

module b17_C_SARLock_k_128_6 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9726,
         n9727, n9729, n9730, n9731, n9732, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088;

  AOI211_X1 U11160 ( .C1(n10756), .C2(n16282), .A(n15068), .B(n15067), .ZN(
        n15069) );
  INV_X1 U11161 ( .A(n17898), .ZN(n17888) );
  XNOR2_X1 U11162 ( .A(n15270), .B(n14370), .ZN(n15258) );
  AND2_X1 U11163 ( .A1(n10364), .A2(n10365), .ZN(n17666) );
  NAND2_X1 U11164 ( .A1(n13954), .A2(n13953), .ZN(n14021) );
  NAND2_X1 U11165 ( .A1(n13765), .A2(n10977), .ZN(n15404) );
  OAI21_X1 U11166 ( .B1(n11236), .B2(n11621), .A(n19175), .ZN(n11007) );
  XNOR2_X1 U11167 ( .A(n10976), .B(n13785), .ZN(n13766) );
  NAND2_X1 U11168 ( .A1(n10975), .A2(n19193), .ZN(n10976) );
  AOI21_X1 U11169 ( .B1(n9940), .B2(n9780), .A(n9857), .ZN(n10933) );
  INV_X1 U11170 ( .A(n13463), .ZN(n14410) );
  INV_X2 U11171 ( .A(n9729), .ZN(n16879) );
  OR2_X1 U11172 ( .A1(n10770), .A2(n10761), .ZN(n19474) );
  AND2_X1 U11173 ( .A1(n13580), .A2(n10750), .ZN(n10943) );
  NAND2_X1 U11174 ( .A1(n10763), .A2(n10762), .ZN(n19711) );
  AND2_X1 U11175 ( .A1(n10756), .A2(n10748), .ZN(n10751) );
  AND2_X2 U11176 ( .A1(n11370), .A2(n11377), .ZN(n11520) );
  NOR2_X1 U11177 ( .A1(n17992), .A2(n17987), .ZN(n17986) );
  AND2_X1 U11178 ( .A1(n16677), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16507) );
  CLKBUF_X2 U11179 ( .A(n10884), .Z(n11375) );
  NOR2_X1 U11180 ( .A1(n16679), .A2(n17634), .ZN(n16677) );
  NOR2_X1 U11181 ( .A1(n17701), .A2(n17702), .ZN(n17673) );
  NOR2_X4 U11182 ( .A1(n10240), .A2(n10234), .ZN(n10331) );
  AND2_X1 U11183 ( .A1(n17786), .A2(n9861), .ZN(n17714) );
  INV_X2 U11184 ( .A(n10253), .ZN(n17185) );
  AND2_X1 U11185 ( .A1(n12429), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10834) );
  NOR3_X2 U11186 ( .A1(n17828), .A2(n17830), .A3(n17810), .ZN(n17786) );
  BUF_X1 U11187 ( .A(n10780), .Z(n12591) );
  NAND2_X2 U11188 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18795) );
  CLKBUF_X2 U11190 ( .A(n11759), .Z(n14221) );
  CLKBUF_X1 U11191 ( .A(n11703), .Z(n14023) );
  CLKBUF_X2 U11192 ( .A(n11948), .Z(n14006) );
  CLKBUF_X2 U11193 ( .A(n11754), .Z(n14105) );
  INV_X2 U11194 ( .A(n12181), .ZN(n12179) );
  INV_X1 U11195 ( .A(n9721), .ZN(n10706) );
  NAND2_X1 U11196 ( .A1(n10662), .A2(n10653), .ZN(n11385) );
  NAND2_X1 U11197 ( .A1(n10652), .A2(n13590), .ZN(n10106) );
  NAND2_X1 U11198 ( .A1(n10047), .A2(n10568), .ZN(n15732) );
  NAND2_X2 U11199 ( .A1(n10231), .A2(n9818), .ZN(n11737) );
  AND2_X2 U11200 ( .A1(n11161), .A2(n10559), .ZN(n10646) );
  BUF_X2 U11201 ( .A(n14265), .Z(n9767) );
  AND2_X1 U11202 ( .A1(n13220), .A2(n13229), .ZN(n11754) );
  CLKBUF_X1 U11203 ( .A(n9757), .Z(n9730) );
  CLKBUF_X2 U11204 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15720) );
  AND2_X1 U11205 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10795) );
  NOR2_X2 U11206 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13592) );
  CLKBUF_X1 U11207 ( .A(n19613), .Z(n9715) );
  AOI22_X1 U11208 ( .A1(n19309), .A2(n15714), .B1(n13655), .B2(n13654), .ZN(
        n19613) );
  NAND2_X1 U11209 ( .A1(n9946), .A2(n9926), .ZN(n9716) );
  NAND2_X1 U11210 ( .A1(n9932), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U11211 ( .A1(n9946), .A2(n9926), .ZN(n15666) );
  NAND2_X1 U11212 ( .A1(n9932), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9727) );
  NOR2_X2 U11213 ( .A1(n13746), .A2(n19414), .ZN(n19886) );
  NAND2_X1 U11214 ( .A1(n15402), .A2(n9794), .ZN(n9718) );
  NAND2_X1 U11215 ( .A1(n15494), .A2(n11112), .ZN(n9719) );
  NAND2_X1 U11216 ( .A1(n15402), .A2(n9794), .ZN(n10209) );
  NAND2_X1 U11217 ( .A1(n15404), .A2(n15403), .ZN(n15402) );
  NAND2_X1 U11218 ( .A1(n15494), .A2(n11112), .ZN(n15304) );
  AND2_X2 U11219 ( .A1(n14621), .A2(n14620), .ZN(n14538) );
  AND2_X1 U11220 ( .A1(n9882), .A2(n13785), .ZN(n9720) );
  XNOR2_X1 U11221 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n10494), .ZN(
        n17987) );
  INV_X1 U11222 ( .A(n10494), .ZN(n17512) );
  NAND2_X1 U11223 ( .A1(n11385), .A2(n10676), .ZN(n9721) );
  AND4_X1 U11225 ( .A1(n10752), .A2(n10754), .A3(n10753), .A4(n10755), .ZN(
        n10775) );
  AND2_X2 U11226 ( .A1(n11675), .A2(n13206), .ZN(n11703) );
  NAND2_X1 U11227 ( .A1(n12880), .A2(n12181), .ZN(n12959) );
  OAI21_X1 U11228 ( .B1(n12911), .B2(n12912), .A(n11891), .ZN(n12003) );
  NAND3_X1 U11229 ( .A1(n10639), .A2(n9928), .A3(n10680), .ZN(n11201) );
  NAND2_X1 U11230 ( .A1(n10733), .A2(n10732), .ZN(n11260) );
  AND2_X1 U11231 ( .A1(n10789), .A2(n12424), .ZN(n10840) );
  AND2_X1 U11232 ( .A1(n12456), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10839) );
  NAND4_X1 U11233 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n12797) );
  XNOR2_X1 U11234 ( .A(n11260), .B(n11259), .ZN(n11261) );
  INV_X1 U11236 ( .A(n14361), .ZN(n11555) );
  INV_X1 U11237 ( .A(n13584), .ZN(n10786) );
  INV_X2 U11238 ( .A(n10404), .ZN(n17202) );
  INV_X2 U11239 ( .A(n17187), .ZN(n10289) );
  NAND2_X1 U11240 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10238) );
  OR2_X1 U11242 ( .A1(n11747), .A2(n11746), .ZN(n12836) );
  INV_X1 U11243 ( .A(n12797), .ZN(n13449) );
  NAND2_X1 U11244 ( .A1(n10181), .A2(n9825), .ZN(n10180) );
  OR2_X1 U11245 ( .A1(n15007), .A2(n15006), .ZN(n15210) );
  NAND3_X2 U11246 ( .A1(n11384), .A2(n11375), .A3(n11377), .ZN(n14361) );
  NAND2_X1 U11247 ( .A1(n11579), .A2(n19387), .ZN(n16479) );
  OR3_X1 U11248 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18795), .ZN(n9813) );
  NAND2_X1 U11249 ( .A1(n18324), .A2(n18218), .ZN(n18279) );
  NAND4_X2 U11250 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n13073) );
  INV_X1 U11251 ( .A(n9736), .ZN(n16241) );
  CLKBUF_X3 U11252 ( .A(n12327), .Z(n9774) );
  INV_X1 U11253 ( .A(n17300), .ZN(n9726) );
  INV_X2 U11254 ( .A(n9814), .ZN(n17205) );
  INV_X2 U11255 ( .A(n17263), .ZN(n10327) );
  XNOR2_X1 U11256 ( .A(n12277), .B(n12276), .ZN(n14553) );
  NAND2_X1 U11257 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17991), .ZN(n17843) );
  AND2_X1 U11258 ( .A1(n11673), .A2(n13220), .ZN(n9757) );
  AND2_X1 U11259 ( .A1(n19431), .A2(n11565), .ZN(n9722) );
  OAI22_X2 U11260 ( .A1(n9787), .A2(n15117), .B1(n15128), .B2(n10177), .ZN(
        n9746) );
  NAND2_X1 U11261 ( .A1(n9882), .A2(n13785), .ZN(n13770) );
  INV_X4 U11262 ( .A(n17313), .ZN(n17334) );
  NAND4_X1 U11263 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n9723) );
  XNOR2_X2 U11264 ( .A(n12011), .B(n13046), .ZN(n13039) );
  INV_X2 U11265 ( .A(n16090), .ZN(n14894) );
  NAND2_X2 U11266 ( .A1(n12001), .A2(n12000), .ZN(n12011) );
  NAND2_X2 U11267 ( .A1(n18944), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10239) );
  NAND2_X2 U11268 ( .A1(n10645), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10105) );
  INV_X1 U11269 ( .A(n10662), .ZN(n10884) );
  NAND2_X2 U11270 ( .A1(n11856), .A2(n11855), .ZN(n11989) );
  NAND2_X2 U11271 ( .A1(n10180), .A2(n10179), .ZN(n13057) );
  AOI21_X4 U11274 ( .B1(n13620), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10673), 
        .ZN(n10674) );
  AND2_X4 U11275 ( .A1(n10789), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9772) );
  AND2_X4 U11276 ( .A1(n10789), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12456) );
  NOR2_X4 U11277 ( .A1(n11377), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11380) );
  INV_X4 U11278 ( .A(n11369), .ZN(n11377) );
  NAND2_X2 U11279 ( .A1(n10712), .A2(n10711), .ZN(n10728) );
  OAI21_X2 U11280 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18976), .A(n16652), 
        .ZN(n17996) );
  AND2_X2 U11281 ( .A1(n10009), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10794) );
  AND2_X4 U11282 ( .A1(n11161), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10781) );
  AND2_X4 U11283 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11161) );
  XNOR2_X2 U11284 ( .A(n12854), .B(n11998), .ZN(n12909) );
  OAI21_X2 U11285 ( .B1(n12912), .B2(n11809), .A(n11997), .ZN(n11998) );
  AND2_X4 U11286 ( .A1(n10796), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10849) );
  AND2_X2 U11288 ( .A1(n11666), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11672) );
  NAND2_X2 U11289 ( .A1(n11239), .A2(n11238), .ZN(n11242) );
  NOR2_X4 U11291 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13229) );
  NOR2_X2 U11292 ( .A1(n17532), .A2(n17401), .ZN(n17397) );
  AND2_X2 U11293 ( .A1(n15343), .A2(n9811), .ZN(n11652) );
  OR2_X1 U11294 ( .A1(n12086), .A2(n14863), .ZN(n14732) );
  AND2_X1 U11295 ( .A1(n16063), .A2(n10135), .ZN(n9777) );
  NAND2_X1 U11296 ( .A1(n13278), .A2(n11221), .ZN(n13373) );
  NAND2_X1 U11297 ( .A1(n13280), .A2(n13279), .ZN(n13278) );
  NOR2_X1 U11298 ( .A1(n15596), .A2(n9856), .ZN(n15525) );
  BUF_X2 U11299 ( .A(n17985), .Z(n9775) );
  CLKBUF_X2 U11300 ( .A(n20266), .Z(n9769) );
  OR2_X1 U11301 ( .A1(n9816), .A2(n14596), .ZN(n14598) );
  NAND2_X1 U11302 ( .A1(n15673), .A2(n15674), .ZN(n15659) );
  XNOR2_X1 U11303 ( .A(n12002), .B(n12003), .ZN(n20266) );
  OR2_X1 U11304 ( .A1(n18776), .A2(n18832), .ZN(n16652) );
  AND2_X1 U11305 ( .A1(n11053), .A2(n11048), .ZN(n11055) );
  CLKBUF_X2 U11306 ( .A(n12318), .Z(n16438) );
  XNOR2_X1 U11307 ( .A(n11919), .B(n11918), .ZN(n12002) );
  NOR2_X1 U11308 ( .A1(n13981), .A2(n13982), .ZN(n14621) );
  NAND2_X1 U11309 ( .A1(n11861), .A2(n9826), .ZN(n11891) );
  OAI21_X1 U11310 ( .B1(n12767), .B2(n12335), .A(n12325), .ZN(n15705) );
  AND2_X1 U11312 ( .A1(n10153), .A2(n9832), .ZN(n17936) );
  OR2_X1 U11313 ( .A1(n11630), .A2(n13269), .ZN(n10733) );
  INV_X1 U11314 ( .A(n10719), .ZN(n11630) );
  NOR2_X1 U11315 ( .A1(n13095), .A2(n13094), .ZN(n13111) );
  CLKBUF_X3 U11316 ( .A(n11278), .Z(n11357) );
  INV_X1 U11317 ( .A(n16865), .ZN(n9729) );
  AND2_X2 U11318 ( .A1(n11574), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11278) );
  BUF_X2 U11319 ( .A(n10720), .Z(n11627) );
  AND3_X1 U11320 ( .A1(n9913), .A2(n9908), .A3(n9914), .ZN(n12170) );
  AND3_X1 U11321 ( .A1(n11716), .A2(n11715), .A3(n9732), .ZN(n9908) );
  NAND2_X4 U11322 ( .A1(n13144), .A2(n12797), .ZN(n12205) );
  NAND2_X1 U11323 ( .A1(n10776), .A2(n20077), .ZN(n10893) );
  NAND2_X1 U11324 ( .A1(n13671), .A2(n12129), .ZN(n11804) );
  NAND2_X2 U11325 ( .A1(n13073), .A2(n11737), .ZN(n11797) );
  INV_X1 U11326 ( .A(n12863), .ZN(n13158) );
  INV_X2 U11327 ( .A(n20077), .ZN(n13746) );
  CLKBUF_X2 U11328 ( .A(n10656), .Z(n12312) );
  NAND2_X1 U11329 ( .A1(n10638), .A2(n10637), .ZN(n10676) );
  INV_X2 U11330 ( .A(n10288), .ZN(n9734) );
  INV_X2 U11331 ( .A(n17322), .ZN(n17237) );
  AND4_X1 U11332 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .ZN(
        n10632) );
  INV_X4 U11333 ( .A(n17204), .ZN(n15818) );
  INV_X1 U11334 ( .A(n10330), .ZN(n10288) );
  INV_X4 U11335 ( .A(n17275), .ZN(n10286) );
  INV_X1 U11336 ( .A(n10265), .ZN(n17322) );
  BUF_X2 U11337 ( .A(n11840), .Z(n14313) );
  CLKBUF_X2 U11338 ( .A(n11934), .Z(n14308) );
  CLKBUF_X2 U11339 ( .A(n11777), .Z(n14284) );
  CLKBUF_X2 U11340 ( .A(n14056), .Z(n14192) );
  INV_X4 U11341 ( .A(n9813), .ZN(n17306) );
  AND2_X1 U11342 ( .A1(n11673), .A2(n11675), .ZN(n11840) );
  AND2_X2 U11343 ( .A1(n13220), .A2(n13206), .ZN(n14265) );
  CLKBUF_X1 U11344 ( .A(n10647), .Z(n9738) );
  INV_X2 U11345 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13602) );
  NAND3_X4 U11346 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15854) );
  NOR2_X1 U11347 ( .A1(n10115), .A2(n10002), .ZN(n10001) );
  NOR2_X1 U11348 ( .A1(n15483), .A2(n9923), .ZN(n16359) );
  NOR2_X1 U11349 ( .A1(n15570), .A2(n10193), .ZN(n15590) );
  AND2_X1 U11350 ( .A1(n15484), .A2(n15486), .ZN(n9923) );
  NAND2_X1 U11351 ( .A1(n14757), .A2(n14773), .ZN(n14766) );
  XNOR2_X1 U11352 ( .A(n11647), .B(n11645), .ZN(n15277) );
  AOI21_X1 U11353 ( .B1(n9855), .B2(n14430), .A(n14429), .ZN(n14738) );
  XNOR2_X1 U11354 ( .A(n14334), .B(n14333), .ZN(n14384) );
  OR2_X1 U11355 ( .A1(n15351), .A2(n15352), .ZN(n10036) );
  AOI211_X1 U11356 ( .C1(n15428), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        n15429) );
  NAND2_X1 U11357 ( .A1(n9919), .A2(n10129), .ZN(n14800) );
  AND2_X1 U11358 ( .A1(n15328), .A2(n15610), .ZN(n16379) );
  XNOR2_X1 U11359 ( .A(n12523), .B(n10227), .ZN(n15107) );
  NAND2_X1 U11360 ( .A1(n15111), .A2(n12503), .ZN(n12523) );
  NOR2_X1 U11361 ( .A1(n9948), .A2(n11253), .ZN(n9947) );
  NOR3_X1 U11362 ( .A1(n15100), .A2(n15099), .A3(n9865), .ZN(n11626) );
  NOR2_X1 U11363 ( .A1(n15863), .A2(n16528), .ZN(n15923) );
  OR2_X1 U11364 ( .A1(n15023), .A2(n15005), .ZN(n15100) );
  XNOR2_X1 U11365 ( .A(n11007), .B(n11604), .ZN(n15403) );
  AND2_X1 U11366 ( .A1(n12062), .A2(n9824), .ZN(n9782) );
  NAND3_X1 U11367 ( .A1(n13770), .A2(n11229), .A3(n11228), .ZN(n13768) );
  INV_X1 U11368 ( .A(n18004), .ZN(n17637) );
  NOR2_X1 U11369 ( .A1(n14812), .A2(n12071), .ZN(n12072) );
  NAND2_X1 U11370 ( .A1(n15146), .A2(n12413), .ZN(n15140) );
  AOI211_X1 U11371 ( .C1(n14849), .C2(n9897), .A(n9896), .B(n9895), .ZN(n9894)
         );
  AND2_X2 U11372 ( .A1(n13835), .A2(n12402), .ZN(n15146) );
  NAND2_X1 U11373 ( .A1(n13255), .A2(n13254), .ZN(n13514) );
  OR2_X1 U11374 ( .A1(n15039), .A2(n15131), .ZN(n15133) );
  NOR2_X2 U11375 ( .A1(n15183), .A2(n15172), .ZN(n15171) );
  AND2_X1 U11376 ( .A1(n13088), .A2(n13089), .ZN(n13109) );
  NAND2_X2 U11377 ( .A1(n12055), .A2(n11983), .ZN(n16090) );
  NAND2_X1 U11378 ( .A1(n11980), .A2(n11979), .ZN(n12055) );
  NOR2_X1 U11379 ( .A1(n18143), .A2(n17819), .ZN(n17804) );
  INV_X1 U11380 ( .A(n17996), .ZN(n17941) );
  NAND2_X1 U11381 ( .A1(n11004), .A2(n11003), .ZN(n11240) );
  NAND2_X1 U11382 ( .A1(n12022), .A2(n12014), .ZN(n20268) );
  NOR2_X1 U11383 ( .A1(n13060), .A2(n10116), .ZN(n13421) );
  NAND2_X1 U11384 ( .A1(n16447), .A2(n15597), .ZN(n15596) );
  OAI22_X1 U11385 ( .A1(n19711), .A2(n10766), .B1(n19640), .B2(n10765), .ZN(
        n10767) );
  NOR2_X1 U11386 ( .A1(n15659), .A2(n10082), .ZN(n16447) );
  NOR2_X1 U11387 ( .A1(n13055), .A2(n13054), .ZN(n13062) );
  OAI21_X1 U11388 ( .B1(n12823), .B2(n12822), .A(n12341), .ZN(n12826) );
  NAND2_X1 U11389 ( .A1(n10763), .A2(n10222), .ZN(n19640) );
  OR2_X1 U11390 ( .A1(n11078), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11079) );
  AND2_X1 U11391 ( .A1(n16438), .A2(n10746), .ZN(n19506) );
  AND2_X1 U11392 ( .A1(n16438), .A2(n10750), .ZN(n19441) );
  INV_X2 U11393 ( .A(n16044), .ZN(n9731) );
  AND2_X1 U11394 ( .A1(n13124), .A2(n12021), .ZN(n10147) );
  OR2_X1 U11395 ( .A1(n11262), .A2(n11261), .ZN(n10108) );
  INV_X2 U11396 ( .A(n19317), .ZN(n19362) );
  NOR2_X2 U11397 ( .A1(n14724), .A2(n13074), .ZN(n13075) );
  NAND2_X1 U11398 ( .A1(n11942), .A2(n11941), .ZN(n13124) );
  NAND2_X1 U11399 ( .A1(n10515), .A2(n17921), .ZN(n17915) );
  NAND2_X1 U11400 ( .A1(n11891), .A2(n11875), .ZN(n12911) );
  NAND2_X1 U11401 ( .A1(n12855), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12854) );
  NAND2_X1 U11402 ( .A1(n11125), .A2(n11038), .ZN(n11036) );
  NAND2_X1 U11403 ( .A1(n12329), .A2(n12328), .ZN(n12793) );
  NAND2_X2 U11404 ( .A1(n13071), .A2(n14413), .ZN(n14724) );
  OR2_X1 U11405 ( .A1(n16219), .A2(n13863), .ZN(n13981) );
  INV_X2 U11406 ( .A(n15159), .ZN(n12766) );
  AND2_X1 U11407 ( .A1(n10745), .A2(n19231), .ZN(n10748) );
  INV_X2 U11408 ( .A(n17366), .ZN(n17355) );
  OR2_X1 U11409 ( .A1(n13070), .A2(n13069), .ZN(n13071) );
  XNOR2_X1 U11410 ( .A(n15705), .B(n12330), .ZN(n12794) );
  OAI21_X1 U11411 ( .B1(n12848), .B2(n12115), .A(n11992), .ZN(n12855) );
  NAND2_X1 U11412 ( .A1(n11989), .A2(n11990), .ZN(n11861) );
  AND2_X1 U11413 ( .A1(n10724), .A2(n10723), .ZN(n10738) );
  AOI21_X1 U11414 ( .B1(n18250), .B2(n17947), .A(n10511), .ZN(n17933) );
  OR2_X1 U11415 ( .A1(n17954), .A2(n17955), .ZN(n10153) );
  NAND2_X1 U11416 ( .A1(n11125), .A2(n11020), .ZN(n11024) );
  AND2_X1 U11417 ( .A1(n11882), .A2(n11881), .ZN(n11885) );
  NAND2_X1 U11418 ( .A1(n10737), .A2(n10736), .ZN(n11259) );
  OR2_X1 U11419 ( .A1(n11019), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11020) );
  AOI21_X1 U11420 ( .B1(n11897), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11898), .ZN(n11903) );
  CLKBUF_X1 U11421 ( .A(n11896), .Z(n11897) );
  AND2_X1 U11422 ( .A1(n10731), .A2(n10730), .ZN(n10732) );
  AOI22_X1 U11423 ( .A1(n10698), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n10735), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10699) );
  AND2_X1 U11424 ( .A1(n10722), .A2(n10721), .ZN(n10723) );
  OR2_X1 U11425 ( .A1(n13035), .A2(n13034), .ZN(n13095) );
  AND2_X1 U11426 ( .A1(n10705), .A2(n10704), .ZN(n10710) );
  AND2_X1 U11427 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  NOR4_X2 U11428 ( .A1(n18319), .A2(n10527), .A3(n17377), .A4(n10533), .ZN(
        n17580) );
  NAND2_X1 U11429 ( .A1(n11827), .A2(n11826), .ZN(n11881) );
  NAND2_X1 U11430 ( .A1(n12979), .A2(n13463), .ZN(n13455) );
  INV_X1 U11431 ( .A(n11278), .ZN(n11263) );
  AOI211_X2 U11432 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n10382), .B(n10381), .ZN(n18335) );
  NOR2_X1 U11433 ( .A1(n10684), .A2(n9930), .ZN(n9929) );
  NAND2_X1 U11434 ( .A1(n12775), .A2(n10671), .ZN(n10677) );
  NAND2_X1 U11435 ( .A1(n18319), .A2(n18970), .ZN(n10529) );
  AOI211_X1 U11436 ( .C1(n10327), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n10313), .B(n10312), .ZN(n17495) );
  AOI211_X2 U11437 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n10392), .B(n10391), .ZN(n18341) );
  CLKBUF_X1 U11438 ( .A(n18347), .Z(n9752) );
  NOR2_X1 U11439 ( .A1(n9912), .A2(n11798), .ZN(n9911) );
  OR2_X1 U11440 ( .A1(n11804), .A2(n11805), .ZN(n14944) );
  AND2_X1 U11441 ( .A1(n13158), .A2(n12836), .ZN(n11800) );
  INV_X1 U11442 ( .A(n12790), .ZN(n19431) );
  AND2_X1 U11443 ( .A1(n10605), .A2(n10669), .ZN(n10198) );
  OR2_X1 U11444 ( .A1(n10860), .A2(n10859), .ZN(n11390) );
  AND4_X1 U11445 ( .A1(n10283), .A2(n10217), .A3(n10158), .A4(n10284), .ZN(
        n17507) );
  AND2_X2 U11446 ( .A1(n9723), .A2(n12180), .ZN(n13463) );
  INV_X1 U11447 ( .A(n10657), .ZN(n12790) );
  INV_X1 U11448 ( .A(n12180), .ZN(n11809) );
  INV_X2 U11449 ( .A(U212), .ZN(n16600) );
  INV_X2 U11450 ( .A(n16601), .ZN(n16605) );
  INV_X1 U11451 ( .A(n11737), .ZN(n13671) );
  NAND3_X1 U11452 ( .A1(n17714), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17701) );
  NAND2_X2 U11453 ( .A1(n11699), .A2(n11698), .ZN(n12129) );
  INV_X1 U11454 ( .A(n12180), .ZN(n9732) );
  NAND2_X2 U11455 ( .A1(n10617), .A2(n10616), .ZN(n10668) );
  NAND3_X1 U11456 ( .A1(n10615), .A2(n10614), .A3(n10613), .ZN(n10616) );
  NAND4_X1 U11457 ( .A1(n9836), .A2(n10556), .A3(n10555), .A4(n9792), .ZN(
        n10047) );
  CLKBUF_X1 U11458 ( .A(n17322), .Z(n9771) );
  NAND2_X1 U11459 ( .A1(n10610), .A2(n13590), .ZN(n10617) );
  AND4_X1 U11460 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11734) );
  AND4_X1 U11461 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11736) );
  AND4_X1 U11462 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n11770) );
  AND4_X1 U11463 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11794) );
  AND4_X1 U11464 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11771) );
  AND4_X1 U11465 ( .A1(n11697), .A2(n11696), .A3(n11695), .A4(n11694), .ZN(
        n11698) );
  AND4_X1 U11466 ( .A1(n11693), .A2(n11692), .A3(n11691), .A4(n11690), .ZN(
        n11699) );
  AND4_X1 U11467 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n11792) );
  AND4_X1 U11468 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11733) );
  NAND2_X2 U11469 ( .A1(n18983), .A2(n18857), .ZN(n18908) );
  INV_X2 U11470 ( .A(n16638), .ZN(U215) );
  INV_X2 U11471 ( .A(n15789), .ZN(n17327) );
  AND4_X1 U11472 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11791) );
  AND4_X1 U11473 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n11735) );
  AND4_X1 U11474 ( .A1(n11709), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n11714) );
  AND4_X1 U11475 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11793) );
  NAND2_X2 U11476 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20088), .ZN(n20017) );
  AND4_X1 U11477 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10610) );
  INV_X2 U11478 ( .A(n20717), .ZN(n9735) );
  AND4_X1 U11479 ( .A1(n11767), .A2(n11766), .A3(n11765), .A4(n11764), .ZN(
        n11768) );
  AND4_X1 U11480 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n11769) );
  CLKBUF_X2 U11481 ( .A(n17563), .Z(n18980) );
  INV_X2 U11482 ( .A(n10329), .ZN(n15789) );
  INV_X1 U11483 ( .A(n10242), .ZN(n10243) );
  NAND2_X2 U11484 ( .A1(n18933), .A2(n10242), .ZN(n17263) );
  BUF_X4 U11485 ( .A(n14265), .Z(n9768) );
  AND2_X1 U11486 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  AND3_X1 U11487 ( .A1(n10563), .A2(n10562), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10567) );
  OR2_X1 U11488 ( .A1(n17027), .A2(n10240), .ZN(n17300) );
  INV_X2 U11489 ( .A(n20177), .ZN(n9736) );
  INV_X2 U11490 ( .A(n10256), .ZN(n17326) );
  INV_X2 U11491 ( .A(n18984), .ZN(n18983) );
  OR2_X2 U11492 ( .A1(n20089), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20020) );
  INV_X2 U11493 ( .A(n20089), .ZN(n20088) );
  INV_X2 U11494 ( .A(n16642), .ZN(n9737) );
  OR2_X2 U11495 ( .A1(n17027), .A2(n10241), .ZN(n10253) );
  AND2_X2 U11496 ( .A1(n13592), .A2(n10559), .ZN(n10778) );
  INV_X1 U11497 ( .A(n17967), .ZN(n9964) );
  OR2_X2 U11498 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15854), .ZN(
        n10404) );
  NAND2_X1 U11499 ( .A1(n18933), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10240) );
  NAND2_X1 U11500 ( .A1(n20969), .A2(n18951), .ZN(n17027) );
  AND2_X2 U11501 ( .A1(n9985), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13220) );
  NOR2_X2 U11502 ( .A1(n9985), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13217) );
  NAND2_X1 U11503 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11674), .ZN(
        n11667) );
  NOR2_X2 U11504 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11675) );
  NOR2_X2 U11505 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10789) );
  INV_X2 U11506 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12842) );
  NAND2_X1 U11507 ( .A1(n19608), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10807) );
  AND2_X1 U11508 ( .A1(n10367), .A2(n18009), .ZN(n17651) );
  NOR3_X4 U11509 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n17870), .ZN(n17814) );
  NAND2_X1 U11510 ( .A1(n9977), .A2(n9978), .ZN(n17692) );
  NAND2_X1 U11511 ( .A1(n11564), .A2(n9722), .ZN(n10685) );
  NAND2_X1 U11512 ( .A1(n10893), .A2(n10679), .ZN(n11564) );
  OAI21_X1 U11513 ( .B1(n12318), .B2(n12335), .A(n12317), .ZN(n12344) );
  OR2_X1 U11514 ( .A1(n13284), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11890) );
  XNOR2_X1 U11515 ( .A(n14766), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9739) );
  INV_X1 U11516 ( .A(n9739), .ZN(n16122) );
  NOR2_X4 U11517 ( .A1(n14465), .A2(n14467), .ZN(n14451) );
  INV_X1 U11518 ( .A(n9717), .ZN(n10719) );
  NOR2_X2 U11519 ( .A1(n17986), .A2(n10340), .ZN(n17978) );
  NOR2_X2 U11520 ( .A1(n17978), .A2(n17977), .ZN(n17976) );
  NAND3_X1 U11521 ( .A1(n9907), .A2(n12174), .A3(n9906), .ZN(n11799) );
  NAND2_X2 U11522 ( .A1(n10675), .A2(n10674), .ZN(n9740) );
  NAND2_X1 U11523 ( .A1(n10675), .A2(n10674), .ZN(n10725) );
  AOI21_X2 U11524 ( .B1(n15393), .B2(n9947), .A(n9830), .ZN(n9946) );
  MUX2_X1 U11525 ( .A(n10662), .B(n15732), .S(n10653), .Z(n10660) );
  NAND2_X1 U11526 ( .A1(n15624), .A2(n15327), .ZN(n9741) );
  AND2_X1 U11527 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U11528 ( .A1(n15624), .A2(n15327), .ZN(n11042) );
  INV_X1 U11529 ( .A(n12349), .ZN(n9743) );
  AND2_X1 U11530 ( .A1(n9744), .A2(n13116), .ZN(n13835) );
  NOR2_X1 U11531 ( .A1(n10186), .A2(n9743), .ZN(n9744) );
  BUF_X1 U11532 ( .A(n12547), .Z(n9745) );
  NOR2_X1 U11533 ( .A1(n12544), .A2(n12543), .ZN(n12547) );
  OR2_X2 U11534 ( .A1(n15304), .A2(n15306), .ZN(n9747) );
  AND2_X2 U11535 ( .A1(n10937), .A2(n9881), .ZN(n9748) );
  INV_X1 U11536 ( .A(n9748), .ZN(n11222) );
  AND2_X1 U11537 ( .A1(n13206), .A2(n11674), .ZN(n9749) );
  AND2_X1 U11538 ( .A1(n13206), .A2(n11674), .ZN(n9750) );
  INV_X1 U11539 ( .A(n9750), .ZN(n9751) );
  AND2_X1 U11540 ( .A1(n19421), .A2(n10668), .ZN(n9928) );
  AND2_X1 U11541 ( .A1(n13592), .A2(n10559), .ZN(n9753) );
  NOR2_X2 U11542 ( .A1(n15107), .A2(n15106), .ZN(n15105) );
  NOR3_X2 U11543 ( .A1(n17450), .A2(n17416), .A3(n17373), .ZN(n17412) );
  AND2_X1 U11544 ( .A1(n13592), .A2(n10559), .ZN(n9754) );
  AND2_X1 U11545 ( .A1(n12544), .A2(n12543), .ZN(n12545) );
  OAI211_X1 U11546 ( .C1(n10660), .C2(n10659), .A(n10665), .B(n13746), .ZN(
        n11569) );
  AND2_X2 U11547 ( .A1(n15637), .A2(n9808), .ZN(n16375) );
  NOR2_X4 U11548 ( .A1(n9925), .A2(n15638), .ZN(n15637) );
  NOR2_X4 U11549 ( .A1(n13514), .A2(n13562), .ZN(n13522) );
  AND2_X2 U11550 ( .A1(n13580), .A2(n10751), .ZN(n10942) );
  AND2_X2 U11551 ( .A1(n16438), .A2(n10751), .ZN(n10941) );
  OR2_X1 U11552 ( .A1(n11241), .A2(n11240), .ZN(n11246) );
  OAI21_X2 U11553 ( .B1(n16375), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15591), .ZN(n16369) );
  NOR2_X4 U11554 ( .A1(n15140), .A2(n15134), .ZN(n12455) );
  NAND2_X2 U11555 ( .A1(n10209), .A2(n9862), .ZN(n15624) );
  INV_X2 U11556 ( .A(n13891), .ZN(n12073) );
  NAND2_X1 U11557 ( .A1(n10726), .A2(n10744), .ZN(n12767) );
  XNOR2_X2 U11558 ( .A(n12455), .B(n12478), .ZN(n15128) );
  OR2_X2 U11559 ( .A1(n10770), .A2(n10769), .ZN(n10771) );
  NOR2_X2 U11560 ( .A1(n10234), .A2(n10239), .ZN(n10330) );
  AND2_X1 U11561 ( .A1(n11672), .A2(n13220), .ZN(n9755) );
  AND2_X1 U11562 ( .A1(n11672), .A2(n13220), .ZN(n9756) );
  AND2_X1 U11563 ( .A1(n11672), .A2(n13220), .ZN(n11948) );
  AND3_X4 U11564 ( .A1(n13602), .A2(n10009), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10647) );
  NAND2_X2 U11565 ( .A1(n11799), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U11566 ( .A1(n10592), .A2(n10591), .ZN(n10657) );
  INV_X2 U11567 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10559) );
  AND2_X1 U11568 ( .A1(n11673), .A2(n13220), .ZN(n9758) );
  CLKBUF_X1 U11569 ( .A(n11833), .Z(n9759) );
  CLKBUF_X1 U11570 ( .A(n11833), .Z(n9760) );
  CLKBUF_X1 U11571 ( .A(n11833), .Z(n9761) );
  AND2_X1 U11574 ( .A1(n11673), .A2(n13220), .ZN(n11833) );
  AND2_X2 U11575 ( .A1(n10559), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10788) );
  NAND4_X1 U11576 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n9765) );
  NAND4_X1 U11577 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n9766) );
  AND2_X1 U11578 ( .A1(n15343), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15314) );
  AND2_X4 U11579 ( .A1(n15359), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15343) );
  NAND2_X2 U11580 ( .A1(n15493), .A2(n15492), .ZN(n15494) );
  NAND2_X1 U11581 ( .A1(n12339), .A2(n12338), .ZN(n12341) );
  AND2_X2 U11582 ( .A1(n11652), .A2(n10213), .ZN(n15270) );
  OAI21_X1 U11583 ( .B1(n10708), .B2(n11560), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10709) );
  NAND2_X2 U11584 ( .A1(n13880), .A2(n12065), .ZN(n14833) );
  OAI21_X2 U11585 ( .B1(n13816), .B2(n12063), .A(n12064), .ZN(n13880) );
  AND2_X2 U11586 ( .A1(n13580), .A2(n10749), .ZN(n10944) );
  INV_X1 U11587 ( .A(n11278), .ZN(n9770) );
  AND2_X2 U11588 ( .A1(n12318), .A2(n10749), .ZN(n19608) );
  OAI21_X1 U11589 ( .B1(n12336), .B2(n12335), .A(n12334), .ZN(n12339) );
  NAND2_X2 U11590 ( .A1(n12758), .A2(n12637), .ZN(n11366) );
  NAND2_X1 U11591 ( .A1(n13116), .A2(n12349), .ZN(n13200) );
  NOR2_X4 U11592 ( .A1(n13057), .A2(n12348), .ZN(n13116) );
  NOR2_X2 U11593 ( .A1(n9746), .A2(n12479), .ZN(n12500) );
  XNOR2_X1 U11594 ( .A(n10726), .B(n10758), .ZN(n12327) );
  BUF_X4 U11595 ( .A(n12336), .Z(n10769) );
  XNOR2_X2 U11596 ( .A(n10739), .B(n10738), .ZN(n12336) );
  NAND2_X1 U11597 ( .A1(n10707), .A2(n9790), .ZN(n10020) );
  NOR2_X1 U11598 ( .A1(n14894), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10136) );
  NOR2_X1 U11599 ( .A1(n10131), .A2(n9921), .ZN(n9920) );
  INV_X1 U11600 ( .A(n12072), .ZN(n9921) );
  NAND2_X1 U11601 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  INV_X1 U11602 ( .A(n12309), .ZN(n10132) );
  INV_X1 U11603 ( .A(n14732), .ZN(n9996) );
  NAND2_X1 U11604 ( .A1(n15211), .A2(n10088), .ZN(n14363) );
  AND2_X1 U11605 ( .A1(n10090), .A2(n10089), .ZN(n10088) );
  INV_X1 U11606 ( .A(n11558), .ZN(n10089) );
  AND2_X1 U11607 ( .A1(n11211), .A2(n19304), .ZN(n11578) );
  NAND2_X1 U11608 ( .A1(n11968), .A2(n11967), .ZN(n12044) );
  INV_X1 U11609 ( .A(n12032), .ZN(n11967) );
  NAND2_X1 U11610 ( .A1(n11815), .A2(n11814), .ZN(n11882) );
  NAND2_X1 U11611 ( .A1(n11803), .A2(n11821), .ZN(n12161) );
  NOR2_X1 U11612 ( .A1(n10908), .A2(n10907), .ZN(n10926) );
  NAND2_X1 U11613 ( .A1(n10890), .A2(n10889), .ZN(n10922) );
  AND2_X1 U11614 ( .A1(n14587), .A2(n14088), .ZN(n14578) );
  OR2_X1 U11615 ( .A1(n13073), .A2(n12842), .ZN(n14294) );
  INV_X1 U11616 ( .A(n14733), .ZN(n9989) );
  AND2_X1 U11617 ( .A1(n9777), .A2(n9878), .ZN(n9998) );
  INV_X1 U11618 ( .A(n14808), .ZN(n10134) );
  INV_X1 U11619 ( .A(n12057), .ZN(n11981) );
  NAND2_X1 U11620 ( .A1(n13463), .A2(n12179), .ZN(n12265) );
  OR2_X1 U11621 ( .A1(n11982), .A2(n11981), .ZN(n11860) );
  OR2_X1 U11622 ( .A1(n11050), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U11623 ( .A1(n11369), .A2(n12319), .ZN(n12518) );
  INV_X1 U11624 ( .A(n15150), .ZN(n10121) );
  AND2_X1 U11625 ( .A1(n15592), .A2(n16382), .ZN(n10058) );
  NAND2_X1 U11626 ( .A1(n10706), .A2(n13746), .ZN(n10654) );
  AND2_X1 U11627 ( .A1(n10201), .A2(n10005), .ZN(n9945) );
  INV_X1 U11628 ( .A(n11608), .ZN(n10005) );
  INV_X1 U11629 ( .A(n13607), .ZN(n12742) );
  AND2_X1 U11630 ( .A1(n12781), .A2(n12782), .ZN(n12780) );
  AND2_X1 U11631 ( .A1(n19431), .A2(n20037), .ZN(n11384) );
  AND2_X1 U11632 ( .A1(n10662), .A2(n20037), .ZN(n11370) );
  OR2_X1 U11633 ( .A1(n12780), .A2(n11389), .ZN(n11395) );
  AND2_X2 U11634 ( .A1(n10668), .A2(n10667), .ZN(n11566) );
  MUX2_X1 U11635 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11188), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11191) );
  NAND2_X1 U11636 ( .A1(n10157), .A2(n17897), .ZN(n9977) );
  AND2_X1 U11637 ( .A1(n13507), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13516) );
  NOR2_X1 U11638 ( .A1(n14894), .A2(n14856), .ZN(n9995) );
  NAND2_X1 U11639 ( .A1(n14756), .A2(n14773), .ZN(n9922) );
  AND2_X1 U11640 ( .A1(n12169), .A2(n14413), .ZN(n12299) );
  NAND2_X1 U11641 ( .A1(n12168), .A2(n9899), .ZN(n12169) );
  AOI211_X1 U11642 ( .C1(n15907), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9899)
         );
  AND2_X1 U11643 ( .A1(n11125), .A2(n11642), .ZN(n11620) );
  INV_X1 U11644 ( .A(n10058), .ZN(n10057) );
  NOR2_X1 U11645 ( .A1(n9822), .A2(n11614), .ZN(n11615) );
  INV_X1 U11646 ( .A(n15266), .ZN(n11614) );
  NAND2_X1 U11647 ( .A1(n10199), .A2(n10200), .ZN(n11647) );
  AOI21_X1 U11648 ( .B1(n10201), .B2(n15306), .A(n9829), .ZN(n10200) );
  CLKBUF_X1 U11649 ( .A(n11369), .Z(n13331) );
  NAND2_X1 U11650 ( .A1(n17650), .A2(n10225), .ZN(n15863) );
  AND2_X1 U11651 ( .A1(n17679), .A2(n9869), .ZN(n10152) );
  NAND2_X1 U11652 ( .A1(n14398), .A2(n14399), .ZN(n20745) );
  AND2_X1 U11653 ( .A1(n14369), .A2(n14368), .ZN(n14371) );
  NAND2_X1 U11654 ( .A1(n15590), .A2(n10192), .ZN(n10191) );
  NAND2_X1 U11655 ( .A1(n16479), .A2(n15589), .ZN(n10192) );
  AND2_X1 U11656 ( .A1(n11825), .A2(n11824), .ZN(n11826) );
  NAND2_X1 U11657 ( .A1(n9911), .A2(n12862), .ZN(n9906) );
  AOI22_X1 U11658 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U11659 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U11660 ( .A1(n9951), .A2(n10664), .ZN(n10707) );
  NAND2_X1 U11661 ( .A1(n11374), .A2(n11373), .ZN(n12781) );
  NAND2_X1 U11662 ( .A1(n10663), .A2(n11199), .ZN(n11561) );
  AND2_X1 U11663 ( .A1(n11193), .A2(n19431), .ZN(n10663) );
  NAND2_X1 U11664 ( .A1(n12773), .A2(n10667), .ZN(n10664) );
  AND2_X1 U11665 ( .A1(n15732), .A2(n10662), .ZN(n10605) );
  NAND2_X1 U11666 ( .A1(n10343), .A2(n10492), .ZN(n10324) );
  AOI21_X1 U11667 ( .B1(n18809), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10466), .ZN(n10475) );
  NOR2_X1 U11668 ( .A1(n11857), .A2(n12129), .ZN(n12837) );
  NOR2_X1 U11669 ( .A1(n9855), .A2(n10150), .ZN(n10149) );
  NAND2_X1 U11670 ( .A1(n10151), .A2(n14258), .ZN(n10150) );
  INV_X1 U11671 ( .A(n14440), .ZN(n10151) );
  INV_X1 U11672 ( .A(n14453), .ZN(n14258) );
  AND2_X1 U11673 ( .A1(n10139), .A2(n14482), .ZN(n10138) );
  OR2_X1 U11674 ( .A1(n10144), .A2(n14593), .ZN(n10143) );
  NAND2_X1 U11675 ( .A1(n14022), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14297) );
  AND2_X1 U11676 ( .A1(n9802), .A2(n13861), .ZN(n10137) );
  INV_X1 U11677 ( .A(n13862), .ZN(n13861) );
  AND2_X1 U11678 ( .A1(n12044), .A2(n12034), .ZN(n13253) );
  NOR2_X1 U11679 ( .A1(n16090), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9993) );
  NAND2_X1 U11680 ( .A1(n14800), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12081) );
  INV_X1 U11681 ( .A(n10136), .ZN(n10000) );
  NOR2_X1 U11682 ( .A1(n10071), .A2(n14613), .ZN(n10070) );
  INV_X1 U11683 ( .A(n10072), .ZN(n10071) );
  NOR2_X1 U11684 ( .A1(n13898), .A2(n10073), .ZN(n10072) );
  INV_X1 U11685 ( .A(n14539), .ZN(n10073) );
  INV_X1 U11686 ( .A(n16105), .ZN(n9918) );
  XNOR2_X1 U11687 ( .A(n12055), .B(n12054), .ZN(n13515) );
  NAND2_X1 U11688 ( .A1(n12181), .A2(n13463), .ZN(n12243) );
  AND2_X1 U11689 ( .A1(n12284), .A2(n12283), .ZN(n12294) );
  INV_X1 U11690 ( .A(n12305), .ZN(n12297) );
  INV_X1 U11691 ( .A(n11874), .ZN(n10127) );
  NAND2_X1 U11692 ( .A1(n11819), .A2(n11796), .ZN(n12960) );
  INV_X1 U11693 ( .A(n12848), .ZN(n13395) );
  NOR2_X1 U11694 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13135), .ZN(n13393) );
  NAND2_X1 U11695 ( .A1(n20271), .A2(n11886), .ZN(n11942) );
  NAND2_X1 U11696 ( .A1(n12129), .A2(n12180), .ZN(n12115) );
  NAND3_X1 U11697 ( .A1(n11857), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n9766), 
        .ZN(n12116) );
  OR2_X1 U11698 ( .A1(n9765), .A2(n11886), .ZN(n11928) );
  NAND2_X1 U11699 ( .A1(n13679), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11982) );
  NOR2_X1 U11700 ( .A1(n11644), .A2(n11136), .ZN(n11137) );
  NOR2_X1 U11701 ( .A1(n10015), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10014) );
  INV_X1 U11702 ( .A(n10016), .ZN(n10015) );
  OR2_X1 U11703 ( .A1(n9815), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11064) );
  NOR2_X1 U11704 ( .A1(n10011), .A2(n11009), .ZN(n10010) );
  INV_X1 U11705 ( .A(n11005), .ZN(n10011) );
  OR2_X1 U11706 ( .A1(n10924), .A2(n10801), .ZN(n10006) );
  AND2_X1 U11707 ( .A1(n12478), .A2(n12477), .ZN(n12479) );
  INV_X1 U11708 ( .A(n15158), .ZN(n10122) );
  AND2_X1 U11709 ( .A1(n10104), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10102) );
  NOR2_X1 U11710 ( .A1(n16432), .A2(n10101), .ZN(n10104) );
  NOR2_X1 U11711 ( .A1(n15287), .A2(n15296), .ZN(n11130) );
  OR2_X1 U11712 ( .A1(n15017), .A2(n9870), .ZN(n11134) );
  OR2_X1 U11713 ( .A1(n16322), .A2(n11023), .ZN(n11120) );
  AND2_X1 U11714 ( .A1(n10203), .A2(n9937), .ZN(n9936) );
  NAND2_X1 U11715 ( .A1(n11093), .A2(n9938), .ZN(n9937) );
  AOI21_X1 U11716 ( .B1(n10205), .B2(n11093), .A(n10204), .ZN(n10203) );
  INV_X1 U11717 ( .A(n15319), .ZN(n10204) );
  INV_X1 U11718 ( .A(n11093), .ZN(n9939) );
  OR2_X1 U11719 ( .A1(n11100), .A2(n15529), .ZN(n15334) );
  AND4_X1 U11720 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10878) );
  NAND2_X1 U11721 ( .A1(n10087), .A2(n13838), .ZN(n10086) );
  INV_X1 U11722 ( .A(n15579), .ZN(n10087) );
  INV_X1 U11723 ( .A(n15647), .ZN(n10085) );
  NAND2_X1 U11724 ( .A1(n11235), .A2(n11237), .ZN(n11238) );
  NOR2_X1 U11725 ( .A1(n11002), .A2(n11001), .ZN(n11410) );
  INV_X1 U11726 ( .A(n11230), .ZN(n9882) );
  INV_X1 U11727 ( .A(n11259), .ZN(n10112) );
  INV_X1 U11728 ( .A(n11260), .ZN(n10113) );
  OR2_X1 U11729 ( .A1(n10847), .A2(n10846), .ZN(n11386) );
  OR2_X1 U11730 ( .A1(n11400), .A2(n11396), .ZN(n12928) );
  NAND2_X1 U11731 ( .A1(n10757), .A2(n10756), .ZN(n10019) );
  AOI21_X1 U11732 ( .B1(n11156), .B2(n11155), .A(n11154), .ZN(n11186) );
  AND2_X1 U11733 ( .A1(n15937), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11154) );
  AOI21_X1 U11734 ( .B1(n17323), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n10162), .ZN(n10161) );
  AND2_X1 U11735 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10162) );
  NAND2_X1 U11736 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10160) );
  NOR2_X1 U11737 ( .A1(n9983), .A2(n20969), .ZN(n10242) );
  NAND2_X1 U11738 ( .A1(n18951), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9983) );
  NOR2_X1 U11739 ( .A1(n10529), .A2(n10528), .ZN(n15845) );
  INV_X1 U11740 ( .A(n17993), .ZN(n10493) );
  NAND2_X1 U11741 ( .A1(n18335), .A2(n18330), .ZN(n18783) );
  INV_X1 U11742 ( .A(n16650), .ZN(n10528) );
  NOR2_X1 U11743 ( .A1(n15740), .A2(n15739), .ZN(n15847) );
  OR3_X1 U11744 ( .A1(n10067), .A2(n12267), .A3(n14442), .ZN(n10066) );
  OR2_X1 U11745 ( .A1(n13207), .A2(n14408), .ZN(n12868) );
  NOR2_X1 U11746 ( .A1(n14724), .A2(n11797), .ZN(n14354) );
  AND2_X1 U11747 ( .A1(n12636), .A2(n12635), .ZN(n20205) );
  INV_X1 U11748 ( .A(n14294), .ZN(n14331) );
  AND2_X1 U11749 ( .A1(n12842), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14330) );
  NAND2_X1 U11750 ( .A1(n14299), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14327) );
  NAND2_X1 U11751 ( .A1(n14252), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14276) );
  NAND2_X1 U11752 ( .A1(n13432), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14187) );
  NOR2_X1 U11753 ( .A1(n14102), .A2(n15971), .ZN(n14119) );
  NAND2_X1 U11754 ( .A1(n14119), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14136) );
  NAND2_X1 U11755 ( .A1(n14894), .A2(n9873), .ZN(n10135) );
  NOR2_X1 U11756 ( .A1(n13249), .A2(n13248), .ZN(n13507) );
  AND2_X1 U11757 ( .A1(n15905), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14413) );
  AND2_X1 U11758 ( .A1(n14949), .A2(n11886), .ZN(n12882) );
  NAND2_X1 U11759 ( .A1(n12916), .A2(n12915), .ZN(n12923) );
  NOR2_X1 U11760 ( .A1(n14441), .A2(n14425), .ZN(n14426) );
  OAI21_X1 U11761 ( .B1(n9922), .B2(n14742), .A(n14743), .ZN(n14758) );
  INV_X1 U11762 ( .A(n16216), .ZN(n10062) );
  OR2_X1 U11763 ( .A1(n13814), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12064) );
  NOR2_X1 U11764 ( .A1(n16254), .A2(n12209), .ZN(n16231) );
  AND2_X1 U11765 ( .A1(n9885), .A2(n9884), .ZN(n14919) );
  NAND2_X1 U11766 ( .A1(n12305), .A2(n20984), .ZN(n9885) );
  AND2_X1 U11767 ( .A1(n12297), .A2(n13045), .ZN(n13901) );
  OR2_X1 U11768 ( .A1(n12299), .A2(n16241), .ZN(n9884) );
  INV_X1 U11769 ( .A(n15907), .ZN(n14408) );
  NAND2_X1 U11770 ( .A1(n9769), .A2(n13261), .ZN(n20423) );
  NAND2_X1 U11771 ( .A1(n13130), .A2(n13395), .ZN(n20510) );
  NAND2_X1 U11772 ( .A1(n11982), .A2(n11928), .ZN(n12131) );
  AND2_X1 U11773 ( .A1(n12098), .A2(n12102), .ZN(n12117) );
  OR2_X1 U11774 ( .A1(n12103), .A2(n12097), .ZN(n12098) );
  AOI21_X1 U11775 ( .B1(n9891), .B2(n9890), .A(n9888), .ZN(n12154) );
  INV_X1 U11776 ( .A(n12153), .ZN(n9890) );
  OAI21_X1 U11777 ( .B1(n12152), .B2(n12151), .A(n9889), .ZN(n9888) );
  OAI21_X1 U11778 ( .B1(n12140), .B2(n12141), .A(n9892), .ZN(n9891) );
  NOR2_X1 U11779 ( .A1(n10017), .A2(n11113), .ZN(n10016) );
  INV_X1 U11780 ( .A(n11103), .ZN(n10017) );
  AND2_X1 U11781 ( .A1(n11052), .A2(n11051), .ZN(n15043) );
  AND2_X1 U11782 ( .A1(n11309), .A2(n11308), .ZN(n15172) );
  XNOR2_X1 U11783 ( .A(n12500), .B(n12497), .ZN(n15113) );
  NOR2_X1 U11784 ( .A1(n15243), .A2(n10081), .ZN(n10080) );
  INV_X1 U11785 ( .A(n15036), .ZN(n10081) );
  INV_X1 U11786 ( .A(n10679), .ZN(n10678) );
  INV_X1 U11787 ( .A(n14968), .ZN(n10124) );
  AND2_X1 U11788 ( .A1(n10125), .A2(n10123), .ZN(n14969) );
  INV_X1 U11789 ( .A(n11654), .ZN(n10123) );
  AOI21_X1 U11790 ( .B1(n10058), .B2(n10056), .A(n10055), .ZN(n10054) );
  INV_X1 U11791 ( .A(n16380), .ZN(n10056) );
  INV_X1 U11792 ( .A(n15593), .ZN(n10055) );
  NOR2_X1 U11793 ( .A1(n19139), .A2(n13319), .ZN(n13322) );
  AND2_X1 U11794 ( .A1(n15034), .A2(n10079), .ZN(n15230) );
  AND2_X1 U11795 ( .A1(n9866), .A2(n15227), .ZN(n10079) );
  AND2_X1 U11796 ( .A1(n15353), .A2(n15550), .ZN(n10035) );
  NAND2_X1 U11797 ( .A1(n10050), .A2(n10048), .ZN(n15363) );
  AOI21_X1 U11798 ( .B1(n10051), .B2(n10057), .A(n10049), .ZN(n10048) );
  INV_X1 U11799 ( .A(n15330), .ZN(n10049) );
  NAND2_X1 U11800 ( .A1(n16379), .A2(n16380), .ZN(n16378) );
  AND3_X1 U11801 ( .A1(n11494), .A2(n11493), .A3(n11492), .ZN(n13312) );
  NOR2_X1 U11802 ( .A1(n15670), .A2(n10208), .ZN(n10207) );
  INV_X1 U11803 ( .A(n11018), .ZN(n10208) );
  NOR2_X1 U11804 ( .A1(n15657), .A2(n15667), .ZN(n9924) );
  NAND2_X1 U11805 ( .A1(n11416), .A2(n11415), .ZN(n15686) );
  NOR2_X1 U11806 ( .A1(n12929), .A2(n10075), .ZN(n13776) );
  NAND2_X1 U11807 ( .A1(n10077), .A2(n10076), .ZN(n10075) );
  INV_X1 U11808 ( .A(n13183), .ZN(n10076) );
  INV_X1 U11809 ( .A(n13272), .ZN(n9940) );
  AND2_X1 U11810 ( .A1(n11554), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10007) );
  AOI21_X1 U11811 ( .B1(n11393), .B2(n11395), .A(n11394), .ZN(n11400) );
  OR2_X1 U11812 ( .A1(n12929), .A2(n10074), .ZN(n13184) );
  INV_X1 U11813 ( .A(n10077), .ZN(n10074) );
  CLKBUF_X1 U11814 ( .A(n10662), .Z(n13659) );
  NAND2_X1 U11815 ( .A1(n19672), .A2(n20059), .ZN(n19579) );
  OR2_X1 U11816 ( .A1(n19672), .A2(n20059), .ZN(n19737) );
  NAND2_X1 U11817 ( .A1(n15715), .A2(n20053), .ZN(n19893) );
  NOR3_X1 U11818 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n10234), .ZN(n10235) );
  INV_X1 U11819 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20824) );
  INV_X1 U11820 ( .A(n17290), .ZN(n17325) );
  NOR2_X1 U11821 ( .A1(n17027), .A2(n10239), .ZN(n10265) );
  AOI21_X1 U11822 ( .B1(n10289), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n10332), .ZN(n10333) );
  NOR2_X1 U11823 ( .A1(n17275), .A2(n18570), .ZN(n10332) );
  AOI21_X1 U11824 ( .B1(n17185), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(n9982), .ZN(n9981) );
  NOR2_X1 U11825 ( .A1(n17300), .A2(n17203), .ZN(n9982) );
  NAND2_X1 U11826 ( .A1(n17673), .A2(n9803), .ZN(n16679) );
  NOR2_X1 U11827 ( .A1(n9798), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9970) );
  NAND2_X1 U11828 ( .A1(n17666), .A2(n18013), .ZN(n17665) );
  NOR2_X1 U11829 ( .A1(n10363), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9978) );
  INV_X1 U11830 ( .A(n9977), .ZN(n17743) );
  NAND2_X1 U11831 ( .A1(n9784), .A2(n9975), .ZN(n9971) );
  NAND2_X1 U11832 ( .A1(n10521), .A2(n17894), .ZN(n17820) );
  AND2_X1 U11833 ( .A1(n15994), .A2(n13445), .ZN(n20126) );
  AND2_X1 U11834 ( .A1(n14379), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13437) );
  AND2_X1 U11835 ( .A1(n15895), .A2(n14413), .ZN(n16116) );
  AND2_X1 U11836 ( .A1(n12311), .A2(n16256), .ZN(n9896) );
  NAND2_X1 U11837 ( .A1(n9986), .A2(n9992), .ZN(n12088) );
  NAND2_X1 U11838 ( .A1(n9996), .A2(n9988), .ZN(n9992) );
  NAND2_X1 U11839 ( .A1(n9994), .A2(n9987), .ZN(n9986) );
  AND2_X1 U11840 ( .A1(n12299), .A2(n12177), .ZN(n16244) );
  CLKBUF_X1 U11841 ( .A(n13284), .Z(n20551) );
  INV_X1 U11842 ( .A(n15416), .ZN(n15090) );
  AND2_X1 U11843 ( .A1(n10183), .A2(n13174), .ZN(n10179) );
  AND2_X1 U11844 ( .A1(n10226), .A2(n10184), .ZN(n10183) );
  AND2_X1 U11845 ( .A1(n15159), .A2(n19431), .ZN(n15149) );
  XNOR2_X1 U11846 ( .A(n14363), .B(n14362), .ZN(n19241) );
  INV_X1 U11847 ( .A(n20059), .ZN(n19638) );
  AND2_X1 U11848 ( .A1(n16445), .A2(n20049), .ZN(n16421) );
  INV_X1 U11849 ( .A(n16435), .ZN(n16427) );
  INV_X1 U11850 ( .A(n16425), .ZN(n16441) );
  NAND2_X1 U11851 ( .A1(n14372), .A2(n10230), .ZN(n10115) );
  XNOR2_X1 U11852 ( .A(n9943), .B(n11623), .ZN(n14373) );
  AOI21_X1 U11853 ( .B1(n15277), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11648), .ZN(n11651) );
  AND2_X1 U11854 ( .A1(n11647), .A2(n11646), .ZN(n11648) );
  NAND2_X1 U11855 ( .A1(n10195), .A2(n10194), .ZN(n10193) );
  NAND2_X1 U11856 ( .A1(n19384), .A2(n15601), .ZN(n10194) );
  AND2_X1 U11857 ( .A1(n11578), .A2(n11368), .ZN(n16474) );
  AND2_X1 U11858 ( .A1(n11252), .A2(n11377), .ZN(n19391) );
  XNOR2_X1 U11859 ( .A(n12794), .B(n12793), .ZN(n20053) );
  INV_X1 U11860 ( .A(n20043), .ZN(n15715) );
  AND2_X1 U11861 ( .A1(n13643), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15714) );
  NAND2_X1 U11862 ( .A1(n16496), .A2(n18212), .ZN(n10551) );
  XNOR2_X1 U11863 ( .A(n10164), .B(n16518), .ZN(n16515) );
  NAND2_X1 U11864 ( .A1(n10166), .A2(n10165), .ZN(n10164) );
  NOR2_X1 U11865 ( .A1(n18279), .A2(n18289), .ZN(n18287) );
  INV_X1 U11866 ( .A(n10232), .ZN(n9912) );
  AND4_X1 U11867 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n10990) );
  AND4_X1 U11868 ( .A1(n10948), .A2(n10947), .A3(n10946), .A4(n10945), .ZN(
        n10955) );
  INV_X1 U11869 ( .A(n12122), .ZN(n12104) );
  AND2_X2 U11870 ( .A1(n11675), .A2(n13229), .ZN(n11782) );
  NAND2_X1 U11871 ( .A1(n11943), .A2(n10147), .ZN(n12033) );
  AND2_X2 U11872 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U11873 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U11874 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11777), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U11875 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9750), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U11877 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10633) );
  AND2_X1 U11878 ( .A1(n11036), .A2(n9860), .ZN(n11053) );
  NOR2_X1 U11879 ( .A1(n11067), .A2(n10013), .ZN(n10012) );
  NAND2_X1 U11880 ( .A1(n11566), .A2(n10688), .ZN(n10692) );
  AND4_X1 U11881 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10879) );
  NOR2_X1 U11882 ( .A1(n10662), .A2(n10656), .ZN(n10680) );
  AOI21_X1 U11883 ( .B1(n13738), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n10808), .ZN(n10819) );
  AOI21_X1 U11884 ( .B1(n10943), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n11377), .ZN(n10806) );
  AOI22_X1 U11885 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10940), .B1(
        n10938), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10774) );
  INV_X1 U11886 ( .A(n10668), .ZN(n11563) );
  AOI22_X1 U11887 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10574) );
  AOI21_X1 U11888 ( .B1(n10922), .B2(n10921), .A(n10920), .ZN(n11153) );
  AND2_X1 U11889 ( .A1(n10529), .A2(n18330), .ZN(n10459) );
  AOI22_X1 U11890 ( .A1(n11833), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11745) );
  NOR2_X1 U11891 ( .A1(n12103), .A2(n12102), .ZN(n12149) );
  AND2_X1 U11892 ( .A1(n14784), .A2(n14188), .ZN(n14189) );
  NOR2_X1 U11893 ( .A1(n10142), .A2(n10140), .ZN(n10139) );
  INV_X1 U11894 ( .A(n10141), .ZN(n10140) );
  NOR2_X1 U11895 ( .A1(n14563), .A2(n14503), .ZN(n10141) );
  INV_X1 U11896 ( .A(n14297), .ZN(n14324) );
  OR2_X1 U11897 ( .A1(n10146), .A2(n10145), .ZN(n10144) );
  INV_X1 U11898 ( .A(n14519), .ZN(n10145) );
  OR2_X1 U11899 ( .A1(n14020), .A2(n14602), .ZN(n10146) );
  OR2_X1 U11900 ( .A1(n13923), .A2(n14548), .ZN(n13955) );
  OR2_X1 U11901 ( .A1(n14477), .A2(n10069), .ZN(n10067) );
  OR2_X1 U11902 ( .A1(n14814), .A2(n16073), .ZN(n12071) );
  NOR2_X1 U11903 ( .A1(n12209), .A2(n10065), .ZN(n10064) );
  INV_X1 U11904 ( .A(n13572), .ZN(n10065) );
  INV_X1 U11905 ( .A(n12866), .ZN(n9900) );
  AND2_X1 U11906 ( .A1(n12158), .A2(n13158), .ZN(n9902) );
  NOR2_X1 U11907 ( .A1(n12159), .A2(n13158), .ZN(n9901) );
  AND2_X1 U11908 ( .A1(n12299), .A2(n12291), .ZN(n12305) );
  OR2_X1 U11909 ( .A1(n11852), .A2(n11851), .ZN(n11993) );
  OR2_X1 U11910 ( .A1(n11839), .A2(n11838), .ZN(n12057) );
  INV_X1 U11911 ( .A(n11881), .ZN(n11828) );
  OR2_X1 U11912 ( .A1(n11871), .A2(n11870), .ZN(n11994) );
  INV_X1 U11913 ( .A(n11928), .ZN(n11917) );
  INV_X1 U11914 ( .A(n12116), .ZN(n12150) );
  NAND2_X1 U11915 ( .A1(n13158), .A2(n11700), .ZN(n11716) );
  NOR2_X1 U11916 ( .A1(n11802), .A2(n9766), .ZN(n9914) );
  NAND2_X1 U11917 ( .A1(n9904), .A2(n11885), .ZN(n11904) );
  AOI221_X1 U11918 ( .B1(n20661), .B2(P1_STATE2_REG_2__SCAN_IN), .C1(
        P1_STATE2_REG_1__SCAN_IN), .C2(n12842), .A(n14957), .ZN(n13135) );
  OR2_X1 U11919 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20263), .ZN(
        n12102) );
  NOR2_X1 U11920 ( .A1(n12145), .A2(n9893), .ZN(n9892) );
  AND2_X1 U11921 ( .A1(n12163), .A2(n12146), .ZN(n9893) );
  NAND2_X1 U11922 ( .A1(n11886), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9889) );
  INV_X1 U11923 ( .A(n11802), .ZN(n12880) );
  AND2_X1 U11924 ( .A1(n12279), .A2(n12162), .ZN(n12881) );
  INV_X1 U11925 ( .A(n10688), .ZN(n10924) );
  NAND2_X1 U11926 ( .A1(n11055), .A2(n11049), .ZN(n11050) );
  NAND2_X1 U11927 ( .A1(n11036), .A2(n10012), .ZN(n11082) );
  NAND2_X1 U11928 ( .A1(n11036), .A2(n11037), .ZN(n11068) );
  NAND2_X1 U11929 ( .A1(n11029), .A2(n19113), .ZN(n11038) );
  NOR2_X1 U11930 ( .A1(n11027), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11029) );
  NAND2_X1 U11931 ( .A1(n11024), .A2(n11021), .ZN(n11027) );
  AND2_X1 U11932 ( .A1(n15201), .A2(n14996), .ZN(n10090) );
  OAI21_X1 U11933 ( .B1(n10583), .B2(n10582), .A(n13590), .ZN(n10592) );
  OAI21_X1 U11934 ( .B1(n10590), .B2(n10589), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10591) );
  NOR2_X1 U11935 ( .A1(n15029), .A2(n10093), .ZN(n10092) );
  NOR2_X1 U11936 ( .A1(n15358), .A2(n10100), .ZN(n10099) );
  INV_X1 U11937 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10100) );
  NOR2_X1 U11938 ( .A1(n19114), .A2(n10097), .ZN(n10096) );
  NAND2_X1 U11939 ( .A1(n10118), .A2(n10229), .ZN(n10117) );
  INV_X1 U11940 ( .A(n13162), .ZN(n10118) );
  OR2_X1 U11941 ( .A1(n11630), .A2(n19408), .ZN(n10724) );
  NAND2_X1 U11942 ( .A1(n10023), .A2(n10022), .ZN(n10696) );
  NOR2_X1 U11943 ( .A1(n15271), .A2(n10214), .ZN(n10213) );
  AND2_X1 U11944 ( .A1(n9810), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10212) );
  OR2_X1 U11945 ( .A1(n15873), .A2(n11023), .ZN(n11107) );
  INV_X1 U11946 ( .A(n15345), .ZN(n10034) );
  AND2_X1 U11947 ( .A1(n11250), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10211) );
  NOR2_X1 U11948 ( .A1(n10052), .A2(n15375), .ZN(n10051) );
  INV_X1 U11949 ( .A(n10054), .ZN(n10052) );
  AND2_X1 U11950 ( .A1(n9808), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10197) );
  INV_X1 U11951 ( .A(n13270), .ZN(n10210) );
  OR2_X1 U11952 ( .A1(n10802), .A2(n10801), .ZN(n10008) );
  INV_X1 U11953 ( .A(n13181), .ZN(n10078) );
  NOR2_X1 U11954 ( .A1(n12518), .A2(n19413), .ZN(n12330) );
  XNOR2_X1 U11955 ( .A(n10740), .B(n9740), .ZN(n10758) );
  OAI21_X1 U11956 ( .B1(n10664), .B2(n10706), .A(n9952), .ZN(n11560) );
  NAND2_X1 U11957 ( .A1(n9950), .A2(n11561), .ZN(n9952) );
  AND2_X1 U11958 ( .A1(n9721), .A2(n19421), .ZN(n9950) );
  NOR2_X1 U11959 ( .A1(n19421), .A2(n10668), .ZN(n10658) );
  NAND2_X1 U11960 ( .A1(n10222), .A2(n10759), .ZN(n10986) );
  INV_X1 U11961 ( .A(n10770), .ZN(n10759) );
  NAND2_X1 U11962 ( .A1(n12318), .A2(n12767), .ZN(n10770) );
  NOR2_X2 U11963 ( .A1(n10771), .A2(n9774), .ZN(n13738) );
  AOI22_X1 U11964 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U11965 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10622) );
  NAND2_X1 U11966 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10562) );
  NAND2_X1 U11967 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U11968 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U11969 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10558) );
  NAND3_X1 U11970 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20029), .A3(n19889), 
        .ZN(n13658) );
  NAND2_X1 U11971 ( .A1(n10882), .A2(n10881), .ZN(n10888) );
  INV_X1 U11972 ( .A(n11201), .ZN(n10687) );
  AOI21_X1 U11973 ( .B1(n17205), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n10273), .ZN(n10274) );
  NOR2_X1 U11974 ( .A1(n17674), .A2(n9966), .ZN(n9965) );
  NOR2_X1 U11975 ( .A1(n17923), .A2(n10351), .ZN(n10353) );
  AND2_X1 U11976 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10350), .ZN(
        n10351) );
  OAI21_X1 U11977 ( .B1(n16548), .B2(n16536), .A(n17897), .ZN(n10352) );
  NOR2_X1 U11978 ( .A1(n17499), .A2(n10324), .ZN(n10347) );
  XNOR2_X1 U11979 ( .A(n17507), .B(n10494), .ZN(n10341) );
  NOR2_X1 U11980 ( .A1(n10494), .A2(n17507), .ZN(n10343) );
  AOI21_X1 U11981 ( .B1(n10537), .B2(n18970), .A(n10538), .ZN(n18782) );
  OR2_X1 U11982 ( .A1(n18783), .A2(n10526), .ZN(n15741) );
  MUX2_X1 U11983 ( .A(n12243), .B(n12205), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12192) );
  AND2_X1 U11984 ( .A1(n14214), .A2(n14213), .ZN(n14482) );
  OR2_X1 U11985 ( .A1(n14777), .A2(n14303), .ZN(n14213) );
  OR2_X1 U11986 ( .A1(n14736), .A2(n14303), .ZN(n14304) );
  INV_X1 U11987 ( .A(n10150), .ZN(n10148) );
  AND2_X1 U11988 ( .A1(n13434), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14252) );
  OR2_X1 U11989 ( .A1(n14761), .A2(n14303), .ZN(n14256) );
  INV_X1 U11990 ( .A(n14136), .ZN(n13431) );
  AND2_X1 U11991 ( .A1(n14121), .A2(n14120), .ZN(n14572) );
  AND2_X1 U11992 ( .A1(n14104), .A2(n14103), .ZN(n14577) );
  AND2_X1 U11993 ( .A1(n14055), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14085) );
  NAND2_X1 U11994 ( .A1(n14085), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14102) );
  CLKBUF_X1 U11995 ( .A(n14578), .Z(n14579) );
  INV_X1 U11996 ( .A(n14587), .ZN(n14595) );
  OR2_X1 U11997 ( .A1(n14037), .A2(n14816), .ZN(n14040) );
  NAND2_X1 U11998 ( .A1(n14014), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14037) );
  NOR2_X1 U11999 ( .A1(n21042), .A2(n13955), .ZN(n14014) );
  OR2_X1 U12000 ( .A1(n13948), .A2(n16028), .ZN(n13923) );
  NAND2_X1 U12001 ( .A1(n13978), .A2(n13922), .ZN(n13954) );
  AND2_X1 U12002 ( .A1(n13846), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13908) );
  NAND2_X1 U12003 ( .A1(n13908), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13948) );
  NOR2_X1 U12004 ( .A1(n13793), .A2(n20122), .ZN(n13846) );
  NAND2_X1 U12005 ( .A1(n13551), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13793) );
  AND2_X1 U12006 ( .A1(n13516), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13551) );
  AND2_X1 U12007 ( .A1(n13522), .A2(n13523), .ZN(n13556) );
  AOI21_X1 U12008 ( .B1(n13513), .B2(n14011), .A(n13512), .ZN(n13562) );
  AOI21_X1 U12009 ( .B1(n13253), .B2(n14011), .A(n13252), .ZN(n13256) );
  AND2_X1 U12010 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13083) );
  NAND2_X1 U12011 ( .A1(n20266), .A2(n14011), .ZN(n13027) );
  NAND2_X1 U12012 ( .A1(n13031), .A2(n13030), .ZN(n13082) );
  INV_X1 U12013 ( .A(n13029), .ZN(n13030) );
  INV_X1 U12014 ( .A(n13033), .ZN(n13031) );
  NAND2_X1 U12015 ( .A1(n9989), .A2(n9851), .ZN(n9987) );
  NOR2_X1 U12016 ( .A1(n14498), .A2(n10067), .ZN(n14464) );
  NOR2_X1 U12017 ( .A1(n14498), .A2(n14477), .ZN(n14478) );
  NAND2_X1 U12018 ( .A1(n14591), .A2(n9867), .ZN(n14512) );
  INV_X1 U12019 ( .A(n14510), .ZN(n10060) );
  NAND2_X1 U12020 ( .A1(n14591), .A2(n9776), .ZN(n14567) );
  AOI21_X1 U12021 ( .B1(n10133), .B2(n10130), .A(n14894), .ZN(n10129) );
  NOR2_X1 U12022 ( .A1(n9777), .A2(n12309), .ZN(n10130) );
  NAND2_X1 U12023 ( .A1(n9999), .A2(n9997), .ZN(n12080) );
  AND2_X1 U12024 ( .A1(n9998), .A2(n12079), .ZN(n9997) );
  NAND2_X1 U12025 ( .A1(n14591), .A2(n14582), .ZN(n14585) );
  AND2_X1 U12026 ( .A1(n9999), .A2(n9998), .ZN(n14895) );
  NAND2_X1 U12027 ( .A1(n10128), .A2(n10133), .ZN(n14807) );
  NAND2_X1 U12028 ( .A1(n16064), .A2(n9777), .ZN(n10128) );
  NAND2_X1 U12029 ( .A1(n12073), .A2(n12072), .ZN(n16064) );
  NAND2_X1 U12030 ( .A1(n14538), .A2(n9850), .ZN(n14605) );
  AND2_X1 U12031 ( .A1(n14538), .A2(n10070), .ZN(n14611) );
  AND2_X1 U12032 ( .A1(n12231), .A2(n12230), .ZN(n13898) );
  NAND2_X1 U12033 ( .A1(n14538), .A2(n10072), .ZN(n14612) );
  AND2_X1 U12034 ( .A1(n12226), .A2(n12225), .ZN(n14539) );
  NAND2_X1 U12035 ( .A1(n14538), .A2(n14539), .ZN(n14541) );
  AND2_X1 U12036 ( .A1(n12219), .A2(n12218), .ZN(n13863) );
  CLKBUF_X1 U12037 ( .A(n13891), .Z(n14834) );
  NAND2_X1 U12038 ( .A1(n10063), .A2(n10064), .ZN(n16217) );
  NAND2_X1 U12039 ( .A1(n16108), .A2(n9782), .ZN(n9916) );
  INV_X1 U12040 ( .A(n16251), .ZN(n12199) );
  INV_X1 U12041 ( .A(n11797), .ZN(n9909) );
  NAND2_X1 U12042 ( .A1(n12205), .A2(n12179), .ZN(n12833) );
  CLKBUF_X1 U12043 ( .A(n12840), .Z(n12841) );
  NAND2_X1 U12044 ( .A1(n10126), .A2(n11874), .ZN(n11875) );
  NAND2_X1 U12045 ( .A1(n11927), .A2(n11926), .ZN(n13343) );
  NOR2_X1 U12046 ( .A1(n12870), .A2(n13070), .ZN(n15881) );
  NOR2_X1 U12047 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20518) );
  INV_X1 U12048 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20599) );
  INV_X1 U12049 ( .A(n12129), .ZN(n13139) );
  INV_X1 U12050 ( .A(n13156), .ZN(n13681) );
  INV_X1 U12051 ( .A(n13155), .ZN(n13682) );
  AOI21_X1 U12052 ( .B1(n20449), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n13676), 
        .ZN(n20607) );
  INV_X1 U12053 ( .A(n11167), .ZN(n11212) );
  OR2_X1 U12054 ( .A1(n11577), .A2(n11576), .ZN(n13607) );
  NAND2_X1 U12055 ( .A1(n11132), .A2(n11131), .ZN(n11644) );
  INV_X1 U12056 ( .A(n11620), .ZN(n11132) );
  AND2_X1 U12057 ( .A1(n11104), .A2(n9807), .ZN(n11129) );
  NAND2_X1 U12058 ( .A1(n11104), .A2(n11103), .ZN(n11114) );
  AND2_X1 U12059 ( .A1(n11065), .A2(n11064), .ZN(n19072) );
  AND2_X1 U12060 ( .A1(n11006), .A2(n10010), .ZN(n11015) );
  NAND2_X1 U12061 ( .A1(n11006), .A2(n11005), .ZN(n11010) );
  INV_X1 U12062 ( .A(n13200), .ZN(n10188) );
  OR2_X1 U12063 ( .A1(n11479), .A2(n11478), .ZN(n12350) );
  AND2_X1 U12064 ( .A1(n11289), .A2(n11288), .ZN(n13196) );
  OR2_X1 U12065 ( .A1(n10117), .A2(n13196), .ZN(n10116) );
  OR2_X1 U12066 ( .A1(n11455), .A2(n11454), .ZN(n12347) );
  AND2_X1 U12067 ( .A1(n11273), .A2(n11272), .ZN(n13054) );
  NOR2_X1 U12068 ( .A1(n12346), .A2(n10185), .ZN(n10184) );
  NOR2_X1 U12069 ( .A1(n10171), .A2(n10174), .ZN(n10169) );
  NAND2_X1 U12070 ( .A1(n9745), .A2(n10170), .ZN(n10167) );
  NOR2_X1 U12071 ( .A1(n10171), .A2(n15092), .ZN(n10170) );
  NAND2_X1 U12072 ( .A1(n10172), .A2(n10175), .ZN(n15086) );
  NAND2_X1 U12073 ( .A1(n9745), .A2(n10176), .ZN(n10175) );
  NAND2_X1 U12074 ( .A1(n15096), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U12075 ( .A1(n15230), .A2(n15026), .ZN(n15007) );
  OR2_X1 U12076 ( .A1(n15117), .A2(n15127), .ZN(n10177) );
  OR2_X1 U12077 ( .A1(n15128), .A2(n15127), .ZN(n10178) );
  NAND2_X1 U12078 ( .A1(n9796), .A2(n15178), .ZN(n10186) );
  INV_X1 U12079 ( .A(n13604), .ZN(n13610) );
  INV_X1 U12080 ( .A(n12631), .ZN(n13840) );
  XNOR2_X1 U12081 ( .A(n11635), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13313) );
  NAND2_X1 U12082 ( .A1(n15259), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11635) );
  AND2_X1 U12083 ( .A1(n9811), .A2(n9879), .ZN(n9956) );
  NOR2_X1 U12084 ( .A1(n14973), .A2(n11634), .ZN(n14992) );
  AND2_X1 U12085 ( .A1(n14992), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15259) );
  NAND2_X1 U12086 ( .A1(n14978), .A2(n10091), .ZN(n14973) );
  AND2_X1 U12087 ( .A1(n9805), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10091) );
  INV_X1 U12088 ( .A(n10125), .ZN(n15102) );
  NAND2_X1 U12089 ( .A1(n14978), .A2(n9805), .ZN(n14975) );
  NAND2_X1 U12090 ( .A1(n14978), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14977) );
  NAND2_X1 U12091 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n14980), .ZN(
        n14979) );
  NOR2_X1 U12092 ( .A1(n16362), .A2(n14979), .ZN(n14978) );
  NOR2_X1 U12093 ( .A1(n15133), .A2(n15123), .ZN(n15124) );
  AND2_X1 U12094 ( .A1(n11329), .A2(n11328), .ZN(n15131) );
  AND2_X1 U12095 ( .A1(n14990), .A2(n10098), .ZN(n14980) );
  AND2_X1 U12096 ( .A1(n9806), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10098) );
  AND2_X1 U12097 ( .A1(n9849), .A2(n15040), .ZN(n10120) );
  NAND2_X1 U12098 ( .A1(n14990), .A2(n9806), .ZN(n14991) );
  AND2_X1 U12099 ( .A1(n11321), .A2(n11320), .ZN(n15150) );
  AND2_X1 U12100 ( .A1(n15171), .A2(n9849), .ZN(n15152) );
  NAND2_X1 U12101 ( .A1(n15171), .A2(n9842), .ZN(n15156) );
  NOR2_X1 U12102 ( .A1(n15369), .A2(n14987), .ZN(n14990) );
  NAND2_X1 U12103 ( .A1(n14990), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14989) );
  NAND2_X1 U12104 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14988), .ZN(
        n14987) );
  NOR2_X1 U12105 ( .A1(n19090), .A2(n14985), .ZN(n14988) );
  AND2_X1 U12106 ( .A1(n11301), .A2(n11300), .ZN(n13732) );
  NAND2_X1 U12107 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n14986), .ZN(
        n14985) );
  NAND2_X1 U12108 ( .A1(n13419), .A2(n13477), .ZN(n13731) );
  AND2_X1 U12109 ( .A1(n13322), .A2(n10095), .ZN(n14986) );
  AND2_X1 U12110 ( .A1(n9797), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10095) );
  NAND2_X1 U12111 ( .A1(n13322), .A2(n9797), .ZN(n14983) );
  OR2_X1 U12112 ( .A1(n13060), .A2(n10117), .ZN(n13197) );
  NAND2_X1 U12113 ( .A1(n13322), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13321) );
  NAND2_X1 U12114 ( .A1(n10103), .A2(n9854), .ZN(n13319) );
  AND2_X1 U12115 ( .A1(n10103), .A2(n10102), .ZN(n13320) );
  NAND2_X1 U12116 ( .A1(n10103), .A2(n10104), .ZN(n13317) );
  NAND2_X1 U12117 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n13316), .ZN(
        n13315) );
  NOR2_X1 U12118 ( .A1(n13315), .A2(n16432), .ZN(n13318) );
  NOR2_X1 U12119 ( .A1(n13314), .A2(n16446), .ZN(n13316) );
  NAND2_X1 U12120 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13314) );
  AOI21_X1 U12121 ( .B1(n9747), .B2(n9945), .A(n9829), .ZN(n9944) );
  OAI21_X1 U12122 ( .B1(n10202), .B2(n9876), .A(n11649), .ZN(n10004) );
  OR2_X1 U12123 ( .A1(n14999), .A2(n11143), .ZN(n15266) );
  AND2_X1 U12124 ( .A1(n16295), .A2(n11621), .ZN(n11649) );
  OR2_X1 U12125 ( .A1(n15203), .A2(n15202), .ZN(n16296) );
  INV_X1 U12126 ( .A(n11646), .ZN(n11645) );
  NAND2_X1 U12127 ( .A1(n11124), .A2(n11134), .ZN(n15287) );
  NAND2_X1 U12128 ( .A1(n15020), .A2(n15021), .ZN(n15023) );
  NAND2_X1 U12129 ( .A1(n9935), .A2(n9933), .ZN(n15493) );
  AOI21_X1 U12130 ( .B1(n9936), .B2(n9939), .A(n9934), .ZN(n9933) );
  INV_X1 U12131 ( .A(n15320), .ZN(n9934) );
  NOR2_X1 U12132 ( .A1(n9821), .A2(n10206), .ZN(n10205) );
  INV_X1 U12133 ( .A(n15335), .ZN(n10206) );
  NAND2_X1 U12134 ( .A1(n15343), .A2(n9880), .ZN(n15484) );
  NAND2_X1 U12135 ( .A1(n10030), .A2(n10027), .ZN(n10026) );
  NAND2_X1 U12136 ( .A1(n10033), .A2(n10029), .ZN(n10027) );
  AOI21_X1 U12137 ( .B1(n10032), .B2(n15352), .A(n10031), .ZN(n10030) );
  INV_X1 U12138 ( .A(n15334), .ZN(n10031) );
  INV_X1 U12139 ( .A(n15336), .ZN(n10029) );
  OAI21_X1 U12140 ( .B1(n15363), .B2(n15364), .A(n15332), .ZN(n15552) );
  OR2_X1 U12141 ( .A1(n15596), .A2(n9844), .ZN(n15559) );
  OR2_X1 U12142 ( .A1(n15596), .A2(n10086), .ZN(n15557) );
  AND2_X1 U12143 ( .A1(n15637), .A2(n10196), .ZN(n15569) );
  AND2_X1 U12144 ( .A1(n10197), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10196) );
  INV_X1 U12145 ( .A(n15604), .ZN(n10195) );
  OR2_X1 U12146 ( .A1(n13731), .A2(n13732), .ZN(n15181) );
  AND2_X1 U12147 ( .A1(n11305), .A2(n11304), .ZN(n15180) );
  OR2_X1 U12148 ( .A1(n15181), .A2(n15180), .ZN(n15183) );
  AND2_X1 U12149 ( .A1(n11524), .A2(n11523), .ZN(n15579) );
  NAND2_X1 U12150 ( .A1(n15637), .A2(n10197), .ZN(n15591) );
  NAND2_X1 U12151 ( .A1(n10084), .A2(n10083), .ZN(n10082) );
  NOR2_X1 U12152 ( .A1(n9838), .A2(n16448), .ZN(n10083) );
  NAND2_X1 U12153 ( .A1(n15637), .A2(n16450), .ZN(n16376) );
  OR3_X1 U12154 ( .A1(n15659), .A2(n11496), .A3(n9838), .ZN(n16449) );
  INV_X1 U12155 ( .A(n15637), .ZN(n15621) );
  OR2_X1 U12156 ( .A1(n16479), .A2(n16464), .ZN(n15646) );
  NAND2_X1 U12157 ( .A1(n9927), .A2(n16411), .ZN(n9926) );
  INV_X1 U12158 ( .A(n11245), .ZN(n9927) );
  AND3_X1 U12159 ( .A1(n11433), .A2(n11432), .A3(n11431), .ZN(n16463) );
  NAND2_X1 U12160 ( .A1(n15393), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9949) );
  NAND2_X1 U12161 ( .A1(n15686), .A2(n15685), .ZN(n16462) );
  OR2_X1 U12162 ( .A1(n13782), .A2(n13781), .ZN(n11603) );
  NAND2_X1 U12163 ( .A1(n13774), .A2(n11412), .ZN(n15694) );
  AND2_X1 U12164 ( .A1(n10108), .A2(n9789), .ZN(n12985) );
  INV_X1 U12165 ( .A(n12986), .ZN(n10109) );
  INV_X1 U12166 ( .A(n13378), .ZN(n10107) );
  OR2_X1 U12167 ( .A1(n13379), .A2(n9868), .ZN(n13779) );
  NOR2_X1 U12168 ( .A1(n13769), .A2(n11231), .ZN(n11232) );
  AND3_X1 U12169 ( .A1(n11406), .A2(n11405), .A3(n11404), .ZN(n13183) );
  INV_X1 U12170 ( .A(n11566), .ZN(n9930) );
  AND2_X1 U12171 ( .A1(n11585), .A2(n16479), .ZN(n13273) );
  NAND2_X1 U12172 ( .A1(n13280), .A2(n11023), .ZN(n10896) );
  NAND2_X1 U12173 ( .A1(n11578), .A2(n12742), .ZN(n19387) );
  XNOR2_X1 U12174 ( .A(n12780), .B(n11383), .ZN(n12813) );
  AND2_X1 U12175 ( .A1(n11388), .A2(n11387), .ZN(n12812) );
  OAI22_X1 U12176 ( .A1(n12794), .A2(n12793), .B1(n12330), .B2(n15705), .ZN(
        n12823) );
  OR2_X1 U12177 ( .A1(n12339), .A2(n12338), .ZN(n12340) );
  NAND2_X1 U12178 ( .A1(n12313), .A2(n20037), .ZN(n12333) );
  OAI22_X2 U12179 ( .A1(n19309), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n13313), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19206) );
  NAND2_X1 U12180 ( .A1(n11191), .A2(n11190), .ZN(n13643) );
  NAND2_X1 U12181 ( .A1(n20043), .A2(n20053), .ZN(n20030) );
  OR2_X1 U12182 ( .A1(n19672), .A2(n19638), .ZN(n19769) );
  NAND2_X1 U12183 ( .A1(n15715), .A2(n20050), .ZN(n19817) );
  INV_X1 U12184 ( .A(n19737), .ZN(n19819) );
  INV_X1 U12185 ( .A(n19434), .ZN(n19420) );
  INV_X1 U12186 ( .A(n19435), .ZN(n19418) );
  NAND2_X1 U12187 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19889), .ZN(n19414) );
  INV_X1 U12188 ( .A(n19769), .ZN(n19847) );
  NOR2_X2 U12189 ( .A1(n13840), .A2(n13658), .ZN(n19435) );
  INV_X1 U12190 ( .A(n19414), .ZN(n19430) );
  NAND2_X1 U12191 ( .A1(n10687), .A2(n20081), .ZN(n13639) );
  NOR2_X1 U12192 ( .A1(n17580), .A2(n15845), .ZN(n18766) );
  OR2_X1 U12193 ( .A1(n9729), .A2(n9958), .ZN(n16832) );
  NOR2_X1 U12194 ( .A1(n16845), .A2(n17790), .ZN(n9958) );
  NAND2_X1 U12195 ( .A1(n16832), .A2(n17782), .ZN(n16831) );
  NOR2_X1 U12196 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16920), .ZN(n16904) );
  NAND2_X1 U12197 ( .A1(n16507), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16506) );
  INV_X1 U12198 ( .A(n16671), .ZN(n16670) );
  OAI211_X1 U12199 ( .C1(n10253), .C2(n18355), .A(n10433), .B(n10432), .ZN(
        n17374) );
  NOR3_X1 U12200 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n20969), .ZN(n10244) );
  NAND2_X1 U12201 ( .A1(n10302), .A2(n10301), .ZN(n10492) );
  NOR2_X1 U12202 ( .A1(n10300), .A2(n10299), .ZN(n10301) );
  AND2_X1 U12203 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10299) );
  NOR2_X1 U12204 ( .A1(n10285), .A2(n10159), .ZN(n10158) );
  OAI21_X1 U12205 ( .B1(n15847), .B2(n15743), .A(n18977), .ZN(n15938) );
  NOR3_X1 U12206 ( .A1(n17456), .A2(n15742), .A3(n15741), .ZN(n15743) );
  OAI221_X1 U12207 ( .B1(n15850), .B2(n17580), .C1(n15850), .C2(n18970), .A(
        n15849), .ZN(n15940) );
  INV_X1 U12208 ( .A(n18789), .ZN(n15850) );
  AOI21_X1 U12209 ( .B1(n15846), .B2(n18826), .A(n18850), .ZN(n17522) );
  INV_X1 U12210 ( .A(n17577), .ZN(n17524) );
  INV_X1 U12211 ( .A(n17521), .ZN(n17579) );
  NAND2_X1 U12212 ( .A1(n17673), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16683) );
  NAND2_X1 U12213 ( .A1(n17673), .A2(n9965), .ZN(n17632) );
  NOR2_X1 U12214 ( .A1(n9960), .A2(n9961), .ZN(n9959) );
  INV_X1 U12215 ( .A(n17835), .ZN(n18160) );
  INV_X1 U12216 ( .A(n17820), .ZN(n18162) );
  INV_X1 U12217 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16937) );
  NAND2_X1 U12218 ( .A1(n9964), .A2(n9962), .ZN(n17901) );
  NOR2_X1 U12219 ( .A1(n17939), .A2(n9963), .ZN(n9962) );
  NAND2_X1 U12220 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9963) );
  AND3_X1 U12221 ( .A1(n9964), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17928) );
  NOR2_X1 U12222 ( .A1(n15922), .A2(n17871), .ZN(n10368) );
  AND2_X1 U12223 ( .A1(n10367), .A2(n9968), .ZN(n15922) );
  NOR2_X1 U12224 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n9969), .ZN(
        n9968) );
  INV_X1 U12225 ( .A(n9970), .ZN(n9969) );
  NAND2_X1 U12226 ( .A1(n10347), .A2(n10346), .ZN(n10349) );
  NOR2_X1 U12227 ( .A1(n17670), .A2(n10545), .ZN(n18006) );
  INV_X1 U12228 ( .A(n17692), .ZN(n17680) );
  NOR2_X1 U12229 ( .A1(n18132), .A2(n17684), .ZN(n18041) );
  INV_X1 U12230 ( .A(n17690), .ZN(n18039) );
  INV_X1 U12231 ( .A(n17804), .ZN(n18057) );
  INV_X1 U12232 ( .A(n18279), .ZN(n18767) );
  NOR2_X1 U12233 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17730), .ZN(
        n17710) );
  NAND2_X1 U12234 ( .A1(n18134), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18132) );
  NAND2_X1 U12235 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17896), .ZN(
        n17835) );
  NAND2_X1 U12236 ( .A1(n9973), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17815) );
  XNOR2_X1 U12237 ( .A(n10353), .B(n10352), .ZN(n17912) );
  NOR2_X1 U12238 ( .A1(n17912), .A2(n17913), .ZN(n17911) );
  NAND2_X1 U12239 ( .A1(n9979), .A2(n17935), .ZN(n17925) );
  OAI21_X1 U12240 ( .B1(n17936), .B2(n17937), .A(n10348), .ZN(n9979) );
  NOR2_X1 U12241 ( .A1(n17925), .A2(n17924), .ZN(n17923) );
  NAND2_X1 U12242 ( .A1(n17936), .A2(n17937), .ZN(n17935) );
  NOR2_X1 U12243 ( .A1(n10491), .A2(n10490), .ZN(n18274) );
  OAI21_X1 U12244 ( .B1(n18783), .B2(n18794), .A(n18782), .ZN(n18803) );
  NOR2_X1 U12245 ( .A1(n10539), .A2(n10538), .ZN(n15848) );
  AOI21_X1 U12246 ( .B1(n10478), .B2(n10477), .A(n10476), .ZN(n18768) );
  INV_X1 U12247 ( .A(n18794), .ZN(n18792) );
  NAND2_X1 U12248 ( .A1(n18792), .A2(n15848), .ZN(n18789) );
  AOI211_X1 U12249 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n10423), .B(n10422), .ZN(n18347) );
  INV_X1 U12250 ( .A(n17374), .ZN(n18352) );
  AOI22_X1 U12251 ( .A1(n18768), .A2(n18767), .B1(n18772), .B2(n18274), .ZN(
        n18776) );
  NOR2_X1 U12252 ( .A1(n18836), .A2(n18986), .ZN(n18977) );
  INV_X1 U12253 ( .A(n13840), .ZN(n15187) );
  INV_X1 U12254 ( .A(n20159), .ZN(n20175) );
  AND2_X1 U12255 ( .A1(n15994), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20178) );
  NAND2_X1 U12256 ( .A1(n20745), .A2(n13451), .ZN(n20152) );
  OR2_X1 U12257 ( .A1(n14427), .A2(n14426), .ZN(n14855) );
  AND2_X2 U12258 ( .A1(n12839), .A2(n14413), .ZN(n20204) );
  AND2_X1 U12259 ( .A1(n16046), .A2(n13072), .ZN(n16044) );
  NAND2_X1 U12260 ( .A1(n13077), .A2(n13076), .ZN(n16043) );
  INV_X1 U12261 ( .A(n16043), .ZN(n14722) );
  CLKBUF_X1 U12262 ( .A(n20227), .Z(n20748) );
  NOR2_X2 U12263 ( .A1(n20259), .A2(n11809), .ZN(n20244) );
  OR2_X1 U12264 ( .A1(n14327), .A2(n20999), .ZN(n13436) );
  XOR2_X1 U12265 ( .A(n14414), .B(n14429), .Z(n14730) );
  INV_X1 U12266 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21042) );
  INV_X1 U12267 ( .A(n16114), .ZN(n16111) );
  OR2_X1 U12268 ( .A1(n16116), .A2(n12883), .ZN(n16120) );
  INV_X1 U12269 ( .A(n14726), .ZN(n9990) );
  INV_X1 U12270 ( .A(n9922), .ZN(n14744) );
  AND2_X1 U12271 ( .A1(n13900), .A2(n12300), .ZN(n9887) );
  NAND2_X1 U12272 ( .A1(n14885), .A2(n9872), .ZN(n9886) );
  NAND2_X1 U12273 ( .A1(n9917), .A2(n16105), .ZN(n16100) );
  NAND2_X1 U12274 ( .A1(n16108), .A2(n16106), .ZN(n9917) );
  INV_X1 U12275 ( .A(n9884), .ZN(n12991) );
  INV_X1 U12276 ( .A(n20518), .ZN(n20601) );
  NAND2_X1 U12277 ( .A1(n11921), .A2(n11905), .ZN(n13125) );
  INV_X1 U12278 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20263) );
  INV_X1 U12279 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13213) );
  CLKBUF_X1 U12280 ( .A(n12170), .Z(n12171) );
  OAI21_X1 U12281 ( .B1(n20333), .B2(n20337), .A(n20332), .ZN(n20355) );
  INV_X1 U12282 ( .A(n20390), .ZN(n20380) );
  OAI21_X1 U12283 ( .B1(n9874), .B2(n20397), .A(n20553), .ZN(n20415) );
  NOR2_X1 U12284 ( .A1(n20423), .A2(n20447), .ZN(n20442) );
  AND2_X1 U12285 ( .A1(n20512), .A2(n13394), .ZN(n20473) );
  OAI21_X1 U12286 ( .B1(n20488), .B2(n20484), .A(n20483), .ZN(n20506) );
  NAND2_X1 U12287 ( .A1(n12156), .A2(n12157), .ZN(n15907) );
  AND2_X1 U12288 ( .A1(n20661), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15905) );
  INV_X1 U12289 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20554) );
  NAND2_X1 U12290 ( .A1(n11104), .A2(n10016), .ZN(n11118) );
  OR2_X1 U12291 ( .A1(n13327), .A2(n13326), .ZN(n19228) );
  INV_X1 U12292 ( .A(n19224), .ZN(n19213) );
  INV_X1 U12293 ( .A(n19178), .ZN(n19223) );
  AND2_X1 U12294 ( .A1(n19380), .A2(n13637), .ZN(n19224) );
  NAND2_X1 U12295 ( .A1(n10188), .A2(n12351), .ZN(n13475) );
  OR2_X1 U12296 ( .A1(n11491), .A2(n11490), .ZN(n13201) );
  OR2_X1 U12297 ( .A1(n11467), .A2(n11466), .ZN(n13199) );
  INV_X1 U12298 ( .A(n10184), .ZN(n10182) );
  AND2_X1 U12299 ( .A1(n12602), .A2(n19304), .ZN(n15159) );
  INV_X1 U12300 ( .A(n15149), .ZN(n15185) );
  NAND2_X1 U12301 ( .A1(n11559), .A2(n14363), .ZN(n16285) );
  NAND2_X1 U12302 ( .A1(n15086), .A2(n15085), .ZN(n15087) );
  NAND2_X1 U12303 ( .A1(n15096), .A2(n15098), .ZN(n15097) );
  OR2_X1 U12304 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  INV_X1 U12305 ( .A(n19280), .ZN(n19299) );
  INV_X1 U12306 ( .A(n16349), .ZN(n19295) );
  AND2_X1 U12307 ( .A1(n19275), .A2(n12788), .ZN(n19280) );
  AND2_X1 U12308 ( .A1(n19306), .A2(n12650), .ZN(n19381) );
  INV_X1 U12309 ( .A(n19381), .ZN(n12725) );
  OAI211_X1 U12310 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n9953), .ZN(n14358)
         );
  NAND2_X1 U12311 ( .A1(n15343), .A2(n9954), .ZN(n9953) );
  OR2_X1 U12312 ( .A1(n15343), .A2(n9957), .ZN(n9955) );
  AND2_X1 U12313 ( .A1(n9956), .A2(n9957), .ZN(n9954) );
  AND2_X1 U12314 ( .A1(n14971), .A2(n14970), .ZN(n15416) );
  NAND2_X1 U12315 ( .A1(n10053), .A2(n10054), .ZN(n15376) );
  OR2_X1 U12316 ( .A1(n16379), .A2(n10057), .ZN(n10053) );
  INV_X1 U12317 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19114) );
  INV_X1 U12318 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19139) );
  INV_X1 U12319 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16432) );
  NAND2_X1 U12320 ( .A1(n19000), .A2(n11633), .ZN(n16445) );
  NOR2_X2 U12321 ( .A1(n19000), .A2(n13331), .ZN(n16435) );
  INV_X1 U12322 ( .A(n16421), .ZN(n16439) );
  OR2_X1 U12323 ( .A1(n15465), .A2(n15446), .ZN(n15441) );
  AND2_X1 U12324 ( .A1(n15034), .A2(n9866), .ZN(n15228) );
  OAI211_X1 U12325 ( .C1(n15351), .C2(n10028), .A(n10025), .B(n10024), .ZN(
        n15521) );
  NAND2_X1 U12326 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  OAI21_X1 U12327 ( .B1(n10030), .B2(n15336), .A(n10026), .ZN(n10025) );
  NAND2_X1 U12328 ( .A1(n15351), .A2(n9848), .ZN(n10024) );
  NAND2_X1 U12329 ( .A1(n10036), .A2(n10035), .ZN(n15346) );
  NAND2_X1 U12330 ( .A1(n10036), .A2(n10032), .ZN(n15523) );
  NAND2_X1 U12331 ( .A1(n16378), .A2(n16382), .ZN(n15595) );
  NAND2_X1 U12332 ( .A1(n9718), .A2(n9843), .ZN(n15640) );
  AND2_X1 U12333 ( .A1(n9718), .A2(n10207), .ZN(n15387) );
  NAND2_X1 U12334 ( .A1(n9718), .A2(n11018), .ZN(n15672) );
  INV_X1 U12335 ( .A(n16474), .ZN(n19400) );
  NAND2_X1 U12336 ( .A1(n9941), .A2(n13377), .ZN(n13384) );
  INV_X1 U12337 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20922) );
  INV_X1 U12338 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20916) );
  INV_X1 U12339 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21022) );
  OR2_X1 U12340 ( .A1(n15705), .A2(n12765), .ZN(n20059) );
  INV_X1 U12341 ( .A(n20053), .ZN(n20050) );
  XNOR2_X1 U12342 ( .A(n12823), .B(n12822), .ZN(n20043) );
  INV_X1 U12343 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20047) );
  NOR2_X1 U12344 ( .A1(n12929), .A2(n11400), .ZN(n13180) );
  NOR2_X1 U12345 ( .A1(n19673), .A2(n19617), .ZN(n19497) );
  INV_X1 U12346 ( .A(n19541), .ZN(n19546) );
  INV_X1 U12347 ( .A(n19585), .ZN(n19604) );
  INV_X1 U12348 ( .A(n19661), .ZN(n19665) );
  OAI21_X1 U12349 ( .B1(n19715), .B2(n19714), .A(n19713), .ZN(n19732) );
  INV_X1 U12350 ( .A(n19760), .ZN(n19765) );
  OR2_X1 U12351 ( .A1(n19776), .A2(n19775), .ZN(n19806) );
  OAI22_X1 U12352 ( .A1(n18316), .A2(n19418), .B1(n16565), .B2(n19420), .ZN(
        n19820) );
  INV_X1 U12353 ( .A(n19836), .ZN(n19844) );
  OAI22_X1 U12354 ( .A1(n20975), .A2(n19418), .B1(n16559), .B2(n19420), .ZN(
        n19867) );
  OAI21_X1 U12355 ( .B1(n19858), .B2(n19857), .A(n19856), .ZN(n19878) );
  INV_X1 U12356 ( .A(n19873), .ZN(n19877) );
  INV_X1 U12357 ( .A(n19688), .ZN(n19908) );
  NAND2_X1 U12358 ( .A1(n19847), .A2(n19846), .ZN(n19930) );
  INV_X1 U12359 ( .A(n19598), .ZN(n19926) );
  INV_X1 U12360 ( .A(n19458), .ZN(n19924) );
  INV_X1 U12361 ( .A(n19802), .ZN(n19934) );
  INV_X1 U12362 ( .A(n19930), .ZN(n19943) );
  INV_X1 U12363 ( .A(n19845), .ZN(n19942) );
  INV_X1 U12364 ( .A(n19895), .ZN(n19944) );
  AND2_X1 U12365 ( .A1(n19431), .A2(n19430), .ZN(n19938) );
  INV_X1 U12366 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20037) );
  NOR2_X1 U12367 ( .A1(n10539), .A2(n18330), .ZN(n16650) );
  AOI21_X1 U12368 ( .B1(n18766), .B2(n18789), .A(n17521), .ZN(n18989) );
  INV_X1 U12369 ( .A(n16507), .ZN(n16520) );
  NAND2_X1 U12370 ( .A1(n16831), .A2(n16879), .ZN(n16822) );
  NOR2_X1 U12371 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16840), .ZN(n16829) );
  NOR2_X1 U12372 ( .A1(n18825), .A2(n16671), .ZN(n17024) );
  INV_X1 U12373 ( .A(n17024), .ZN(n17034) );
  INV_X1 U12374 ( .A(n16999), .ZN(n17043) );
  INV_X1 U12375 ( .A(n17033), .ZN(n17044) );
  NOR2_X1 U12376 ( .A1(n16757), .A2(n17097), .ZN(n17102) );
  NOR2_X1 U12377 ( .A1(n17152), .A2(n17151), .ZN(n17136) );
  NOR3_X1 U12378 ( .A1(n18324), .A2(n18319), .A3(n15938), .ZN(n17362) );
  INV_X1 U12379 ( .A(n17362), .ZN(n17365) );
  INV_X1 U12380 ( .A(n17383), .ZN(n17379) );
  INV_X1 U12381 ( .A(n17407), .ZN(n17402) );
  NAND2_X1 U12382 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17402), .ZN(n17401) );
  NOR2_X1 U12383 ( .A1(n17456), .A2(n17411), .ZN(n17408) );
  NOR2_X1 U12384 ( .A1(n17630), .A2(n17458), .ZN(n17451) );
  NAND2_X1 U12385 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17451), .ZN(n17450) );
  INV_X1 U12386 ( .A(n17423), .ZN(n17448) );
  AOI211_X1 U12387 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n10323), .B(n10322), .ZN(n17488) );
  INV_X1 U12388 ( .A(n10496), .ZN(n17492) );
  INV_X1 U12389 ( .A(n10492), .ZN(n17502) );
  AND2_X1 U12390 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17505), .ZN(n17510) );
  INV_X1 U12391 ( .A(n17514), .ZN(n17511) );
  OR4_X2 U12392 ( .A1(n10337), .A2(n9980), .A3(n10336), .A4(n10339), .ZN(
        n17993) );
  NAND2_X1 U12393 ( .A1(n10338), .A2(n9981), .ZN(n9980) );
  NOR2_X1 U12394 ( .A1(n17506), .A2(n18804), .ZN(n17514) );
  OAI211_X1 U12395 ( .C1(n18979), .C2(n18324), .A(n17580), .B(n17579), .ZN(
        n17619) );
  INV_X1 U12396 ( .A(n17629), .ZN(n17620) );
  NOR2_X1 U12398 ( .A1(n17626), .A2(n18324), .ZN(n17627) );
  NAND2_X1 U12399 ( .A1(n17786), .A2(n9786), .ZN(n17737) );
  NAND2_X1 U12400 ( .A1(n17786), .A2(n9783), .ZN(n17773) );
  NAND2_X1 U12401 ( .A1(n16536), .A2(n17994), .ZN(n17898) );
  INV_X1 U12402 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17810) );
  OAI22_X1 U12403 ( .A1(n17691), .A2(n17835), .B1(n18000), .B2(n18162), .ZN(
        n17841) );
  INV_X1 U12404 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17909) );
  NAND2_X1 U12405 ( .A1(n9964), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17940) );
  NOR2_X1 U12406 ( .A1(n18970), .A2(n16652), .ZN(n17985) );
  NOR2_X2 U12407 ( .A1(n16652), .A2(n18324), .ZN(n17994) );
  INV_X1 U12408 ( .A(n9775), .ZN(n18000) );
  NAND2_X1 U12409 ( .A1(n10367), .A2(n9970), .ZN(n15862) );
  NOR2_X1 U12410 ( .A1(n17492), .A2(n10349), .ZN(n16548) );
  NOR2_X1 U12411 ( .A1(n17743), .A2(n10363), .ZN(n17694) );
  NOR2_X1 U12412 ( .A1(n18780), .A2(n18803), .ZN(n18290) );
  INV_X1 U12413 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18986) );
  INV_X1 U12414 ( .A(n10157), .ZN(n17775) );
  NAND2_X1 U12415 ( .A1(n17783), .A2(n9778), .ZN(n17776) );
  NAND2_X1 U12416 ( .A1(n18290), .A2(n18805), .ZN(n18145) );
  AND2_X1 U12417 ( .A1(n17815), .A2(n17870), .ZN(n18213) );
  INV_X1 U12418 ( .A(n10153), .ZN(n17953) );
  NOR2_X1 U12419 ( .A1(n18301), .A2(n18298), .ZN(n18291) );
  NOR2_X1 U12420 ( .A1(n15848), .A2(n18794), .ZN(n18805) );
  INV_X1 U12421 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18565) );
  INV_X1 U12422 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18818) );
  INV_X1 U12423 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18327) );
  INV_X1 U12424 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20925) );
  INV_X1 U12425 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18355) );
  INV_X1 U12426 ( .A(n18977), .ZN(n18832) );
  OAI21_X1 U12429 ( .B1(n14386), .B2(n16259), .A(n9894), .ZN(P1_U3000) );
  NOR2_X1 U12430 ( .A1(n9898), .A2(n12087), .ZN(n9897) );
  NAND2_X1 U12431 ( .A1(n12310), .A2(n14380), .ZN(n9895) );
  AOI21_X1 U12432 ( .B1(n16274), .B2(n16282), .A(n16281), .ZN(n16283) );
  OAI21_X1 U12433 ( .B1(n12604), .B2(n12766), .A(n12603), .ZN(n12605) );
  NOR2_X1 U12434 ( .A1(n12982), .A2(n10182), .ZN(n10218) );
  OAI21_X1 U12435 ( .B1(n15431), .B2(n16427), .A(n11662), .ZN(n11663) );
  NAND2_X1 U12436 ( .A1(n14371), .A2(n10114), .ZN(n10002) );
  AND2_X1 U12437 ( .A1(n11611), .A2(n11610), .ZN(n11612) );
  OR2_X1 U12438 ( .A1(n15578), .A2(n16477), .ZN(n10189) );
  NAND2_X1 U12439 ( .A1(n10191), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10190) );
  OAI211_X1 U12440 ( .C1(n16502), .C2(n18305), .A(n10551), .B(n10550), .ZN(
        n10552) );
  OR2_X1 U12441 ( .A1(n15925), .A2(n16508), .ZN(n10163) );
  AND2_X1 U12442 ( .A1(n10647), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10833) );
  NAND2_X1 U12443 ( .A1(n15343), .A2(n9810), .ZN(n15308) );
  NAND2_X1 U12444 ( .A1(n15343), .A2(n9809), .ZN(n15278) );
  AND2_X1 U12445 ( .A1(n9800), .A2(n14565), .ZN(n9776) );
  AND2_X2 U12446 ( .A1(n10786), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10863) );
  AND2_X1 U12447 ( .A1(n9976), .A2(n9859), .ZN(n9778) );
  NOR2_X1 U12448 ( .A1(n14021), .A2(n10146), .ZN(n14518) );
  AND2_X1 U12449 ( .A1(n11795), .A2(n13158), .ZN(n11819) );
  NAND2_X1 U12450 ( .A1(n14141), .A2(n10141), .ZN(n9779) );
  OR2_X1 U12451 ( .A1(n13270), .A2(n13269), .ZN(n9780) );
  AND2_X1 U12452 ( .A1(n9716), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9781) );
  AND2_X1 U12453 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9783) );
  NOR2_X1 U12454 ( .A1(n10353), .A2(n10352), .ZN(n9784) );
  AND4_X1 U12455 ( .A1(n11748), .A2(n11816), .A3(n11715), .A4(n11716), .ZN(
        n11808) );
  INV_X1 U12456 ( .A(n19421), .ZN(n10667) );
  AND2_X1 U12457 ( .A1(n9783), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9785) );
  AND2_X1 U12458 ( .A1(n9785), .A2(n9959), .ZN(n9786) );
  NAND2_X1 U12459 ( .A1(n12455), .A2(n12478), .ZN(n9787) );
  OR3_X1 U12460 ( .A1(n14498), .A2(n10067), .A3(n12267), .ZN(n9788) );
  AND4_X1 U12461 ( .A1(n10107), .A2(n10109), .A3(n10111), .A4(n13778), .ZN(
        n9789) );
  AND2_X1 U12462 ( .A1(n10688), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9790) );
  AND2_X1 U12463 ( .A1(n10010), .A2(n11013), .ZN(n9791) );
  AND3_X1 U12464 ( .A1(n10558), .A2(n10557), .A3(n13590), .ZN(n9792) );
  AND2_X1 U12465 ( .A1(n10064), .A2(n10062), .ZN(n9793) );
  AND2_X1 U12466 ( .A1(n11008), .A2(n9841), .ZN(n9794) );
  NOR2_X1 U12467 ( .A1(n15659), .A2(n15660), .ZN(n9795) );
  AND2_X1 U12468 ( .A1(n12351), .A2(n10187), .ZN(n9796) );
  NOR2_X1 U12469 ( .A1(n10685), .A2(n10684), .ZN(n11364) );
  AND2_X1 U12470 ( .A1(n10096), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9797) );
  OR2_X1 U12471 ( .A1(n17871), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9798) );
  AND2_X1 U12472 ( .A1(n9965), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9799) );
  NOR2_X1 U12473 ( .A1(n10061), .A2(n14574), .ZN(n9800) );
  AND2_X1 U12474 ( .A1(n10188), .A2(n9796), .ZN(n9801) );
  AND2_X1 U12475 ( .A1(n13807), .A2(n13557), .ZN(n9802) );
  AND2_X1 U12476 ( .A1(n9799), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9803) );
  AND2_X1 U12477 ( .A1(n10012), .A2(n9853), .ZN(n9804) );
  INV_X1 U12478 ( .A(n15085), .ZN(n10171) );
  OR2_X1 U12479 ( .A1(n11495), .A2(n13312), .ZN(n11496) );
  AND2_X1 U12480 ( .A1(n10092), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9805) );
  AND2_X1 U12481 ( .A1(n10099), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9806) );
  AND2_X1 U12482 ( .A1(n10014), .A2(n15114), .ZN(n9807) );
  AND2_X1 U12483 ( .A1(n16450), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9808) );
  AND2_X2 U12484 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13206) );
  AND2_X1 U12485 ( .A1(n10212), .A2(n11251), .ZN(n9809) );
  AND2_X1 U12486 ( .A1(n15473), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9810) );
  AND2_X1 U12487 ( .A1(n9809), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9811) );
  INV_X1 U12488 ( .A(n10676), .ZN(n10776) );
  AND2_X1 U12489 ( .A1(n10974), .A2(n10973), .ZN(n9812) );
  OR2_X2 U12490 ( .A1(n10240), .A2(n18795), .ZN(n9814) );
  NAND2_X1 U12491 ( .A1(n11036), .A2(n9804), .ZN(n9815) );
  OR2_X1 U12492 ( .A1(n14605), .A2(n14522), .ZN(n9816) );
  BUF_X1 U12493 ( .A(n11702), .Z(n14126) );
  AND2_X2 U12494 ( .A1(n9772), .A2(n13590), .ZN(n10779) );
  AND2_X1 U12495 ( .A1(n10202), .A2(n15305), .ZN(n15285) );
  NOR2_X1 U12496 ( .A1(n14021), .A2(n14020), .ZN(n14601) );
  AND2_X1 U12497 ( .A1(n15343), .A2(n10212), .ZN(n15284) );
  OR2_X1 U12498 ( .A1(n14021), .A2(n10144), .ZN(n9817) );
  INV_X1 U12499 ( .A(n10726), .ZN(n10741) );
  INV_X1 U12500 ( .A(n9925), .ZN(n15383) );
  AND4_X1 U12501 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n9818) );
  NOR2_X1 U12502 ( .A1(n14021), .A2(n10143), .ZN(n14587) );
  AND2_X1 U12503 ( .A1(n14578), .A2(n14577), .ZN(n14571) );
  OR2_X1 U12504 ( .A1(n12318), .A2(n19231), .ZN(n10764) );
  OAI21_X1 U12505 ( .B1(n10004), .B2(n10003), .A(n9944), .ZN(n15268) );
  NAND2_X1 U12506 ( .A1(n9741), .A2(n15326), .ZN(n15611) );
  NOR2_X1 U12507 ( .A1(n11129), .A2(n11128), .ZN(n9819) );
  NOR2_X1 U12508 ( .A1(n10357), .A2(n9974), .ZN(n9820) );
  INV_X2 U12509 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U12510 ( .A1(n9949), .A2(n11245), .ZN(n16410) );
  AND4_X1 U12511 ( .A1(n11102), .A2(n15329), .A3(n15333), .A4(n15550), .ZN(
        n9821) );
  NOR3_X1 U12512 ( .A1(n11145), .A2(n11023), .A3(n14370), .ZN(n9822) );
  NAND2_X1 U12513 ( .A1(n9999), .A2(n9777), .ZN(n14806) );
  INV_X4 U12514 ( .A(n17300), .ZN(n17323) );
  NAND2_X1 U12515 ( .A1(n10021), .A2(n10020), .ZN(n10734) );
  XNOR2_X1 U12516 ( .A(n11247), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16411) );
  INV_X1 U12517 ( .A(n16411), .ZN(n9948) );
  AND2_X1 U12518 ( .A1(n9778), .A2(n18106), .ZN(n9823) );
  OR2_X1 U12519 ( .A1(n16106), .A2(n9918), .ZN(n9824) );
  NAND2_X1 U12520 ( .A1(n12344), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9825) );
  INV_X1 U12521 ( .A(n10229), .ZN(n10119) );
  AND2_X1 U12522 ( .A1(n10127), .A2(n11860), .ZN(n9826) );
  XNOR2_X1 U12523 ( .A(n11632), .B(n11631), .ZN(n16274) );
  AND2_X1 U12524 ( .A1(n16098), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9827) );
  OR2_X1 U12525 ( .A1(n19474), .A2(n10805), .ZN(n9828) );
  NAND2_X1 U12526 ( .A1(n11134), .A2(n15294), .ZN(n9829) );
  AND2_X1 U12527 ( .A1(n10657), .A2(n10656), .ZN(n10669) );
  AND2_X1 U12528 ( .A1(n14141), .A2(n10139), .ZN(n14480) );
  AND3_X1 U12529 ( .A1(n11248), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11621), .ZN(n9830) );
  NAND2_X1 U12530 ( .A1(n14141), .A2(n14140), .ZN(n14504) );
  AND2_X1 U12531 ( .A1(n12072), .A2(n10000), .ZN(n9831) );
  NAND2_X1 U12532 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10325), .ZN(
        n9832) );
  OR2_X1 U12533 ( .A1(n12005), .A2(n11982), .ZN(n9833) );
  AND2_X1 U12534 ( .A1(n11130), .A2(n15305), .ZN(n10201) );
  AND2_X1 U12535 ( .A1(n9990), .A2(n9988), .ZN(n9834) );
  AND2_X1 U12536 ( .A1(n9791), .A2(n13659), .ZN(n9835) );
  AND2_X1 U12537 ( .A1(n10561), .A2(n10560), .ZN(n9836) );
  INV_X1 U12538 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10009) );
  INV_X1 U12539 ( .A(n12243), .ZN(n10059) );
  XNOR2_X1 U12540 ( .A(n16506), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16865) );
  NAND2_X1 U12541 ( .A1(n16548), .A2(n16536), .ZN(n17897) );
  NAND2_X1 U12542 ( .A1(n17786), .A2(n9785), .ZN(n9837) );
  INV_X1 U12543 ( .A(n13315), .ZN(n10103) );
  INV_X1 U12544 ( .A(n12170), .ZN(n9907) );
  OR2_X1 U12545 ( .A1(n15660), .A2(n10085), .ZN(n9838) );
  NOR2_X1 U12546 ( .A1(n15596), .A2(n15579), .ZN(n13837) );
  NAND3_X1 U12547 ( .A1(n13522), .A2(n13523), .A3(n9802), .ZN(n9839) );
  AND2_X1 U12548 ( .A1(n13322), .A2(n10096), .ZN(n9840) );
  AND2_X1 U12549 ( .A1(n16413), .A2(n16414), .ZN(n9841) );
  AND2_X1 U12550 ( .A1(n15167), .A2(n10122), .ZN(n9842) );
  AND2_X1 U12551 ( .A1(n15385), .A2(n10207), .ZN(n9843) );
  OR2_X1 U12552 ( .A1(n10086), .A2(n15556), .ZN(n9844) );
  AND2_X1 U12553 ( .A1(n13421), .A2(n13420), .ZN(n13419) );
  AND2_X1 U12554 ( .A1(n15124), .A2(n15120), .ZN(n15020) );
  NAND2_X1 U12555 ( .A1(n15034), .A2(n10080), .ZN(n9845) );
  AND2_X1 U12556 ( .A1(n14591), .A2(n9800), .ZN(n9846) );
  INV_X1 U12557 ( .A(n15326), .ZN(n9938) );
  OR2_X1 U12558 ( .A1(n15659), .A2(n9838), .ZN(n13311) );
  NOR2_X1 U12559 ( .A1(n14498), .A2(n10066), .ZN(n10068) );
  NAND2_X1 U12560 ( .A1(n13082), .A2(n13081), .ZN(n13088) );
  AND2_X1 U12561 ( .A1(n10178), .A2(n9787), .ZN(n9847) );
  NAND2_X1 U12562 ( .A1(n15113), .A2(n15112), .ZN(n15111) );
  AND2_X1 U12563 ( .A1(n10032), .A2(n15336), .ZN(n9848) );
  NAND2_X1 U12564 ( .A1(n11229), .A2(n11228), .ZN(n13771) );
  AND2_X1 U12565 ( .A1(n9842), .A2(n10121), .ZN(n9849) );
  NAND2_X1 U12566 ( .A1(n15034), .A2(n15036), .ZN(n15035) );
  NAND2_X1 U12567 ( .A1(n10198), .A2(n9928), .ZN(n11167) );
  AND2_X1 U12568 ( .A1(n10070), .A2(n14603), .ZN(n9850) );
  AND2_X1 U12569 ( .A1(n9993), .A2(n9988), .ZN(n9851) );
  NAND2_X1 U12570 ( .A1(n11375), .A2(n11045), .ZN(n9852) );
  OR2_X1 U12571 ( .A1(n13659), .A2(n11043), .ZN(n9853) );
  NAND2_X1 U12572 ( .A1(n15171), .A2(n15167), .ZN(n15155) );
  INV_X1 U12573 ( .A(n14563), .ZN(n14140) );
  AND2_X1 U12574 ( .A1(n10102), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9854) );
  NAND2_X1 U12575 ( .A1(n14305), .A2(n14304), .ZN(n9855) );
  OR2_X1 U12576 ( .A1(n9844), .A2(n13886), .ZN(n9856) );
  NOR2_X1 U12577 ( .A1(n10210), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9857) );
  NAND2_X1 U12578 ( .A1(n11104), .A2(n10014), .ZN(n10018) );
  INV_X1 U12579 ( .A(n10033), .ZN(n10032) );
  NAND2_X1 U12580 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  INV_X1 U12581 ( .A(n11496), .ZN(n10084) );
  AND2_X1 U12582 ( .A1(n10149), .A2(n14414), .ZN(n9858) );
  OR2_X1 U12583 ( .A1(n17897), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9859) );
  AND2_X1 U12584 ( .A1(n9804), .A2(n9852), .ZN(n9860) );
  AND2_X1 U12585 ( .A1(n9786), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9861) );
  AND2_X1 U12586 ( .A1(n9843), .A2(n10215), .ZN(n9862) );
  INV_X1 U12587 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15396) );
  INV_X1 U12588 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U12589 ( .A1(n10180), .A2(n13174), .ZN(n12982) );
  NOR2_X1 U12590 ( .A1(n12982), .A2(n12346), .ZN(n12968) );
  NAND2_X1 U12591 ( .A1(n12200), .A2(n12199), .ZN(n16254) );
  INV_X1 U12592 ( .A(n16254), .ZN(n10063) );
  NOR2_X1 U12593 ( .A1(n16462), .A2(n16463), .ZN(n15673) );
  OR2_X1 U12594 ( .A1(n13060), .A2(n10119), .ZN(n13114) );
  INV_X1 U12595 ( .A(n9883), .ZN(n14898) );
  OAI211_X1 U12596 ( .C1(n13901), .C2(n9887), .A(n9886), .B(n14919), .ZN(n9883) );
  INV_X1 U12597 ( .A(n11023), .ZN(n11621) );
  AND2_X1 U12598 ( .A1(n14990), .A2(n10099), .ZN(n9863) );
  INV_X1 U12599 ( .A(n13730), .ZN(n10187) );
  INV_X1 U12600 ( .A(n14492), .ZN(n10142) );
  INV_X1 U12601 ( .A(n9975), .ZN(n9974) );
  NOR2_X1 U12602 ( .A1(n18110), .A2(n18221), .ZN(n9975) );
  INV_X1 U12603 ( .A(n11037), .ZN(n10013) );
  AND2_X1 U12604 ( .A1(n14978), .A2(n10092), .ZN(n9864) );
  OR2_X1 U12605 ( .A1(n11654), .A2(n10124), .ZN(n9865) );
  AND2_X1 U12606 ( .A1(n10080), .A2(n15238), .ZN(n9866) );
  INV_X1 U12607 ( .A(n16477), .ZN(n19395) );
  AND2_X1 U12608 ( .A1(n9776), .A2(n10060), .ZN(n9867) );
  OR2_X1 U12609 ( .A1(n13378), .A2(n10110), .ZN(n9868) );
  OR2_X1 U12610 ( .A1(n17897), .A2(n18002), .ZN(n9869) );
  NAND2_X1 U12611 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9870) );
  NAND2_X1 U12612 ( .A1(n9910), .A2(n9909), .ZN(n12174) );
  AND2_X1 U12613 ( .A1(n17673), .A2(n9799), .ZN(n9871) );
  INV_X1 U12614 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n9961) );
  INV_X1 U12615 ( .A(n14582), .ZN(n10061) );
  OR2_X1 U12616 ( .A1(n13902), .A2(n16159), .ZN(n9872) );
  INV_X1 U12617 ( .A(n15092), .ZN(n10176) );
  INV_X1 U12618 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14525) );
  OR2_X1 U12619 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9873) );
  INV_X1 U12620 ( .A(n10174), .ZN(n10173) );
  NAND2_X1 U12621 ( .A1(n15098), .A2(n10176), .ZN(n10174) );
  NOR2_X1 U12622 ( .A1(n20545), .A2(n20419), .ZN(n9874) );
  NOR2_X1 U12623 ( .A1(n20545), .A2(n20598), .ZN(n9875) );
  OR2_X1 U12624 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U12625 ( .A1(n10211), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9877) );
  AND2_X1 U12626 ( .A1(n16160), .A2(n16164), .ZN(n9878) );
  AND2_X1 U12627 ( .A1(n10213), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9879) );
  INV_X1 U12628 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17939) );
  INV_X1 U12629 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10214) );
  INV_X1 U12630 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9967) );
  INV_X1 U12631 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10101) );
  INV_X1 U12632 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10097) );
  AND2_X1 U12633 ( .A1(n15316), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9880) );
  INV_X1 U12634 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9988) );
  INV_X1 U12635 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10093) );
  INV_X1 U12636 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9960) );
  INV_X1 U12637 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10094) );
  INV_X1 U12638 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9957) );
  INV_X1 U12639 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10185) );
  NAND3_X2 U12640 ( .A1(n18987), .A2(n18974), .A3(n18986), .ZN(n18199) );
  AOI22_X2 U12641 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19435), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19434), .ZN(n19948) );
  NOR3_X2 U12642 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20599), .A3(
        n20598), .ZN(n13712) );
  AOI22_X2 U12643 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19435), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19434), .ZN(n19931) );
  NOR2_X2 U12644 ( .A1(n15187), .A2(n13658), .ZN(n19434) );
  NOR2_X4 U12645 ( .A1(n18808), .A2(n18643), .ZN(n18761) );
  NOR2_X2 U12646 ( .A1(n13680), .A2(n13671), .ZN(n20644) );
  XNOR2_X2 U12647 ( .A(n9881), .B(n10936), .ZN(n13280) );
  NAND2_X1 U12648 ( .A1(n10804), .A2(n10803), .ZN(n9881) );
  INV_X1 U12649 ( .A(n13768), .ZN(n11233) );
  NAND2_X1 U12650 ( .A1(n11242), .A2(n11244), .ZN(n11245) );
  NOR2_X1 U12651 ( .A1(n12304), .A2(n14910), .ZN(n9898) );
  NAND2_X2 U12652 ( .A1(n13679), .A2(n12129), .ZN(n11802) );
  INV_X2 U12653 ( .A(n11857), .ZN(n13679) );
  NAND2_X2 U12654 ( .A1(n11714), .A2(n10233), .ZN(n11857) );
  NAND2_X1 U12655 ( .A1(n13080), .A2(n13079), .ZN(n12020) );
  XNOR2_X1 U12656 ( .A(n12018), .B(n13239), .ZN(n13080) );
  NAND2_X1 U12657 ( .A1(n9903), .A2(n12012), .ZN(n12018) );
  NAND2_X1 U12658 ( .A1(n13038), .A2(n13039), .ZN(n9903) );
  INV_X1 U12659 ( .A(n9904), .ZN(n11884) );
  XNOR2_X2 U12660 ( .A(n11880), .B(n11876), .ZN(n9904) );
  NAND2_X1 U12661 ( .A1(n12841), .A2(n9904), .ZN(n20513) );
  NAND3_X1 U12662 ( .A1(n11921), .A2(n11905), .A3(n11886), .ZN(n9905) );
  NAND2_X1 U12663 ( .A1(n9905), .A2(n9833), .ZN(n11919) );
  NAND2_X1 U12664 ( .A1(n12862), .A2(n10232), .ZN(n12173) );
  INV_X1 U12665 ( .A(n12960), .ZN(n9910) );
  INV_X1 U12666 ( .A(n12112), .ZN(n12862) );
  AND2_X1 U12667 ( .A1(n11748), .A2(n11816), .ZN(n9913) );
  NAND2_X1 U12668 ( .A1(n11808), .A2(n9914), .ZN(n12166) );
  NAND2_X2 U12669 ( .A1(n9916), .A2(n9915), .ZN(n13816) );
  AOI21_X2 U12670 ( .B1(n9782), .B2(n9918), .A(n9827), .ZN(n9915) );
  NAND2_X1 U12671 ( .A1(n12073), .A2(n9920), .ZN(n9919) );
  NAND2_X2 U12672 ( .A1(n12081), .A2(n14801), .ZN(n14741) );
  NAND2_X2 U12673 ( .A1(n15666), .A2(n9924), .ZN(n9925) );
  NOR2_X2 U12674 ( .A1(n9925), .A2(n9877), .ZN(n15359) );
  NAND2_X1 U12675 ( .A1(n9931), .A2(n9929), .ZN(n10697) );
  INV_X1 U12676 ( .A(n10685), .ZN(n9931) );
  NAND4_X1 U12677 ( .A1(n10697), .A2(n10677), .A3(n13639), .A4(n12758), .ZN(
        n9932) );
  NAND2_X2 U12678 ( .A1(n10666), .A2(n13746), .ZN(n12758) );
  NAND2_X1 U12679 ( .A1(n11042), .A2(n9936), .ZN(n9935) );
  INV_X1 U12680 ( .A(n10933), .ZN(n9941) );
  NAND2_X1 U12681 ( .A1(n9942), .A2(n10001), .ZN(P2_U3015) );
  OR2_X2 U12682 ( .A1(n14373), .A2(n16477), .ZN(n9942) );
  OAI21_X2 U12683 ( .B1(n11617), .B2(n11616), .A(n11615), .ZN(n9943) );
  NAND2_X2 U12684 ( .A1(n10862), .A2(n10861), .ZN(n10936) );
  NAND2_X1 U12685 ( .A1(n11561), .A2(n19421), .ZN(n9951) );
  NOR2_X2 U12686 ( .A1(n17911), .A2(n9784), .ZN(n10357) );
  NAND3_X1 U12687 ( .A1(n9972), .A2(n9971), .A3(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12688 ( .A1(n17911), .A2(n9975), .ZN(n9972) );
  INV_X1 U12689 ( .A(n10357), .ZN(n9973) );
  INV_X2 U12690 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18944) );
  NAND2_X2 U12691 ( .A1(n9984), .A2(n12042), .ZN(n16108) );
  NAND2_X1 U12692 ( .A1(n16113), .A2(n16112), .ZN(n9984) );
  INV_X2 U12693 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U12694 ( .A1(n12165), .A2(n14944), .ZN(n11806) );
  NAND3_X1 U12695 ( .A1(n11821), .A2(n11803), .A3(n13679), .ZN(n12165) );
  XNOR2_X2 U12696 ( .A(n11989), .B(n11990), .ZN(n12848) );
  NAND2_X1 U12697 ( .A1(n9989), .A2(n9993), .ZN(n9991) );
  NAND2_X2 U12698 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  AND2_X2 U12699 ( .A1(n9994), .A2(n9991), .ZN(n14726) );
  NAND2_X1 U12700 ( .A1(n12073), .A2(n9831), .ZN(n9999) );
  NOR2_X1 U12701 ( .A1(n10201), .A2(n9876), .ZN(n10003) );
  OAI21_X1 U12702 ( .B1(n10802), .B2(n10006), .A(n10894), .ZN(n10895) );
  AOI21_X1 U12703 ( .B1(n10008), .B2(n11520), .A(n10007), .ZN(n11401) );
  NAND2_X1 U12704 ( .A1(n11377), .A2(n10008), .ZN(n10803) );
  NAND2_X1 U12705 ( .A1(n11006), .A2(n9791), .ZN(n11019) );
  NAND2_X1 U12706 ( .A1(n9835), .A2(n11006), .ZN(n11125) );
  INV_X1 U12707 ( .A(n10018), .ZN(n11127) );
  NAND2_X1 U12708 ( .A1(n11365), .A2(n20077), .ZN(n10655) );
  NAND2_X1 U12709 ( .A1(n10640), .A2(n11201), .ZN(n11365) );
  NOR2_X2 U12710 ( .A1(n10019), .A2(n15080), .ZN(n10938) );
  NOR2_X2 U12711 ( .A1(n10019), .A2(n9774), .ZN(n10940) );
  NAND2_X1 U12712 ( .A1(n10708), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10021) );
  NAND2_X1 U12713 ( .A1(n10707), .A2(n10688), .ZN(n10022) );
  INV_X1 U12714 ( .A(n10708), .ZN(n10023) );
  NAND2_X1 U12715 ( .A1(n10734), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10675) );
  OAI211_X1 U12716 ( .C1(n10714), .C2(n9740), .A(n10741), .B(n10728), .ZN(
        n10718) );
  OAI211_X1 U12717 ( .C1(n10727), .C2(n10726), .A(n10715), .B(n10037), .ZN(
        n10041) );
  INV_X1 U12718 ( .A(n10038), .ZN(n10037) );
  OAI21_X1 U12719 ( .B1(n10740), .B2(n10726), .A(n10729), .ZN(n10038) );
  NAND2_X1 U12720 ( .A1(n10040), .A2(n10039), .ZN(n10717) );
  OAI21_X1 U12721 ( .B1(n10728), .B2(n10725), .A(n10740), .ZN(n10039) );
  NAND2_X1 U12722 ( .A1(n10713), .A2(n10714), .ZN(n10040) );
  NAND2_X1 U12723 ( .A1(n10042), .A2(n10041), .ZN(n11258) );
  NAND4_X1 U12724 ( .A1(n10738), .A2(n10716), .A3(n10717), .A4(n10718), .ZN(
        n10042) );
  NAND2_X2 U12725 ( .A1(n10045), .A2(n10043), .ZN(n10662) );
  NAND2_X1 U12726 ( .A1(n10044), .A2(n13590), .ZN(n10043) );
  NAND4_X1 U12727 ( .A1(n10576), .A2(n10575), .A3(n10573), .A4(n10574), .ZN(
        n10044) );
  NAND2_X1 U12728 ( .A1(n10046), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10045) );
  NAND4_X1 U12729 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10046) );
  NAND2_X1 U12730 ( .A1(n16379), .A2(n10051), .ZN(n10050) );
  NAND2_X2 U12731 ( .A1(n9748), .A2(n11403), .ZN(n11225) );
  INV_X1 U12732 ( .A(n11225), .ZN(n10978) );
  NAND3_X1 U12733 ( .A1(n12181), .A2(n13463), .A3(n12182), .ZN(n12186) );
  NAND2_X1 U12734 ( .A1(n10059), .A2(n15983), .ZN(n12241) );
  NAND2_X1 U12735 ( .A1(n10059), .A2(n12255), .ZN(n12259) );
  NAND2_X1 U12736 ( .A1(n10059), .A2(n12269), .ZN(n12273) );
  NAND2_X1 U12737 ( .A1(n10059), .A2(n13870), .ZN(n12219) );
  NAND2_X1 U12738 ( .A1(n10059), .A2(n16017), .ZN(n12231) );
  NAND2_X1 U12739 ( .A1(n10059), .A2(n14568), .ZN(n12253) );
  NAND2_X1 U12740 ( .A1(n10059), .A2(n14558), .ZN(n12264) );
  NAND2_X1 U12741 ( .A1(n10063), .A2(n9793), .ZN(n16219) );
  INV_X1 U12742 ( .A(n10068), .ZN(n14441) );
  INV_X1 U12743 ( .A(n14462), .ZN(n10069) );
  NOR2_X1 U12744 ( .A1(n12928), .A2(n12927), .ZN(n12929) );
  NOR2_X1 U12745 ( .A1(n11400), .A2(n10078), .ZN(n10077) );
  NAND2_X1 U12746 ( .A1(n15211), .A2(n10090), .ZN(n14995) );
  AND2_X1 U12747 ( .A1(n15211), .A2(n15201), .ZN(n15203) );
  INV_X1 U12748 ( .A(n10676), .ZN(n11369) );
  NAND2_X1 U12749 ( .A1(n13746), .A2(n10676), .ZN(n10679) );
  NAND2_X4 U12750 ( .A1(n10106), .A2(n10105), .ZN(n20077) );
  INV_X1 U12751 ( .A(n13778), .ZN(n10110) );
  NAND2_X1 U12752 ( .A1(n10108), .A2(n10111), .ZN(n13379) );
  NOR2_X1 U12753 ( .A1(n13379), .A2(n13378), .ZN(n13777) );
  NAND2_X1 U12754 ( .A1(n10113), .A2(n10112), .ZN(n10111) );
  NAND2_X1 U12755 ( .A1(n16274), .A2(n16475), .ZN(n10114) );
  NAND2_X1 U12756 ( .A1(n15171), .A2(n10120), .ZN(n15039) );
  NOR2_X1 U12757 ( .A1(n15100), .A2(n15099), .ZN(n10125) );
  INV_X1 U12758 ( .A(n11626), .ZN(n14970) );
  NAND2_X1 U12759 ( .A1(n11861), .A2(n11860), .ZN(n10126) );
  AOI21_X2 U12760 ( .B1(n9777), .B2(n10136), .A(n10134), .ZN(n10133) );
  AND3_X2 U12761 ( .A1(n13522), .A2(n13523), .A3(n10137), .ZN(n13921) );
  NAND3_X1 U12762 ( .A1(n13522), .A2(n13523), .A3(n13557), .ZN(n13808) );
  NAND2_X1 U12763 ( .A1(n14141), .A2(n10138), .ZN(n14465) );
  NAND2_X1 U12764 ( .A1(n11943), .A2(n13124), .ZN(n12022) );
  INV_X1 U12765 ( .A(n12033), .ZN(n11968) );
  AND2_X1 U12766 ( .A1(n14451), .A2(n10148), .ZN(n14428) );
  AND2_X1 U12767 ( .A1(n14451), .A2(n10149), .ZN(n14429) );
  NAND2_X1 U12768 ( .A1(n14451), .A2(n9858), .ZN(n14334) );
  NAND2_X1 U12769 ( .A1(n14451), .A2(n14258), .ZN(n14439) );
  NOR2_X2 U12770 ( .A1(n10367), .A2(n18009), .ZN(n17650) );
  NAND2_X2 U12771 ( .A1(n17665), .A2(n10152), .ZN(n10367) );
  NAND2_X1 U12772 ( .A1(n10155), .A2(n10154), .ZN(n17729) );
  OR2_X1 U12773 ( .A1(n17728), .A2(n17897), .ZN(n10154) );
  NAND3_X1 U12774 ( .A1(n10156), .A2(n9823), .A3(n17783), .ZN(n10155) );
  INV_X1 U12775 ( .A(n17728), .ZN(n10156) );
  NAND2_X1 U12776 ( .A1(n9823), .A2(n17783), .ZN(n10157) );
  NAND3_X1 U12777 ( .A1(n10282), .A2(n10161), .A3(n10160), .ZN(n10159) );
  AOI21_X1 U12778 ( .B1(n16515), .B2(n18203), .A(n10163), .ZN(n15926) );
  INV_X1 U12779 ( .A(n15923), .ZN(n10165) );
  INV_X1 U12780 ( .A(n15922), .ZN(n10166) );
  INV_X2 U12781 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18951) );
  INV_X2 U12782 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20969) );
  XNOR2_X2 U12783 ( .A(n11258), .B(n11261), .ZN(n12318) );
  NAND3_X1 U12784 ( .A1(n10718), .A2(n10716), .A3(n10717), .ZN(n10739) );
  NAND2_X1 U12785 ( .A1(n15096), .A2(n10169), .ZN(n10168) );
  NAND3_X1 U12786 ( .A1(n10168), .A2(n10167), .A3(n12582), .ZN(n12600) );
  INV_X1 U12787 ( .A(n10178), .ZN(n15126) );
  INV_X1 U12788 ( .A(n13178), .ZN(n10181) );
  NAND3_X1 U12789 ( .A1(n10190), .A2(n15577), .A3(n10189), .ZN(P2_U3029) );
  INV_X1 U12790 ( .A(n13373), .ZN(n11227) );
  NAND2_X1 U12791 ( .A1(n13373), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11226) );
  NAND2_X1 U12792 ( .A1(n10658), .A2(n10198), .ZN(n10665) );
  NAND2_X1 U12793 ( .A1(n9719), .A2(n10201), .ZN(n10199) );
  OR2_X2 U12794 ( .A1(n15304), .A2(n15306), .ZN(n10202) );
  OAI21_X1 U12795 ( .B1(n15611), .B2(n10205), .A(n11093), .ZN(n15318) );
  NAND2_X1 U12796 ( .A1(n15402), .A2(n11008), .ZN(n15394) );
  NAND2_X1 U12797 ( .A1(n15383), .A2(n10211), .ZN(n15365) );
  NAND2_X1 U12798 ( .A1(n11652), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11653) );
  INV_X1 U12799 ( .A(n13256), .ZN(n13254) );
  INV_X1 U12800 ( .A(n13246), .ZN(n13255) );
  NAND2_X1 U12801 ( .A1(n13921), .A2(n13979), .ZN(n13978) );
  INV_X1 U12803 ( .A(n15146), .ZN(n15138) );
  NAND2_X1 U12804 ( .A1(n12840), .A2(n11886), .ZN(n11856) );
  XNOR2_X1 U12805 ( .A(n11882), .B(n11828), .ZN(n12840) );
  NAND2_X1 U12806 ( .A1(n15258), .A2(n19391), .ZN(n11613) );
  AND4_X1 U12807 ( .A1(n10815), .A2(n10813), .A3(n10814), .A4(n10812), .ZN(
        n10816) );
  XNOR2_X1 U12808 ( .A(n12088), .B(n12087), .ZN(n14386) );
  AOI21_X1 U12809 ( .B1(n14384), .B2(n16069), .A(n14383), .ZN(n14385) );
  NAND2_X1 U12810 ( .A1(n14384), .A2(n14352), .ZN(n14356) );
  NAND2_X1 U12811 ( .A1(n9740), .A2(n10714), .ZN(n10715) );
  AND2_X1 U12812 ( .A1(n13580), .A2(n10746), .ZN(n19742) );
  INV_X1 U12813 ( .A(n17506), .ZN(n17432) );
  INV_X1 U12814 ( .A(n12918), .ZN(n14303) );
  INV_X1 U12815 ( .A(n14303), .ZN(n14188) );
  NAND2_X1 U12816 ( .A1(n11032), .A2(n15638), .ZN(n10215) );
  NOR2_X1 U12817 ( .A1(n20545), .A2(n20514), .ZN(n10216) );
  AND2_X1 U12818 ( .A1(n10287), .A2(n10219), .ZN(n10217) );
  INV_X1 U12819 ( .A(n15305), .ZN(n11121) );
  INV_X1 U12820 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10354) );
  INV_X1 U12821 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10344) );
  OR2_X1 U12822 ( .A1(n17263), .A2(n17299), .ZN(n10219) );
  NOR2_X1 U12823 ( .A1(n15034), .A2(n15526), .ZN(n10220) );
  AND2_X1 U12824 ( .A1(n10776), .A2(n10668), .ZN(n10221) );
  INV_X1 U12825 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19309) );
  AND2_X1 U12826 ( .A1(n10769), .A2(n15080), .ZN(n10222) );
  INV_X1 U12827 ( .A(n17897), .ZN(n17871) );
  AND2_X1 U12828 ( .A1(n10633), .A2(n13590), .ZN(n10223) );
  NAND2_X1 U12829 ( .A1(n11361), .A2(n11360), .ZN(n10224) );
  AND2_X1 U12830 ( .A1(n17871), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10225) );
  INV_X1 U12831 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12087) );
  INV_X1 U12832 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14548) );
  INV_X1 U12833 ( .A(n11380), .ZN(n11534) );
  OR2_X1 U12834 ( .A1(n11430), .A2(n11429), .ZN(n10226) );
  INV_X1 U12835 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n12754) );
  INV_X1 U12836 ( .A(n11397), .ZN(n11535) );
  INV_X1 U12837 ( .A(n17691), .ZN(n17900) );
  NAND2_X1 U12838 ( .A1(n17488), .A2(n17994), .ZN(n17691) );
  INV_X1 U12839 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10880) );
  AND2_X1 U12840 ( .A1(n12520), .A2(n12539), .ZN(n10227) );
  INV_X1 U12841 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12315) );
  NOR2_X1 U12842 ( .A1(n17995), .A2(n17941), .ZN(n17738) );
  INV_X1 U12843 ( .A(n17738), .ZN(n17770) );
  INV_X1 U12844 ( .A(n15284), .ZN(n15309) );
  AND2_X1 U12845 ( .A1(n15327), .A2(n15609), .ZN(n10228) );
  INV_X1 U12846 ( .A(n11600), .ZN(n19210) );
  NAND2_X1 U12847 ( .A1(n11282), .A2(n11281), .ZN(n10229) );
  INV_X1 U12848 ( .A(n10728), .ZN(n10729) );
  INV_X1 U12849 ( .A(n10714), .ZN(n10740) );
  OR4_X1 U12850 ( .A1(n15418), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14370), .A4(n15271), .ZN(n10230) );
  AND2_X1 U12851 ( .A1(n11578), .A2(n11363), .ZN(n16475) );
  AND4_X1 U12852 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n10231) );
  INV_X1 U12853 ( .A(n14451), .ZN(n14466) );
  NAND2_X2 U12854 ( .A1(n9732), .A2(n12797), .ZN(n11818) );
  AND2_X1 U12855 ( .A1(n9766), .A2(n13073), .ZN(n10232) );
  AND4_X1 U12856 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n10233) );
  NAND2_X1 U12857 ( .A1(n20204), .A2(n14351), .ZN(n20194) );
  NAND3_X1 U12858 ( .A1(n11800), .A2(n13671), .A3(n12837), .ZN(n12112) );
  AOI22_X1 U12859 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19441), .B1(
        n10942), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10813) );
  OR2_X1 U12860 ( .A1(n11966), .A2(n11965), .ZN(n12035) );
  AOI22_X1 U12861 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U12862 ( .A1(n11804), .A2(n12836), .ZN(n11816) );
  NAND2_X1 U12863 ( .A1(n11802), .A2(n12863), .ZN(n11715) );
  INV_X1 U12864 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11666) );
  OR2_X1 U12865 ( .A1(n11978), .A2(n11977), .ZN(n12047) );
  AOI22_X1 U12866 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10628) );
  INV_X1 U12867 ( .A(n15528), .ZN(n11250) );
  AND4_X1 U12868 ( .A1(n10875), .A2(n10874), .A3(n10873), .A4(n10872), .ZN(
        n10877) );
  AND2_X1 U12869 ( .A1(n10735), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10673) );
  NOR2_X1 U12870 ( .A1(n10256), .A2(n18327), .ZN(n10273) );
  OR2_X1 U12871 ( .A1(n14610), .A2(n14019), .ZN(n14020) );
  INV_X1 U12873 ( .A(n14167), .ZN(n13432) );
  INV_X1 U12874 ( .A(n14588), .ZN(n14088) );
  INV_X1 U12875 ( .A(n11800), .ZN(n12160) );
  OR2_X1 U12876 ( .A1(n11954), .A2(n11953), .ZN(n12023) );
  OR2_X1 U12877 ( .A1(n11915), .A2(n11914), .ZN(n11916) );
  AND2_X1 U12878 ( .A1(n21022), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11151) );
  AND2_X1 U12879 ( .A1(n12523), .A2(n10227), .ZN(n12524) );
  NOR2_X1 U12880 ( .A1(n15720), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12424) );
  AND3_X1 U12881 ( .A1(n10612), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10611), .ZN(n10615) );
  NAND2_X1 U12882 ( .A1(n10597), .A2(n13590), .ZN(n10604) );
  OR2_X1 U12883 ( .A1(n10474), .A2(n10475), .ZN(n10467) );
  NAND2_X1 U12884 ( .A1(n18319), .A2(n17456), .ZN(n10463) );
  AND2_X1 U12885 ( .A1(n13435), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14299) );
  NOR2_X1 U12886 ( .A1(n14187), .A2(n13433), .ZN(n14209) );
  INV_X1 U12887 ( .A(n11916), .ZN(n12005) );
  NOR2_X1 U12888 ( .A1(n13474), .A2(n13473), .ZN(n12351) );
  OAI211_X1 U12889 ( .C1(n12542), .C2(n12541), .A(n12577), .B(n12540), .ZN(
        n12543) );
  NAND2_X1 U12890 ( .A1(n12502), .A2(n12497), .ZN(n12503) );
  NAND2_X1 U12891 ( .A1(n10578), .A2(n10577), .ZN(n10583) );
  OR2_X1 U12892 ( .A1(n10919), .A2(n10918), .ZN(n11403) );
  INV_X1 U12893 ( .A(n15446), .ZN(n11251) );
  INV_X1 U12894 ( .A(n10677), .ZN(n10672) );
  OAI21_X1 U12895 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18944), .A(
        n10467), .ZN(n10468) );
  NAND2_X1 U12896 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20969), .ZN(
        n10234) );
  AND2_X1 U12897 ( .A1(n18143), .A2(n10354), .ZN(n10355) );
  INV_X1 U12898 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10348) );
  OR2_X1 U12899 ( .A1(n15939), .A2(n18361), .ZN(n10530) );
  OAI21_X1 U12900 ( .B1(n12869), .B2(n9907), .A(n12868), .ZN(n13070) );
  OR2_X1 U12901 ( .A1(n9751), .A2(n11749), .ZN(n11750) );
  XNOR2_X1 U12902 ( .A(n13436), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14379) );
  NAND2_X1 U12903 ( .A1(n14209), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14232) );
  OR2_X1 U12904 ( .A1(n11940), .A2(n11939), .ZN(n12015) );
  INV_X1 U12905 ( .A(n12115), .ZN(n12163) );
  INV_X1 U12906 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11892) );
  INV_X1 U12907 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20272) );
  INV_X1 U12908 ( .A(n12318), .ZN(n13580) );
  OR2_X1 U12909 ( .A1(n10971), .A2(n10970), .ZN(n11407) );
  NAND2_X1 U12910 ( .A1(n10687), .A2(n20077), .ZN(n12637) );
  NOR2_X1 U12911 ( .A1(n15543), .A2(n11606), .ZN(n15515) );
  AND2_X1 U12912 ( .A1(n11080), .A2(n11079), .ZN(n19047) );
  INV_X1 U12913 ( .A(n11390), .ZN(n11214) );
  OAI21_X1 U12914 ( .B1(n18335), .B2(n10536), .A(n10535), .ZN(n10538) );
  NOR2_X1 U12915 ( .A1(n18361), .A2(n18335), .ZN(n10531) );
  INV_X1 U12916 ( .A(n10362), .ZN(n10363) );
  NOR2_X1 U12917 ( .A1(n17914), .A2(n17913), .ZN(n10516) );
  NOR2_X1 U12918 ( .A1(n17916), .A2(n17915), .ZN(n17914) );
  OAI21_X1 U12919 ( .B1(n15741), .B2(n10530), .A(n18766), .ZN(n18794) );
  AND2_X1 U12920 ( .A1(n12294), .A2(n12293), .ZN(n14403) );
  NAND2_X1 U12921 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13248) );
  OR3_X1 U12922 ( .A1(n20745), .A2(n13430), .A3(n13429), .ZN(n15994) );
  OAI21_X1 U12923 ( .B1(n20268), .B2(n13971), .A(n13087), .ZN(n13089) );
  INV_X1 U12924 ( .A(n14332), .ZN(n14333) );
  NAND2_X1 U12925 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n13431), .ZN(
        n14167) );
  NOR2_X1 U12926 ( .A1(n14040), .A2(n14525), .ZN(n14055) );
  AND3_X1 U12927 ( .A1(n14018), .A2(n14017), .A3(n14016), .ZN(n14610) );
  INV_X1 U12928 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16028) );
  INV_X1 U12929 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20122) );
  AND3_X1 U12930 ( .A1(n12881), .A2(n12880), .A3(n15907), .ZN(n15895) );
  AND2_X1 U12931 ( .A1(n16077), .A2(n12077), .ZN(n16063) );
  AND2_X1 U12932 ( .A1(n13892), .A2(n12074), .ZN(n16077) );
  NAND2_X1 U12933 ( .A1(n12299), .A2(n14403), .ZN(n14920) );
  AND2_X1 U12934 ( .A1(n12297), .A2(n14920), .ZN(n12856) );
  NOR2_X1 U12935 ( .A1(n20554), .A2(n14408), .ZN(n14957) );
  OR2_X1 U12936 ( .A1(n20423), .A2(n20477), .ZN(n13683) );
  NOR2_X1 U12937 ( .A1(n13287), .A2(n13676), .ZN(n20553) );
  OR3_X1 U12938 ( .A1(n20554), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13135), 
        .ZN(n13680) );
  NAND2_X1 U12939 ( .A1(n19241), .A2(n19224), .ZN(n16280) );
  INV_X1 U12940 ( .A(n19222), .ZN(n19197) );
  AND2_X1 U12941 ( .A1(n11333), .A2(n11332), .ZN(n15123) );
  NAND2_X1 U12942 ( .A1(n12340), .A2(n12341), .ZN(n12822) );
  INV_X1 U12943 ( .A(n12501), .ZN(n12497) );
  INV_X1 U12944 ( .A(n19246), .ZN(n15250) );
  AND2_X1 U12945 ( .A1(n11317), .A2(n11316), .ZN(n15158) );
  OR2_X1 U12946 ( .A1(n15441), .A2(n11608), .ZN(n15418) );
  NAND2_X1 U12947 ( .A1(n20043), .A2(n20050), .ZN(n19673) );
  INV_X1 U12948 ( .A(n9715), .ZN(n19889) );
  NOR2_X2 U12949 ( .A1(n18988), .A2(n15739), .ZN(n18780) );
  NOR2_X1 U12950 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16868), .ZN(n16855) );
  NOR2_X1 U12951 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16893), .ZN(n16874) );
  INV_X1 U12952 ( .A(n17042), .ZN(n16913) );
  NAND2_X1 U12953 ( .A1(n18989), .A2(n17523), .ZN(n16671) );
  NOR2_X1 U12954 ( .A1(n17684), .A2(n18057), .ZN(n17690) );
  NAND2_X1 U12955 ( .A1(n18160), .A2(n18131), .ZN(n17805) );
  NAND2_X1 U12956 ( .A1(n18213), .A2(n17897), .ZN(n17896) );
  NOR2_X1 U12957 ( .A1(n17693), .A2(n18039), .ZN(n17678) );
  NAND2_X1 U12958 ( .A1(n10356), .A2(n17897), .ZN(n17783) );
  INV_X1 U12959 ( .A(n17805), .ZN(n18134) );
  NAND2_X1 U12960 ( .A1(n10357), .A2(n18221), .ZN(n17870) );
  INV_X1 U12961 ( .A(n18145), .ZN(n18218) );
  INV_X1 U12962 ( .A(n18298), .ZN(n18289) );
  INV_X1 U12963 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18809) );
  INV_X1 U12964 ( .A(n10485), .ZN(n18330) );
  INV_X1 U12965 ( .A(n20601), .ZN(n20548) );
  INV_X1 U12966 ( .A(n20136), .ZN(n20170) );
  AND2_X1 U12967 ( .A1(n13464), .A2(n13463), .ZN(n20159) );
  AND2_X1 U12968 ( .A1(n15994), .A2(n13437), .ZN(n20154) );
  NAND2_X1 U12969 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13083), .ZN(
        n13249) );
  INV_X1 U12970 ( .A(n20194), .ZN(n20199) );
  AND2_X1 U12971 ( .A1(n14354), .A2(n14353), .ZN(n14713) );
  INV_X1 U12972 ( .A(n14642), .ZN(n14353) );
  AND2_X1 U12973 ( .A1(n14609), .A2(n13973), .ZN(n16021) );
  INV_X1 U12974 ( .A(n16120), .ZN(n16104) );
  AND2_X1 U12975 ( .A1(n16120), .A2(n12910), .ZN(n16114) );
  AOI21_X1 U12976 ( .B1(n14900), .B2(n12307), .A(n14899), .ZN(n16189) );
  AND2_X1 U12977 ( .A1(n12882), .A2(n12842), .ZN(n20177) );
  NOR2_X1 U12978 ( .A1(n16189), .A2(n16195), .ZN(n16140) );
  INV_X1 U12979 ( .A(n14920), .ZN(n14885) );
  OAI21_X1 U12980 ( .B1(n13171), .B2(n14920), .A(n14926), .ZN(n16250) );
  INV_X1 U12981 ( .A(n16220), .ZN(n16256) );
  INV_X1 U12982 ( .A(n13393), .ZN(n13676) );
  NOR2_X1 U12983 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14949) );
  INV_X1 U12984 ( .A(n20659), .ZN(n20295) );
  INV_X1 U12985 ( .A(n20326), .ZN(n20316) );
  INV_X1 U12986 ( .A(n20358), .ZN(n20350) );
  INV_X1 U12987 ( .A(n20418), .ZN(n20410) );
  NAND2_X1 U12988 ( .A1(n20268), .A2(n20267), .ZN(n20360) );
  OR2_X1 U12989 ( .A1(n13130), .A2(n13395), .ZN(n20394) );
  INV_X1 U12990 ( .A(n13683), .ZN(n13758) );
  INV_X1 U12991 ( .A(n20509), .ZN(n20501) );
  INV_X1 U12992 ( .A(n20530), .ZN(n20541) );
  NOR2_X1 U12993 ( .A1(n20268), .A2(n9769), .ZN(n20512) );
  INV_X1 U12994 ( .A(n20547), .ZN(n20588) );
  NAND2_X1 U12995 ( .A1(n16280), .A2(n16279), .ZN(n16281) );
  INV_X1 U12996 ( .A(n19200), .ZN(n16282) );
  INV_X1 U12997 ( .A(n19228), .ZN(n19194) );
  AND2_X1 U12998 ( .A1(n13333), .A2(n13332), .ZN(n19222) );
  INV_X1 U12999 ( .A(n19174), .ZN(n19236) );
  OR2_X1 U13000 ( .A1(n11443), .A2(n11442), .ZN(n13117) );
  NOR2_X1 U13001 ( .A1(n15164), .A2(n15163), .ZN(n15166) );
  AND2_X1 U13002 ( .A1(n19275), .A2(n12779), .ZN(n19246) );
  INV_X1 U13003 ( .A(n19275), .ZN(n19294) );
  AND2_X1 U13004 ( .A1(n12649), .A2(n13610), .ZN(n19380) );
  AND2_X1 U13005 ( .A1(n16445), .A2(n12731), .ZN(n16434) );
  INV_X1 U13006 ( .A(n16445), .ZN(n16409) );
  NOR2_X1 U13007 ( .A1(n11604), .A2(n11603), .ZN(n16469) );
  OAI21_X1 U13008 ( .B1(n13666), .B2(n13665), .A(n13664), .ZN(n19436) );
  INV_X1 U13009 ( .A(n19524), .ZN(n19526) );
  INV_X1 U13010 ( .A(n19578), .ZN(n19564) );
  INV_X1 U13011 ( .A(n19567), .ZN(n19603) );
  NOR2_X1 U13012 ( .A1(n19893), .A2(n19579), .ZN(n19630) );
  NAND2_X1 U13013 ( .A1(n19672), .A2(n19638), .ZN(n19617) );
  INV_X1 U13014 ( .A(n19697), .ZN(n19699) );
  INV_X1 U13015 ( .A(n19673), .ZN(n19670) );
  NOR2_X1 U13016 ( .A1(n19737), .A2(n20030), .ZN(n19805) );
  INV_X1 U13017 ( .A(n19835), .ZN(n19841) );
  NOR2_X1 U13018 ( .A1(n19769), .A2(n19817), .ZN(n19836) );
  INV_X1 U13019 ( .A(n19749), .ZN(n19896) );
  NOR2_X1 U13020 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n13648), .ZN(n19304) );
  INV_X1 U13021 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n21085) );
  OR2_X1 U13022 ( .A1(n16726), .A2(P3_EBX_REG_28__SCAN_IN), .ZN(n16717) );
  INV_X2 U13023 ( .A(n18324), .ZN(n18970) );
  NAND2_X1 U13024 ( .A1(n17041), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17031) );
  NOR2_X1 U13025 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16823), .ZN(n16811) );
  NOR2_X1 U13026 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16939), .ZN(n16928) );
  INV_X1 U13027 ( .A(n17031), .ZN(n16997) );
  INV_X1 U13028 ( .A(n17030), .ZN(n17041) );
  OR2_X1 U13029 ( .A1(n17343), .A2(n17346), .ZN(n17339) );
  NOR3_X1 U13030 ( .A1(n17456), .A2(n17450), .A3(n17583), .ZN(n17442) );
  INV_X1 U13031 ( .A(n17508), .ZN(n17513) );
  INV_X1 U13032 ( .A(n18319), .ZN(n17523) );
  NOR2_X1 U13033 ( .A1(n16497), .A2(n17691), .ZN(n16498) );
  INV_X1 U13034 ( .A(n17795), .ZN(n17779) );
  INV_X1 U13035 ( .A(n17488), .ZN(n16536) );
  NAND2_X1 U13036 ( .A1(n18131), .A2(n17820), .ZN(n17819) );
  NOR2_X2 U13037 ( .A1(n18289), .A2(n18137), .ZN(n18203) );
  INV_X1 U13038 ( .A(n18036), .ZN(n18212) );
  AOI21_X2 U13039 ( .B1(n15852), .B2(n10489), .A(n18832), .ZN(n18298) );
  NOR2_X1 U13040 ( .A1(n18773), .A2(n18289), .ZN(n18297) );
  NAND2_X1 U13041 ( .A1(n18974), .A2(n18317), .ZN(n18367) );
  INV_X1 U13042 ( .A(n18829), .ZN(n18952) );
  INV_X1 U13043 ( .A(n18704), .ZN(n18358) );
  CLKBUF_X1 U13044 ( .A(n18427), .Z(n18423) );
  INV_X1 U13045 ( .A(n18407), .ZN(n18470) );
  INV_X1 U13046 ( .A(n18588), .ZN(n18666) );
  NAND3_X1 U13047 ( .A1(n12860), .A2(n14413), .A3(n15907), .ZN(n14399) );
  INV_X1 U13048 ( .A(n20738), .ZN(n20751) );
  INV_X1 U13049 ( .A(n20178), .ZN(n20162) );
  INV_X1 U13050 ( .A(n20154), .ZN(n20141) );
  INV_X1 U13051 ( .A(n20126), .ZN(n20186) );
  NAND2_X1 U13052 ( .A1(n14354), .A2(n14642), .ZN(n14717) );
  OAI21_X1 U13053 ( .B1(n14506), .B2(n14505), .A(n9779), .ZN(n14791) );
  INV_X1 U13054 ( .A(n14724), .ZN(n16046) );
  INV_X1 U13055 ( .A(n20205), .ZN(n20229) );
  NOR2_X1 U13056 ( .A1(n14399), .A2(n12940), .ZN(n12975) );
  INV_X1 U13057 ( .A(n15949), .ZN(n14805) );
  INV_X1 U13058 ( .A(n16069), .ZN(n14832) );
  INV_X1 U13059 ( .A(n16116), .ZN(n20100) );
  NAND2_X1 U13060 ( .A1(n12299), .A2(n12178), .ZN(n16220) );
  INV_X1 U13061 ( .A(n16244), .ZN(n16259) );
  INV_X1 U13062 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20449) );
  OR2_X1 U13063 ( .A1(n20360), .A2(n20394), .ZN(n20326) );
  OR2_X1 U13064 ( .A1(n20360), .A2(n20447), .ZN(n20358) );
  OR2_X1 U13065 ( .A1(n20360), .A2(n20477), .ZN(n20390) );
  OR2_X1 U13066 ( .A1(n20360), .A2(n20510), .ZN(n20418) );
  OR2_X1 U13067 ( .A1(n20423), .A2(n20394), .ZN(n20446) );
  INV_X1 U13068 ( .A(n13398), .ZN(n13729) );
  NAND2_X1 U13069 ( .A1(n20512), .A2(n20448), .ZN(n20509) );
  NAND2_X1 U13070 ( .A1(n20512), .A2(n20511), .ZN(n20593) );
  INV_X1 U13071 ( .A(n13129), .ZN(n13724) );
  INV_X1 U13072 ( .A(n13289), .ZN(n13717) );
  OR2_X1 U13073 ( .A1(n20606), .A2(n20510), .ZN(n20659) );
  INV_X1 U13074 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20661) );
  INV_X1 U13075 ( .A(n20736), .ZN(n20738) );
  AND2_X1 U13076 ( .A1(n11366), .A2(n12642), .ZN(n20074) );
  OR2_X1 U13077 ( .A1(n13327), .A2(n13329), .ZN(n19200) );
  OR2_X1 U13078 ( .A1(n20074), .A2(n13335), .ZN(n19178) );
  INV_X1 U13079 ( .A(n12605), .ZN(n12606) );
  NAND2_X1 U13080 ( .A1(n12830), .A2(n12829), .ZN(n19672) );
  AND2_X1 U13081 ( .A1(n12778), .A2(n19304), .ZN(n19275) );
  NOR2_X1 U13082 ( .A1(n19295), .A2(n19280), .ZN(n19286) );
  INV_X1 U13083 ( .A(n19278), .ZN(n19303) );
  OR2_X1 U13084 ( .A1(n19376), .A2(n19312), .ZN(n19344) );
  NAND2_X1 U13085 ( .A1(n19308), .A2(n20082), .ZN(n19376) );
  INV_X1 U13086 ( .A(n19380), .ZN(n19306) );
  INV_X1 U13087 ( .A(n11663), .ZN(n11664) );
  INV_X1 U13088 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19102) );
  INV_X1 U13089 ( .A(n16434), .ZN(n16424) );
  INV_X1 U13090 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16446) );
  INV_X1 U13091 ( .A(n19391), .ZN(n15702) );
  INV_X1 U13092 ( .A(n16475), .ZN(n19404) );
  INV_X1 U13093 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15937) );
  AOI211_X2 U13094 ( .C1(n13657), .C2(n13665), .A(n9715), .B(n13656), .ZN(
        n19439) );
  INV_X1 U13095 ( .A(n19497), .ZN(n19492) );
  OR2_X1 U13096 ( .A1(n19579), .A2(n20030), .ZN(n19524) );
  OR2_X1 U13097 ( .A1(n19617), .A2(n20030), .ZN(n19541) );
  OR2_X1 U13098 ( .A1(n19617), .A2(n19817), .ZN(n19567) );
  OR2_X1 U13099 ( .A1(n19579), .A2(n19817), .ZN(n19578) );
  INV_X1 U13100 ( .A(n19630), .ZN(n19637) );
  OR2_X1 U13101 ( .A1(n19617), .A2(n19893), .ZN(n19661) );
  NAND2_X1 U13102 ( .A1(n19847), .A2(n19670), .ZN(n19697) );
  NAND2_X1 U13103 ( .A1(n19819), .A2(n19670), .ZN(n19736) );
  NAND2_X1 U13104 ( .A1(n19847), .A2(n19704), .ZN(n19760) );
  INV_X1 U13105 ( .A(n19805), .ZN(n19801) );
  AND2_X1 U13106 ( .A1(n19813), .A2(n19812), .ZN(n19835) );
  NAND2_X1 U13107 ( .A1(n19819), .A2(n19818), .ZN(n19873) );
  INV_X1 U13108 ( .A(n19820), .ZN(n19899) );
  INV_X1 U13109 ( .A(n19867), .ZN(n19923) );
  INV_X1 U13110 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18974) );
  NAND4_X1 U13111 ( .A1(n16670), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n18970), 
        .A4(n16669), .ZN(n16999) );
  INV_X2 U13112 ( .A(n18361), .ZN(n17456) );
  AND2_X1 U13113 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17102), .ZN(n17096) );
  NOR2_X1 U13114 ( .A1(n17154), .A2(n17181), .ZN(n17169) );
  NOR2_X1 U13115 ( .A1(n17456), .A2(n17484), .ZN(n17490) );
  NAND2_X1 U13116 ( .A1(n18804), .A2(n17369), .ZN(n17508) );
  NAND2_X1 U13117 ( .A1(n17524), .A2(n17523), .ZN(n17548) );
  NAND2_X1 U13118 ( .A1(n17579), .A2(n17522), .ZN(n17577) );
  INV_X1 U13119 ( .A(n17627), .ZN(n17622) );
  AOI21_X1 U13120 ( .B1(n16499), .B2(n17888), .A(n16498), .ZN(n16500) );
  NAND2_X1 U13121 ( .A1(n17841), .A2(n16538), .ZN(n17795) );
  INV_X1 U13122 ( .A(n17988), .ZN(n17975) );
  NOR2_X1 U13123 ( .A1(n17968), .A2(n17941), .ZN(n17991) );
  INV_X1 U13124 ( .A(n18291), .ZN(n18285) );
  INV_X1 U13125 ( .A(n18287), .ZN(n18305) );
  INV_X1 U13126 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18814) );
  AOI211_X1 U13127 ( .C1(n18977), .C2(n18802), .A(n18318), .B(n15853), .ZN(
        n18957) );
  INV_X1 U13128 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18338) );
  INV_X1 U13129 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18365) );
  INV_X1 U13130 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18593) );
  INV_X1 U13131 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18650) );
  INV_X1 U13132 ( .A(n18709), .ZN(n18679) );
  INV_X1 U13133 ( .A(n18722), .ZN(n18684) );
  INV_X1 U13134 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18713) );
  INV_X1 U13135 ( .A(n18581), .ZN(n18746) );
  INV_X1 U13136 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21062) );
  INV_X1 U13137 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18852) );
  CLKBUF_X1 U13138 ( .A(n16641), .Z(n16642) );
  NAND2_X1 U13139 ( .A1(n10554), .A2(n10553), .ZN(P3_U2831) );
  INV_X1 U13140 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16528) );
  OR2_X2 U13141 ( .A1(n18795), .A2(n10238), .ZN(n10256) );
  AOI22_X1 U13142 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10252) );
  NAND4_X1 U13143 ( .A1(n18944), .A2(n18951), .A3(n18933), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17187) );
  INV_X1 U13144 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20886) );
  AOI22_X1 U13145 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10237) );
  INV_X2 U13146 ( .A(n10235), .ZN(n17204) );
  AOI22_X1 U13147 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10236) );
  OAI211_X1 U13148 ( .C1(n10404), .C2(n20886), .A(n10237), .B(n10236), .ZN(
        n10250) );
  NOR2_X2 U13149 ( .A1(n17027), .A2(n10238), .ZN(n10329) );
  NOR2_X4 U13150 ( .A1(n18795), .A2(n10239), .ZN(n17290) );
  AOI22_X1 U13151 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10248) );
  NAND2_X1 U13152 ( .A1(n18944), .A2(n18933), .ZN(n10241) );
  AOI22_X1 U13153 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10247) );
  NOR2_X4 U13154 ( .A1(n18933), .A2(n10243), .ZN(n17313) );
  AOI22_X1 U13155 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10246) );
  NAND2_X1 U13157 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10245) );
  NAND4_X1 U13158 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10249) );
  AOI211_X1 U13159 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n10250), .B(n10249), .ZN(n10251) );
  OAI211_X1 U13160 ( .C1(n10256), .C2(n18355), .A(n10252), .B(n10251), .ZN(
        n10496) );
  INV_X1 U13161 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U13162 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10264) );
  INV_X1 U13163 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18739) );
  AOI22_X1 U13164 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13165 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17327), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10254) );
  OAI211_X1 U13166 ( .C1(n10404), .C2(n18739), .A(n10255), .B(n10254), .ZN(
        n10262) );
  AOI22_X1 U13167 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13168 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U13169 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U13170 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10257) );
  NAND4_X1 U13171 ( .A1(n10260), .A2(n10259), .A3(n10258), .A4(n10257), .ZN(
        n10261) );
  AOI211_X1 U13172 ( .C1(n10286), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n10262), .B(n10261), .ZN(n10263) );
  OAI211_X1 U13173 ( .C1(n10253), .C2(n17141), .A(n10264), .B(n10263), .ZN(
        n10502) );
  INV_X1 U13174 ( .A(n10502), .ZN(n17499) );
  AOI22_X1 U13175 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10265), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10266) );
  OAI21_X1 U13176 ( .B1(n17263), .B2(n21085), .A(n10266), .ZN(n10270) );
  INV_X1 U13177 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18573) );
  AOI22_X1 U13178 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10330), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U13179 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10267) );
  OAI211_X1 U13180 ( .C1(n17275), .C2(n18573), .A(n10268), .B(n10267), .ZN(
        n10269) );
  AOI211_X1 U13181 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n10270), .B(n10269), .ZN(n10279) );
  INV_X2 U13182 ( .A(n17204), .ZN(n17270) );
  AOI22_X1 U13183 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10271) );
  OAI21_X1 U13184 ( .B1(n15789), .B2(n18650), .A(n10271), .ZN(n10272) );
  INV_X1 U13185 ( .A(n10272), .ZN(n10276) );
  AOI22_X1 U13186 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10275) );
  AND2_X2 U13189 ( .A1(n10279), .A2(n21088), .ZN(n10494) );
  INV_X1 U13190 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18726) );
  AOI22_X1 U13191 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10330), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13192 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10329), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10280) );
  OAI211_X1 U13193 ( .C1(n10404), .C2(n18726), .A(n10281), .B(n10280), .ZN(
        n10285) );
  AOI22_X1 U13194 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13195 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10265), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U13196 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10282) );
  AOI22_X1 U13197 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10287) );
  INV_X1 U13198 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17299) );
  INV_X1 U13199 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U13200 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10296) );
  INV_X1 U13201 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18578) );
  INV_X1 U13202 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17157) );
  OAI22_X1 U13203 ( .A1(n17275), .A2(n18578), .B1(n17334), .B2(n17157), .ZN(
        n10294) );
  AOI22_X1 U13204 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13205 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13206 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10290) );
  NAND3_X1 U13207 ( .A1(n10292), .A2(n10291), .A3(n10290), .ZN(n10293) );
  AOI211_X1 U13208 ( .C1(n9734), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n10294), .B(n10293), .ZN(n10295) );
  OAI211_X1 U13209 ( .C1(n9814), .C2(n17165), .A(n10296), .B(n10295), .ZN(
        n10297) );
  INV_X1 U13210 ( .A(n10297), .ZN(n10302) );
  AOI22_X1 U13211 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10298) );
  OAI21_X1 U13212 ( .B1(n10256), .B2(n18338), .A(n10298), .ZN(n10300) );
  AOI22_X1 U13213 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10303) );
  INV_X1 U13214 ( .A(n10303), .ZN(n10313) );
  INV_X1 U13215 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18584) );
  AOI22_X1 U13216 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13217 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10304) );
  OAI21_X1 U13218 ( .B1(n17325), .B2(n20824), .A(n10304), .ZN(n10309) );
  AOI22_X1 U13219 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13220 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13221 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10305) );
  NAND3_X1 U13222 ( .A1(n10307), .A2(n10306), .A3(n10305), .ZN(n10308) );
  AOI211_X1 U13223 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n10309), .B(n10308), .ZN(n10310) );
  OAI211_X1 U13224 ( .C1(n17275), .C2(n18584), .A(n10311), .B(n10310), .ZN(
        n10312) );
  INV_X1 U13225 ( .A(n17495), .ZN(n10346) );
  INV_X1 U13226 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18670) );
  AOI22_X1 U13227 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10314) );
  OAI21_X1 U13228 ( .B1(n15789), .B2(n18670), .A(n10314), .ZN(n10323) );
  INV_X1 U13229 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21050) );
  AOI22_X1 U13230 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10321) );
  INV_X1 U13231 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17225) );
  OAI22_X1 U13232 ( .A1(n17275), .A2(n18593), .B1(n17334), .B2(n17225), .ZN(
        n10319) );
  AOI22_X1 U13233 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13234 ( .A1(n17290), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13235 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10315) );
  NAND3_X1 U13236 ( .A1(n10317), .A2(n10316), .A3(n10315), .ZN(n10318) );
  AOI211_X1 U13237 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n10319), .B(n10318), .ZN(n10320) );
  OAI211_X1 U13238 ( .C1(n21050), .C2(n17263), .A(n10321), .B(n10320), .ZN(
        n10322) );
  INV_X1 U13239 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17913) );
  XOR2_X1 U13240 ( .A(n10324), .B(n17499), .Z(n10325) );
  INV_X1 U13241 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18250) );
  XOR2_X1 U13242 ( .A(n18250), .B(n10325), .Z(n17955) );
  INV_X1 U13243 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20943) );
  NOR2_X1 U13244 ( .A1(n20943), .A2(n10341), .ZN(n10342) );
  INV_X1 U13245 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15787) );
  AOI22_X1 U13246 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10326) );
  OAI21_X1 U13247 ( .B1(n9771), .B2(n15787), .A(n10326), .ZN(n10339) );
  INV_X1 U13248 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U13249 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10338) );
  INV_X1 U13250 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18322) );
  AOI22_X1 U13251 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10328) );
  OAI21_X1 U13252 ( .B1(n10256), .B2(n18322), .A(n10328), .ZN(n10337) );
  AOI22_X1 U13253 ( .A1(n10329), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13254 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10330), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10334) );
  INV_X1 U13255 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18570) );
  NAND3_X1 U13256 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n10336) );
  NAND2_X1 U13257 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17993), .ZN(
        n17992) );
  INV_X1 U13258 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18938) );
  NOR2_X1 U13259 ( .A1(n17512), .A2(n18938), .ZN(n10340) );
  XOR2_X1 U13260 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10341), .Z(
        n17977) );
  NOR2_X1 U13261 ( .A1(n10342), .A2(n17976), .ZN(n17961) );
  XNOR2_X1 U13262 ( .A(n10343), .B(n10492), .ZN(n17962) );
  NAND2_X1 U13263 ( .A1(n17961), .A2(n17962), .ZN(n17960) );
  OAI21_X1 U13264 ( .B1(n17961), .B2(n17962), .A(n10344), .ZN(n10345) );
  NAND2_X1 U13265 ( .A1(n17960), .A2(n10345), .ZN(n17954) );
  XNOR2_X1 U13266 ( .A(n10347), .B(n10346), .ZN(n17937) );
  INV_X1 U13267 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18220) );
  XOR2_X1 U13268 ( .A(n10349), .B(n17492), .Z(n10350) );
  XOR2_X1 U13269 ( .A(n18220), .B(n10350), .Z(n17924) );
  INV_X1 U13270 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18221) );
  NOR3_X1 U13271 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17817) );
  INV_X1 U13272 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18143) );
  NAND3_X1 U13273 ( .A1(n17814), .A2(n17817), .A3(n10355), .ZN(n10356) );
  INV_X1 U13274 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18178) );
  INV_X1 U13275 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21002) );
  INV_X1 U13276 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18206) );
  NOR2_X1 U13277 ( .A1(n21002), .A2(n18206), .ZN(n18180) );
  NAND2_X1 U13278 ( .A1(n18180), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18172) );
  INV_X1 U13279 ( .A(n18172), .ZN(n18187) );
  NAND3_X1 U13280 ( .A1(n18187), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17796) );
  NOR2_X1 U13281 ( .A1(n18178), .A2(n17796), .ZN(n18131) );
  NAND2_X1 U13282 ( .A1(n18131), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18110) );
  INV_X1 U13283 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18125) );
  INV_X1 U13284 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18106) );
  NOR2_X1 U13285 ( .A1(n18125), .A2(n18106), .ZN(n18105) );
  INV_X1 U13286 ( .A(n18105), .ZN(n18062) );
  INV_X1 U13287 ( .A(n9820), .ZN(n10361) );
  NOR2_X1 U13288 ( .A1(n18062), .A2(n10361), .ZN(n17728) );
  INV_X1 U13289 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18058) );
  NAND2_X1 U13290 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18060) );
  INV_X1 U13291 ( .A(n18060), .ZN(n18082) );
  NAND3_X1 U13292 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18082), .ZN(n10358) );
  NOR3_X1 U13293 ( .A1(n17729), .A2(n18058), .A3(n10358), .ZN(n17697) );
  NOR2_X1 U13294 ( .A1(n18062), .A2(n10358), .ZN(n18066) );
  INV_X1 U13295 ( .A(n18066), .ZN(n18055) );
  NOR2_X1 U13296 ( .A1(n18055), .A2(n18058), .ZN(n18021) );
  NAND2_X1 U13297 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18021), .ZN(
        n17684) );
  INV_X1 U13298 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17769) );
  NAND2_X1 U13299 ( .A1(n17897), .A2(n17769), .ZN(n17764) );
  NOR2_X1 U13300 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17764), .ZN(
        n10359) );
  INV_X1 U13301 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17735) );
  NAND2_X1 U13302 ( .A1(n10359), .A2(n17735), .ZN(n17730) );
  INV_X1 U13303 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20822) );
  NAND3_X1 U13304 ( .A1(n17710), .A2(n20822), .A3(n18058), .ZN(n10360) );
  OAI21_X1 U13305 ( .B1(n10361), .B2(n17684), .A(n10360), .ZN(n10362) );
  INV_X1 U13306 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17693) );
  NAND3_X1 U13307 ( .A1(n17697), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17692), .ZN(n10366) );
  NAND2_X1 U13308 ( .A1(n10366), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10365) );
  INV_X1 U13309 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18022) );
  MUX2_X1 U13310 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17680), .S(
        n17897), .Z(n10364) );
  INV_X1 U13311 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18013) );
  NAND2_X1 U13312 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10545) );
  INV_X1 U13313 ( .A(n10545), .ZN(n18002) );
  NAND2_X1 U13314 ( .A1(n10366), .A2(n17871), .ZN(n17679) );
  INV_X1 U13315 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18009) );
  AOI221_X1 U13316 ( .B1(n15923), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), 
        .C1(n17897), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n10368), .ZN(
        n10372) );
  INV_X1 U13317 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18939) );
  AOI22_X1 U13318 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17897), .B1(
        n17871), .B2(n18939), .ZN(n10371) );
  NOR2_X1 U13319 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18939), .ZN(
        n10549) );
  AOI211_X1 U13320 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18939), .A(
        n15923), .B(n10368), .ZN(n10369) );
  OAI21_X1 U13321 ( .B1(n10549), .B2(n10369), .A(n10371), .ZN(n10370) );
  OAI21_X1 U13322 ( .B1(n10372), .B2(n10371), .A(n10370), .ZN(n16499) );
  INV_X1 U13323 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U13324 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10373) );
  OAI21_X1 U13325 ( .B1(n17325), .B2(n17274), .A(n10373), .ZN(n10382) );
  AOI22_X1 U13326 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10380) );
  INV_X1 U13327 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18656) );
  AOI22_X1 U13328 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10374) );
  OAI21_X1 U13329 ( .B1(n17334), .B2(n18656), .A(n10374), .ZN(n10378) );
  INV_X1 U13330 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U13331 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10330), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13332 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10375) );
  OAI211_X1 U13333 ( .C1(n17187), .C2(n17283), .A(n10376), .B(n10375), .ZN(
        n10377) );
  AOI211_X1 U13334 ( .C1(n10286), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n10378), .B(n10377), .ZN(n10379) );
  OAI211_X1 U13335 ( .C1(n10253), .C2(n18338), .A(n10380), .B(n10379), .ZN(
        n10381) );
  INV_X1 U13336 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18344) );
  AOI22_X1 U13337 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10383) );
  OAI21_X1 U13338 ( .B1(n10253), .B2(n18344), .A(n10383), .ZN(n10392) );
  INV_X1 U13339 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17262) );
  AOI22_X1 U13340 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10327), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10390) );
  INV_X1 U13341 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18659) );
  AOI22_X1 U13342 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10384) );
  OAI21_X1 U13343 ( .B1(n17334), .B2(n18659), .A(n10384), .ZN(n10388) );
  INV_X1 U13344 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15810) );
  AOI22_X1 U13345 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13346 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10385) );
  OAI211_X1 U13347 ( .C1(n17275), .C2(n15810), .A(n10386), .B(n10385), .ZN(
        n10387) );
  AOI211_X1 U13348 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n10388), .B(n10387), .ZN(n10389) );
  OAI211_X1 U13349 ( .C1(n9814), .C2(n17262), .A(n10390), .B(n10389), .ZN(
        n10391) );
  AOI22_X1 U13350 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10393) );
  OAI21_X1 U13351 ( .B1(n10256), .B2(n18713), .A(n10393), .ZN(n10402) );
  INV_X1 U13352 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18646) );
  AOI22_X1 U13353 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13354 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10394) );
  OAI21_X1 U13355 ( .B1(n10253), .B2(n18322), .A(n10394), .ZN(n10398) );
  AOI22_X1 U13356 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13357 ( .A1(n10330), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10395) );
  OAI211_X1 U13358 ( .C1(n17275), .C2(n15787), .A(n10396), .B(n10395), .ZN(
        n10397) );
  AOI211_X1 U13359 ( .C1(n17202), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n10398), .B(n10397), .ZN(n10399) );
  OAI211_X1 U13360 ( .C1(n17334), .C2(n18646), .A(n10400), .B(n10399), .ZN(
        n10401) );
  AOI211_X4 U13361 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n10402), .B(n10401), .ZN(n18319) );
  AOI22_X1 U13362 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17290), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17270), .ZN(n10403) );
  OAI21_X1 U13363 ( .B1(n10288), .B2(n18593), .A(n10403), .ZN(n10413) );
  AOI22_X1 U13364 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17313), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10411) );
  INV_X1 U13365 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18765) );
  OAI22_X1 U13366 ( .A1(n17225), .A2(n10404), .B1(n18765), .B2(n10256), .ZN(
        n10409) );
  AOI22_X1 U13367 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17237), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13368 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13369 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10289), .B1(
        n10286), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10405) );
  NAND3_X1 U13370 ( .A1(n10407), .A2(n10406), .A3(n10405), .ZN(n10408) );
  AOI211_X1 U13371 ( .C1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n10327), .A(
        n10409), .B(n10408), .ZN(n10410) );
  OAI211_X1 U13372 ( .C1(n10253), .C2(n18365), .A(n10411), .B(n10410), .ZN(
        n10412) );
  AOI211_X4 U13373 ( .C1(n10329), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n10413), .B(n10412), .ZN(n18361) );
  INV_X1 U13374 ( .A(n10463), .ZN(n10434) );
  INV_X1 U13375 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U13376 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10414) );
  OAI21_X1 U13377 ( .B1(n9771), .B2(n17123), .A(n10414), .ZN(n10423) );
  AOI22_X1 U13378 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13379 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10415) );
  OAI21_X1 U13380 ( .B1(n10253), .B2(n20925), .A(n10415), .ZN(n10419) );
  INV_X1 U13381 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15826) );
  AOI22_X1 U13382 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13383 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10416) );
  OAI211_X1 U13384 ( .C1(n17275), .C2(n15826), .A(n10417), .B(n10416), .ZN(
        n10418) );
  AOI211_X1 U13385 ( .C1(n17202), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n10419), .B(n10418), .ZN(n10420) );
  OAI211_X1 U13386 ( .C1(n15789), .C2(n20824), .A(n10421), .B(n10420), .ZN(
        n10422) );
  AOI22_X1 U13387 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10327), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10433) );
  INV_X1 U13388 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U13389 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13390 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10424) );
  OAI211_X1 U13391 ( .C1(n17187), .C2(n17111), .A(n10425), .B(n10424), .ZN(
        n10431) );
  AOI22_X1 U13392 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13393 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13394 ( .A1(n10330), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10427) );
  NAND2_X1 U13395 ( .A1(n17202), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10426) );
  NAND4_X1 U13396 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  AOI211_X1 U13397 ( .C1(n10286), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n10431), .B(n10430), .ZN(n10432) );
  NOR2_X1 U13398 ( .A1(n9752), .A2(n18352), .ZN(n10460) );
  NAND4_X1 U13399 ( .A1(n18335), .A2(n18341), .A3(n10434), .A4(n10460), .ZN(
        n10539) );
  AOI22_X1 U13400 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13401 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13402 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10442) );
  INV_X1 U13403 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18333) );
  INV_X1 U13404 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17171) );
  OAI22_X1 U13405 ( .A1(n10253), .A2(n18333), .B1(n17204), .B2(n17171), .ZN(
        n10440) );
  AOI22_X1 U13406 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13407 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13408 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U13409 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10435) );
  NAND4_X1 U13410 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n10439) );
  AOI211_X1 U13411 ( .C1(n10327), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n10440), .B(n10439), .ZN(n10441) );
  NAND4_X1 U13412 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10485) );
  AOI22_X1 U13413 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10445) );
  OAI21_X1 U13414 ( .B1(n10253), .B2(n18327), .A(n10445), .ZN(n10454) );
  INV_X1 U13415 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U13416 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10452) );
  INV_X1 U13417 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17316) );
  OAI22_X1 U13418 ( .A1(n17275), .A2(n17316), .B1(n17334), .B2(n18650), .ZN(
        n10450) );
  AOI22_X1 U13419 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13420 ( .A1(n10330), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13421 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10446) );
  NAND3_X1 U13422 ( .A1(n10448), .A2(n10447), .A3(n10446), .ZN(n10449) );
  AOI211_X1 U13423 ( .C1(n17205), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n10450), .B(n10449), .ZN(n10451) );
  OAI211_X1 U13424 ( .C1(n17300), .C2(n17186), .A(n10452), .B(n10451), .ZN(
        n10453) );
  AOI211_X4 U13425 ( .C1(n10329), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n10454), .B(n10453), .ZN(n18324) );
  NOR2_X1 U13426 ( .A1(n17374), .A2(n9752), .ZN(n18804) );
  NAND2_X1 U13427 ( .A1(n17374), .A2(n9752), .ZN(n10526) );
  OAI211_X1 U13428 ( .C1(n18341), .C2(n18804), .A(n10526), .B(n10531), .ZN(
        n10455) );
  INV_X1 U13429 ( .A(n10455), .ZN(n10456) );
  NAND2_X1 U13430 ( .A1(n10459), .A2(n10456), .ZN(n10490) );
  INV_X1 U13431 ( .A(n18804), .ZN(n10464) );
  NAND3_X1 U13432 ( .A1(n18330), .A2(n18319), .A3(n10526), .ZN(n10457) );
  INV_X1 U13433 ( .A(n18341), .ZN(n15742) );
  NAND2_X1 U13434 ( .A1(n15742), .A2(n18352), .ZN(n18784) );
  INV_X1 U13435 ( .A(n18784), .ZN(n10524) );
  AOI21_X1 U13436 ( .B1(n10464), .B2(n10457), .A(n10524), .ZN(n10462) );
  OAI21_X1 U13437 ( .B1(n10460), .B2(n18361), .A(n15742), .ZN(n10458) );
  OAI21_X1 U13438 ( .B1(n10460), .B2(n10459), .A(n10458), .ZN(n10461) );
  AOI211_X2 U13439 ( .C1(n18335), .C2(n10463), .A(n10462), .B(n10461), .ZN(
        n10535) );
  INV_X1 U13440 ( .A(n10535), .ZN(n10465) );
  NAND2_X1 U13441 ( .A1(n18324), .A2(n17523), .ZN(n10523) );
  AOI21_X1 U13442 ( .B1(n17456), .B2(n10464), .A(n10523), .ZN(n10532) );
  AOI211_X1 U13443 ( .C1(n10528), .C2(n10490), .A(n10465), .B(n10532), .ZN(
        n15852) );
  NAND2_X1 U13444 ( .A1(n18565), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10480) );
  OAI21_X1 U13445 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18565), .A(
        n10480), .ZN(n10483) );
  OAI22_X1 U13446 ( .A1(n18951), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18809), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10479) );
  NOR2_X1 U13447 ( .A1(n10483), .A2(n10479), .ZN(n10478) );
  OAI22_X1 U13448 ( .A1(n18944), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18814), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10474) );
  NOR2_X1 U13449 ( .A1(n10479), .A2(n10480), .ZN(n10466) );
  OAI22_X1 U13450 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18818), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10468), .ZN(n10470) );
  NOR2_X1 U13451 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18818), .ZN(
        n10469) );
  NAND2_X1 U13452 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10468), .ZN(
        n10471) );
  AOI22_X1 U13453 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10470), .B1(
        n10469), .B2(n10471), .ZN(n10477) );
  AOI21_X1 U13454 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n10471), .A(
        n10470), .ZN(n10472) );
  AOI21_X1 U13455 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18818), .A(
        n10472), .ZN(n10481) );
  NAND2_X1 U13456 ( .A1(n10475), .A2(n10474), .ZN(n10473) );
  OAI211_X1 U13457 ( .C1(n10475), .C2(n10474), .A(n10477), .B(n10473), .ZN(
        n10484) );
  NAND2_X1 U13458 ( .A1(n10481), .A2(n10484), .ZN(n10476) );
  INV_X1 U13459 ( .A(n9752), .ZN(n17377) );
  NAND2_X1 U13460 ( .A1(n17377), .A2(n18330), .ZN(n10534) );
  INV_X1 U13461 ( .A(n10534), .ZN(n10525) );
  XNOR2_X1 U13462 ( .A(n10480), .B(n10479), .ZN(n10482) );
  OAI21_X1 U13463 ( .B1(n10482), .B2(n10484), .A(n10481), .ZN(n16489) );
  INV_X1 U13464 ( .A(n16489), .ZN(n18771) );
  NOR2_X1 U13465 ( .A1(n10484), .A2(n10483), .ZN(n16488) );
  NOR2_X1 U13466 ( .A1(n18324), .A2(n10485), .ZN(n10487) );
  NAND2_X1 U13467 ( .A1(n10487), .A2(n17374), .ZN(n10491) );
  NAND2_X1 U13468 ( .A1(n18852), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18984) );
  NAND2_X1 U13469 ( .A1(n18983), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18917) );
  OAI211_X1 U13470 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18852), .B(n18910), .ZN(n18850) );
  OAI21_X1 U13471 ( .B1(n18330), .B2(n18970), .A(n18850), .ZN(n10486) );
  NAND2_X1 U13472 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18979) );
  OAI21_X1 U13473 ( .B1(n10487), .B2(n10486), .A(n18979), .ZN(n16649) );
  OAI22_X1 U13474 ( .A1(n16488), .A2(n10491), .B1(n10525), .B2(n16649), .ZN(
        n10488) );
  AOI22_X1 U13475 ( .A1(n18768), .A2(n10525), .B1(n18771), .B2(n10488), .ZN(
        n10489) );
  INV_X1 U13476 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18937) );
  NAND2_X1 U13477 ( .A1(n18937), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18836) );
  NAND2_X1 U13478 ( .A1(n18274), .A2(n16536), .ZN(n18137) );
  NAND2_X1 U13479 ( .A1(n16499), .A2(n18203), .ZN(n10554) );
  INV_X1 U13480 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17638) );
  NOR2_X1 U13481 ( .A1(n18009), .A2(n17638), .ZN(n15856) );
  NAND2_X1 U13482 ( .A1(n15856), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10544) );
  INV_X1 U13483 ( .A(n10544), .ZN(n16504) );
  NOR2_X1 U13484 ( .A1(n10494), .A2(n10493), .ZN(n10505) );
  INV_X1 U13485 ( .A(n17507), .ZN(n10495) );
  NOR2_X1 U13486 ( .A1(n10505), .A2(n10495), .ZN(n10503) );
  NOR2_X1 U13487 ( .A1(n17502), .A2(n10503), .ZN(n10501) );
  NAND2_X1 U13488 ( .A1(n10501), .A2(n10502), .ZN(n10499) );
  NOR2_X1 U13489 ( .A1(n17495), .A2(n10499), .ZN(n10498) );
  NAND2_X1 U13490 ( .A1(n10498), .A2(n10496), .ZN(n10497) );
  NOR2_X1 U13491 ( .A1(n17488), .A2(n10497), .ZN(n10520) );
  XOR2_X1 U13492 ( .A(n17488), .B(n10497), .Z(n17916) );
  XNOR2_X1 U13493 ( .A(n17492), .B(n10498), .ZN(n10513) );
  XOR2_X1 U13494 ( .A(n17495), .B(n10499), .Z(n10500) );
  NAND2_X1 U13495 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10500), .ZN(
        n10512) );
  XOR2_X1 U13496 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n10500), .Z(
        n17934) );
  XOR2_X1 U13497 ( .A(n10502), .B(n10501), .Z(n17948) );
  XOR2_X1 U13498 ( .A(n10503), .B(n17502), .Z(n10504) );
  NAND2_X1 U13499 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10504), .ZN(
        n10510) );
  XOR2_X1 U13500 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n10504), .Z(
        n17966) );
  XNOR2_X1 U13501 ( .A(n17507), .B(n10505), .ZN(n10506) );
  OR2_X1 U13502 ( .A1(n20943), .A2(n10506), .ZN(n10509) );
  XOR2_X1 U13503 ( .A(n20943), .B(n10506), .Z(n18272) );
  AOI21_X1 U13504 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17512), .A(
        n17993), .ZN(n10508) );
  INV_X1 U13505 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18954) );
  NOR2_X1 U13506 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17512), .ZN(
        n10507) );
  AOI221_X1 U13507 ( .B1(n17993), .B2(n17512), .C1(n10508), .C2(n18954), .A(
        n10507), .ZN(n18271) );
  NAND2_X1 U13508 ( .A1(n18272), .A2(n18271), .ZN(n18270) );
  NAND2_X1 U13509 ( .A1(n10509), .A2(n18270), .ZN(n17965) );
  NAND2_X1 U13510 ( .A1(n17966), .A2(n17965), .ZN(n17964) );
  NAND2_X1 U13511 ( .A1(n10510), .A2(n17964), .ZN(n17949) );
  NAND2_X1 U13512 ( .A1(n17948), .A2(n17949), .ZN(n17947) );
  NOR2_X1 U13513 ( .A1(n17948), .A2(n17949), .ZN(n10511) );
  NAND2_X1 U13514 ( .A1(n17934), .A2(n17933), .ZN(n17932) );
  NAND2_X1 U13515 ( .A1(n10512), .A2(n17932), .ZN(n10514) );
  NAND2_X1 U13516 ( .A1(n10513), .A2(n10514), .ZN(n10515) );
  XOR2_X1 U13517 ( .A(n10514), .B(n10513), .Z(n17922) );
  NAND2_X1 U13518 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17922), .ZN(
        n17921) );
  NAND2_X1 U13519 ( .A1(n10520), .A2(n10516), .ZN(n10521) );
  INV_X1 U13520 ( .A(n10516), .ZN(n10519) );
  NAND2_X1 U13521 ( .A1(n17916), .A2(n17915), .ZN(n10518) );
  NAND2_X1 U13522 ( .A1(n10520), .A2(n10519), .ZN(n10517) );
  OAI211_X1 U13523 ( .C1(n10520), .C2(n10519), .A(n10518), .B(n10517), .ZN(
        n17895) );
  NAND2_X1 U13524 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17895), .ZN(
        n17894) );
  NAND2_X1 U13525 ( .A1(n18002), .A2(n17678), .ZN(n18004) );
  NAND2_X1 U13526 ( .A1(n16504), .A2(n17637), .ZN(n16505) );
  INV_X1 U13527 ( .A(n16505), .ZN(n16527) );
  NAND2_X1 U13528 ( .A1(n16527), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10522) );
  XNOR2_X1 U13529 ( .A(n18939), .B(n10522), .ZN(n16502) );
  NAND2_X1 U13530 ( .A1(n10529), .A2(n10523), .ZN(n18988) );
  NAND3_X1 U13531 ( .A1(n10531), .A2(n10525), .A3(n10524), .ZN(n15739) );
  NAND2_X1 U13532 ( .A1(n18324), .A2(n18319), .ZN(n15939) );
  INV_X1 U13533 ( .A(n10531), .ZN(n10527) );
  NAND3_X1 U13534 ( .A1(n18330), .A2(n18341), .A3(n18352), .ZN(n10533) );
  NOR2_X1 U13535 ( .A1(n10531), .A2(n15845), .ZN(n10537) );
  AOI21_X1 U13536 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(n10536) );
  NAND2_X1 U13537 ( .A1(n18041), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17670) );
  NAND2_X1 U13538 ( .A1(n18006), .A2(n15856), .ZN(n16541) );
  NAND3_X1 U13539 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n18939), .ZN(n10547) );
  INV_X1 U13540 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16518) );
  NAND2_X1 U13541 ( .A1(n18006), .A2(n16504), .ZN(n16525) );
  OAI21_X1 U13542 ( .B1(n16518), .B2(n16525), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10540) );
  OAI21_X1 U13543 ( .B1(n16541), .B2(n10547), .A(n10540), .ZN(n16496) );
  INV_X1 U13544 ( .A(n18274), .ZN(n18773) );
  NAND2_X1 U13545 ( .A1(n17488), .A2(n18297), .ZN(n18036) );
  NOR2_X1 U13546 ( .A1(n18218), .A2(n18289), .ZN(n18292) );
  INV_X1 U13547 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18914) );
  NOR2_X1 U13548 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18987) );
  NOR2_X1 U13549 ( .A1(n18914), .A2(n18199), .ZN(n16495) );
  INV_X2 U13550 ( .A(n18199), .ZN(n18301) );
  NAND3_X1 U13551 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18107) );
  AOI21_X1 U13552 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18275) );
  OR2_X1 U13553 ( .A1(n18107), .A2(n18275), .ZN(n18217) );
  NAND3_X1 U13554 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18109) );
  OR2_X1 U13555 ( .A1(n18217), .A2(n18109), .ZN(n18121) );
  NOR2_X1 U13556 ( .A1(n18110), .A2(n18121), .ZN(n18020) );
  INV_X1 U13557 ( .A(n18020), .ZN(n18061) );
  INV_X1 U13558 ( .A(n18021), .ZN(n18049) );
  NAND2_X1 U13559 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18023) );
  NOR3_X1 U13560 ( .A1(n18049), .A2(n10545), .A3(n18023), .ZN(n16503) );
  INV_X1 U13561 ( .A(n16503), .ZN(n18007) );
  OAI21_X1 U13562 ( .B1(n18061), .B2(n18007), .A(n18780), .ZN(n18001) );
  INV_X1 U13563 ( .A(n18110), .ZN(n16538) );
  INV_X1 U13564 ( .A(n18109), .ZN(n10541) );
  NAND2_X1 U13565 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18248) );
  NOR2_X1 U13566 ( .A1(n18107), .A2(n18248), .ZN(n18215) );
  NAND2_X1 U13567 ( .A1(n10541), .A2(n18215), .ZN(n18120) );
  NOR2_X1 U13568 ( .A1(n18954), .A2(n18120), .ZN(n18185) );
  NAND2_X1 U13569 ( .A1(n16538), .A2(n18185), .ZN(n18122) );
  NAND2_X1 U13570 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16503), .ZN(
        n16539) );
  OAI21_X1 U13571 ( .B1(n18122), .B2(n16539), .A(n9773), .ZN(n10543) );
  NOR2_X1 U13572 ( .A1(n18110), .A2(n18120), .ZN(n18100) );
  INV_X1 U13573 ( .A(n18100), .ZN(n18064) );
  INV_X1 U13574 ( .A(n18805), .ZN(n18778) );
  OAI21_X1 U13575 ( .B1(n18007), .B2(n18064), .A(n18778), .ZN(n10542) );
  NAND4_X1 U13576 ( .A1(n18285), .A2(n18001), .A3(n10543), .A4(n10542), .ZN(
        n15860) );
  AOI22_X1 U13577 ( .A1(n18292), .A2(n10544), .B1(n18199), .B2(n15860), .ZN(
        n15928) );
  NOR2_X1 U13578 ( .A1(n10545), .A2(n18023), .ZN(n10546) );
  INV_X1 U13579 ( .A(n18780), .ZN(n18798) );
  AOI21_X1 U13580 ( .B1(n9773), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18778), .ZN(n18276) );
  OAI22_X1 U13581 ( .A1(n18798), .A2(n18061), .B1(n18064), .B2(n18276), .ZN(
        n16537) );
  AND2_X1 U13582 ( .A1(n16537), .A2(n18021), .ZN(n18024) );
  NAND4_X1 U13583 ( .A1(n15856), .A2(n18298), .A3(n10546), .A4(n18024), .ZN(
        n15857) );
  OAI22_X1 U13584 ( .A1(n15928), .A2(n18939), .B1(n10547), .B2(n15857), .ZN(
        n10548) );
  AOI211_X1 U13585 ( .C1(n10549), .C2(n18292), .A(n16495), .B(n10548), .ZN(
        n10550) );
  INV_X1 U13586 ( .A(n10552), .ZN(n10553) );
  AND2_X4 U13587 ( .A1(n10795), .A2(n13602), .ZN(n12429) );
  AOI22_X1 U13588 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10556) );
  AND2_X4 U13589 ( .A1(n10794), .A2(n15720), .ZN(n12430) );
  AOI22_X1 U13590 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10778), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10555) );
  NAND2_X1 U13591 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10557) );
  NAND2_X1 U13592 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10561) );
  AND2_X4 U13593 ( .A1(n10788), .A2(n13602), .ZN(n10780) );
  AOI22_X1 U13594 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13595 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13596 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10564) );
  NAND4_X1 U13597 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10568) );
  AOI22_X1 U13598 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10778), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13599 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12456), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13600 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13601 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13602 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12430), .B1(
        n10778), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13603 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13604 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13605 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13606 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13607 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10581) );
  NAND2_X1 U13608 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10580) );
  NAND2_X1 U13609 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10579) );
  NAND3_X1 U13610 ( .A1(n10581), .A2(n10580), .A3(n10579), .ZN(n10582) );
  AOI22_X1 U13611 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12456), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13612 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10585) );
  NAND2_X1 U13613 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10584) );
  NAND3_X1 U13614 ( .A1(n10586), .A2(n10585), .A3(n10584), .ZN(n10590) );
  NAND2_X1 U13615 ( .A1(n10588), .A2(n10587), .ZN(n10589) );
  AOI22_X1 U13616 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U13617 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12456), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13618 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13619 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10593) );
  NAND4_X1 U13620 ( .A1(n10596), .A2(n10595), .A3(n10594), .A4(n10593), .ZN(
        n10597) );
  AOI22_X1 U13621 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9753), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13622 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13623 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10598) );
  NAND4_X1 U13624 ( .A1(n10601), .A2(n10600), .A3(n10599), .A4(n10598), .ZN(
        n10602) );
  NAND2_X1 U13625 ( .A1(n10602), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10603) );
  NAND2_X2 U13626 ( .A1(n10604), .A2(n10603), .ZN(n10656) );
  AOI22_X1 U13627 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13628 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13629 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13630 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13631 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13632 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12456), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13633 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13634 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13635 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13636 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13637 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13638 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10627) );
  AOI22_X1 U13639 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13640 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13641 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10623) );
  NAND4_X1 U13642 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10626) );
  MUX2_X2 U13643 ( .A(n10627), .B(n10626), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19421) );
  AOI22_X1 U13644 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U13645 ( .A1(n10778), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12456), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U13646 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10629) );
  NAND2_X1 U13647 ( .A1(n10632), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10638) );
  AOI22_X1 U13648 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13649 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12456), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13650 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10634) );
  NAND4_X1 U13651 ( .A1(n10223), .A2(n10636), .A3(n10635), .A4(n10634), .ZN(
        n10637) );
  NAND2_X1 U13652 ( .A1(n11167), .A2(n10221), .ZN(n10640) );
  AND2_X1 U13653 ( .A1(n10657), .A2(n15732), .ZN(n10639) );
  AOI22_X1 U13654 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13655 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9772), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13656 ( .A1(n9753), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13657 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10641) );
  NAND4_X1 U13658 ( .A1(n10644), .A2(n10643), .A3(n10642), .A4(n10641), .ZN(
        n10645) );
  AOI22_X1 U13659 ( .A1(n12430), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10778), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13660 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12456), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13661 ( .A1(n10781), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10646), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13662 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10648) );
  NAND4_X1 U13663 ( .A1(n10651), .A2(n10650), .A3(n10649), .A4(n10648), .ZN(
        n10652) );
  INV_X1 U13664 ( .A(n10656), .ZN(n10653) );
  NAND2_X1 U13665 ( .A1(n10655), .A2(n10654), .ZN(n10661) );
  NAND2_X1 U13666 ( .A1(n11385), .A2(n19421), .ZN(n10682) );
  NAND3_X1 U13667 ( .A1(n10682), .A2(n10668), .A3(n19431), .ZN(n10659) );
  NAND2_X1 U13668 ( .A1(n10661), .A2(n11569), .ZN(n10708) );
  INV_X1 U13669 ( .A(n15732), .ZN(n11565) );
  NAND2_X1 U13670 ( .A1(n11385), .A2(n11565), .ZN(n11193) );
  XNOR2_X1 U13671 ( .A(n12312), .B(n10884), .ZN(n11195) );
  NAND2_X1 U13672 ( .A1(n11195), .A2(n15732), .ZN(n11199) );
  NAND4_X1 U13673 ( .A1(n10884), .A2(n12790), .A3(n15732), .A4(n12312), .ZN(
        n12773) );
  INV_X1 U13674 ( .A(n10665), .ZN(n10666) );
  AND2_X1 U13675 ( .A1(n11566), .A2(n10678), .ZN(n12775) );
  INV_X1 U13676 ( .A(n10669), .ZN(n10670) );
  NOR2_X1 U13677 ( .A1(n10670), .A2(n10662), .ZN(n10671) );
  OR2_X2 U13678 ( .A1(n11366), .A2(n10672), .ZN(n13620) );
  NOR2_X1 U13679 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10735) );
  AND2_X1 U13680 ( .A1(n10676), .A2(n20077), .ZN(n20081) );
  NAND2_X1 U13681 ( .A1(n10680), .A2(n13746), .ZN(n10681) );
  NAND2_X1 U13682 ( .A1(n10681), .A2(n10667), .ZN(n10683) );
  NAND2_X1 U13683 ( .A1(n10683), .A2(n10682), .ZN(n10684) );
  NOR2_X1 U13684 ( .A1(n10893), .A2(n19309), .ZN(n10686) );
  AND2_X2 U13685 ( .A1(n10687), .A2(n10686), .ZN(n10720) );
  AOI22_X1 U13686 ( .A1(n10720), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10690) );
  INV_X2 U13687 ( .A(n10893), .ZN(n10688) );
  NOR2_X2 U13688 ( .A1(n10692), .A2(n12773), .ZN(n11574) );
  NAND2_X1 U13689 ( .A1(n11278), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10689) );
  OAI21_X2 U13690 ( .B1(n9717), .B2(n20922), .A(n10691), .ZN(n10714) );
  INV_X1 U13691 ( .A(n10692), .ZN(n10695) );
  NAND2_X1 U13692 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U13693 ( .A1(n9770), .A2(n10693), .ZN(n10694) );
  OAI21_X1 U13694 ( .B1(n10696), .B2(n10695), .A(n10694), .ZN(n10700) );
  INV_X1 U13695 ( .A(n10697), .ZN(n10698) );
  NAND2_X1 U13696 ( .A1(n10700), .A2(n10699), .ZN(n10743) );
  NAND2_X1 U13697 ( .A1(n11278), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10705) );
  INV_X1 U13698 ( .A(n10735), .ZN(n10702) );
  NAND2_X1 U13699 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U13700 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  AOI21_X1 U13701 ( .B1(n10720), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10703), .ZN(
        n10704) );
  OAI211_X2 U13702 ( .C1(n9727), .C2(n20916), .A(n10710), .B(n10709), .ZN(
        n10742) );
  NAND2_X2 U13703 ( .A1(n10743), .A2(n10742), .ZN(n10726) );
  NAND2_X1 U13704 ( .A1(n10734), .A2(n15720), .ZN(n10712) );
  AOI21_X1 U13705 ( .B1(n19309), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U13706 ( .A1(n10728), .A2(n10725), .ZN(n10713) );
  NAND3_X1 U13707 ( .A1(n10715), .A2(n10726), .A3(n10729), .ZN(n10716) );
  INV_X1 U13708 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19408) );
  AOI22_X1 U13709 ( .A1(n10720), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U13710 ( .A1(n11357), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10721) );
  INV_X1 U13711 ( .A(n9740), .ZN(n10727) );
  INV_X1 U13712 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13269) );
  AOI22_X1 U13713 ( .A1(n10720), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10731) );
  NAND2_X1 U13714 ( .A1(n11357), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13715 ( .A1(n10734), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13716 ( .A1(n10735), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10736) );
  OR2_X1 U13717 ( .A1(n10743), .A2(n10742), .ZN(n10744) );
  INV_X1 U13718 ( .A(n12767), .ZN(n19231) );
  AND2_X1 U13719 ( .A1(n10758), .A2(n19231), .ZN(n10747) );
  AND2_X1 U13720 ( .A1(n10769), .A2(n10747), .ZN(n10746) );
  INV_X1 U13721 ( .A(n10758), .ZN(n10745) );
  AOI22_X1 U13722 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19742), .B1(
        n10942), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13724 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19506), .B1(
        n19608), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10754) );
  AND2_X1 U13725 ( .A1(n10769), .A2(n10748), .ZN(n10750) );
  AOI22_X1 U13726 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19441), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13727 ( .A1(n10943), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10941), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10752) );
  INV_X1 U13728 ( .A(n10764), .ZN(n10757) );
  INV_X1 U13729 ( .A(n10769), .ZN(n10756) );
  INV_X2 U13730 ( .A(n9774), .ZN(n15080) );
  INV_X1 U13731 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U13732 ( .A1(n10769), .A2(n9774), .ZN(n10761) );
  INV_X1 U13733 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10760) );
  OAI22_X1 U13734 ( .A1(n12320), .A2(n10986), .B1(n19474), .B2(n10760), .ZN(
        n10768) );
  INV_X1 U13735 ( .A(n10764), .ZN(n10763) );
  INV_X1 U13736 ( .A(n10761), .ZN(n10762) );
  INV_X1 U13737 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10766) );
  INV_X1 U13738 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10765) );
  NOR2_X1 U13739 ( .A1(n10768), .A2(n10767), .ZN(n10773) );
  NOR2_X4 U13740 ( .A1(n10771), .A2(n15080), .ZN(n10939) );
  AOI22_X1 U13741 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13738), .B1(
        n10939), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10772) );
  NAND4_X1 U13742 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(
        n10777) );
  NAND2_X1 U13743 ( .A1(n10777), .A2(n13331), .ZN(n10804) );
  AND2_X2 U13744 ( .A1(n9754), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10909) );
  INV_X1 U13745 ( .A(n10779), .ZN(n10963) );
  AOI22_X1 U13746 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10909), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10785) );
  BUF_X1 U13747 ( .A(n12430), .Z(n10796) );
  AOI22_X1 U13748 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10849), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10784) );
  AND2_X2 U13749 ( .A1(n12591), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10850) );
  AOI22_X1 U13750 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10783) );
  INV_X1 U13751 ( .A(n10781), .ZN(n13584) );
  AND2_X2 U13752 ( .A1(n10786), .A2(n13590), .ZN(n10820) );
  INV_X1 U13753 ( .A(n10646), .ZN(n12426) );
  INV_X1 U13754 ( .A(n12426), .ZN(n10787) );
  AND2_X2 U13755 ( .A1(n10787), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11419) );
  AOI22_X1 U13756 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10820), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10782) );
  NAND4_X1 U13757 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10802) );
  AND2_X2 U13758 ( .A1(n10787), .A2(n13590), .ZN(n11420) );
  AOI22_X1 U13759 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10863), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10800) );
  INV_X1 U13760 ( .A(n10839), .ZN(n10964) );
  INV_X1 U13761 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10792) );
  AND2_X2 U13762 ( .A1(n10788), .A2(n12424), .ZN(n12447) );
  NAND2_X1 U13763 ( .A1(n12447), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10791) );
  NAND2_X1 U13764 ( .A1(n10840), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10790) );
  OAI211_X1 U13765 ( .C1(n10964), .C2(n10792), .A(n10791), .B(n10790), .ZN(
        n10793) );
  INV_X1 U13766 ( .A(n10793), .ZN(n10799) );
  AND2_X1 U13767 ( .A1(n10794), .A2(n12424), .ZN(n10825) );
  AND2_X1 U13768 ( .A1(n12424), .A2(n9742), .ZN(n10841) );
  AOI22_X1 U13769 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10798) );
  AND2_X2 U13770 ( .A1(n10796), .A2(n13590), .ZN(n10832) );
  NAND2_X1 U13771 ( .A1(n10832), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10797) );
  NAND4_X1 U13772 ( .A1(n10800), .A2(n10799), .A3(n10798), .A4(n10797), .ZN(
        n10801) );
  INV_X1 U13773 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10805) );
  NAND3_X1 U13774 ( .A1(n9828), .A2(n10807), .A3(n10806), .ZN(n10808) );
  INV_X1 U13775 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10810) );
  INV_X1 U13776 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10809) );
  OAI22_X1 U13777 ( .A1(n10810), .A2(n19640), .B1(n19711), .B2(n10809), .ZN(
        n10811) );
  AOI21_X1 U13778 ( .B1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n10940), .A(
        n10811), .ZN(n10818) );
  AOI22_X1 U13779 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10939), .B1(
        n10938), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13780 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19506), .B1(
        n10941), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13781 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19742), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10814) );
  INV_X1 U13782 ( .A(n10986), .ZN(n13663) );
  NAND2_X1 U13783 ( .A1(n13663), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10812) );
  NAND4_X1 U13784 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10862) );
  AOI22_X1 U13785 ( .A1(n10909), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13786 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13787 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13788 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n10833), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10821) );
  NAND4_X1 U13789 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n10831) );
  AOI22_X1 U13790 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13791 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13792 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13793 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U13794 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10830) );
  NOR2_X1 U13795 ( .A1(n10831), .A2(n10830), .ZN(n12727) );
  AOI22_X1 U13796 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13797 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13798 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10836) );
  INV_X1 U13799 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19413) );
  AOI22_X1 U13800 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10820), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10835) );
  NAND4_X1 U13801 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10847) );
  AOI22_X1 U13802 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13803 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13804 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13805 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10842) );
  NAND4_X1 U13806 ( .A1(n10845), .A2(n10844), .A3(n10843), .A4(n10842), .ZN(
        n10846) );
  NAND2_X1 U13807 ( .A1(n11377), .A2(n11386), .ZN(n10848) );
  OR2_X1 U13808 ( .A1(n12727), .A2(n10848), .ZN(n11213) );
  AOI22_X1 U13809 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13810 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13811 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13812 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10851) );
  NAND4_X1 U13813 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10860) );
  AOI22_X1 U13814 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13815 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13816 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13817 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10855) );
  NAND4_X1 U13818 ( .A1(n10858), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(
        n10859) );
  NAND2_X1 U13819 ( .A1(n11213), .A2(n11214), .ZN(n10861) );
  NAND2_X1 U13820 ( .A1(n10832), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10867) );
  NAND2_X1 U13821 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10866) );
  NAND2_X1 U13822 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10865) );
  NAND2_X1 U13823 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10864) );
  AOI22_X1 U13824 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13825 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U13826 ( .A1(n10839), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10869) );
  NAND2_X1 U13827 ( .A1(n10779), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10868) );
  NAND2_X1 U13828 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10875) );
  NAND2_X1 U13829 ( .A1(n10909), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10874) );
  NAND2_X1 U13830 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10873) );
  NAND2_X1 U13831 ( .A1(n10834), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10872) );
  AOI22_X1 U13832 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10876) );
  NAND4_X1 U13833 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(
        n11011) );
  INV_X1 U13834 ( .A(n11011), .ZN(n11023) );
  MUX2_X1 U13835 ( .A(n10880), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11150) );
  NAND2_X1 U13836 ( .A1(n11150), .A2(n11151), .ZN(n10882) );
  NAND2_X1 U13837 ( .A1(n10880), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10881) );
  XNOR2_X1 U13838 ( .A(n15720), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10887) );
  INV_X1 U13839 ( .A(n10887), .ZN(n10883) );
  XNOR2_X1 U13840 ( .A(n10888), .B(n10883), .ZN(n11177) );
  NAND2_X1 U13841 ( .A1(n10924), .A2(n11177), .ZN(n11179) );
  OAI21_X1 U13842 ( .B1(n11214), .B2(n10924), .A(n11179), .ZN(n10885) );
  INV_X1 U13843 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12824) );
  MUX2_X1 U13844 ( .A(n10885), .B(n12824), .S(n11375), .Z(n10904) );
  NOR2_X1 U13845 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10886) );
  MUX2_X1 U13846 ( .A(n11386), .B(n10886), .S(n11375), .Z(n10903) );
  NAND2_X1 U13847 ( .A1(n10904), .A2(n10903), .ZN(n10908) );
  NAND2_X1 U13848 ( .A1(n10888), .A2(n10887), .ZN(n10890) );
  NAND2_X1 U13849 ( .A1(n20047), .A2(n15720), .ZN(n10889) );
  MUX2_X1 U13850 ( .A(n12315), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10921) );
  INV_X1 U13851 ( .A(n10921), .ZN(n10891) );
  XNOR2_X1 U13852 ( .A(n10922), .B(n10891), .ZN(n11148) );
  INV_X1 U13853 ( .A(n11148), .ZN(n10892) );
  NAND2_X1 U13854 ( .A1(n10893), .A2(n10892), .ZN(n10894) );
  MUX2_X1 U13855 ( .A(n10895), .B(P2_EBX_REG_3__SCAN_IN), .S(n11375), .Z(
        n10907) );
  XNOR2_X1 U13856 ( .A(n10908), .B(n10907), .ZN(n15055) );
  NAND2_X1 U13857 ( .A1(n10896), .A2(n15055), .ZN(n13272) );
  INV_X1 U13858 ( .A(n11151), .ZN(n10898) );
  NAND2_X1 U13859 ( .A1(n10559), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10897) );
  AND2_X1 U13860 ( .A1(n10898), .A2(n10897), .ZN(n11158) );
  INV_X1 U13861 ( .A(n11158), .ZN(n11173) );
  MUX2_X1 U13862 ( .A(n12727), .B(n11173), .S(n10924), .Z(n11164) );
  INV_X1 U13863 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10899) );
  MUX2_X1 U13864 ( .A(n11164), .B(n10899), .S(n11375), .Z(n19229) );
  NOR2_X1 U13865 ( .A1(n19229), .A2(n20916), .ZN(n12737) );
  INV_X1 U13866 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10900) );
  NOR3_X1 U13867 ( .A1(n13659), .A2(n10899), .A3(n10900), .ZN(n10901) );
  NOR2_X1 U13868 ( .A1(n10903), .A2(n10901), .ZN(n15077) );
  NAND2_X1 U13869 ( .A1(n12737), .A2(n15077), .ZN(n12736) );
  NOR2_X1 U13870 ( .A1(n12737), .A2(n15077), .ZN(n10902) );
  AOI21_X1 U13871 ( .B1(n20922), .B2(n12736), .A(n10902), .ZN(n14389) );
  XNOR2_X1 U13872 ( .A(n10904), .B(n10903), .ZN(n15066) );
  XNOR2_X1 U13873 ( .A(n15066), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14387) );
  INV_X1 U13874 ( .A(n15066), .ZN(n10905) );
  AND2_X1 U13875 ( .A1(n10905), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10906) );
  AOI21_X1 U13876 ( .B1(n14389), .B2(n14387), .A(n10906), .ZN(n13270) );
  INV_X1 U13877 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U13878 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10850), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13879 ( .A1(n10909), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13880 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10832), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13881 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11420), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10910) );
  NAND4_X1 U13882 ( .A1(n10913), .A2(n10912), .A3(n10911), .A4(n10910), .ZN(
        n10919) );
  AOI22_X1 U13883 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13884 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10863), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13885 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13886 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10914) );
  NAND4_X1 U13887 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10918) );
  NOR2_X1 U13888 ( .A1(n13590), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10920) );
  NOR2_X1 U13889 ( .A1(n15937), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10923) );
  NAND2_X1 U13890 ( .A1(n11153), .A2(n10923), .ZN(n11149) );
  MUX2_X1 U13891 ( .A(n11403), .B(n11149), .S(n10924), .Z(n10925) );
  MUX2_X1 U13892 ( .A(n14377), .B(n10925), .S(n13659), .Z(n10927) );
  AND2_X2 U13893 ( .A1(n10926), .A2(n10927), .ZN(n11006) );
  INV_X1 U13894 ( .A(n11006), .ZN(n10931) );
  INV_X1 U13895 ( .A(n10926), .ZN(n10929) );
  INV_X1 U13896 ( .A(n10927), .ZN(n10928) );
  NAND2_X1 U13897 ( .A1(n10929), .A2(n10928), .ZN(n10930) );
  NAND2_X1 U13898 ( .A1(n10931), .A2(n10930), .ZN(n19209) );
  INV_X1 U13899 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21003) );
  XNOR2_X1 U13900 ( .A(n19209), .B(n21003), .ZN(n13377) );
  INV_X1 U13901 ( .A(n13377), .ZN(n10932) );
  NAND2_X1 U13902 ( .A1(n10933), .A2(n10932), .ZN(n13376) );
  INV_X1 U13903 ( .A(n19209), .ZN(n10934) );
  NAND2_X1 U13904 ( .A1(n10934), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10935) );
  NAND2_X1 U13905 ( .A1(n13376), .A2(n10935), .ZN(n13767) );
  INV_X1 U13906 ( .A(n10936), .ZN(n10937) );
  INV_X1 U13907 ( .A(n11403), .ZN(n11223) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n13738), .B1(
        n10938), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13909 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10939), .B1(
        n10940), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U13910 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10941), .B1(
        n19742), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13911 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19441), .B1(
        n19506), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13912 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n10942), .B1(
        n10943), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13913 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19608), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10945) );
  INV_X1 U13914 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13669) );
  INV_X1 U13915 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10949) );
  OAI22_X1 U13916 ( .A1(n13669), .A2(n10986), .B1(n19640), .B2(n10949), .ZN(
        n10953) );
  INV_X1 U13917 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10951) );
  INV_X1 U13918 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10950) );
  OAI22_X1 U13919 ( .A1(n10951), .A2(n19474), .B1(n19711), .B2(n10950), .ZN(
        n10952) );
  NOR2_X1 U13920 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  NAND4_X1 U13921 ( .A1(n10957), .A2(n10956), .A3(n10955), .A4(n10954), .ZN(
        n10974) );
  AOI22_X1 U13922 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13923 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13924 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13925 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10958) );
  NAND4_X1 U13926 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10971) );
  INV_X1 U13927 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20860) );
  INV_X1 U13928 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10962) );
  OAI22_X1 U13929 ( .A1(n20860), .A2(n10964), .B1(n10963), .B2(n10962), .ZN(
        n10965) );
  INV_X1 U13930 ( .A(n10965), .ZN(n10969) );
  AOI22_X1 U13931 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13932 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13933 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10966) );
  NAND4_X1 U13934 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10970) );
  INV_X1 U13935 ( .A(n11407), .ZN(n10972) );
  NAND2_X1 U13936 ( .A1(n10972), .A2(n11377), .ZN(n10973) );
  XNOR2_X2 U13937 ( .A(n11225), .B(n9812), .ZN(n11230) );
  NAND2_X1 U13938 ( .A1(n11230), .A2(n11023), .ZN(n10975) );
  INV_X1 U13939 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19198) );
  MUX2_X1 U13940 ( .A(n11407), .B(n19198), .S(n11375), .Z(n11005) );
  XNOR2_X1 U13941 ( .A(n11006), .B(n11005), .ZN(n19193) );
  INV_X1 U13942 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13785) );
  NAND2_X1 U13943 ( .A1(n13766), .A2(n13767), .ZN(n13765) );
  NAND2_X1 U13944 ( .A1(n10976), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10977) );
  NAND2_X2 U13945 ( .A1(n10978), .A2(n9812), .ZN(n11241) );
  AOI22_X1 U13946 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10940), .B1(
        n10938), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13947 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13738), .B1(
        n10939), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13948 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10941), .B1(
        n10943), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U13949 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19441), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U13950 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19742), .B1(
        n10942), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U13951 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19506), .B1(
        n19608), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10979) );
  INV_X1 U13952 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10984) );
  INV_X1 U13953 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10983) );
  OAI22_X1 U13954 ( .A1(n10984), .A2(n19711), .B1(n19640), .B2(n10983), .ZN(
        n10988) );
  INV_X1 U13955 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19429) );
  INV_X1 U13956 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10985) );
  OAI22_X1 U13957 ( .A1(n19429), .A2(n10986), .B1(n19474), .B2(n10985), .ZN(
        n10987) );
  NOR2_X1 U13958 ( .A1(n10988), .A2(n10987), .ZN(n10989) );
  NAND4_X1 U13959 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n11004) );
  AOI22_X1 U13960 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U13961 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U13962 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13963 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10863), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U13964 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n11002) );
  AOI22_X1 U13965 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13966 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11420), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U13967 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10841), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13968 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10825), .B1(
        n12447), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10997) );
  NAND4_X1 U13969 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11001) );
  NAND2_X1 U13970 ( .A1(n11410), .A2(n11377), .ZN(n11003) );
  XNOR2_X2 U13971 ( .A(n11241), .B(n11240), .ZN(n11236) );
  MUX2_X1 U13972 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11410), .S(n13659), .Z(
        n11009) );
  XNOR2_X1 U13973 ( .A(n11010), .B(n11009), .ZN(n19175) );
  INV_X1 U13974 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U13975 ( .A1(n11007), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11008) );
  INV_X1 U13976 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n19168) );
  MUX2_X1 U13977 ( .A(n19168), .B(n11011), .S(n13659), .Z(n11013) );
  NAND2_X1 U13978 ( .A1(n11375), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11012) );
  XNOR2_X1 U13979 ( .A(n11019), .B(n11012), .ZN(n19154) );
  NAND2_X1 U13980 ( .A1(n19154), .A2(n11011), .ZN(n11016) );
  INV_X1 U13981 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20987) );
  OR2_X1 U13982 ( .A1(n11016), .A2(n20987), .ZN(n16413) );
  INV_X1 U13983 ( .A(n11013), .ZN(n11014) );
  XNOR2_X1 U13984 ( .A(n11015), .B(n11014), .ZN(n19166) );
  NAND2_X1 U13985 ( .A1(n19166), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16414) );
  NAND2_X1 U13986 ( .A1(n11016), .A2(n20987), .ZN(n16412) );
  INV_X1 U13987 ( .A(n19166), .ZN(n11017) );
  INV_X1 U13988 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U13989 ( .A1(n11017), .A2(n11253), .ZN(n16416) );
  AND2_X1 U13990 ( .A1(n16412), .A2(n16416), .ZN(n11018) );
  INV_X1 U13991 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11021) );
  NOR2_X1 U13992 ( .A1(n13659), .A2(n11021), .ZN(n11022) );
  XNOR2_X1 U13993 ( .A(n11024), .B(n11022), .ZN(n19138) );
  AOI21_X1 U13994 ( .B1(n19138), .B2(n11621), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15670) );
  NAND2_X1 U13995 ( .A1(n11375), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11025) );
  MUX2_X1 U13996 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11025), .S(n11027), .Z(
        n11026) );
  AND2_X1 U13997 ( .A1(n11026), .A2(n11125), .ZN(n19128) );
  NAND2_X1 U13998 ( .A1(n19128), .A2(n11621), .ZN(n11035) );
  INV_X1 U13999 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15657) );
  NAND2_X1 U14000 ( .A1(n11035), .A2(n15657), .ZN(n15385) );
  NAND2_X1 U14001 ( .A1(n11375), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11028) );
  OR2_X1 U14002 ( .A1(n11029), .A2(n11028), .ZN(n11031) );
  INV_X1 U14003 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19113) );
  INV_X1 U14004 ( .A(n11036), .ZN(n11030) );
  NAND2_X1 U14005 ( .A1(n11031), .A2(n11030), .ZN(n19115) );
  OR2_X1 U14006 ( .A1(n19115), .A2(n11023), .ZN(n11032) );
  INV_X1 U14007 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15638) );
  NAND2_X1 U14008 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11033) );
  OR2_X1 U14009 ( .A1(n19115), .A2(n11033), .ZN(n15641) );
  AND2_X1 U14010 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U14011 ( .A1(n19138), .A2(n11034), .ZN(n15386) );
  OR2_X1 U14012 ( .A1(n15657), .A2(n11035), .ZN(n15384) );
  AND2_X1 U14013 ( .A1(n15386), .A2(n15384), .ZN(n15639) );
  NAND2_X1 U14014 ( .A1(n15641), .A2(n15639), .ZN(n15622) );
  NAND2_X1 U14015 ( .A1(n11375), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11037) );
  NAND2_X1 U14016 ( .A1(n10013), .A2(n11038), .ZN(n11039) );
  NAND2_X1 U14017 ( .A1(n11068), .A2(n11039), .ZN(n13328) );
  NAND2_X1 U14018 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11040) );
  NOR2_X1 U14019 ( .A1(n13328), .A2(n11040), .ZN(n15625) );
  NOR2_X1 U14020 ( .A1(n15622), .A2(n15625), .ZN(n15327) );
  OR2_X1 U14021 ( .A1(n13328), .A2(n11023), .ZN(n11041) );
  NAND2_X1 U14022 ( .A1(n11041), .A2(n20891), .ZN(n15326) );
  INV_X1 U14023 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11293) );
  NOR2_X1 U14024 ( .A1(n13659), .A2(n11293), .ZN(n11067) );
  NOR2_X1 U14025 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n11043) );
  INV_X1 U14026 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11062) );
  INV_X1 U14027 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U14028 ( .A1(n11062), .A2(n11044), .ZN(n11045) );
  INV_X1 U14029 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15169) );
  INV_X1 U14030 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11046) );
  NAND2_X1 U14031 ( .A1(n15169), .A2(n11046), .ZN(n11047) );
  NAND2_X1 U14032 ( .A1(n11375), .A2(n11047), .ZN(n11048) );
  INV_X1 U14033 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11049) );
  NAND2_X2 U14034 ( .A1(n11105), .A2(n11125), .ZN(n11104) );
  INV_X1 U14035 ( .A(n11104), .ZN(n11052) );
  NAND3_X1 U14036 ( .A1(n11050), .A2(n11375), .A3(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n11051) );
  NAND2_X1 U14037 ( .A1(n15043), .A2(n11011), .ZN(n15335) );
  NAND3_X1 U14038 ( .A1(n15043), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n11621), .ZN(n11089) );
  INV_X1 U14039 ( .A(n11053), .ZN(n11078) );
  NOR2_X1 U14040 ( .A1(n13659), .A2(n11046), .ZN(n11054) );
  NAND2_X1 U14041 ( .A1(n11079), .A2(n11054), .ZN(n11056) );
  INV_X1 U14042 ( .A(n11055), .ZN(n11091) );
  NAND2_X1 U14043 ( .A1(n11056), .A2(n11091), .ZN(n19037) );
  NAND2_X1 U14044 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11057) );
  NOR2_X1 U14045 ( .A1(n19037), .A2(n11057), .ZN(n15352) );
  NOR2_X1 U14046 ( .A1(n13659), .A2(n11044), .ZN(n11058) );
  NAND2_X1 U14047 ( .A1(n11064), .A2(n11058), .ZN(n11059) );
  NAND2_X1 U14048 ( .A1(n11059), .A2(n11078), .ZN(n19061) );
  INV_X1 U14049 ( .A(n19061), .ZN(n11061) );
  AND2_X1 U14050 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11060) );
  NAND2_X1 U14051 ( .A1(n11061), .A2(n11060), .ZN(n15331) );
  NOR2_X1 U14052 ( .A1(n13659), .A2(n11062), .ZN(n11063) );
  INV_X1 U14053 ( .A(n11125), .ZN(n11116) );
  AOI21_X1 U14054 ( .B1(n9815), .B2(n11063), .A(n11116), .ZN(n11065) );
  AND2_X1 U14055 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11066) );
  NAND2_X1 U14056 ( .A1(n19072), .A2(n11066), .ZN(n15330) );
  NAND2_X1 U14057 ( .A1(n11068), .A2(n11067), .ZN(n11069) );
  AND2_X1 U14058 ( .A1(n11082), .A2(n11069), .ZN(n19101) );
  AND2_X1 U14059 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11070) );
  NAND2_X1 U14060 ( .A1(n19101), .A2(n11070), .ZN(n15609) );
  INV_X1 U14061 ( .A(n11082), .ZN(n11071) );
  INV_X1 U14062 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U14063 ( .A1(n11071), .A2(n13481), .ZN(n11084) );
  INV_X1 U14064 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11072) );
  NOR2_X1 U14065 ( .A1(n13659), .A2(n11072), .ZN(n11073) );
  NAND2_X1 U14066 ( .A1(n11084), .A2(n11073), .ZN(n11074) );
  NAND2_X1 U14067 ( .A1(n11074), .A2(n9815), .ZN(n19080) );
  NAND2_X1 U14068 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11075) );
  OR2_X1 U14069 ( .A1(n19080), .A2(n11075), .ZN(n15592) );
  NAND4_X1 U14070 ( .A1(n15331), .A2(n15330), .A3(n15609), .A4(n15592), .ZN(
        n11076) );
  NOR2_X1 U14071 ( .A1(n15352), .A2(n11076), .ZN(n11088) );
  NAND2_X1 U14072 ( .A1(n11078), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11077) );
  MUX2_X1 U14073 ( .A(n11078), .B(n11077), .S(n11375), .Z(n11080) );
  AND2_X1 U14074 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11081) );
  NAND2_X1 U14075 ( .A1(n19047), .A2(n11081), .ZN(n15549) );
  NAND2_X1 U14076 ( .A1(n11082), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11083) );
  MUX2_X1 U14077 ( .A(n11083), .B(n11082), .S(n13659), .Z(n11085) );
  NAND2_X1 U14078 ( .A1(n11085), .A2(n11084), .ZN(n19095) );
  INV_X1 U14079 ( .A(n19095), .ZN(n11086) );
  NAND2_X1 U14080 ( .A1(n11086), .A2(n11621), .ZN(n11097) );
  INV_X1 U14081 ( .A(n11097), .ZN(n11087) );
  NAND2_X1 U14082 ( .A1(n11087), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16382) );
  AND4_X1 U14083 ( .A1(n11089), .A2(n11088), .A3(n15549), .A4(n16382), .ZN(
        n11092) );
  NAND2_X1 U14084 ( .A1(n11375), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11090) );
  XNOR2_X1 U14085 ( .A(n11091), .B(n11090), .ZN(n19023) );
  NAND2_X1 U14086 ( .A1(n19023), .A2(n11011), .ZN(n11100) );
  INV_X1 U14087 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15529) );
  AND2_X2 U14088 ( .A1(n11092), .A2(n15334), .ZN(n11093) );
  OR2_X1 U14089 ( .A1(n19037), .A2(n11023), .ZN(n11094) );
  INV_X1 U14090 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15539) );
  NAND2_X1 U14091 ( .A1(n11094), .A2(n15539), .ZN(n15353) );
  OR2_X1 U14092 ( .A1(n19080), .A2(n11023), .ZN(n11095) );
  INV_X1 U14093 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U14094 ( .A1(n11095), .A2(n15601), .ZN(n15593) );
  NAND2_X1 U14095 ( .A1(n19101), .A2(n11621), .ZN(n11096) );
  INV_X1 U14096 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11290) );
  NAND2_X1 U14097 ( .A1(n11096), .A2(n11290), .ZN(n15610) );
  AND3_X1 U14098 ( .A1(n15593), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15610), .ZN(n11098) );
  INV_X1 U14099 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16377) );
  NAND2_X1 U14100 ( .A1(n11097), .A2(n16377), .ZN(n16380) );
  INV_X1 U14101 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15367) );
  OAI21_X1 U14102 ( .B1(n19061), .B2(n11023), .A(n15367), .ZN(n15332) );
  AND4_X1 U14103 ( .A1(n15353), .A2(n11098), .A3(n16380), .A4(n15332), .ZN(
        n11102) );
  NAND2_X1 U14104 ( .A1(n19072), .A2(n11011), .ZN(n11099) );
  XNOR2_X1 U14105 ( .A(n11099), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15329) );
  NAND2_X1 U14106 ( .A1(n11100), .A2(n15529), .ZN(n15333) );
  NAND2_X1 U14107 ( .A1(n19047), .A2(n11011), .ZN(n11101) );
  INV_X1 U14108 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15553) );
  NAND2_X1 U14109 ( .A1(n11101), .A2(n15553), .ZN(n15550) );
  NAND2_X1 U14110 ( .A1(n11375), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11103) );
  NAND3_X1 U14111 ( .A1(n11105), .A2(n11375), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n11106) );
  NAND2_X1 U14112 ( .A1(n11114), .A2(n11106), .ZN(n15873) );
  INV_X1 U14113 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15487) );
  NAND2_X1 U14114 ( .A1(n11107), .A2(n15487), .ZN(n15319) );
  INV_X1 U14115 ( .A(n11107), .ZN(n11108) );
  NAND2_X1 U14116 ( .A1(n11108), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15320) );
  INV_X1 U14117 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11109) );
  NOR2_X1 U14118 ( .A1(n13659), .A2(n11109), .ZN(n11113) );
  INV_X1 U14119 ( .A(n11113), .ZN(n11110) );
  XNOR2_X1 U14120 ( .A(n11114), .B(n11110), .ZN(n16331) );
  NAND2_X1 U14121 ( .A1(n16331), .A2(n11011), .ZN(n11111) );
  XNOR2_X1 U14122 ( .A(n11111), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15492) );
  INV_X1 U14123 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15486) );
  OR2_X1 U14124 ( .A1(n11111), .A2(n15486), .ZN(n11112) );
  INV_X1 U14125 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11115) );
  NOR2_X1 U14126 ( .A1(n13659), .A2(n11115), .ZN(n11117) );
  AOI21_X1 U14127 ( .B1(n11118), .B2(n11117), .A(n11116), .ZN(n11119) );
  NAND2_X1 U14128 ( .A1(n10018), .A2(n11119), .ZN(n16322) );
  INV_X1 U14129 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15474) );
  NOR2_X1 U14130 ( .A1(n11120), .A2(n15474), .ZN(n15306) );
  NAND2_X1 U14131 ( .A1(n11120), .A2(n15474), .ZN(n15305) );
  INV_X1 U14132 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15114) );
  NAND2_X1 U14133 ( .A1(n11375), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11122) );
  OR2_X1 U14134 ( .A1(n11129), .A2(n11122), .ZN(n11123) );
  INV_X1 U14135 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15009) );
  NAND2_X1 U14136 ( .A1(n11129), .A2(n15009), .ZN(n11642) );
  NAND2_X1 U14137 ( .A1(n11123), .A2(n11620), .ZN(n15017) );
  INV_X1 U14138 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15452) );
  OAI21_X1 U14139 ( .B1(n15017), .B2(n11023), .A(n15452), .ZN(n11124) );
  NAND2_X1 U14140 ( .A1(n11375), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11126) );
  OAI21_X1 U14141 ( .B1(n11127), .B2(n11126), .A(n11125), .ZN(n11128) );
  AOI21_X1 U14142 ( .B1(n9819), .B2(n11621), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15296) );
  NAND2_X1 U14143 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11608) );
  NAND2_X1 U14144 ( .A1(n11375), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11131) );
  NAND2_X1 U14145 ( .A1(n11375), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11135) );
  XNOR2_X1 U14146 ( .A(n11644), .B(n11135), .ZN(n16295) );
  AND2_X1 U14147 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14148 ( .A1(n9819), .A2(n11133), .ZN(n15294) );
  INV_X1 U14149 ( .A(n11135), .ZN(n11136) );
  NAND2_X1 U14150 ( .A1(n11375), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U14151 ( .A1(n11137), .A2(n11138), .ZN(n11618) );
  INV_X1 U14152 ( .A(n11137), .ZN(n11140) );
  INV_X1 U14153 ( .A(n11138), .ZN(n11139) );
  NAND2_X1 U14154 ( .A1(n11140), .A2(n11139), .ZN(n11141) );
  NAND2_X1 U14155 ( .A1(n11618), .A2(n11141), .ZN(n14999) );
  OR2_X1 U14156 ( .A1(n14999), .A2(n11023), .ZN(n11142) );
  INV_X1 U14157 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15271) );
  NAND2_X1 U14158 ( .A1(n11142), .A2(n15271), .ZN(n15267) );
  NAND2_X1 U14159 ( .A1(n15268), .A2(n15267), .ZN(n11617) );
  NAND2_X1 U14160 ( .A1(n11621), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U14161 ( .A1(n11617), .A2(n15266), .ZN(n11147) );
  NAND2_X1 U14162 ( .A1(n11375), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11144) );
  XNOR2_X1 U14163 ( .A(n11618), .B(n11144), .ZN(n16284) );
  AOI21_X1 U14164 ( .B1(n16284), .B2(n11621), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11616) );
  INV_X1 U14165 ( .A(n16284), .ZN(n11145) );
  INV_X1 U14166 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14370) );
  NOR2_X1 U14167 ( .A1(n11616), .A2(n9822), .ZN(n11146) );
  XNOR2_X1 U14168 ( .A(n11147), .B(n11146), .ZN(n15265) );
  NAND2_X1 U14169 ( .A1(n11149), .A2(n11148), .ZN(n11184) );
  INV_X1 U14170 ( .A(n11150), .ZN(n11174) );
  XNOR2_X1 U14171 ( .A(n11174), .B(n11151), .ZN(n11168) );
  NAND2_X1 U14172 ( .A1(n11177), .A2(n11168), .ZN(n11152) );
  OR2_X1 U14173 ( .A1(n11184), .A2(n11152), .ZN(n11157) );
  INV_X1 U14174 ( .A(n11153), .ZN(n11156) );
  INV_X1 U14175 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12760) );
  NAND2_X1 U14176 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12760), .ZN(
        n11155) );
  NAND2_X1 U14177 ( .A1(n11157), .A2(n11186), .ZN(n13604) );
  NAND2_X1 U14178 ( .A1(n11177), .A2(n11158), .ZN(n11159) );
  NOR2_X1 U14179 ( .A1(n11184), .A2(n11159), .ZN(n11160) );
  OAI21_X1 U14180 ( .B1(n13604), .B2(n11160), .A(n19950), .ZN(n11163) );
  NAND2_X1 U14181 ( .A1(n11161), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11162) );
  NAND2_X1 U14182 ( .A1(n11162), .A2(n12760), .ZN(n12756) );
  INV_X1 U14183 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19001) );
  OAI211_X1 U14184 ( .C1(n10849), .C2(n12756), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n19001), .ZN(n20061) );
  NAND2_X1 U14185 ( .A1(n11163), .A2(n20061), .ZN(n13636) );
  INV_X1 U14186 ( .A(n13636), .ZN(n15936) );
  OAI21_X1 U14187 ( .B1(n11164), .B2(n11174), .A(n11179), .ZN(n11165) );
  INV_X1 U14188 ( .A(n11184), .ZN(n11182) );
  INV_X1 U14189 ( .A(n11186), .ZN(n11189) );
  AOI21_X1 U14190 ( .B1(n11165), .B2(n11182), .A(n11189), .ZN(n11166) );
  MUX2_X1 U14191 ( .A(n15936), .B(n11166), .S(n11377), .Z(n20069) );
  NAND2_X1 U14192 ( .A1(n20069), .A2(n11212), .ZN(n11210) );
  NOR2_X1 U14193 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20753) );
  AOI211_X1 U14194 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n20753), .ZN(n20082) );
  NAND2_X1 U14195 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20756) );
  NAND2_X1 U14196 ( .A1(n20082), .A2(n20756), .ZN(n13310) );
  INV_X1 U14197 ( .A(n13310), .ZN(n13608) );
  NAND2_X1 U14198 ( .A1(n11563), .A2(n13608), .ZN(n11207) );
  NAND2_X1 U14199 ( .A1(n11377), .A2(n11173), .ZN(n11169) );
  NAND2_X1 U14200 ( .A1(n11169), .A2(n11168), .ZN(n11171) );
  NAND2_X1 U14201 ( .A1(n11377), .A2(n11177), .ZN(n11170) );
  NAND2_X1 U14202 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  NAND2_X1 U14203 ( .A1(n11172), .A2(n13746), .ZN(n11176) );
  OAI21_X1 U14204 ( .B1(n11174), .B2(n11173), .A(n10688), .ZN(n11175) );
  NAND2_X1 U14205 ( .A1(n11176), .A2(n11175), .ZN(n11183) );
  AND2_X1 U14206 ( .A1(n20077), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19311) );
  INV_X1 U14207 ( .A(n11177), .ZN(n11178) );
  OAI21_X1 U14208 ( .B1(n19311), .B2(n11377), .A(n11178), .ZN(n11180) );
  NAND2_X1 U14209 ( .A1(n11180), .A2(n11179), .ZN(n11181) );
  NAND3_X1 U14210 ( .A1(n11183), .A2(n11182), .A3(n11181), .ZN(n11187) );
  NAND2_X1 U14211 ( .A1(n10688), .A2(n11184), .ZN(n11185) );
  NAND3_X1 U14212 ( .A1(n11187), .A2(n11186), .A3(n11185), .ZN(n11188) );
  NAND2_X1 U14213 ( .A1(n11189), .A2(n19311), .ZN(n11190) );
  NAND2_X1 U14214 ( .A1(n13643), .A2(n13331), .ZN(n12751) );
  INV_X1 U14215 ( .A(n11191), .ZN(n11192) );
  OAI211_X1 U14216 ( .C1(n11192), .C2(n20077), .A(n12751), .B(n11565), .ZN(
        n11206) );
  NAND2_X1 U14217 ( .A1(n11193), .A2(n10668), .ZN(n11194) );
  NAND2_X1 U14218 ( .A1(n12758), .A2(n11194), .ZN(n11200) );
  OAI21_X1 U14219 ( .B1(n11195), .B2(n12790), .A(n20081), .ZN(n11562) );
  NAND2_X1 U14220 ( .A1(n11565), .A2(n11377), .ZN(n11576) );
  NAND2_X1 U14221 ( .A1(n11576), .A2(n13746), .ZN(n11196) );
  NAND3_X1 U14222 ( .A1(n11196), .A2(n19421), .A3(n19431), .ZN(n11197) );
  NAND2_X1 U14223 ( .A1(n11197), .A2(n10668), .ZN(n11198) );
  NAND4_X1 U14224 ( .A1(n11200), .A2(n11199), .A3(n11562), .A4(n11198), .ZN(
        n11577) );
  NOR3_X1 U14225 ( .A1(n11201), .A2(n13604), .A3(n13310), .ZN(n11202) );
  OR2_X1 U14226 ( .A1(n11577), .A2(n11202), .ZN(n12747) );
  MUX2_X1 U14227 ( .A(n11201), .B(n10668), .S(n11377), .Z(n11203) );
  NAND2_X1 U14228 ( .A1(n13610), .A2(n20756), .ZN(n12743) );
  NOR2_X1 U14229 ( .A1(n11203), .A2(n12743), .ZN(n11204) );
  NOR2_X1 U14230 ( .A1(n12747), .A2(n11204), .ZN(n11205) );
  OAI211_X1 U14231 ( .C1(n11207), .C2(n12751), .A(n11206), .B(n11205), .ZN(
        n11208) );
  INV_X1 U14232 ( .A(n11208), .ZN(n11209) );
  NAND2_X1 U14233 ( .A1(n11210), .A2(n11209), .ZN(n11211) );
  NOR2_X1 U14234 ( .A1(n19309), .A2(n12754), .ZN(n20073) );
  INV_X1 U14235 ( .A(n20073), .ZN(n13648) );
  INV_X1 U14236 ( .A(n11578), .ZN(n11581) );
  NAND2_X1 U14237 ( .A1(n11212), .A2(n20077), .ZN(n20068) );
  NOR2_X1 U14238 ( .A1(n11581), .A2(n20068), .ZN(n11252) );
  NAND2_X1 U14239 ( .A1(n11252), .A2(n13331), .ZN(n16477) );
  XOR2_X1 U14240 ( .A(n11214), .B(n11213), .Z(n14392) );
  OR2_X1 U14241 ( .A1(n12727), .A2(n13331), .ZN(n11215) );
  NAND2_X1 U14242 ( .A1(n11215), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12729) );
  XOR2_X1 U14243 ( .A(n12727), .B(n11386), .Z(n11216) );
  NOR2_X1 U14244 ( .A1(n12729), .A2(n11216), .ZN(n11217) );
  XNOR2_X1 U14245 ( .A(n12729), .B(n11216), .ZN(n12735) );
  NOR2_X1 U14246 ( .A1(n20922), .A2(n12735), .ZN(n12734) );
  NOR2_X1 U14247 ( .A1(n11217), .A2(n12734), .ZN(n11218) );
  XOR2_X1 U14248 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11218), .Z(
        n14391) );
  NOR2_X1 U14249 ( .A1(n14392), .A2(n14391), .ZN(n14390) );
  NOR2_X1 U14250 ( .A1(n11218), .A2(n19408), .ZN(n11219) );
  OR2_X1 U14251 ( .A1(n14390), .A2(n11219), .ZN(n11220) );
  XNOR2_X1 U14252 ( .A(n11220), .B(n13269), .ZN(n13279) );
  NAND2_X1 U14253 ( .A1(n11220), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11221) );
  NAND2_X1 U14254 ( .A1(n11222), .A2(n11223), .ZN(n11224) );
  NAND2_X1 U14255 ( .A1(n11225), .A2(n11224), .ZN(n13374) );
  NAND2_X1 U14256 ( .A1(n11226), .A2(n13374), .ZN(n11229) );
  NAND2_X1 U14257 ( .A1(n11227), .A2(n21003), .ZN(n11228) );
  NAND2_X1 U14258 ( .A1(n11230), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13769) );
  NAND2_X1 U14259 ( .A1(n13768), .A2(n13769), .ZN(n11235) );
  INV_X1 U14260 ( .A(n11240), .ZN(n11231) );
  AOI21_X1 U14261 ( .B1(n11233), .B2(n11236), .A(n11232), .ZN(n11234) );
  OAI21_X1 U14262 ( .B1(n11235), .B2(n11236), .A(n11234), .ZN(n15401) );
  NAND2_X1 U14263 ( .A1(n15401), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11239) );
  INV_X1 U14264 ( .A(n11236), .ZN(n11237) );
  XNOR2_X1 U14265 ( .A(n11246), .B(n11023), .ZN(n11243) );
  XNOR2_X2 U14266 ( .A(n11242), .B(n11243), .ZN(n15393) );
  INV_X1 U14267 ( .A(n11243), .ZN(n11244) );
  INV_X1 U14268 ( .A(n11246), .ZN(n11248) );
  NAND2_X1 U14269 ( .A1(n11248), .A2(n11621), .ZN(n11247) );
  AND2_X1 U14270 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16450) );
  NAND2_X1 U14271 ( .A1(n16450), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15598) );
  NAND2_X1 U14272 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15574) );
  NOR2_X1 U14273 ( .A1(n15574), .A2(n15367), .ZN(n11249) );
  NAND2_X1 U14274 ( .A1(n9808), .A2(n11249), .ZN(n15528) );
  AND2_X1 U14275 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15316) );
  AND2_X1 U14276 ( .A1(n15316), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15473) );
  NAND2_X1 U14277 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15446) );
  INV_X1 U14278 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15437) );
  OR2_X1 U14279 ( .A1(n9764), .A2(n11253), .ZN(n11257) );
  AOI22_X1 U14280 ( .A1(n11627), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11255) );
  NAND2_X1 U14281 ( .A1(n11357), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11254) );
  AND2_X1 U14282 ( .A1(n11255), .A2(n11254), .ZN(n11256) );
  NAND2_X1 U14283 ( .A1(n11257), .A2(n11256), .ZN(n12969) );
  INV_X1 U14284 ( .A(n11258), .ZN(n11262) );
  INV_X1 U14285 ( .A(n9764), .ZN(n11352) );
  AOI22_X1 U14286 ( .A1(n10720), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11264) );
  OAI21_X1 U14287 ( .B1(n11263), .B2(n14377), .A(n11264), .ZN(n11265) );
  AOI21_X1 U14288 ( .B1(n10719), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11265), .ZN(n13378) );
  OR2_X1 U14289 ( .A1(n11630), .A2(n13785), .ZN(n11267) );
  AOI22_X1 U14290 ( .A1(n10720), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11266) );
  OAI211_X1 U14291 ( .C1(n11263), .C2(n19198), .A(n11267), .B(n11266), .ZN(
        n13778) );
  INV_X1 U14292 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U14293 ( .A1(n11627), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11268) );
  OAI21_X1 U14294 ( .B1(n11263), .B2(n12989), .A(n11268), .ZN(n11269) );
  AOI21_X1 U14295 ( .B1(n10719), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11269), .ZN(n12986) );
  NAND2_X1 U14296 ( .A1(n12969), .A2(n12985), .ZN(n13055) );
  OR2_X1 U14297 ( .A1(n9764), .A2(n20987), .ZN(n11273) );
  AOI22_X1 U14298 ( .A1(n11627), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14299 ( .A1(n11357), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11270) );
  AND2_X1 U14300 ( .A1(n11271), .A2(n11270), .ZN(n11272) );
  INV_X1 U14301 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15667) );
  OR2_X1 U14302 ( .A1(n9764), .A2(n15667), .ZN(n11277) );
  AOI22_X1 U14303 ( .A1(n11627), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11275) );
  NAND2_X1 U14304 ( .A1(n11357), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11274) );
  AND2_X1 U14305 ( .A1(n11275), .A2(n11274), .ZN(n11276) );
  NAND2_X1 U14306 ( .A1(n11277), .A2(n11276), .ZN(n13061) );
  NAND2_X1 U14307 ( .A1(n13062), .A2(n13061), .ZN(n13060) );
  OR2_X1 U14308 ( .A1(n9764), .A2(n15657), .ZN(n11282) );
  AOI22_X1 U14309 ( .A1(n11627), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11280) );
  NAND2_X1 U14310 ( .A1(n11357), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11279) );
  AND2_X1 U14311 ( .A1(n11280), .A2(n11279), .ZN(n11281) );
  NAND2_X1 U14312 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11284) );
  NAND2_X1 U14313 ( .A1(n11627), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11283) );
  OAI211_X1 U14314 ( .C1(n11263), .C2(n19113), .A(n11284), .B(n11283), .ZN(
        n11285) );
  AOI21_X1 U14315 ( .B1(n11352), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11285), .ZN(n13162) );
  INV_X1 U14316 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20891) );
  OR2_X1 U14317 ( .A1(n9764), .A2(n20891), .ZN(n11289) );
  AOI22_X1 U14318 ( .A1(n11627), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11287) );
  NAND2_X1 U14319 ( .A1(n11357), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11286) );
  AND2_X1 U14320 ( .A1(n11287), .A2(n11286), .ZN(n11288) );
  OR2_X1 U14321 ( .A1(n9764), .A2(n11290), .ZN(n11292) );
  AOI22_X1 U14322 ( .A1(n11627), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11291) );
  OAI211_X1 U14323 ( .C1(n11293), .C2(n11263), .A(n11292), .B(n11291), .ZN(
        n13420) );
  OR2_X1 U14324 ( .A1(n9764), .A2(n16377), .ZN(n11297) );
  AOI22_X1 U14325 ( .A1(n11627), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11295) );
  NAND2_X1 U14326 ( .A1(n11357), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11294) );
  AND2_X1 U14327 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  NAND2_X1 U14328 ( .A1(n11297), .A2(n11296), .ZN(n13477) );
  OR2_X1 U14329 ( .A1(n9764), .A2(n15601), .ZN(n11301) );
  AOI22_X1 U14330 ( .A1(n11627), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11299) );
  NAND2_X1 U14331 ( .A1(n11357), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11298) );
  AND2_X1 U14332 ( .A1(n11299), .A2(n11298), .ZN(n11300) );
  INV_X1 U14333 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15589) );
  OR2_X1 U14334 ( .A1(n9764), .A2(n15589), .ZN(n11305) );
  AOI22_X1 U14335 ( .A1(n11627), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11303) );
  NAND2_X1 U14336 ( .A1(n11357), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11302) );
  AND2_X1 U14337 ( .A1(n11303), .A2(n11302), .ZN(n11304) );
  OR2_X1 U14338 ( .A1(n9764), .A2(n15367), .ZN(n11309) );
  AOI22_X1 U14339 ( .A1(n11627), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11307) );
  NAND2_X1 U14340 ( .A1(n11357), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11306) );
  AND2_X1 U14341 ( .A1(n11307), .A2(n11306), .ZN(n11308) );
  OR2_X1 U14342 ( .A1(n9764), .A2(n15553), .ZN(n11313) );
  AOI22_X1 U14343 ( .A1(n11627), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11311) );
  NAND2_X1 U14344 ( .A1(n11357), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11310) );
  AND2_X1 U14345 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  NAND2_X1 U14346 ( .A1(n11313), .A2(n11312), .ZN(n15167) );
  OR2_X1 U14347 ( .A1(n9764), .A2(n15539), .ZN(n11317) );
  AOI22_X1 U14348 ( .A1(n11627), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11315) );
  NAND2_X1 U14349 ( .A1(n11357), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11314) );
  AND2_X1 U14350 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  OR2_X1 U14351 ( .A1(n9764), .A2(n15529), .ZN(n11321) );
  AOI22_X1 U14352 ( .A1(n11627), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11319) );
  NAND2_X1 U14353 ( .A1(n11357), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11318) );
  AND2_X1 U14354 ( .A1(n11319), .A2(n11318), .ZN(n11320) );
  INV_X1 U14355 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15514) );
  OR2_X1 U14356 ( .A1(n9764), .A2(n15514), .ZN(n11325) );
  AOI22_X1 U14357 ( .A1(n11627), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11323) );
  NAND2_X1 U14358 ( .A1(n11357), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11322) );
  AND2_X1 U14359 ( .A1(n11323), .A2(n11322), .ZN(n11324) );
  NAND2_X1 U14360 ( .A1(n11325), .A2(n11324), .ZN(n15040) );
  OR2_X1 U14361 ( .A1(n9764), .A2(n15487), .ZN(n11329) );
  AOI22_X1 U14362 ( .A1(n11627), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11327) );
  NAND2_X1 U14363 ( .A1(n11357), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11326) );
  AND2_X1 U14364 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  OR2_X1 U14365 ( .A1(n9764), .A2(n15486), .ZN(n11333) );
  AOI22_X1 U14366 ( .A1(n11627), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11331) );
  NAND2_X1 U14367 ( .A1(n11357), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11330) );
  AND2_X1 U14368 ( .A1(n11331), .A2(n11330), .ZN(n11332) );
  OR2_X1 U14369 ( .A1(n9764), .A2(n15474), .ZN(n11337) );
  AOI22_X1 U14370 ( .A1(n11627), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11335) );
  NAND2_X1 U14371 ( .A1(n11357), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11334) );
  AND2_X1 U14372 ( .A1(n11335), .A2(n11334), .ZN(n11336) );
  NAND2_X1 U14373 ( .A1(n11337), .A2(n11336), .ZN(n15120) );
  INV_X1 U14374 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15463) );
  OR2_X1 U14375 ( .A1(n9764), .A2(n15463), .ZN(n11341) );
  AOI22_X1 U14376 ( .A1(n11627), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11339) );
  NAND2_X1 U14377 ( .A1(n11357), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11338) );
  AND2_X1 U14378 ( .A1(n11339), .A2(n11338), .ZN(n11340) );
  NAND2_X1 U14379 ( .A1(n11341), .A2(n11340), .ZN(n15021) );
  NAND2_X1 U14380 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11343) );
  NAND2_X1 U14381 ( .A1(n11627), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11342) );
  OAI211_X1 U14382 ( .C1(n11263), .C2(n15009), .A(n11343), .B(n11342), .ZN(
        n11344) );
  AOI21_X1 U14383 ( .B1(n11352), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11344), .ZN(n15005) );
  INV_X1 U14384 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16307) );
  NAND2_X1 U14385 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11346) );
  NAND2_X1 U14386 ( .A1(n11627), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11345) );
  OAI211_X1 U14387 ( .C1(n11263), .C2(n16307), .A(n11346), .B(n11345), .ZN(
        n11347) );
  AOI21_X1 U14388 ( .B1(n11352), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11347), .ZN(n15099) );
  INV_X1 U14389 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11350) );
  NAND2_X1 U14390 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U14391 ( .A1(n11627), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11348) );
  OAI211_X1 U14392 ( .C1(n11263), .C2(n11350), .A(n11349), .B(n11348), .ZN(
        n11351) );
  AOI21_X1 U14393 ( .B1(n11352), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11351), .ZN(n11654) );
  OR2_X1 U14394 ( .A1(n9764), .A2(n15271), .ZN(n11356) );
  AOI22_X1 U14395 ( .A1(n11627), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11354) );
  NAND2_X1 U14396 ( .A1(n11357), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11353) );
  AND2_X1 U14397 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  NAND2_X1 U14398 ( .A1(n11356), .A2(n11355), .ZN(n14968) );
  OR2_X1 U14399 ( .A1(n9764), .A2(n14370), .ZN(n11361) );
  AOI22_X1 U14400 ( .A1(n11627), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11359) );
  NAND2_X1 U14401 ( .A1(n11357), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11358) );
  AND2_X1 U14402 ( .A1(n11359), .A2(n11358), .ZN(n11360) );
  XNOR2_X1 U14403 ( .A(n14970), .B(n10224), .ZN(n16287) );
  NAND2_X1 U14404 ( .A1(n13620), .A2(n11377), .ZN(n11362) );
  NAND2_X1 U14405 ( .A1(n11362), .A2(n10697), .ZN(n11363) );
  NAND2_X1 U14406 ( .A1(n11364), .A2(n11365), .ZN(n13581) );
  NAND2_X1 U14407 ( .A1(n11366), .A2(n13331), .ZN(n11367) );
  NAND2_X1 U14408 ( .A1(n13581), .A2(n11367), .ZN(n11368) );
  INV_X1 U14409 ( .A(n11520), .ZN(n11508) );
  OR2_X1 U14410 ( .A1(n12727), .A2(n11508), .ZN(n11374) );
  INV_X1 U14411 ( .A(n11385), .ZN(n12788) );
  NAND2_X1 U14412 ( .A1(n11380), .A2(n12788), .ZN(n11392) );
  INV_X1 U14413 ( .A(n11384), .ZN(n11371) );
  NAND2_X1 U14414 ( .A1(n21022), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20057) );
  NAND2_X1 U14415 ( .A1(n11371), .A2(n20057), .ZN(n11372) );
  AND2_X1 U14416 ( .A1(n11392), .A2(n11372), .ZN(n11373) );
  INV_X1 U14417 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20901) );
  NAND2_X1 U14418 ( .A1(n12790), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11376) );
  OAI211_X1 U14419 ( .C1(n11377), .C2(n20916), .A(n11376), .B(n20037), .ZN(
        n11378) );
  INV_X1 U14420 ( .A(n11378), .ZN(n11379) );
  OAI21_X1 U14421 ( .B1(n14361), .B2(n20901), .A(n11379), .ZN(n12782) );
  INV_X1 U14422 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19970) );
  INV_X2 U14423 ( .A(n11534), .ZN(n11525) );
  NAND2_X1 U14424 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11382) );
  NOR2_X1 U14425 ( .A1(n19431), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U14426 ( .A1(n11397), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n11381) );
  OAI211_X1 U14427 ( .C1(n14361), .C2(n19970), .A(n11382), .B(n11381), .ZN(
        n11389) );
  INV_X1 U14428 ( .A(n11389), .ZN(n11383) );
  AOI22_X1 U14429 ( .A1(n11385), .A2(n11384), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U14430 ( .A1(n11520), .A2(n11386), .ZN(n11387) );
  NAND2_X1 U14431 ( .A1(n12813), .A2(n12812), .ZN(n11393) );
  NAND2_X1 U14432 ( .A1(n11520), .A2(n11390), .ZN(n11391) );
  OAI211_X1 U14433 ( .C1(n20037), .C2(n20047), .A(n11392), .B(n11391), .ZN(
        n11394) );
  AND3_X1 U14434 ( .A1(n11393), .A2(n11395), .A3(n11394), .ZN(n11396) );
  INV_X1 U14435 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19973) );
  NAND2_X1 U14436 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11399) );
  INV_X2 U14437 ( .A(n11535), .ZN(n11554) );
  NAND2_X1 U14438 ( .A1(n11554), .A2(P2_EAX_REG_2__SCAN_IN), .ZN(n11398) );
  OAI211_X1 U14439 ( .C1(n14361), .C2(n19973), .A(n11399), .B(n11398), .ZN(
        n12927) );
  AOI22_X1 U14440 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11402) );
  OAI211_X1 U14441 ( .C1(n19975), .C2(n14361), .A(n11402), .B(n11401), .ZN(
        n13181) );
  AOI22_X1 U14442 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11406) );
  NAND2_X1 U14443 ( .A1(n11555), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U14444 ( .A1(n11520), .A2(n11403), .ZN(n11404) );
  AOI22_X1 U14445 ( .A1(n11555), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11554), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14446 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n11520), .B2(n11407), .ZN(n11408) );
  NAND2_X1 U14447 ( .A1(n11409), .A2(n11408), .ZN(n13775) );
  NAND2_X1 U14448 ( .A1(n13776), .A2(n13775), .ZN(n13774) );
  INV_X1 U14449 ( .A(n11410), .ZN(n11411) );
  NAND2_X1 U14450 ( .A1(n11520), .A2(n11411), .ZN(n11412) );
  INV_X1 U14451 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19980) );
  NAND2_X1 U14452 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11414) );
  NAND2_X1 U14453 ( .A1(n11554), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n11413) );
  OAI211_X1 U14454 ( .C1(n14361), .C2(n19980), .A(n11414), .B(n11413), .ZN(
        n15693) );
  NAND2_X1 U14455 ( .A1(n15694), .A2(n15693), .ZN(n11416) );
  NAND2_X1 U14456 ( .A1(n11520), .A2(n11621), .ZN(n11415) );
  INV_X1 U14457 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19982) );
  NAND2_X1 U14458 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11418) );
  NAND2_X1 U14459 ( .A1(n11554), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n11417) );
  OAI211_X1 U14460 ( .C1(n14361), .C2(n19982), .A(n11418), .B(n11417), .ZN(
        n15685) );
  AOI22_X1 U14461 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n11433) );
  NAND2_X1 U14462 ( .A1(n11555), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14463 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n10850), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14464 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n10833), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14465 ( .A1(n10832), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14466 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11421) );
  NAND4_X1 U14467 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11430) );
  AOI22_X1 U14468 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14469 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14470 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10840), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14471 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12447), .B1(
        n10825), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11425) );
  NAND4_X1 U14472 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11429) );
  NAND2_X1 U14473 ( .A1(n11520), .A2(n10226), .ZN(n11431) );
  AOI22_X1 U14474 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14475 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14476 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14477 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11434) );
  NAND4_X1 U14478 ( .A1(n11437), .A2(n11436), .A3(n11435), .A4(n11434), .ZN(
        n11443) );
  AOI22_X1 U14479 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14480 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14481 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14482 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U14483 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11442) );
  AOI22_X1 U14484 ( .A1(n11555), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n11520), 
        .B2(n13117), .ZN(n11445) );
  AOI22_X1 U14485 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U14486 ( .A1(n11445), .A2(n11444), .ZN(n15674) );
  AOI22_X1 U14487 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10849), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14488 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14489 ( .A1(n10832), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14490 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11446) );
  NAND4_X1 U14491 ( .A1(n11449), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11455) );
  AOI22_X1 U14492 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14493 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14494 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10840), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14495 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12447), .B1(
        n10825), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11450) );
  NAND4_X1 U14496 ( .A1(n11453), .A2(n11452), .A3(n11451), .A4(n11450), .ZN(
        n11454) );
  INV_X1 U14497 ( .A(n12347), .ZN(n13118) );
  AOI22_X1 U14498 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11456) );
  OAI21_X1 U14499 ( .B1(n13118), .B2(n11508), .A(n11456), .ZN(n11457) );
  AOI21_X1 U14500 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n11555), .A(n11457), 
        .ZN(n15660) );
  AOI22_X1 U14501 ( .A1(n11555), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11554), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14502 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14503 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14504 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14505 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11458) );
  NAND4_X1 U14506 ( .A1(n11461), .A2(n11460), .A3(n11459), .A4(n11458), .ZN(
        n11467) );
  AOI22_X1 U14507 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14508 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14509 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14510 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11462) );
  NAND4_X1 U14511 ( .A1(n11465), .A2(n11464), .A3(n11463), .A4(n11462), .ZN(
        n11466) );
  AOI22_X1 U14512 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n11525), .B1(
        n11520), .B2(n13199), .ZN(n11468) );
  NAND2_X1 U14513 ( .A1(n11469), .A2(n11468), .ZN(n15647) );
  AOI22_X1 U14514 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14515 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14516 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14517 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11470) );
  NAND4_X1 U14518 ( .A1(n11473), .A2(n11472), .A3(n11471), .A4(n11470), .ZN(
        n11479) );
  AOI22_X1 U14519 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14520 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14521 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14522 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11474) );
  NAND4_X1 U14523 ( .A1(n11477), .A2(n11476), .A3(n11475), .A4(n11474), .ZN(
        n11478) );
  AOI22_X1 U14524 ( .A1(n11555), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11520), 
        .B2(n12350), .ZN(n11481) );
  AOI22_X1 U14525 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11480) );
  NAND2_X1 U14526 ( .A1(n11481), .A2(n11480), .ZN(n15613) );
  INV_X1 U14527 ( .A(n15613), .ZN(n11495) );
  AOI22_X1 U14528 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U14529 ( .A1(n11555), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14530 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14531 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14532 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14533 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11420), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14534 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11491) );
  AOI22_X1 U14535 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14536 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10863), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14537 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10840), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14538 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12447), .B1(
        n10825), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14539 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  NAND2_X1 U14540 ( .A1(n11520), .A2(n13201), .ZN(n11492) );
  AOI22_X1 U14541 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10832), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14542 ( .A1(n10849), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14543 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10833), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14544 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11497) );
  NAND4_X1 U14545 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11506) );
  AOI22_X1 U14546 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14547 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14548 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10840), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14549 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12447), .B1(
        n10825), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11501) );
  NAND4_X1 U14550 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  NOR2_X1 U14551 ( .A1(n11506), .A2(n11505), .ZN(n13473) );
  AOI22_X1 U14552 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11507) );
  OAI21_X1 U14553 ( .B1(n13473), .B2(n11508), .A(n11507), .ZN(n11509) );
  AOI21_X1 U14554 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n11555), .A(n11509), 
        .ZN(n16448) );
  AOI22_X1 U14555 ( .A1(n11555), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11554), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14556 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14557 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14558 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14559 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11510) );
  NAND4_X1 U14560 ( .A1(n11513), .A2(n11512), .A3(n11511), .A4(n11510), .ZN(
        n11519) );
  AOI22_X1 U14561 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14562 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14563 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14564 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11514) );
  NAND4_X1 U14565 ( .A1(n11517), .A2(n11516), .A3(n11515), .A4(n11514), .ZN(
        n11518) );
  NOR2_X1 U14566 ( .A1(n11519), .A2(n11518), .ZN(n13730) );
  AOI22_X1 U14567 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n11380), .B1(
        n11520), .B2(n10187), .ZN(n11521) );
  NAND2_X1 U14568 ( .A1(n11522), .A2(n11521), .ZN(n15597) );
  AOI22_X1 U14569 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14570 ( .A1(n11555), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11523) );
  INV_X1 U14571 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19999) );
  NAND2_X1 U14572 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U14573 ( .A1(n11554), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n11526) );
  OAI211_X1 U14574 ( .C1(n14361), .C2(n19999), .A(n11527), .B(n11526), .ZN(
        n13838) );
  AOI22_X1 U14575 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11529) );
  NAND2_X1 U14576 ( .A1(n11555), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11528) );
  AND2_X1 U14577 ( .A1(n11529), .A2(n11528), .ZN(n15556) );
  AOI22_X1 U14578 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11531) );
  NAND2_X1 U14579 ( .A1(n11555), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11530) );
  AND2_X1 U14580 ( .A1(n11531), .A2(n11530), .ZN(n13886) );
  INV_X1 U14581 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20002) );
  NAND2_X1 U14582 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11533) );
  NAND2_X1 U14583 ( .A1(n11554), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n11532) );
  OAI211_X1 U14584 ( .C1(n14361), .C2(n20002), .A(n11533), .B(n11532), .ZN(
        n15524) );
  AND2_X2 U14585 ( .A1(n15525), .A2(n15524), .ZN(n15034) );
  INV_X1 U14586 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n21000) );
  INV_X1 U14587 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n20873) );
  OAI222_X1 U14588 ( .A1(n14361), .A2(n21000), .B1(n11535), .B2(n20873), .C1(
        n15514), .C2(n11534), .ZN(n15036) );
  AOI22_X1 U14589 ( .A1(n11380), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14590 ( .A1(n11555), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11536) );
  AND2_X1 U14591 ( .A1(n11537), .A2(n11536), .ZN(n15243) );
  INV_X1 U14592 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21070) );
  NAND2_X1 U14593 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11539) );
  NAND2_X1 U14594 ( .A1(n11554), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n11538) );
  OAI211_X1 U14595 ( .C1(n14361), .C2(n21070), .A(n11539), .B(n11538), .ZN(
        n15238) );
  INV_X1 U14596 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U14597 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11541) );
  NAND2_X1 U14598 ( .A1(n11554), .A2(P2_EAX_REG_24__SCAN_IN), .ZN(n11540) );
  OAI211_X1 U14599 ( .C1(n14361), .C2(n11542), .A(n11541), .B(n11540), .ZN(
        n15227) );
  INV_X1 U14600 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20009) );
  NAND2_X1 U14601 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11544) );
  NAND2_X1 U14602 ( .A1(n11554), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n11543) );
  OAI211_X1 U14603 ( .C1(n14361), .C2(n20009), .A(n11544), .B(n11543), .ZN(
        n15026) );
  AOI22_X1 U14604 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11546) );
  NAND2_X1 U14605 ( .A1(n11555), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11545) );
  AND2_X1 U14606 ( .A1(n11546), .A2(n11545), .ZN(n15006) );
  AOI22_X1 U14607 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U14608 ( .A1(n11555), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11547) );
  AND2_X1 U14609 ( .A1(n11548), .A2(n11547), .ZN(n15209) );
  NOR2_X2 U14610 ( .A1(n15210), .A2(n15209), .ZN(n15211) );
  INV_X1 U14611 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U14612 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11550) );
  NAND2_X1 U14613 ( .A1(n11554), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n11549) );
  OAI211_X1 U14614 ( .C1(n14361), .C2(n11551), .A(n11550), .B(n11549), .ZN(
        n15201) );
  INV_X1 U14615 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20015) );
  NAND2_X1 U14616 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11553) );
  NAND2_X1 U14617 ( .A1(n11554), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n11552) );
  OAI211_X1 U14618 ( .C1(n14361), .C2(n20015), .A(n11553), .B(n11552), .ZN(
        n14996) );
  AOI22_X1 U14619 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n11554), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U14620 ( .A1(n11555), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11556) );
  AND2_X1 U14621 ( .A1(n11557), .A2(n11556), .ZN(n11558) );
  NAND2_X1 U14622 ( .A1(n14995), .A2(n11558), .ZN(n11559) );
  NAND2_X1 U14623 ( .A1(n11560), .A2(n11566), .ZN(n11573) );
  NAND2_X1 U14624 ( .A1(n11561), .A2(n13331), .ZN(n13615) );
  NAND2_X1 U14625 ( .A1(n13615), .A2(n11562), .ZN(n11571) );
  NAND2_X1 U14626 ( .A1(n11563), .A2(n20077), .ZN(n11568) );
  INV_X1 U14627 ( .A(n11564), .ZN(n12643) );
  OAI21_X1 U14628 ( .B1(n11566), .B2(n11565), .A(n12643), .ZN(n11567) );
  NAND3_X1 U14629 ( .A1(n11569), .A2(n11568), .A3(n11567), .ZN(n11570) );
  AOI21_X1 U14630 ( .B1(n19421), .B2(n11571), .A(n11570), .ZN(n11572) );
  AND2_X1 U14631 ( .A1(n11573), .A2(n11572), .ZN(n13600) );
  INV_X1 U14632 ( .A(n11574), .ZN(n13583) );
  NAND2_X1 U14633 ( .A1(n13600), .A2(n13583), .ZN(n11575) );
  NAND2_X1 U14634 ( .A1(n11578), .A2(n11575), .ZN(n11579) );
  INV_X1 U14635 ( .A(n16479), .ZN(n15571) );
  NAND2_X1 U14636 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13781) );
  INV_X1 U14637 ( .A(n13781), .ZN(n11582) );
  INV_X1 U14638 ( .A(n11579), .ZN(n19384) );
  NAND2_X1 U14639 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19388) );
  INV_X1 U14640 ( .A(n19388), .ZN(n19393) );
  NAND2_X1 U14641 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19393), .ZN(
        n11584) );
  NAND2_X1 U14642 ( .A1(n19384), .A2(n11584), .ZN(n19390) );
  INV_X1 U14643 ( .A(n19387), .ZN(n11580) );
  NOR2_X1 U14644 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19393), .ZN(
        n11583) );
  NAND2_X1 U14645 ( .A1(n11580), .A2(n11583), .ZN(n19398) );
  NOR2_X1 U14646 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15718) );
  NOR2_X1 U14647 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15935) );
  AND2_X1 U14648 ( .A1(n15718), .A2(n15935), .ZN(n11600) );
  INV_X1 U14649 ( .A(n11600), .ZN(n15581) );
  NAND2_X1 U14650 ( .A1(n11581), .A2(n15581), .ZN(n19385) );
  AND3_X1 U14651 ( .A1(n19390), .A2(n19398), .A3(n19385), .ZN(n13274) );
  OAI21_X1 U14652 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15571), .A(
        n13274), .ZN(n13387) );
  INV_X1 U14653 ( .A(n13387), .ZN(n13784) );
  OAI21_X1 U14654 ( .B1(n15571), .B2(n11582), .A(n13784), .ZN(n15695) );
  AOI21_X1 U14655 ( .B1(n19387), .B2(n11584), .A(n11583), .ZN(n11585) );
  NAND2_X1 U14656 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13273), .ZN(
        n13782) );
  NOR2_X1 U14657 ( .A1(n11603), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15699) );
  NOR2_X1 U14658 ( .A1(n15695), .A2(n15699), .ZN(n11586) );
  INV_X1 U14659 ( .A(n11586), .ZN(n16464) );
  NAND2_X1 U14660 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11606) );
  INV_X1 U14661 ( .A(n11606), .ZN(n11592) );
  NAND2_X1 U14662 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16468) );
  NAND2_X1 U14663 ( .A1(n16479), .A2(n16468), .ZN(n11588) );
  AND2_X1 U14664 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n11586), .ZN(
        n11587) );
  NAND2_X1 U14665 ( .A1(n11588), .A2(n11587), .ZN(n15676) );
  NOR2_X1 U14666 ( .A1(n15657), .A2(n15638), .ZN(n15645) );
  INV_X1 U14667 ( .A(n15645), .ZN(n11589) );
  OR2_X1 U14668 ( .A1(n15676), .A2(n11589), .ZN(n11590) );
  NAND2_X1 U14669 ( .A1(n11590), .A2(n15646), .ZN(n15630) );
  NAND2_X1 U14670 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15630), .ZN(
        n15527) );
  INV_X1 U14671 ( .A(n15527), .ZN(n11591) );
  NAND2_X1 U14672 ( .A1(n11592), .A2(n11591), .ZN(n11593) );
  OR2_X1 U14673 ( .A1(n15528), .A2(n11593), .ZN(n11594) );
  NAND2_X1 U14674 ( .A1(n15646), .A2(n11594), .ZN(n15511) );
  INV_X1 U14675 ( .A(n15473), .ZN(n11595) );
  NAND2_X1 U14676 ( .A1(n15646), .A2(n11595), .ZN(n11596) );
  NAND2_X1 U14677 ( .A1(n15511), .A2(n11596), .ZN(n15479) );
  AND2_X1 U14678 ( .A1(n16479), .A2(n15474), .ZN(n11597) );
  NOR2_X1 U14679 ( .A1(n15479), .A2(n11597), .ZN(n15464) );
  NAND2_X1 U14680 ( .A1(n16479), .A2(n15446), .ZN(n11598) );
  AND2_X1 U14681 ( .A1(n15464), .A2(n11598), .ZN(n15438) );
  OAI21_X1 U14682 ( .B1(n11608), .B2(n15271), .A(n16479), .ZN(n11599) );
  NAND2_X1 U14683 ( .A1(n15438), .A2(n11599), .ZN(n14365) );
  NAND2_X1 U14684 ( .A1(n14365), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14685 ( .A1(n19180), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15261) );
  OAI211_X1 U14686 ( .C1(n19400), .C2(n16285), .A(n11601), .B(n15261), .ZN(
        n11602) );
  AOI21_X1 U14687 ( .B1(n16287), .B2(n16475), .A(n11602), .ZN(n11611) );
  INV_X1 U14688 ( .A(n16468), .ZN(n11605) );
  NAND2_X1 U14689 ( .A1(n16469), .A2(n11605), .ZN(n15675) );
  NOR2_X1 U14690 ( .A1(n15667), .A2(n15675), .ZN(n15644) );
  NAND2_X1 U14691 ( .A1(n15644), .A2(n15645), .ZN(n16452) );
  NOR2_X1 U14692 ( .A1(n15528), .A2(n16452), .ZN(n15562) );
  NAND2_X1 U14693 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15562), .ZN(
        n15543) );
  AND2_X1 U14694 ( .A1(n15473), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11607) );
  NAND2_X1 U14695 ( .A1(n15515), .A2(n11607), .ZN(n15465) );
  INV_X1 U14696 ( .A(n15418), .ZN(n11609) );
  NAND3_X1 U14697 ( .A1(n11609), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14370), .ZN(n11610) );
  OAI211_X1 U14698 ( .C1(n15265), .C2(n16477), .A(n11613), .B(n11612), .ZN(
        P2_U3016) );
  NOR2_X1 U14699 ( .A1(n11618), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11619) );
  MUX2_X1 U14700 ( .A(n11620), .B(n11619), .S(n11375), .Z(n16278) );
  NAND2_X1 U14701 ( .A1(n16278), .A2(n11621), .ZN(n11622) );
  XNOR2_X1 U14702 ( .A(n11622), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11623) );
  INV_X1 U14703 ( .A(n19304), .ZN(n12648) );
  NOR2_X1 U14704 ( .A1(n20068), .A2(n12648), .ZN(n11624) );
  NAND2_X1 U14705 ( .A1(n20069), .A2(n11624), .ZN(n19000) );
  INV_X1 U14706 ( .A(n19000), .ZN(n11625) );
  NAND2_X1 U14707 ( .A1(n11625), .A2(n13331), .ZN(n16425) );
  NAND2_X1 U14708 ( .A1(n14358), .A2(n16435), .ZN(n11641) );
  NAND2_X1 U14709 ( .A1(n11626), .A2(n10224), .ZN(n11632) );
  AOI22_X1 U14710 ( .A1(n11627), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11629) );
  NAND2_X1 U14711 ( .A1(n11357), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11628) );
  OAI211_X1 U14712 ( .C1(n9764), .C2(n9957), .A(n11629), .B(n11628), .ZN(
        n11631) );
  NOR2_X2 U14713 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20029) );
  OR2_X1 U14714 ( .A1(n20029), .A2(n15718), .ZN(n20048) );
  NAND2_X1 U14715 ( .A1(n20048), .A2(n19309), .ZN(n11633) );
  AND2_X1 U14716 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20049) );
  INV_X1 U14717 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11638) );
  INV_X1 U14718 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16362) );
  INV_X1 U14719 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15337) );
  INV_X1 U14720 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15358) );
  INV_X1 U14721 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15369) );
  INV_X1 U14722 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19090) );
  INV_X1 U14723 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15029) );
  INV_X1 U14724 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16306) );
  INV_X1 U14725 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14726 ( .A1(n19309), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12335) );
  INV_X1 U14727 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19770) );
  NAND2_X1 U14728 ( .A1(n19770), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11636) );
  NAND2_X1 U14729 ( .A1(n12335), .A2(n11636), .ZN(n12731) );
  NAND2_X1 U14730 ( .A1(n13313), .A2(n16434), .ZN(n11637) );
  INV_X1 U14731 ( .A(n19210), .ZN(n19180) );
  NAND2_X1 U14732 ( .A1(n19180), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14366) );
  OAI211_X1 U14733 ( .C1(n16445), .C2(n11638), .A(n11637), .B(n14366), .ZN(
        n11639) );
  AOI21_X1 U14734 ( .B1(n16274), .B2(n16421), .A(n11639), .ZN(n11640) );
  OAI211_X1 U14735 ( .C1(n14373), .C2(n16425), .A(n11641), .B(n11640), .ZN(
        P2_U2983) );
  NAND3_X1 U14736 ( .A1(n11375), .A2(n11642), .A3(P2_EBX_REG_27__SCAN_IN), 
        .ZN(n11643) );
  NAND2_X1 U14737 ( .A1(n11644), .A2(n11643), .ZN(n16310) );
  NOR2_X1 U14738 ( .A1(n16310), .A2(n11023), .ZN(n11646) );
  XNOR2_X1 U14739 ( .A(n11649), .B(n10214), .ZN(n11650) );
  XNOR2_X1 U14740 ( .A(n11651), .B(n11650), .ZN(n15423) );
  NAND2_X1 U14741 ( .A1(n15423), .A2(n16441), .ZN(n11665) );
  OAI21_X1 U14742 ( .B1(n11652), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11653), .ZN(n15431) );
  INV_X1 U14743 ( .A(n14969), .ZN(n11656) );
  NAND2_X1 U14744 ( .A1(n15102), .A2(n11654), .ZN(n11655) );
  NAND2_X1 U14745 ( .A1(n11656), .A2(n11655), .ZN(n16297) );
  INV_X1 U14746 ( .A(n16297), .ZN(n11661) );
  INV_X1 U14747 ( .A(n14973), .ZN(n11658) );
  INV_X1 U14748 ( .A(n14992), .ZN(n11657) );
  OAI21_X1 U14749 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11658), .A(
        n11657), .ZN(n16301) );
  NAND2_X1 U14750 ( .A1(n19180), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15424) );
  NAND2_X1 U14751 ( .A1(n16409), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11659) );
  OAI211_X1 U14752 ( .C1(n16301), .C2(n16424), .A(n15424), .B(n11659), .ZN(
        n11660) );
  AOI21_X1 U14753 ( .B1(n11661), .B2(n16421), .A(n11660), .ZN(n11662) );
  NAND2_X1 U14754 ( .A1(n11665), .A2(n11664), .ZN(P2_U2986) );
  NOR2_X4 U14755 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n11667), .ZN(
        n11934) );
  AOI22_X1 U14756 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11670) );
  BUF_X8 U14757 ( .A(n11782), .Z(n14314) );
  AOI22_X1 U14758 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11669) );
  AND2_X4 U14759 ( .A1(n13206), .A2(n11674), .ZN(n11772) );
  AOI22_X1 U14760 ( .A1(n9758), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11668) );
  NAND4_X1 U14761 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(
        n11681) );
  AND2_X2 U14762 ( .A1(n11672), .A2(n11675), .ZN(n11777) );
  AOI22_X1 U14763 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11777), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11679) );
  AND2_X2 U14764 ( .A1(n13217), .A2(n13229), .ZN(n11701) );
  AND2_X2 U14765 ( .A1(n13217), .A2(n13206), .ZN(n14056) );
  AOI22_X1 U14766 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11678) );
  AND2_X2 U14767 ( .A1(n11672), .A2(n11674), .ZN(n11702) );
  AOI22_X1 U14768 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11840), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11677) );
  AND2_X2 U14769 ( .A1(n13229), .A2(n11674), .ZN(n11929) );
  AOI22_X1 U14770 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11676) );
  NAND4_X1 U14771 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11680) );
  OR2_X2 U14772 ( .A1(n11681), .A2(n11680), .ZN(n12863) );
  AOI22_X1 U14773 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11777), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14774 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14775 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11840), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14776 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14777 ( .A1(n9755), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14265), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14778 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14779 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14780 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11777), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14781 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14782 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11840), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14783 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14784 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14785 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14786 ( .A1(n9758), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14787 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11694) );
  AND2_X1 U14788 ( .A1(n11737), .A2(n12129), .ZN(n11700) );
  AOI22_X1 U14789 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14790 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11840), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11707) );
  NAND2_X1 U14791 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U14792 ( .A1(n11703), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11704) );
  AOI22_X1 U14793 ( .A1(n9758), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9749), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14794 ( .A1(n9756), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14265), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14795 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11782), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14796 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U14797 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11720) );
  NAND2_X1 U14798 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11719) );
  NAND2_X1 U14799 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U14800 ( .A1(n14314), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11717) );
  NAND2_X1 U14801 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U14802 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U14803 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11722) );
  NAND2_X1 U14804 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14805 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11728) );
  NAND2_X1 U14806 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14807 ( .A1(n11934), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11726) );
  NAND2_X1 U14808 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U14809 ( .A1(n14056), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U14810 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U14811 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11730) );
  NAND2_X1 U14812 ( .A1(n11703), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U14813 ( .A1(n11857), .A2(n13073), .ZN(n11805) );
  NAND2_X1 U14814 ( .A1(n11805), .A2(n11797), .ZN(n11748) );
  AOI22_X1 U14815 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14816 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14817 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11840), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14818 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11738) );
  NAND4_X1 U14819 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11747) );
  AOI22_X1 U14820 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14821 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14822 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11742) );
  NAND4_X1 U14823 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11746) );
  NAND2_X1 U14824 ( .A1(n9758), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11753) );
  NAND2_X1 U14825 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11752) );
  NAND2_X1 U14826 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11751) );
  INV_X1 U14827 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11749) );
  NAND2_X1 U14828 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U14829 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11757) );
  NAND2_X1 U14830 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11756) );
  NAND2_X1 U14831 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U14832 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U14833 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11762) );
  NAND2_X1 U14834 ( .A1(n11934), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11761) );
  NAND2_X1 U14835 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11760) );
  NAND2_X1 U14836 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11767) );
  NAND2_X1 U14837 ( .A1(n14056), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11766) );
  NAND2_X1 U14838 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11765) );
  NAND2_X1 U14839 ( .A1(n11703), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U14840 ( .A1(n11833), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11776) );
  NAND2_X1 U14841 ( .A1(n11948), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11775) );
  NAND2_X1 U14842 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14843 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U14844 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U14845 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U14846 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U14847 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U14848 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11786) );
  NAND2_X1 U14849 ( .A1(n11759), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U14850 ( .A1(n11934), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U14851 ( .A1(n11782), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U14852 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U14853 ( .A1(n14056), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11789) );
  NAND2_X1 U14854 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11788) );
  NAND2_X1 U14855 ( .A1(n11703), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11787) );
  NAND4_X4 U14856 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n12180) );
  INV_X1 U14857 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20091) );
  XNOR2_X1 U14858 ( .A(n20091), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12090) );
  NOR2_X1 U14859 ( .A1(n12180), .A2(n12090), .ZN(n11798) );
  NOR2_X1 U14860 ( .A1(n12836), .A2(n9765), .ZN(n11795) );
  NOR2_X1 U14861 ( .A1(n12129), .A2(n12180), .ZN(n11796) );
  AND2_X2 U14862 ( .A1(n12836), .A2(n12180), .ZN(n12181) );
  NAND2_X1 U14863 ( .A1(n12863), .A2(n9765), .ZN(n12285) );
  OAI211_X1 U14864 ( .C1(n11818), .C2(n13679), .A(n12959), .B(n12285), .ZN(
        n11823) );
  NOR2_X1 U14865 ( .A1(n11823), .A2(n12160), .ZN(n11807) );
  NAND2_X1 U14866 ( .A1(n13139), .A2(n11737), .ZN(n11801) );
  AND2_X1 U14867 ( .A1(n11801), .A2(n13073), .ZN(n11821) );
  OR2_X1 U14868 ( .A1(n11802), .A2(n11737), .ZN(n11803) );
  NAND2_X1 U14869 ( .A1(n11807), .A2(n11806), .ZN(n11811) );
  NAND2_X1 U14870 ( .A1(n11808), .A2(n11809), .ZN(n11810) );
  AOI22_X1 U14871 ( .A1(n11811), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11810), 
        .B2(n11917), .ZN(n11812) );
  NAND2_X1 U14872 ( .A1(n11876), .A2(n11812), .ZN(n11896) );
  NAND2_X1 U14873 ( .A1(n11896), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11815) );
  INV_X1 U14874 ( .A(n12882), .ZN(n11813) );
  MUX2_X1 U14875 ( .A(n15905), .B(n11813), .S(n20449), .Z(n11814) );
  NAND2_X1 U14876 ( .A1(n11816), .A2(n12179), .ZN(n11817) );
  NOR2_X1 U14877 ( .A1(n9766), .A2(n12180), .ZN(n13438) );
  INV_X1 U14878 ( .A(n13438), .ZN(n14411) );
  MUX2_X1 U14879 ( .A(n11808), .B(n11817), .S(n14411), .Z(n11827) );
  NAND2_X1 U14880 ( .A1(n11819), .A2(n13671), .ZN(n12290) );
  NAND2_X1 U14881 ( .A1(n13449), .A2(n12180), .ZN(n13425) );
  AND3_X1 U14882 ( .A1(n13425), .A2(n14949), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11820) );
  OAI211_X1 U14883 ( .C1(n11821), .C2(n11818), .A(n12290), .B(n11820), .ZN(
        n11822) );
  NOR2_X1 U14884 ( .A1(n11823), .A2(n11822), .ZN(n11825) );
  NAND3_X1 U14885 ( .A1(n12165), .A2(n12180), .A3(n14944), .ZN(n11824) );
  INV_X1 U14886 ( .A(n11982), .ZN(n11854) );
  AOI22_X1 U14887 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14888 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14889 ( .A1(n11934), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14890 ( .A1(n14056), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11829) );
  NAND4_X1 U14891 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n11839) );
  AOI22_X1 U14892 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14221), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14893 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14894 ( .A1(n11833), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14895 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11834) );
  NAND4_X1 U14896 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n11834), .ZN(
        n11838) );
  AOI22_X1 U14897 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14898 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14899 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14900 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11841) );
  NAND4_X1 U14901 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .ZN(
        n11852) );
  AOI22_X1 U14902 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14903 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14105), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14905 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11848) );
  BUF_X1 U14906 ( .A(n11929), .Z(n11846) );
  AOI22_X1 U14907 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U14908 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11851) );
  XNOR2_X1 U14909 ( .A(n11981), .B(n11993), .ZN(n11853) );
  NAND2_X1 U14910 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  INV_X1 U14911 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n21006) );
  AOI21_X1 U14912 ( .B1(n13449), .B2(n11993), .A(n11886), .ZN(n11859) );
  NAND2_X1 U14913 ( .A1(n13679), .A2(n12057), .ZN(n11858) );
  OAI211_X1 U14914 ( .C1(n12116), .C2(n21006), .A(n11859), .B(n11858), .ZN(
        n11990) );
  INV_X1 U14915 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20282) );
  OR2_X1 U14916 ( .A1(n11982), .A2(n12057), .ZN(n11873) );
  AOI22_X1 U14917 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14221), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14918 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14126), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14919 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14920 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11862) );
  NAND4_X1 U14921 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11871) );
  AOI22_X1 U14922 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14923 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14924 ( .A1(n11934), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14925 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U14926 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  NAND2_X1 U14927 ( .A1(n11917), .A2(n11994), .ZN(n11872) );
  OAI211_X1 U14928 ( .C1(n20282), .C2(n12116), .A(n11873), .B(n11872), .ZN(
        n11874) );
  NAND2_X1 U14929 ( .A1(n11896), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11879) );
  INV_X1 U14930 ( .A(n15905), .ZN(n11925) );
  NAND2_X1 U14931 ( .A1(n11925), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11893) );
  NAND2_X1 U14932 ( .A1(n20599), .A2(n20449), .ZN(n20545) );
  NAND2_X1 U14933 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20595) );
  AND2_X1 U14934 ( .A1(n20545), .A2(n20595), .ZN(n20264) );
  NAND2_X1 U14935 ( .A1(n12882), .A2(n20264), .ZN(n11877) );
  AND2_X1 U14936 ( .A1(n11893), .A2(n11877), .ZN(n11878) );
  NAND2_X1 U14937 ( .A1(n11879), .A2(n11878), .ZN(n11880) );
  INV_X1 U14938 ( .A(n11885), .ZN(n11883) );
  NAND2_X1 U14939 ( .A1(n11884), .A2(n11883), .ZN(n13127) );
  NAND2_X1 U14940 ( .A1(n13127), .A2(n11904), .ZN(n13284) );
  INV_X1 U14941 ( .A(n13284), .ZN(n11887) );
  INV_X1 U14942 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n11886) );
  INV_X1 U14943 ( .A(n11994), .ZN(n11888) );
  OR2_X1 U14944 ( .A1(n11982), .A2(n11888), .ZN(n11889) );
  NAND2_X2 U14945 ( .A1(n11890), .A2(n11889), .ZN(n12912) );
  INV_X1 U14946 ( .A(n12003), .ZN(n11920) );
  INV_X1 U14947 ( .A(n11876), .ZN(n11895) );
  NAND2_X1 U14948 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  NAND2_X1 U14949 ( .A1(n11895), .A2(n11894), .ZN(n11902) );
  NAND2_X1 U14950 ( .A1(n11904), .A2(n11902), .ZN(n11900) );
  NOR2_X1 U14951 ( .A1(n15905), .A2(n20272), .ZN(n11898) );
  XNOR2_X1 U14952 ( .A(n20595), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13290) );
  NAND2_X1 U14953 ( .A1(n12882), .A2(n13290), .ZN(n11901) );
  NAND2_X1 U14954 ( .A1(n11903), .A2(n11901), .ZN(n11899) );
  NAND2_X2 U14955 ( .A1(n11900), .A2(n11899), .ZN(n11921) );
  NAND4_X1 U14956 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .ZN(
        n11905) );
  AOI22_X1 U14957 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11777), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14958 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14959 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14960 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11906) );
  NAND4_X1 U14961 ( .A1(n11909), .A2(n11908), .A3(n11907), .A4(n11906), .ZN(
        n11915) );
  AOI22_X1 U14962 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14963 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11934), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U14964 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14965 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11910) );
  NAND4_X1 U14966 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n11914) );
  AOI22_X1 U14967 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11917), .B2(n11916), .ZN(n11918) );
  NAND2_X1 U14968 ( .A1(n11920), .A2(n12002), .ZN(n12013) );
  INV_X1 U14969 ( .A(n12013), .ZN(n11943) );
  NAND2_X1 U14970 ( .A1(n11897), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11927) );
  OAI21_X1 U14971 ( .B1(n20595), .B2(n20272), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11924) );
  INV_X1 U14972 ( .A(n20595), .ZN(n11923) );
  INV_X1 U14973 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20273) );
  NAND2_X1 U14974 ( .A1(n20273), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20419) );
  INV_X1 U14975 ( .A(n20419), .ZN(n11922) );
  NAND2_X1 U14976 ( .A1(n11923), .A2(n11922), .ZN(n13488) );
  NAND2_X1 U14977 ( .A1(n11924), .A2(n13488), .ZN(n20265) );
  AOI22_X1 U14978 ( .A1(n12882), .A2(n20265), .B1(n11925), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11926) );
  XNOR2_X2 U14979 ( .A(n11921), .B(n13343), .ZN(n20271) );
  AOI22_X1 U14980 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14981 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14982 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14983 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11930) );
  NAND4_X1 U14984 ( .A1(n11933), .A2(n11932), .A3(n11931), .A4(n11930), .ZN(
        n11940) );
  AOI22_X1 U14985 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U14986 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11937) );
  INV_X1 U14987 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n21027) );
  AOI22_X1 U14988 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U14989 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11935) );
  NAND4_X1 U14990 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11939) );
  AOI22_X1 U14991 ( .A1(n12131), .A2(n12015), .B1(n12150), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U14992 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U14993 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U14994 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U14995 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14023), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11944) );
  NAND4_X1 U14996 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(
        n11954) );
  AOI22_X1 U14997 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14998 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U14999 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n14283), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15000 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11949) );
  NAND4_X1 U15001 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(
        n11953) );
  NAND2_X1 U15002 ( .A1(n12131), .A2(n12023), .ZN(n11956) );
  NAND2_X1 U15003 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11955) );
  NAND2_X1 U15004 ( .A1(n11956), .A2(n11955), .ZN(n12021) );
  AOI22_X1 U15005 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U15006 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15007 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15008 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11957) );
  NAND4_X1 U15009 ( .A1(n11960), .A2(n11959), .A3(n11958), .A4(n11957), .ZN(
        n11966) );
  AOI22_X1 U15010 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15011 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15012 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15013 ( .A1(n11833), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11961) );
  NAND4_X1 U15014 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n11965) );
  AOI22_X1 U15015 ( .A1(n12131), .A2(n12035), .B1(n12150), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12032) );
  INV_X1 U15016 ( .A(n12044), .ZN(n11980) );
  AOI22_X1 U15017 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15018 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11833), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15019 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15020 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U15021 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11978) );
  AOI22_X1 U15022 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15023 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15024 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15025 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U15026 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11977) );
  AOI22_X1 U15027 ( .A1(n12131), .A2(n12047), .B1(n12150), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12043) );
  INV_X1 U15028 ( .A(n12043), .ZN(n11979) );
  NOR3_X1 U15029 ( .A1(n11982), .A2(n12115), .A3(n11981), .ZN(n11983) );
  INV_X1 U15030 ( .A(n12035), .ZN(n11985) );
  NAND2_X1 U15031 ( .A1(n11994), .A2(n11993), .ZN(n12004) );
  NAND2_X1 U15032 ( .A1(n12004), .A2(n12005), .ZN(n12016) );
  NAND2_X1 U15033 ( .A1(n12016), .A2(n12015), .ZN(n12024) );
  INV_X1 U15034 ( .A(n12023), .ZN(n11984) );
  OR2_X1 U15035 ( .A1(n12024), .A2(n11984), .ZN(n12036) );
  NOR2_X1 U15036 ( .A1(n11985), .A2(n12036), .ZN(n12045) );
  NAND2_X1 U15037 ( .A1(n12045), .A2(n12047), .ZN(n12056) );
  INV_X1 U15038 ( .A(n12056), .ZN(n11986) );
  NAND2_X1 U15039 ( .A1(n12057), .A2(n11986), .ZN(n11987) );
  OR2_X1 U15040 ( .A1(n11818), .A2(n11987), .ZN(n11988) );
  NAND2_X1 U15041 ( .A1(n16090), .A2(n11988), .ZN(n13814) );
  AND2_X1 U15042 ( .A1(n13814), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12063) );
  NAND2_X1 U15043 ( .A1(n13449), .A2(n12836), .ZN(n12006) );
  OAI21_X1 U15044 ( .B1(n11818), .B2(n11993), .A(n12006), .ZN(n11991) );
  INV_X1 U15045 ( .A(n11991), .ZN(n11992) );
  XNOR2_X1 U15046 ( .A(n11994), .B(n11993), .ZN(n11995) );
  OAI211_X1 U15047 ( .C1(n11995), .C2(n11818), .A(n13158), .B(n12129), .ZN(
        n11996) );
  INV_X1 U15048 ( .A(n11996), .ZN(n11997) );
  NAND2_X1 U15049 ( .A1(n12909), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12001) );
  INV_X1 U15050 ( .A(n11998), .ZN(n11999) );
  OR2_X1 U15051 ( .A1(n12854), .A2(n11999), .ZN(n12000) );
  INV_X1 U15052 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13046) );
  NAND2_X1 U15053 ( .A1(n9769), .A2(n12163), .ZN(n12010) );
  OAI21_X1 U15054 ( .B1(n12005), .B2(n12004), .A(n12016), .ZN(n12008) );
  INV_X1 U15055 ( .A(n11818), .ZN(n12059) );
  INV_X1 U15056 ( .A(n12006), .ZN(n12007) );
  AOI21_X1 U15057 ( .B1(n12008), .B2(n12059), .A(n12007), .ZN(n12009) );
  NAND2_X1 U15058 ( .A1(n12010), .A2(n12009), .ZN(n13038) );
  NAND2_X1 U15059 ( .A1(n12011), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12012) );
  INV_X1 U15060 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13239) );
  INV_X1 U15061 ( .A(n13124), .ZN(n13261) );
  NAND2_X1 U15062 ( .A1(n12013), .A2(n13261), .ZN(n12014) );
  XNOR2_X1 U15063 ( .A(n12016), .B(n12015), .ZN(n12017) );
  OAI22_X1 U15064 ( .A1(n20268), .A2(n12115), .B1(n11818), .B2(n12017), .ZN(
        n13079) );
  NAND2_X1 U15065 ( .A1(n12018), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12019) );
  NAND2_X1 U15066 ( .A1(n12020), .A2(n12019), .ZN(n13168) );
  XNOR2_X1 U15067 ( .A(n12022), .B(n12021), .ZN(n13099) );
  NAND2_X1 U15068 ( .A1(n13099), .A2(n12163), .ZN(n12027) );
  XNOR2_X1 U15069 ( .A(n12024), .B(n12023), .ZN(n12025) );
  NAND2_X1 U15070 ( .A1(n12025), .A2(n12059), .ZN(n12026) );
  NAND2_X1 U15071 ( .A1(n12027), .A2(n12026), .ZN(n12029) );
  INV_X1 U15072 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12028) );
  XNOR2_X1 U15073 ( .A(n12029), .B(n12028), .ZN(n13167) );
  NAND2_X1 U15074 ( .A1(n13168), .A2(n13167), .ZN(n12031) );
  NAND2_X1 U15075 ( .A1(n12029), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12030) );
  NAND2_X1 U15076 ( .A1(n12031), .A2(n12030), .ZN(n16113) );
  NAND2_X1 U15077 ( .A1(n12033), .A2(n12032), .ZN(n12034) );
  NAND2_X1 U15078 ( .A1(n13253), .A2(n12163), .ZN(n12039) );
  XNOR2_X1 U15079 ( .A(n12036), .B(n12035), .ZN(n12037) );
  NAND2_X1 U15080 ( .A1(n12037), .A2(n12059), .ZN(n12038) );
  NAND2_X1 U15081 ( .A1(n12039), .A2(n12038), .ZN(n12041) );
  INV_X1 U15082 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12040) );
  XNOR2_X1 U15083 ( .A(n12041), .B(n12040), .ZN(n16112) );
  NAND2_X1 U15084 ( .A1(n12041), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12042) );
  NAND2_X1 U15085 ( .A1(n12044), .A2(n12043), .ZN(n13513) );
  NAND3_X1 U15086 ( .A1(n12055), .A2(n12163), .A3(n13513), .ZN(n12050) );
  INV_X1 U15087 ( .A(n12045), .ZN(n12046) );
  XNOR2_X1 U15088 ( .A(n12047), .B(n12046), .ZN(n12048) );
  NAND2_X1 U15089 ( .A1(n12059), .A2(n12048), .ZN(n12049) );
  NAND2_X1 U15090 ( .A1(n12050), .A2(n12049), .ZN(n12051) );
  OR2_X1 U15091 ( .A1(n12051), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16106) );
  NAND2_X1 U15092 ( .A1(n12051), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16105) );
  INV_X1 U15093 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U15094 ( .A1(n12131), .A2(n12057), .ZN(n12052) );
  OAI21_X1 U15095 ( .B1(n12053), .B2(n12116), .A(n12052), .ZN(n12054) );
  NAND2_X1 U15096 ( .A1(n13515), .A2(n12163), .ZN(n12061) );
  XNOR2_X1 U15097 ( .A(n12057), .B(n12056), .ZN(n12058) );
  NAND2_X1 U15098 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  NAND2_X1 U15099 ( .A1(n12061), .A2(n12060), .ZN(n16098) );
  OR2_X1 U15100 ( .A1(n16098), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12062) );
  INV_X1 U15101 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16228) );
  OR2_X1 U15102 ( .A1(n16090), .A2(n16228), .ZN(n12065) );
  NAND2_X1 U15103 ( .A1(n16090), .A2(n16228), .ZN(n12066) );
  NAND2_X1 U15104 ( .A1(n14833), .A2(n12066), .ZN(n13891) );
  INV_X1 U15105 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16195) );
  OR2_X1 U15106 ( .A1(n16090), .A2(n16195), .ZN(n13892) );
  NAND2_X1 U15107 ( .A1(n16090), .A2(n16195), .ZN(n12067) );
  NAND2_X1 U15108 ( .A1(n13892), .A2(n12067), .ZN(n14826) );
  INV_X1 U15109 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12075) );
  NAND2_X1 U15110 ( .A1(n16090), .A2(n12075), .ZN(n14824) );
  NAND2_X1 U15111 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12068) );
  NAND2_X1 U15112 ( .A1(n16090), .A2(n12068), .ZN(n14822) );
  NAND2_X1 U15113 ( .A1(n14824), .A2(n14822), .ZN(n12069) );
  NOR2_X1 U15114 ( .A1(n14826), .A2(n12069), .ZN(n13894) );
  INV_X1 U15115 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12227) );
  NAND2_X1 U15116 ( .A1(n16090), .A2(n12227), .ZN(n12070) );
  NAND2_X1 U15117 ( .A1(n13894), .A2(n12070), .ZN(n14812) );
  INV_X1 U15118 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12296) );
  XNOR2_X1 U15119 ( .A(n16090), .B(n12296), .ZN(n14814) );
  INV_X1 U15120 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14912) );
  AND2_X1 U15121 ( .A1(n16090), .A2(n14912), .ZN(n16073) );
  INV_X1 U15122 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12078) );
  OR2_X1 U15123 ( .A1(n16090), .A2(n12227), .ZN(n12074) );
  NOR2_X1 U15124 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14820) );
  AND2_X1 U15125 ( .A1(n14820), .A2(n12075), .ZN(n12076) );
  OR2_X1 U15126 ( .A1(n16090), .A2(n12076), .ZN(n16076) );
  OR2_X1 U15127 ( .A1(n16090), .A2(n14912), .ZN(n16074) );
  AND2_X1 U15128 ( .A1(n16076), .A2(n16074), .ZN(n12077) );
  XNOR2_X1 U15129 ( .A(n16090), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14808) );
  NAND3_X1 U15130 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12309) );
  INV_X1 U15131 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16160) );
  INV_X1 U15132 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16164) );
  INV_X1 U15133 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14902) );
  INV_X1 U15134 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15917) );
  AND2_X1 U15135 ( .A1(n14902), .A2(n15917), .ZN(n12079) );
  NAND2_X1 U15136 ( .A1(n12080), .A2(n14894), .ZN(n14801) );
  NAND3_X1 U15137 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12301) );
  NAND2_X1 U15138 ( .A1(n14741), .A2(n12301), .ZN(n12082) );
  NAND2_X1 U15139 ( .A1(n12081), .A2(n16090), .ZN(n14772) );
  NAND3_X1 U15140 ( .A1(n12082), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14772), .ZN(n12086) );
  NAND2_X1 U15141 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14863) );
  INV_X1 U15142 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14856) );
  NOR2_X1 U15143 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12083) );
  INV_X1 U15144 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16136) );
  AND2_X1 U15145 ( .A1(n12083), .A2(n16136), .ZN(n14753) );
  NOR2_X1 U15146 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14864) );
  NAND2_X1 U15147 ( .A1(n14753), .A2(n14864), .ZN(n12084) );
  NOR2_X1 U15148 ( .A1(n14741), .A2(n12084), .ZN(n12085) );
  NAND2_X1 U15149 ( .A1(n12086), .A2(n12085), .ZN(n14733) );
  INV_X1 U15150 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12089) );
  NAND2_X1 U15151 ( .A1(n12090), .A2(n12089), .ZN(n15930) );
  NAND2_X1 U15152 ( .A1(n12180), .A2(n15930), .ZN(n12111) );
  XNOR2_X1 U15153 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12105) );
  NAND2_X1 U15154 ( .A1(n20449), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12122) );
  NAND2_X1 U15155 ( .A1(n12105), .A2(n12104), .ZN(n12092) );
  NAND2_X1 U15156 ( .A1(n20599), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12091) );
  NAND2_X1 U15157 ( .A1(n12092), .A2(n12091), .ZN(n12107) );
  XNOR2_X1 U15158 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12106) );
  NAND2_X1 U15159 ( .A1(n12107), .A2(n12106), .ZN(n12094) );
  NAND2_X1 U15160 ( .A1(n20272), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12093) );
  NAND2_X1 U15161 ( .A1(n12094), .A2(n12093), .ZN(n12101) );
  MUX2_X1 U15162 ( .A(n20273), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12099) );
  NAND2_X1 U15163 ( .A1(n12101), .A2(n12099), .ZN(n12096) );
  NAND2_X1 U15164 ( .A1(n20273), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12095) );
  NAND2_X1 U15165 ( .A1(n12096), .A2(n12095), .ZN(n12103) );
  INV_X1 U15166 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12878) );
  NOR2_X1 U15167 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12878), .ZN(
        n12097) );
  INV_X1 U15168 ( .A(n12099), .ZN(n12100) );
  XNOR2_X1 U15169 ( .A(n12101), .B(n12100), .ZN(n12148) );
  XNOR2_X1 U15170 ( .A(n12105), .B(n12104), .ZN(n12134) );
  XNOR2_X1 U15171 ( .A(n12107), .B(n12106), .ZN(n12143) );
  NOR3_X1 U15172 ( .A1(n12149), .A2(n12134), .A3(n12143), .ZN(n12108) );
  AND2_X1 U15173 ( .A1(n12148), .A2(n12108), .ZN(n12109) );
  NOR2_X1 U15174 ( .A1(n12117), .A2(n12109), .ZN(n14406) );
  NAND2_X1 U15175 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20747) );
  NAND2_X1 U15176 ( .A1(n14406), .A2(n20747), .ZN(n12869) );
  INV_X1 U15177 ( .A(n12869), .ZN(n12110) );
  NAND2_X1 U15178 ( .A1(n12111), .A2(n12110), .ZN(n12159) );
  INV_X1 U15179 ( .A(n15930), .ZN(n13442) );
  INV_X1 U15180 ( .A(n20747), .ZN(n15929) );
  OAI21_X1 U15181 ( .B1(n12112), .B2(n15929), .A(n9765), .ZN(n12113) );
  OAI21_X1 U15182 ( .B1(n13442), .B2(n11818), .A(n12113), .ZN(n12114) );
  NAND2_X1 U15183 ( .A1(n12114), .A2(n11797), .ZN(n12158) );
  NOR2_X1 U15184 ( .A1(n12116), .A2(n12115), .ZN(n12121) );
  NAND2_X1 U15185 ( .A1(n12121), .A2(n12117), .ZN(n12157) );
  NAND2_X1 U15186 ( .A1(n12117), .A2(n12131), .ZN(n12155) );
  INV_X1 U15187 ( .A(n12148), .ZN(n12146) );
  NAND2_X1 U15188 ( .A1(n13139), .A2(n9765), .ZN(n12118) );
  NAND2_X1 U15189 ( .A1(n12118), .A2(n11809), .ZN(n12142) );
  INV_X1 U15190 ( .A(n12142), .ZN(n12120) );
  INV_X1 U15191 ( .A(n12131), .ZN(n12144) );
  NOR2_X1 U15192 ( .A1(n12144), .A2(n12143), .ZN(n12119) );
  AOI211_X1 U15193 ( .C1(n12150), .C2(n12143), .A(n12120), .B(n12119), .ZN(
        n12141) );
  INV_X1 U15194 ( .A(n12121), .ZN(n12125) );
  OAI21_X1 U15195 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20449), .A(
        n12122), .ZN(n12123) );
  INV_X1 U15196 ( .A(n12123), .ZN(n12126) );
  NAND2_X1 U15197 ( .A1(n12131), .A2(n12126), .ZN(n12124) );
  NAND2_X1 U15198 ( .A1(n12125), .A2(n12124), .ZN(n12128) );
  OAI211_X1 U15199 ( .C1(n11802), .C2(n13449), .A(n12142), .B(n12126), .ZN(
        n12127) );
  NAND2_X1 U15200 ( .A1(n12128), .A2(n12127), .ZN(n12135) );
  INV_X1 U15201 ( .A(n12135), .ZN(n12139) );
  NOR2_X1 U15202 ( .A1(n12129), .A2(n11886), .ZN(n12130) );
  AOI21_X1 U15203 ( .B1(n12131), .B2(n12180), .A(n12130), .ZN(n12133) );
  NAND2_X1 U15204 ( .A1(n12150), .A2(n12134), .ZN(n12132) );
  AND2_X1 U15205 ( .A1(n12133), .A2(n12132), .ZN(n12136) );
  INV_X1 U15206 ( .A(n12136), .ZN(n12138) );
  NAND2_X1 U15207 ( .A1(n12133), .A2(n12180), .ZN(n12152) );
  AOI22_X1 U15208 ( .A1(n12136), .A2(n12135), .B1(n12134), .B2(n12152), .ZN(
        n12137) );
  AOI21_X1 U15209 ( .B1(n12139), .B2(n12138), .A(n12137), .ZN(n12140) );
  NOR3_X1 U15210 ( .A1(n12144), .A2(n12143), .A3(n12142), .ZN(n12145) );
  INV_X1 U15211 ( .A(n12149), .ZN(n12147) );
  AOI21_X1 U15212 ( .B1(n12148), .B2(n12147), .A(n12150), .ZN(n12153) );
  NAND2_X1 U15213 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  NAND2_X1 U15214 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  NOR2_X1 U15215 ( .A1(n12161), .A2(n12160), .ZN(n12279) );
  NAND2_X1 U15216 ( .A1(n14944), .A2(n13449), .ZN(n12162) );
  NAND2_X1 U15217 ( .A1(n12163), .A2(n13671), .ZN(n12292) );
  AND2_X1 U15218 ( .A1(n12292), .A2(n9766), .ZN(n12164) );
  NAND2_X1 U15219 ( .A1(n12165), .A2(n12164), .ZN(n12286) );
  NAND2_X1 U15220 ( .A1(n12881), .A2(n12286), .ZN(n12167) );
  NAND2_X1 U15221 ( .A1(n12167), .A2(n12166), .ZN(n12866) );
  OR2_X1 U15222 ( .A1(n15907), .A2(n12292), .ZN(n12168) );
  OR2_X1 U15223 ( .A1(n12880), .A2(n13438), .ZN(n12172) );
  NAND2_X1 U15224 ( .A1(n12881), .A2(n12172), .ZN(n14401) );
  OAI22_X1 U15225 ( .A1(n11809), .A2(n12173), .B1(n12174), .B2(n13679), .ZN(
        n12175) );
  INV_X1 U15226 ( .A(n12175), .ZN(n12176) );
  NAND3_X1 U15227 ( .A1(n9907), .A2(n14401), .A3(n12176), .ZN(n12177) );
  INV_X1 U15228 ( .A(n12173), .ZN(n12860) );
  NAND2_X1 U15229 ( .A1(n12860), .A2(n11809), .ZN(n12633) );
  OAI21_X1 U15230 ( .B1(n12174), .B2(n11857), .A(n12633), .ZN(n12178) );
  INV_X1 U15231 ( .A(n12836), .ZN(n13144) );
  AOI22_X1 U15232 ( .A1(n12833), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14410), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14416) );
  INV_X1 U15233 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12182) );
  INV_X1 U15234 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U15235 ( .A1(n12205), .A2(n12996), .ZN(n12184) );
  NAND2_X1 U15236 ( .A1(n13463), .A2(n12182), .ZN(n12183) );
  NAND3_X1 U15237 ( .A1(n12184), .A2(n12179), .A3(n12183), .ZN(n12185) );
  NAND2_X1 U15238 ( .A1(n12186), .A2(n12185), .ZN(n12189) );
  NAND2_X1 U15239 ( .A1(n12205), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12188) );
  INV_X1 U15240 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12852) );
  NAND2_X1 U15241 ( .A1(n12179), .A2(n12852), .ZN(n12187) );
  NAND2_X1 U15242 ( .A1(n12188), .A2(n12187), .ZN(n12834) );
  XNOR2_X1 U15243 ( .A(n12189), .B(n12834), .ZN(n12979) );
  NAND2_X1 U15244 ( .A1(n13455), .A2(n12189), .ZN(n13035) );
  NAND2_X1 U15245 ( .A1(n12213), .A2(n14410), .ZN(n12245) );
  NAND2_X1 U15246 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14410), .ZN(
        n12190) );
  AND2_X1 U15247 ( .A1(n12245), .A2(n12190), .ZN(n12191) );
  AND2_X1 U15248 ( .A1(n12192), .A2(n12191), .ZN(n13034) );
  MUX2_X1 U15249 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12193) );
  OAI21_X1 U15250 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n12833), .A(
        n12193), .ZN(n13094) );
  MUX2_X1 U15251 ( .A(n12243), .B(n12205), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12196) );
  NAND2_X1 U15252 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14410), .ZN(
        n12194) );
  AND2_X1 U15253 ( .A1(n12245), .A2(n12194), .ZN(n12195) );
  NAND2_X1 U15254 ( .A1(n12196), .A2(n12195), .ZN(n13110) );
  NAND2_X1 U15255 ( .A1(n13111), .A2(n13110), .ZN(n16252) );
  INV_X1 U15256 ( .A(n16252), .ZN(n12200) );
  NAND2_X1 U15257 ( .A1(n12179), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12197) );
  OAI211_X1 U15258 ( .C1(n14410), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12205), .B(
        n12197), .ZN(n12198) );
  OAI21_X1 U15259 ( .B1(n12265), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12198), .ZN(
        n16251) );
  MUX2_X1 U15260 ( .A(n12243), .B(n12205), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12203) );
  NAND2_X1 U15261 ( .A1(n14410), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12201) );
  AND2_X1 U15262 ( .A1(n12245), .A2(n12201), .ZN(n12202) );
  NAND2_X1 U15263 ( .A1(n12203), .A2(n12202), .ZN(n16230) );
  INV_X1 U15264 ( .A(n12265), .ZN(n12204) );
  NAND2_X1 U15265 ( .A1(n12204), .A2(n20135), .ZN(n12208) );
  INV_X1 U15266 ( .A(n12205), .ZN(n12213) );
  NAND2_X1 U15267 ( .A1(n12179), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12206) );
  OAI211_X1 U15268 ( .C1(n14410), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12205), .B(
        n12206), .ZN(n12207) );
  AND2_X1 U15269 ( .A1(n12208), .A2(n12207), .ZN(n16229) );
  NAND2_X1 U15270 ( .A1(n16230), .A2(n16229), .ZN(n12209) );
  MUX2_X1 U15271 ( .A(n12243), .B(n12205), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12212) );
  NAND2_X1 U15272 ( .A1(n14410), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12210) );
  AND2_X1 U15273 ( .A1(n12245), .A2(n12210), .ZN(n12211) );
  NAND2_X1 U15274 ( .A1(n12212), .A2(n12211), .ZN(n13572) );
  NAND2_X1 U15275 ( .A1(n12179), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12214) );
  OAI211_X1 U15276 ( .C1(n14410), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12205), .B(
        n12214), .ZN(n12215) );
  OAI21_X1 U15277 ( .B1(n12265), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12215), .ZN(
        n16216) );
  INV_X1 U15278 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13870) );
  INV_X1 U15279 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14837) );
  NAND2_X1 U15280 ( .A1(n12205), .A2(n14837), .ZN(n12217) );
  NAND2_X1 U15281 ( .A1(n13463), .A2(n13870), .ZN(n12216) );
  NAND3_X1 U15282 ( .A1(n12217), .A2(n12179), .A3(n12216), .ZN(n12218) );
  INV_X1 U15283 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16202) );
  INV_X1 U15284 ( .A(n12833), .ZN(n12278) );
  NAND2_X1 U15285 ( .A1(n16202), .A2(n12278), .ZN(n12221) );
  MUX2_X1 U15286 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12220) );
  NAND2_X1 U15287 ( .A1(n12221), .A2(n12220), .ZN(n13982) );
  MUX2_X1 U15288 ( .A(n12243), .B(n12205), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12224) );
  NAND2_X1 U15289 ( .A1(n14410), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12222) );
  AND2_X1 U15290 ( .A1(n12245), .A2(n12222), .ZN(n12223) );
  NAND2_X1 U15291 ( .A1(n12224), .A2(n12223), .ZN(n14620) );
  MUX2_X1 U15292 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12226) );
  OR2_X1 U15293 ( .A1(n12833), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12225) );
  INV_X1 U15294 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n16017) );
  NAND2_X1 U15295 ( .A1(n12205), .A2(n12227), .ZN(n12229) );
  NAND2_X1 U15296 ( .A1(n13463), .A2(n16017), .ZN(n12228) );
  NAND3_X1 U15297 ( .A1(n12229), .A2(n12179), .A3(n12228), .ZN(n12230) );
  MUX2_X1 U15298 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12232) );
  OAI21_X1 U15299 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n12833), .A(
        n12232), .ZN(n14613) );
  NAND2_X1 U15300 ( .A1(n12205), .A2(n12296), .ZN(n12234) );
  INV_X1 U15301 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15999) );
  NAND2_X1 U15302 ( .A1(n13463), .A2(n15999), .ZN(n12233) );
  NAND3_X1 U15303 ( .A1(n12234), .A2(n12179), .A3(n12233), .ZN(n12235) );
  OAI21_X1 U15304 ( .B1(n12243), .B2(P1_EBX_REG_16__SCAN_IN), .A(n12235), .ZN(
        n14603) );
  NAND2_X1 U15305 ( .A1(n12179), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12236) );
  OAI211_X1 U15306 ( .C1(n14410), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12205), .B(
        n12236), .ZN(n12237) );
  OAI21_X1 U15307 ( .B1(n12265), .B2(P1_EBX_REG_17__SCAN_IN), .A(n12237), .ZN(
        n14522) );
  INV_X1 U15308 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U15309 ( .A1(n12205), .A2(n16164), .ZN(n12239) );
  NAND2_X1 U15310 ( .A1(n13463), .A2(n15983), .ZN(n12238) );
  NAND3_X1 U15311 ( .A1(n12239), .A2(n12179), .A3(n12238), .ZN(n12240) );
  AND2_X1 U15312 ( .A1(n12241), .A2(n12240), .ZN(n14596) );
  MUX2_X1 U15313 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12242) );
  OAI21_X1 U15314 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n12833), .A(
        n12242), .ZN(n14589) );
  NOR2_X4 U15315 ( .A1(n14598), .A2(n14589), .ZN(n14591) );
  MUX2_X1 U15316 ( .A(n12243), .B(n12205), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12247) );
  NAND2_X1 U15317 ( .A1(n14410), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12244) );
  AND2_X1 U15318 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  NAND2_X1 U15319 ( .A1(n12247), .A2(n12246), .ZN(n14582) );
  MUX2_X1 U15320 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12248) );
  OAI21_X1 U15321 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n12833), .A(
        n12248), .ZN(n14574) );
  INV_X1 U15322 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14568) );
  INV_X1 U15323 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12249) );
  NAND2_X1 U15324 ( .A1(n12205), .A2(n12249), .ZN(n12251) );
  NAND2_X1 U15325 ( .A1(n13463), .A2(n14568), .ZN(n12250) );
  NAND3_X1 U15326 ( .A1(n12251), .A2(n12179), .A3(n12250), .ZN(n12252) );
  NAND2_X1 U15327 ( .A1(n12253), .A2(n12252), .ZN(n14565) );
  MUX2_X1 U15328 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12254) );
  OAI21_X1 U15329 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n12833), .A(
        n12254), .ZN(n14510) );
  INV_X1 U15330 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n12255) );
  INV_X1 U15331 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14886) );
  NAND2_X1 U15332 ( .A1(n12205), .A2(n14886), .ZN(n12257) );
  NAND2_X1 U15333 ( .A1(n13463), .A2(n12255), .ZN(n12256) );
  NAND3_X1 U15334 ( .A1(n12257), .A2(n12179), .A3(n12256), .ZN(n12258) );
  AND2_X1 U15335 ( .A1(n12259), .A2(n12258), .ZN(n14500) );
  OR2_X2 U15336 ( .A1(n14512), .A2(n14500), .ZN(n14498) );
  MUX2_X1 U15337 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12260) );
  OAI21_X1 U15338 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n12833), .A(
        n12260), .ZN(n14477) );
  INV_X1 U15339 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14558) );
  INV_X1 U15340 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14765) );
  NAND2_X1 U15341 ( .A1(n12205), .A2(n14765), .ZN(n12262) );
  NAND2_X1 U15342 ( .A1(n13463), .A2(n14558), .ZN(n12261) );
  NAND3_X1 U15343 ( .A1(n12262), .A2(n12179), .A3(n12261), .ZN(n12263) );
  NAND2_X1 U15344 ( .A1(n12264), .A2(n12263), .ZN(n14462) );
  MUX2_X1 U15345 ( .A(n12265), .B(n12179), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12266) );
  OAI21_X1 U15346 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n12833), .A(
        n12266), .ZN(n12267) );
  INV_X1 U15347 ( .A(n12267), .ZN(n14449) );
  INV_X1 U15348 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n12269) );
  INV_X1 U15349 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12268) );
  NAND2_X1 U15350 ( .A1(n12205), .A2(n12268), .ZN(n12271) );
  NAND2_X1 U15351 ( .A1(n13463), .A2(n12269), .ZN(n12270) );
  NAND3_X1 U15352 ( .A1(n12271), .A2(n12179), .A3(n12270), .ZN(n12272) );
  AND2_X1 U15353 ( .A1(n12273), .A2(n12272), .ZN(n14442) );
  OR2_X1 U15354 ( .A1(n12833), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12274) );
  INV_X1 U15355 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14556) );
  NAND2_X1 U15356 ( .A1(n13463), .A2(n14556), .ZN(n12275) );
  NAND2_X1 U15357 ( .A1(n12274), .A2(n12275), .ZN(n14415) );
  MUX2_X1 U15358 ( .A(n14415), .B(n12275), .S(n12181), .Z(n14425) );
  MUX2_X1 U15359 ( .A(n12179), .B(n14416), .S(n14426), .Z(n12277) );
  AOI22_X1 U15360 ( .A1(n12833), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14410), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12276) );
  INV_X1 U15361 ( .A(n14553), .ZN(n12311) );
  OR2_X1 U15362 ( .A1(n12279), .A2(n12278), .ZN(n12284) );
  INV_X1 U15363 ( .A(n11819), .ZN(n12281) );
  NAND2_X1 U15364 ( .A1(n11797), .A2(n12863), .ZN(n12280) );
  OAI211_X1 U15365 ( .C1(n12880), .C2(n9723), .A(n12281), .B(n12280), .ZN(
        n12282) );
  NAND2_X1 U15366 ( .A1(n12282), .A2(n12180), .ZN(n12283) );
  AND2_X1 U15367 ( .A1(n12286), .A2(n12285), .ZN(n12289) );
  INV_X1 U15368 ( .A(n11808), .ZN(n12287) );
  NAND2_X1 U15369 ( .A1(n12287), .A2(n13438), .ZN(n12288) );
  AND3_X1 U15370 ( .A1(n12294), .A2(n12289), .A3(n12288), .ZN(n12962) );
  OAI211_X1 U15371 ( .C1(n12959), .C2(n9766), .A(n12962), .B(n12290), .ZN(
        n12291) );
  INV_X1 U15372 ( .A(n12292), .ZN(n12293) );
  NOR2_X1 U15373 ( .A1(n12166), .A2(n11809), .ZN(n14948) );
  NAND2_X1 U15374 ( .A1(n12299), .A2(n14948), .ZN(n13045) );
  NAND2_X1 U15375 ( .A1(n12856), .A2(n13045), .ZN(n14910) );
  AOI21_X1 U15376 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13171) );
  NAND2_X1 U15377 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13825) );
  NOR2_X1 U15378 ( .A1(n12040), .A2(n13825), .ZN(n16239) );
  INV_X1 U15379 ( .A(n16239), .ZN(n14918) );
  NOR2_X1 U15380 ( .A1(n13171), .A2(n14918), .ZN(n16204) );
  INV_X1 U15381 ( .A(n16204), .ZN(n12295) );
  INV_X1 U15382 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13827) );
  NAND2_X1 U15383 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16213) );
  NOR2_X1 U15384 ( .A1(n13827), .A2(n16213), .ZN(n16205) );
  NAND3_X1 U15385 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16205), .ZN(n14924) );
  NOR2_X1 U15386 ( .A1(n16202), .A2(n14924), .ZN(n14927) );
  NAND2_X1 U15387 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14927), .ZN(
        n12298) );
  NOR2_X1 U15388 ( .A1(n12295), .A2(n12298), .ZN(n14907) );
  INV_X1 U15389 ( .A(n14907), .ZN(n13902) );
  NOR3_X1 U15390 ( .A1(n14912), .A2(n12296), .A3(n12078), .ZN(n16166) );
  NAND3_X1 U15391 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n16166), .ZN(n12308) );
  INV_X1 U15392 ( .A(n12308), .ZN(n12300) );
  NAND2_X1 U15393 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12300), .ZN(
        n16159) );
  NAND3_X1 U15394 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n16239), .ZN(n14922) );
  NOR2_X1 U15395 ( .A1(n12298), .A2(n14922), .ZN(n12307) );
  AND2_X1 U15396 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12307), .ZN(
        n13900) );
  INV_X1 U15397 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20984) );
  NAND3_X1 U15398 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n14898), .ZN(n15912) );
  NAND2_X1 U15399 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16153) );
  INV_X1 U15400 ( .A(n14910), .ZN(n16167) );
  NAND2_X1 U15401 ( .A1(n16167), .A2(n14919), .ZN(n16206) );
  OAI21_X1 U15402 ( .B1(n15912), .B2(n16153), .A(n16206), .ZN(n16147) );
  INV_X1 U15403 ( .A(n12301), .ZN(n14740) );
  OR2_X1 U15404 ( .A1(n13045), .A2(n14740), .ZN(n12302) );
  OAI211_X1 U15405 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n12856), .A(
        n16147), .B(n12302), .ZN(n12304) );
  AND2_X1 U15406 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16128) );
  INV_X1 U15407 ( .A(n12856), .ZN(n12303) );
  AOI21_X1 U15408 ( .B1(n14886), .B2(n12303), .A(n12304), .ZN(n16137) );
  OAI21_X1 U15409 ( .B1(n16167), .B2(n16128), .A(n16137), .ZN(n14880) );
  AOI21_X1 U15410 ( .B1(n14863), .B2(n14910), .A(n14880), .ZN(n14857) );
  OAI211_X1 U15411 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16167), .A(
        n14857), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14849) );
  NAND2_X1 U15412 ( .A1(n20177), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14380) );
  INV_X1 U15413 ( .A(n13045), .ZN(n14900) );
  NAND3_X1 U15414 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12305), .A3(
        n12307), .ZN(n12306) );
  OAI21_X1 U15415 ( .B1(n13902), .B2(n14920), .A(n12306), .ZN(n14899) );
  NOR3_X1 U15416 ( .A1(n12249), .A2(n12309), .A3(n12308), .ZN(n16138) );
  NAND3_X1 U15417 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16140), .A3(
        n16138), .ZN(n14883) );
  NOR2_X1 U15418 ( .A1(n14886), .A2(n14883), .ZN(n16129) );
  NAND2_X1 U15419 ( .A1(n16129), .A2(n16128), .ZN(n14866) );
  NOR3_X1 U15420 ( .A1(n14866), .A2(n14863), .A3(n14856), .ZN(n14850) );
  NAND3_X1 U15421 ( .A1(n14850), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12087), .ZN(n12310) );
  NAND2_X1 U15422 ( .A1(n12312), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12313) );
  NOR2_X1 U15423 ( .A1(n20047), .A2(n10880), .ZN(n19883) );
  AND2_X1 U15424 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19883), .ZN(
        n12314) );
  NAND2_X1 U15425 ( .A1(n12314), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19882) );
  INV_X1 U15426 ( .A(n12314), .ZN(n12331) );
  NAND2_X1 U15427 ( .A1(n12315), .A2(n12331), .ZN(n12316) );
  AND3_X1 U15428 ( .A1(n19882), .A2(n20029), .A3(n12316), .ZN(n19777) );
  AOI21_X1 U15429 ( .B1(n12333), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19777), .ZN(n12317) );
  INV_X1 U15430 ( .A(n12344), .ZN(n12322) );
  NOR2_X1 U15431 ( .A1(n12312), .A2(n19309), .ZN(n12319) );
  NOR2_X1 U15432 ( .A1(n12518), .A2(n12320), .ZN(n12323) );
  INV_X1 U15433 ( .A(n12323), .ZN(n12321) );
  NAND2_X1 U15434 ( .A1(n12322), .A2(n12321), .ZN(n12324) );
  NAND2_X1 U15435 ( .A1(n12344), .A2(n12323), .ZN(n13176) );
  NAND2_X1 U15436 ( .A1(n12324), .A2(n13176), .ZN(n12827) );
  INV_X1 U15437 ( .A(n12827), .ZN(n12342) );
  AOI22_X1 U15438 ( .A1(n12333), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20029), .B2(n21022), .ZN(n12325) );
  INV_X1 U15439 ( .A(n12335), .ZN(n12326) );
  NAND2_X1 U15440 ( .A1(n9774), .A2(n12326), .ZN(n12329) );
  NAND2_X1 U15441 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10880), .ZN(
        n19671) );
  NAND2_X1 U15442 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21022), .ZN(
        n19705) );
  NAND2_X1 U15443 ( .A1(n19671), .A2(n19705), .ZN(n19707) );
  AND2_X1 U15444 ( .A1(n20029), .A2(n19707), .ZN(n19471) );
  AOI21_X1 U15445 ( .B1(n12333), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19471), .ZN(n12328) );
  NAND2_X1 U15446 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19739) );
  NAND2_X1 U15447 ( .A1(n19739), .A2(n20047), .ZN(n12332) );
  AND2_X1 U15448 ( .A1(n12332), .A2(n12331), .ZN(n13739) );
  AOI22_X1 U15449 ( .A1(n12333), .A2(n15720), .B1(n20029), .B2(n13739), .ZN(
        n12334) );
  INV_X1 U15450 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12337) );
  NOR2_X1 U15451 ( .A1(n12518), .A2(n12337), .ZN(n12338) );
  NAND2_X1 U15452 ( .A1(n12342), .A2(n12826), .ZN(n12829) );
  NAND2_X1 U15453 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10656), .ZN(
        n12343) );
  NAND2_X1 U15454 ( .A1(n12829), .A2(n12343), .ZN(n13178) );
  INV_X1 U15455 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12345) );
  NOR2_X1 U15456 ( .A1(n12518), .A2(n12345), .ZN(n13174) );
  NAND2_X1 U15457 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12346) );
  NAND2_X1 U15458 ( .A1(n13117), .A2(n12347), .ZN(n12348) );
  AND2_X1 U15459 ( .A1(n13199), .A2(n13201), .ZN(n12349) );
  INV_X1 U15460 ( .A(n12350), .ZN(n13474) );
  AOI22_X1 U15461 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10849), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15462 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15463 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15464 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12352) );
  NAND4_X1 U15465 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12361) );
  AOI22_X1 U15466 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15467 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15468 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15469 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12356) );
  NAND4_X1 U15470 ( .A1(n12359), .A2(n12358), .A3(n12357), .A4(n12356), .ZN(
        n12360) );
  OR2_X1 U15471 ( .A1(n12361), .A2(n12360), .ZN(n15178) );
  AOI22_X1 U15472 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15473 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15474 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15475 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12362) );
  NAND4_X1 U15476 ( .A1(n12365), .A2(n12364), .A3(n12363), .A4(n12362), .ZN(
        n12371) );
  AOI22_X1 U15477 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15478 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15479 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15480 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12366) );
  NAND4_X1 U15481 ( .A1(n12369), .A2(n12368), .A3(n12367), .A4(n12366), .ZN(
        n12370) );
  OR2_X1 U15482 ( .A1(n12371), .A2(n12370), .ZN(n13885) );
  AOI22_X1 U15483 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10832), .B1(
        n10849), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15484 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15485 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U15486 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12372) );
  NAND4_X1 U15487 ( .A1(n12375), .A2(n12374), .A3(n12373), .A4(n12372), .ZN(
        n12381) );
  AOI22_X1 U15488 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15489 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15490 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15491 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12376) );
  NAND4_X1 U15492 ( .A1(n12379), .A2(n12378), .A3(n12377), .A4(n12376), .ZN(
        n12380) );
  OR2_X1 U15493 ( .A1(n12381), .A2(n12380), .ZN(n13836) );
  AOI22_X1 U15494 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10849), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15495 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15496 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15497 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12382) );
  NAND4_X1 U15498 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12391) );
  AOI22_X1 U15499 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15500 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15501 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15502 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12386) );
  NAND4_X1 U15503 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12390) );
  OR2_X1 U15504 ( .A1(n12391), .A2(n12390), .ZN(n13884) );
  AOI22_X1 U15505 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10849), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15506 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15507 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15508 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12392) );
  NAND4_X1 U15509 ( .A1(n12395), .A2(n12394), .A3(n12393), .A4(n12392), .ZN(
        n12401) );
  AOI22_X1 U15510 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15511 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15512 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15513 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12396) );
  NAND4_X1 U15514 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12400) );
  OR2_X1 U15515 ( .A1(n12401), .A2(n12400), .ZN(n15145) );
  AND4_X1 U15516 ( .A1(n13885), .A2(n13836), .A3(n13884), .A4(n15145), .ZN(
        n12402) );
  AOI22_X1 U15517 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10849), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15518 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U15519 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15520 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12403) );
  NAND4_X1 U15521 ( .A1(n12406), .A2(n12405), .A3(n12404), .A4(n12403), .ZN(
        n12412) );
  AOI22_X1 U15522 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15523 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15524 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15525 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12407) );
  NAND4_X1 U15526 ( .A1(n12410), .A2(n12409), .A3(n12408), .A4(n12407), .ZN(
        n12411) );
  NOR2_X1 U15527 ( .A1(n12412), .A2(n12411), .ZN(n15137) );
  INV_X1 U15528 ( .A(n15137), .ZN(n12413) );
  AOI22_X1 U15529 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10849), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15530 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15531 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15532 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10863), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12414) );
  NAND4_X1 U15533 ( .A1(n12417), .A2(n12416), .A3(n12415), .A4(n12414), .ZN(
        n12423) );
  AOI22_X1 U15534 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15535 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11419), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15536 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12447), .B1(
        n10840), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15537 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10825), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12418) );
  NAND4_X1 U15538 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12422) );
  NOR2_X1 U15539 ( .A1(n12423), .A2(n12422), .ZN(n15134) );
  AND2_X1 U15540 ( .A1(n15720), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12425) );
  OR2_X1 U15541 ( .A1(n12425), .A2(n12424), .ZN(n12590) );
  INV_X1 U15542 ( .A(n12590), .ZN(n12564) );
  NAND2_X1 U15543 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12428) );
  NAND2_X1 U15544 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12427) );
  AND3_X1 U15545 ( .A1(n12564), .A2(n12428), .A3(n12427), .ZN(n12434) );
  AOI22_X1 U15546 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15547 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15548 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12431) );
  NAND4_X1 U15549 ( .A1(n12434), .A2(n12433), .A3(n12432), .A4(n12431), .ZN(
        n12442) );
  AOI22_X1 U15550 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12440) );
  NAND2_X1 U15551 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12436) );
  NAND2_X1 U15552 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12435) );
  AND3_X1 U15553 ( .A1(n12436), .A2(n12590), .A3(n12435), .ZN(n12439) );
  AOI22_X1 U15554 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15555 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12437) );
  NAND4_X1 U15556 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12441) );
  NAND2_X1 U15557 ( .A1(n12442), .A2(n12441), .ZN(n12476) );
  NOR2_X1 U15558 ( .A1(n11377), .A2(n12476), .ZN(n12454) );
  AOI22_X1 U15559 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10849), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15560 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15561 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10850), .B1(
        n10909), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15562 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11419), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12443) );
  NAND4_X1 U15563 ( .A1(n12446), .A2(n12445), .A3(n12444), .A4(n12443), .ZN(
        n12453) );
  AOI22_X1 U15564 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10779), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15565 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10863), .B1(
        n11420), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15566 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10840), .B1(
        n10841), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15567 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10825), .B1(
        n12447), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12448) );
  NAND4_X1 U15568 ( .A1(n12451), .A2(n12450), .A3(n12449), .A4(n12448), .ZN(
        n12452) );
  NOR2_X1 U15569 ( .A1(n12453), .A2(n12452), .ZN(n12471) );
  XNOR2_X1 U15570 ( .A(n12454), .B(n12471), .ZN(n12478) );
  INV_X1 U15571 ( .A(n12476), .ZN(n12472) );
  NAND2_X1 U15572 ( .A1(n11377), .A2(n12472), .ZN(n15127) );
  NAND2_X1 U15573 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12458) );
  NAND2_X1 U15574 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12457) );
  AND3_X1 U15575 ( .A1(n12564), .A2(n12458), .A3(n12457), .ZN(n12462) );
  AOI22_X1 U15576 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U15577 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15578 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12459) );
  NAND4_X1 U15579 ( .A1(n12462), .A2(n12461), .A3(n12460), .A4(n12459), .ZN(
        n12470) );
  AOI22_X1 U15580 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U15581 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12464) );
  NAND2_X1 U15582 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12463) );
  AND3_X1 U15583 ( .A1(n12464), .A2(n12590), .A3(n12463), .ZN(n12467) );
  AOI22_X1 U15584 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15585 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12465) );
  NAND4_X1 U15586 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12465), .ZN(
        n12469) );
  NAND2_X1 U15587 ( .A1(n12470), .A2(n12469), .ZN(n12480) );
  INV_X1 U15588 ( .A(n12471), .ZN(n12473) );
  NAND2_X1 U15589 ( .A1(n12473), .A2(n12472), .ZN(n12481) );
  XOR2_X1 U15590 ( .A(n12480), .B(n12481), .Z(n12474) );
  INV_X1 U15591 ( .A(n12518), .ZN(n12540) );
  NAND2_X1 U15592 ( .A1(n12474), .A2(n12540), .ZN(n15117) );
  INV_X1 U15593 ( .A(n12480), .ZN(n12475) );
  NAND2_X1 U15594 ( .A1(n11377), .A2(n12475), .ZN(n15119) );
  NOR2_X1 U15595 ( .A1(n15119), .A2(n12476), .ZN(n12477) );
  NOR2_X1 U15596 ( .A1(n12481), .A2(n12480), .ZN(n12496) );
  AOI22_X1 U15597 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12487) );
  INV_X1 U15598 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n21068) );
  NAND2_X1 U15599 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12483) );
  NAND2_X1 U15600 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12482) );
  AND3_X1 U15601 ( .A1(n12564), .A2(n12483), .A3(n12482), .ZN(n12486) );
  AOI22_X1 U15602 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15603 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15604 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12495) );
  AOI22_X1 U15605 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9738), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12493) );
  NAND2_X1 U15606 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12489) );
  NAND2_X1 U15607 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12488) );
  AND3_X1 U15608 ( .A1(n12489), .A2(n12590), .A3(n12488), .ZN(n12492) );
  AOI22_X1 U15609 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15610 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12490) );
  NAND4_X1 U15611 ( .A1(n12493), .A2(n12492), .A3(n12491), .A4(n12490), .ZN(
        n12494) );
  AND2_X1 U15612 ( .A1(n12495), .A2(n12494), .ZN(n12498) );
  NAND2_X1 U15613 ( .A1(n12496), .A2(n12498), .ZN(n12519) );
  OAI211_X1 U15614 ( .C1(n12496), .C2(n12498), .A(n12540), .B(n12519), .ZN(
        n12501) );
  INV_X1 U15615 ( .A(n12498), .ZN(n12499) );
  NOR2_X1 U15616 ( .A1(n13331), .A2(n12499), .ZN(n15112) );
  INV_X1 U15617 ( .A(n12500), .ZN(n12502) );
  NAND2_X1 U15618 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12505) );
  NAND2_X1 U15619 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12504) );
  AND3_X1 U15620 ( .A1(n12564), .A2(n12505), .A3(n12504), .ZN(n12509) );
  AOI22_X1 U15621 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15622 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U15623 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12506) );
  NAND4_X1 U15624 ( .A1(n12509), .A2(n12508), .A3(n12507), .A4(n12506), .ZN(
        n12517) );
  AOI22_X1 U15625 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12515) );
  NAND2_X1 U15626 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12511) );
  NAND2_X1 U15627 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12510) );
  AND3_X1 U15628 ( .A1(n12511), .A2(n12590), .A3(n12510), .ZN(n12514) );
  AOI22_X1 U15629 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15630 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12512) );
  NAND4_X1 U15631 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12516) );
  NAND2_X1 U15632 ( .A1(n12517), .A2(n12516), .ZN(n12521) );
  AOI21_X1 U15633 ( .B1(n12519), .B2(n12521), .A(n12518), .ZN(n12520) );
  OR2_X1 U15634 ( .A1(n12519), .A2(n12521), .ZN(n12539) );
  INV_X1 U15635 ( .A(n12521), .ZN(n12522) );
  NAND2_X1 U15636 ( .A1(n11377), .A2(n12522), .ZN(n15106) );
  NOR2_X2 U15637 ( .A1(n15105), .A2(n12524), .ZN(n12544) );
  AOI22_X1 U15638 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15639 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9738), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15640 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U15641 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12526) );
  NAND2_X1 U15642 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12525) );
  AND3_X1 U15643 ( .A1(n12526), .A2(n12590), .A3(n12525), .ZN(n12527) );
  NAND4_X1 U15644 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        n12538) );
  AOI22_X1 U15645 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U15646 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12532) );
  NAND2_X1 U15647 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12531) );
  AND3_X1 U15648 ( .A1(n12564), .A2(n12532), .A3(n12531), .ZN(n12535) );
  AOI22_X1 U15649 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15650 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12533) );
  NAND4_X1 U15651 ( .A1(n12536), .A2(n12535), .A3(n12534), .A4(n12533), .ZN(
        n12537) );
  NAND2_X1 U15652 ( .A1(n12538), .A2(n12537), .ZN(n12546) );
  INV_X1 U15653 ( .A(n12546), .ZN(n12542) );
  INV_X1 U15654 ( .A(n12539), .ZN(n12541) );
  OR2_X1 U15655 ( .A1(n12539), .A2(n12546), .ZN(n12577) );
  NOR2_X2 U15656 ( .A1(n12547), .A2(n12545), .ZN(n15096) );
  NOR2_X1 U15657 ( .A1(n13331), .A2(n12546), .ZN(n15098) );
  NAND2_X1 U15658 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12549) );
  NAND2_X1 U15659 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12548) );
  AND3_X1 U15660 ( .A1(n12564), .A2(n12549), .A3(n12548), .ZN(n12553) );
  AOI22_X1 U15661 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15662 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15663 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12550) );
  NAND4_X1 U15664 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12561) );
  AOI22_X1 U15665 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12559) );
  NAND2_X1 U15666 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12555) );
  NAND2_X1 U15667 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12554) );
  AND3_X1 U15668 ( .A1(n12555), .A2(n12590), .A3(n12554), .ZN(n12558) );
  AOI22_X1 U15669 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15670 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12556) );
  NAND4_X1 U15671 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12560) );
  NAND2_X1 U15672 ( .A1(n12561), .A2(n12560), .ZN(n15092) );
  AOI22_X1 U15673 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15674 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U15675 ( .A1(n12456), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12563) );
  NAND2_X1 U15676 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12562) );
  AND3_X1 U15677 ( .A1(n12564), .A2(n12563), .A3(n12562), .ZN(n12566) );
  AOI22_X1 U15678 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12565) );
  NAND4_X1 U15679 ( .A1(n12568), .A2(n12567), .A3(n12566), .A4(n12565), .ZN(
        n12576) );
  AOI22_X1 U15680 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9738), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15681 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15682 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12572) );
  NAND2_X1 U15683 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12570) );
  NAND2_X1 U15684 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12569) );
  AND3_X1 U15685 ( .A1(n12570), .A2(n12590), .A3(n12569), .ZN(n12571) );
  NAND4_X1 U15686 ( .A1(n12574), .A2(n12573), .A3(n12572), .A4(n12571), .ZN(
        n12575) );
  NAND2_X1 U15687 ( .A1(n12576), .A2(n12575), .ZN(n12580) );
  INV_X1 U15688 ( .A(n12577), .ZN(n15091) );
  NOR2_X1 U15689 ( .A1(n11377), .A2(n15092), .ZN(n12578) );
  NAND2_X1 U15690 ( .A1(n15091), .A2(n12578), .ZN(n12579) );
  NOR2_X1 U15691 ( .A1(n12579), .A2(n12580), .ZN(n12581) );
  AOI21_X1 U15692 ( .B1(n12580), .B2(n12579), .A(n12581), .ZN(n15085) );
  INV_X1 U15693 ( .A(n12581), .ZN(n12582) );
  AOI22_X1 U15694 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15695 ( .A1(n9772), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U15696 ( .A1(n10787), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12583) );
  NAND4_X1 U15697 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12590), .ZN(
        n12598) );
  AOI22_X1 U15698 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9754), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15699 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15700 ( .A1(n12587), .A2(n12586), .ZN(n12597) );
  INV_X1 U15701 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12588) );
  NOR2_X1 U15702 ( .A1(n12426), .A2(n12588), .ZN(n12589) );
  AOI211_X1 U15703 ( .C1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n12456), .A(
        n12590), .B(n12589), .ZN(n12595) );
  AOI22_X1 U15704 ( .A1(n9754), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12429), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15705 ( .A1(n12591), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15706 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10786), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12592) );
  NAND4_X1 U15707 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12596) );
  OAI21_X1 U15708 ( .B1(n12598), .B2(n12597), .A(n12596), .ZN(n12599) );
  XNOR2_X1 U15709 ( .A(n12600), .B(n12599), .ZN(n15193) );
  INV_X1 U15710 ( .A(n13643), .ZN(n12601) );
  INV_X1 U15711 ( .A(n13581), .ZN(n13605) );
  NAND2_X1 U15712 ( .A1(n12601), .A2(n13605), .ZN(n12749) );
  NAND2_X1 U15713 ( .A1(n12749), .A2(n13583), .ZN(n12602) );
  NAND2_X1 U15714 ( .A1(n15193), .A2(n15149), .ZN(n12607) );
  INV_X1 U15715 ( .A(n16287), .ZN(n12604) );
  NAND2_X1 U15716 ( .A1(n12766), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U15717 ( .A1(n12607), .A2(n12606), .ZN(P2_U2857) );
  INV_X1 U15718 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20065) );
  NOR2_X1 U15719 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n20065), .ZN(n12609) );
  NOR4_X1 U15720 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_BE_N_REG_3__SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12608) );
  INV_X1 U15721 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n18998) );
  NAND4_X1 U15722 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n12609), .A3(n12608), .A4(
        n18998), .ZN(n12632) );
  NOR2_X1 U15723 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12632), .ZN(n16630)
         );
  NOR4_X1 U15724 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12613) );
  NOR4_X1 U15725 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12612) );
  NOR4_X1 U15726 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12611) );
  NOR4_X1 U15727 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12610) );
  AND4_X1 U15728 ( .A1(n12613), .A2(n12612), .A3(n12611), .A4(n12610), .ZN(
        n12618) );
  NOR4_X1 U15729 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_19__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12616) );
  NOR4_X1 U15730 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12615) );
  NOR4_X1 U15731 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12614) );
  INV_X1 U15732 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20684) );
  AND4_X1 U15733 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n20684), .ZN(
        n12617) );
  NAND2_X1 U15734 ( .A1(n12618), .A2(n12617), .ZN(n12619) );
  AND2_X2 U15735 ( .A1(n12619), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14642)
         );
  INV_X1 U15736 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20737) );
  NOR3_X1 U15737 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20737), .ZN(n12621) );
  NOR4_X1 U15738 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12620) );
  NAND4_X1 U15739 ( .A1(n14642), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12621), .A4(
        n12620), .ZN(U214) );
  NOR4_X1 U15740 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12625) );
  NOR4_X1 U15741 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12624) );
  NOR4_X1 U15742 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12623) );
  NOR4_X1 U15743 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12622) );
  NAND4_X1 U15744 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n12630) );
  NOR4_X1 U15745 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_7__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12628) );
  NOR4_X1 U15746 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12627) );
  NOR4_X1 U15747 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12626) );
  INV_X1 U15748 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19974) );
  NAND4_X1 U15749 ( .A1(n12628), .A2(n12627), .A3(n12626), .A4(n19974), .ZN(
        n12629) );
  OAI21_X1 U15750 ( .B1(n12630), .B2(n12629), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12631) );
  NOR2_X1 U15751 ( .A1(n15187), .A2(n12632), .ZN(n16555) );
  NAND2_X1 U15752 ( .A1(n16555), .A2(U214), .ZN(U212) );
  INV_X1 U15753 ( .A(n12633), .ZN(n15901) );
  OR2_X1 U15754 ( .A1(n14948), .A2(n15901), .ZN(n12636) );
  INV_X1 U15755 ( .A(n14413), .ZN(n20094) );
  NOR2_X1 U15756 ( .A1(n20094), .A2(n15930), .ZN(n12634) );
  AND2_X1 U15757 ( .A1(n15907), .A2(n12634), .ZN(n12635) );
  NAND2_X1 U15758 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16271) );
  NOR2_X1 U15759 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16271), .ZN(n20227) );
  NOR2_X4 U15760 ( .A1(n20205), .A2(n20748), .ZN(n20226) );
  AND2_X1 U15761 ( .A1(n20226), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OR3_X1 U15762 ( .A1(n12758), .A2(n13604), .A3(n12648), .ZN(n19233) );
  INV_X1 U15763 ( .A(n12637), .ZN(n12638) );
  NOR2_X1 U15764 ( .A1(n13604), .A2(n12648), .ZN(n12642) );
  AND2_X1 U15765 ( .A1(n12638), .A2(n12642), .ZN(n13333) );
  NOR2_X1 U15766 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15934) );
  NAND2_X1 U15767 ( .A1(n15934), .A2(n20037), .ZN(n18995) );
  INV_X1 U15768 ( .A(n18995), .ZN(n12639) );
  OR2_X1 U15769 ( .A1(n13333), .A2(n12639), .ZN(n12646) );
  AOI21_X1 U15770 ( .B1(P2_MEMORYFETCH_REG_SCAN_IN), .B2(n19233), .A(n12646), 
        .ZN(n12640) );
  INV_X1 U15771 ( .A(n12640), .ZN(P2_U2814) );
  INV_X1 U15772 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n12641) );
  NAND2_X1 U15773 ( .A1(n19233), .A2(n12641), .ZN(n12645) );
  NAND2_X1 U15774 ( .A1(n20074), .A2(n12643), .ZN(n12644) );
  OAI21_X1 U15775 ( .B1(n12646), .B2(n12645), .A(n12644), .ZN(n12647) );
  INV_X1 U15776 ( .A(n12647), .ZN(P2_U3612) );
  NOR2_X1 U15777 ( .A1(n13639), .A2(n12648), .ZN(n12649) );
  INV_X1 U15778 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19320) );
  NAND2_X1 U15779 ( .A1(n13333), .A2(n20756), .ZN(n12650) );
  NAND2_X1 U15780 ( .A1(n19381), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12652) );
  NAND3_X1 U15781 ( .A1(n13333), .A2(n13331), .A3(n20756), .ZN(n12724) );
  INV_X1 U15782 ( .A(n12724), .ZN(n19378) );
  AOI22_X1 U15783 ( .A1(n13840), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n15187), .ZN(n19262) );
  INV_X1 U15784 ( .A(n19262), .ZN(n12651) );
  NAND2_X1 U15785 ( .A1(n19378), .A2(n12651), .ZN(n12671) );
  OAI211_X1 U15786 ( .C1(n19306), .C2(n19320), .A(n12652), .B(n12671), .ZN(
        P2_U2964) );
  INV_X1 U15787 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19355) );
  NAND2_X1 U15788 ( .A1(n19381), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12655) );
  NAND2_X1 U15789 ( .A1(n15187), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12654) );
  INV_X1 U15790 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16583) );
  OR2_X1 U15791 ( .A1(n15187), .A2(n16583), .ZN(n12653) );
  NAND2_X1 U15792 ( .A1(n12654), .A2(n12653), .ZN(n19266) );
  NAND2_X1 U15793 ( .A1(n19378), .A2(n19266), .ZN(n12664) );
  OAI211_X1 U15794 ( .C1(n19355), .C2(n19306), .A(n12655), .B(n12664), .ZN(
        P2_U2977) );
  INV_X1 U15795 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19357) );
  NAND2_X1 U15796 ( .A1(n19381), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12658) );
  NAND2_X1 U15797 ( .A1(n15187), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12657) );
  INV_X1 U15798 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16585) );
  OR2_X1 U15799 ( .A1(n15187), .A2(n16585), .ZN(n12656) );
  NAND2_X1 U15800 ( .A1(n12657), .A2(n12656), .ZN(n19269) );
  NAND2_X1 U15801 ( .A1(n19378), .A2(n19269), .ZN(n12674) );
  OAI211_X1 U15802 ( .C1(n19357), .C2(n19306), .A(n12658), .B(n12674), .ZN(
        P2_U2976) );
  INV_X1 U15803 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n20903) );
  NAND2_X1 U15804 ( .A1(n19381), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12663) );
  INV_X1 U15805 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n12659) );
  OR2_X1 U15806 ( .A1(n15187), .A2(n12659), .ZN(n12661) );
  NAND2_X1 U15807 ( .A1(n15187), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12660) );
  AND2_X1 U15808 ( .A1(n12661), .A2(n12660), .ZN(n19260) );
  INV_X1 U15809 ( .A(n19260), .ZN(n12662) );
  NAND2_X1 U15810 ( .A1(n19378), .A2(n12662), .ZN(n12676) );
  OAI211_X1 U15811 ( .C1(n19306), .C2(n20903), .A(n12663), .B(n12676), .ZN(
        P2_U2965) );
  INV_X1 U15812 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19324) );
  NAND2_X1 U15813 ( .A1(n19381), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12665) );
  OAI211_X1 U15814 ( .C1(n19324), .C2(n19306), .A(n12665), .B(n12664), .ZN(
        P2_U2962) );
  INV_X1 U15815 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19322) );
  NAND2_X1 U15816 ( .A1(n19381), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12670) );
  INV_X1 U15817 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12666) );
  OR2_X1 U15818 ( .A1(n15187), .A2(n12666), .ZN(n12668) );
  NAND2_X1 U15819 ( .A1(n15187), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12667) );
  AND2_X1 U15820 ( .A1(n12668), .A2(n12667), .ZN(n19264) );
  INV_X1 U15821 ( .A(n19264), .ZN(n12669) );
  NAND2_X1 U15822 ( .A1(n19378), .A2(n12669), .ZN(n12720) );
  OAI211_X1 U15823 ( .C1(n19306), .C2(n19322), .A(n12670), .B(n12720), .ZN(
        P2_U2963) );
  INV_X1 U15824 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n12673) );
  NAND2_X1 U15825 ( .A1(n19381), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12672) );
  OAI211_X1 U15826 ( .C1(n19306), .C2(n12673), .A(n12672), .B(n12671), .ZN(
        P2_U2979) );
  INV_X1 U15827 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19326) );
  NAND2_X1 U15828 ( .A1(n19381), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12675) );
  OAI211_X1 U15829 ( .C1(n19306), .C2(n19326), .A(n12675), .B(n12674), .ZN(
        P2_U2961) );
  INV_X1 U15830 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n12678) );
  NAND2_X1 U15831 ( .A1(n19381), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n12677) );
  OAI211_X1 U15832 ( .C1(n19306), .C2(n12678), .A(n12677), .B(n12676), .ZN(
        P2_U2980) );
  INV_X1 U15833 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n12680) );
  OAI22_X1 U15834 ( .A1(n15187), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13840), .ZN(n15731) );
  NOR2_X1 U15835 ( .A1(n12724), .A2(n15731), .ZN(n12695) );
  AOI21_X1 U15836 ( .B1(n19380), .B2(P2_EAX_REG_20__SCAN_IN), .A(n12695), .ZN(
        n12679) );
  OAI21_X1 U15837 ( .B1(n12725), .B2(n12680), .A(n12679), .ZN(P2_U2956) );
  INV_X1 U15838 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15839 ( .A1(n13840), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15187), .ZN(n19410) );
  NOR2_X1 U15840 ( .A1(n12724), .A2(n19410), .ZN(n12692) );
  AOI21_X1 U15841 ( .B1(n19380), .B2(P2_EAX_REG_17__SCAN_IN), .A(n12692), .ZN(
        n12681) );
  OAI21_X1 U15842 ( .B1(n12725), .B2(n12682), .A(n12681), .ZN(P2_U2953) );
  INV_X1 U15843 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15844 ( .A1(n13840), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15187), .ZN(n19426) );
  NOR2_X1 U15845 ( .A1(n12724), .A2(n19426), .ZN(n12702) );
  AOI21_X1 U15846 ( .B1(n19380), .B2(P2_EAX_REG_6__SCAN_IN), .A(n12702), .ZN(
        n12683) );
  OAI21_X1 U15847 ( .B1(n12725), .B2(n12684), .A(n12683), .ZN(P2_U2973) );
  INV_X1 U15848 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15849 ( .A1(n13840), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15187), .ZN(n19277) );
  NOR2_X1 U15850 ( .A1(n12724), .A2(n19277), .ZN(n12707) );
  AOI21_X1 U15851 ( .B1(n19380), .B2(P2_EAX_REG_5__SCAN_IN), .A(n12707), .ZN(
        n12685) );
  OAI21_X1 U15852 ( .B1(n12725), .B2(n12686), .A(n12685), .ZN(P2_U2972) );
  INV_X1 U15853 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U15854 ( .A1(n13840), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15187), .ZN(n19272) );
  NOR2_X1 U15855 ( .A1(n12724), .A2(n19272), .ZN(n12689) );
  AOI21_X1 U15856 ( .B1(P2_EAX_REG_8__SCAN_IN), .B2(n19380), .A(n12689), .ZN(
        n12687) );
  OAI21_X1 U15857 ( .B1(n12725), .B2(n12688), .A(n12687), .ZN(P2_U2975) );
  INV_X1 U15858 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n12691) );
  AOI21_X1 U15859 ( .B1(n19380), .B2(P2_EAX_REG_24__SCAN_IN), .A(n12689), .ZN(
        n12690) );
  OAI21_X1 U15860 ( .B1(n12725), .B2(n12691), .A(n12690), .ZN(P2_U2960) );
  INV_X1 U15861 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n12694) );
  AOI21_X1 U15862 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n19380), .A(n12692), .ZN(
        n12693) );
  OAI21_X1 U15863 ( .B1(n12725), .B2(n12694), .A(n12693), .ZN(P2_U2968) );
  INV_X1 U15864 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n12697) );
  AOI21_X1 U15865 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n19380), .A(n12695), .ZN(
        n12696) );
  OAI21_X1 U15866 ( .B1(n12725), .B2(n12697), .A(n12696), .ZN(P2_U2971) );
  INV_X1 U15867 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15868 ( .A1(n13840), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15187), .ZN(n19422) );
  NOR2_X1 U15869 ( .A1(n12724), .A2(n19422), .ZN(n12716) );
  AOI21_X1 U15870 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n19380), .A(n12716), .ZN(
        n12698) );
  OAI21_X1 U15871 ( .B1(n12725), .B2(n12699), .A(n12698), .ZN(P2_U2970) );
  INV_X1 U15872 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15873 ( .A1(n13840), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15187), .ZN(n19433) );
  NOR2_X1 U15874 ( .A1(n12724), .A2(n19433), .ZN(n12710) );
  AOI21_X1 U15875 ( .B1(n19380), .B2(P2_EAX_REG_23__SCAN_IN), .A(n12710), .ZN(
        n12700) );
  OAI21_X1 U15876 ( .B1(n12725), .B2(n12701), .A(n12700), .ZN(P2_U2959) );
  INV_X1 U15877 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12704) );
  AOI21_X1 U15878 ( .B1(n19380), .B2(P2_EAX_REG_22__SCAN_IN), .A(n12702), .ZN(
        n12703) );
  OAI21_X1 U15879 ( .B1(n12725), .B2(n12704), .A(n12703), .ZN(P2_U2958) );
  INV_X1 U15880 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12706) );
  OAI22_X1 U15881 ( .A1(n15187), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13840), .ZN(n19415) );
  NOR2_X1 U15882 ( .A1(n12724), .A2(n19415), .ZN(n12713) );
  AOI21_X1 U15883 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n19380), .A(n12713), .ZN(
        n12705) );
  OAI21_X1 U15884 ( .B1(n12725), .B2(n12706), .A(n12705), .ZN(P2_U2969) );
  INV_X1 U15885 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12709) );
  AOI21_X1 U15886 ( .B1(n19380), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12707), .ZN(
        n12708) );
  OAI21_X1 U15887 ( .B1(n12725), .B2(n12709), .A(n12708), .ZN(P2_U2957) );
  INV_X1 U15888 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12712) );
  AOI21_X1 U15889 ( .B1(n19380), .B2(P2_EAX_REG_7__SCAN_IN), .A(n12710), .ZN(
        n12711) );
  OAI21_X1 U15890 ( .B1(n12725), .B2(n12712), .A(n12711), .ZN(P2_U2974) );
  INV_X1 U15891 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n12715) );
  AOI21_X1 U15892 ( .B1(n19380), .B2(P2_EAX_REG_18__SCAN_IN), .A(n12713), .ZN(
        n12714) );
  OAI21_X1 U15893 ( .B1(n12725), .B2(n12715), .A(n12714), .ZN(P2_U2954) );
  INV_X1 U15894 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12718) );
  AOI21_X1 U15895 ( .B1(n19380), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12716), .ZN(
        n12717) );
  OAI21_X1 U15896 ( .B1(n12725), .B2(n12718), .A(n12717), .ZN(P2_U2955) );
  INV_X1 U15897 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n12721) );
  NAND2_X1 U15898 ( .A1(n19380), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n12719) );
  OAI211_X1 U15899 ( .C1(n12725), .C2(n12721), .A(n12720), .B(n12719), .ZN(
        P2_U2978) );
  INV_X1 U15900 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n20917) );
  AOI22_X1 U15901 ( .A1(n13840), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15187), .ZN(n19255) );
  INV_X1 U15902 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19347) );
  OAI222_X1 U15903 ( .A1(n12725), .A2(n20917), .B1(n12724), .B2(n19255), .C1(
        n19306), .C2(n19347), .ZN(P2_U2982) );
  INV_X1 U15904 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12722) );
  INV_X1 U15905 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19345) );
  OAI22_X1 U15906 ( .A1(n15187), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13840), .ZN(n19244) );
  OAI222_X1 U15907 ( .A1(n12722), .A2(n12725), .B1(n19306), .B2(n19345), .C1(
        n19244), .C2(n12724), .ZN(P2_U2952) );
  INV_X1 U15908 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12726) );
  INV_X1 U15909 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12723) );
  OAI222_X1 U15910 ( .A1(n12726), .A2(n12725), .B1(n12724), .B2(n19244), .C1(
        n19306), .C2(n12723), .ZN(P2_U2967) );
  OR2_X1 U15911 ( .A1(n12727), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12728) );
  AND2_X1 U15912 ( .A1(n12729), .A2(n12728), .ZN(n16478) );
  XNOR2_X1 U15913 ( .A(n19229), .B(n20916), .ZN(n16476) );
  NAND2_X1 U15914 ( .A1(n11600), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16484) );
  OAI21_X1 U15915 ( .B1(n16425), .B2(n16476), .A(n16484), .ZN(n12730) );
  AOI21_X1 U15916 ( .B1(n16435), .B2(n16478), .A(n12730), .ZN(n12733) );
  OAI21_X1 U15917 ( .B1(n16409), .B2(n12731), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12732) );
  OAI211_X1 U15918 ( .C1(n16439), .C2(n12767), .A(n12733), .B(n12732), .ZN(
        P2_U3014) );
  AOI21_X1 U15919 ( .B1(n20922), .B2(n12735), .A(n12734), .ZN(n12820) );
  AND2_X1 U15920 ( .A1(n19180), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12814) );
  OAI21_X1 U15921 ( .B1(n12737), .B2(n15077), .A(n12736), .ZN(n12738) );
  XOR2_X1 U15922 ( .A(n12738), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n12817) );
  NOR2_X1 U15923 ( .A1(n12817), .A2(n16425), .ZN(n12739) );
  AOI211_X1 U15924 ( .C1(n16435), .C2(n12820), .A(n12814), .B(n12739), .ZN(
        n12741) );
  MUX2_X1 U15925 ( .A(n16424), .B(n16445), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n12740) );
  OAI211_X1 U15926 ( .C1(n16439), .C2(n15080), .A(n12741), .B(n12740), .ZN(
        P2_U3013) );
  NAND2_X1 U15927 ( .A1(n12742), .A2(n13643), .ZN(n12746) );
  INV_X1 U15928 ( .A(n12743), .ZN(n12744) );
  NAND3_X1 U15929 ( .A1(n11366), .A2(n12744), .A3(n11564), .ZN(n12745) );
  NAND2_X1 U15930 ( .A1(n12746), .A2(n12745), .ZN(n12777) );
  INV_X1 U15931 ( .A(n12747), .ZN(n12748) );
  NAND2_X1 U15932 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  NOR2_X1 U15933 ( .A1(n12777), .A2(n12750), .ZN(n12753) );
  NOR2_X1 U15934 ( .A1(n12751), .A2(n12758), .ZN(n19305) );
  NAND2_X1 U15935 ( .A1(n19305), .A2(n13608), .ZN(n12752) );
  NAND2_X1 U15936 ( .A1(n12753), .A2(n12752), .ZN(n13601) );
  INV_X1 U15937 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19950) );
  NOR2_X1 U15938 ( .A1(n19950), .A2(n12754), .ZN(n20072) );
  NAND2_X1 U15939 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20072), .ZN(n16486) );
  OAI22_X1 U15940 ( .A1(n16486), .A2(n19001), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n20037), .ZN(n12755) );
  AOI21_X1 U15941 ( .B1(n13601), .B2(n19304), .A(n12755), .ZN(n15725) );
  INV_X1 U15942 ( .A(n15725), .ZN(n12761) );
  INV_X1 U15943 ( .A(n12756), .ZN(n12757) );
  NOR3_X1 U15944 ( .A1(n12758), .A2(n12757), .A3(n13331), .ZN(n13611) );
  NAND3_X1 U15945 ( .A1(n12761), .A2(n15718), .A3(n13611), .ZN(n12759) );
  OAI21_X1 U15946 ( .B1(n12761), .B2(n12760), .A(n12759), .ZN(P2_U3595) );
  INV_X1 U15947 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12763) );
  NAND2_X1 U15948 ( .A1(n20037), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19949) );
  NOR2_X1 U15949 ( .A1(n10656), .A2(n19949), .ZN(n12762) );
  OAI21_X1 U15950 ( .B1(n11377), .B2(n12763), .A(n12762), .ZN(n12764) );
  INV_X1 U15951 ( .A(n12764), .ZN(n12765) );
  MUX2_X1 U15952 ( .A(n12767), .B(n10899), .S(n12766), .Z(n12768) );
  OAI21_X1 U15953 ( .B1(n20059), .B2(n15185), .A(n12768), .ZN(P2_U2887) );
  NAND2_X1 U15954 ( .A1(n20548), .A2(n20661), .ZN(n20097) );
  INV_X1 U15955 ( .A(n20097), .ZN(n12769) );
  NOR2_X1 U15956 ( .A1(n12769), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12772)
         );
  INV_X1 U15957 ( .A(n14406), .ZN(n12770) );
  NOR2_X1 U15958 ( .A1(n12166), .A2(n12770), .ZN(n14407) );
  NAND2_X1 U15959 ( .A1(n14407), .A2(n14413), .ZN(n14398) );
  OAI21_X1 U15960 ( .B1(n12181), .B2(n13438), .A(n20745), .ZN(n12771) );
  OAI21_X1 U15961 ( .B1(n12772), .B2(n20745), .A(n12771), .ZN(P1_U3487) );
  INV_X1 U15962 ( .A(n12773), .ZN(n12774) );
  AND2_X1 U15963 ( .A1(n12775), .A2(n12774), .ZN(n12776) );
  AND2_X1 U15964 ( .A1(n11375), .A2(n19431), .ZN(n12779) );
  NAND2_X1 U15965 ( .A1(n19275), .A2(n10669), .ZN(n13841) );
  NAND2_X1 U15966 ( .A1(n15250), .A2(n13841), .ZN(n19278) );
  INV_X1 U15967 ( .A(n12780), .ZN(n12786) );
  INV_X1 U15968 ( .A(n12781), .ZN(n12784) );
  INV_X1 U15969 ( .A(n12782), .ZN(n12783) );
  NAND2_X1 U15970 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  NAND2_X1 U15971 ( .A1(n12786), .A2(n12785), .ZN(n12787) );
  INV_X1 U15972 ( .A(n12787), .ZN(n19225) );
  NOR2_X1 U15973 ( .A1(n20059), .A2(n12787), .ZN(n19298) );
  INV_X1 U15974 ( .A(n19298), .ZN(n12789) );
  OAI211_X1 U15975 ( .C1(n19638), .C2(n19225), .A(n12789), .B(n19280), .ZN(
        n12792) );
  NAND2_X1 U15976 ( .A1(n19275), .A2(n12790), .ZN(n16349) );
  AOI22_X1 U15977 ( .A1(n19295), .A2(n19225), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19294), .ZN(n12791) );
  OAI211_X1 U15978 ( .C1(n19303), .C2(n19244), .A(n12792), .B(n12791), .ZN(
        P2_U2919) );
  NOR2_X1 U15979 ( .A1(n15080), .A2(n12766), .ZN(n12795) );
  AOI21_X1 U15980 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n12766), .A(n12795), .ZN(
        n12796) );
  OAI21_X1 U15981 ( .B1(n20050), .B2(n15185), .A(n12796), .ZN(P2_U2886) );
  INV_X1 U15982 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U15983 ( .A1(n20205), .A2(n9723), .ZN(n12907) );
  AOI22_X1 U15984 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12798) );
  OAI21_X1 U15985 ( .B1(n12799), .B2(n12907), .A(n12798), .ZN(P1_U2907) );
  INV_X1 U15986 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U15987 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12800) );
  OAI21_X1 U15988 ( .B1(n12801), .B2(n12907), .A(n12800), .ZN(P1_U2908) );
  INV_X1 U15989 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U15990 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12802) );
  OAI21_X1 U15991 ( .B1(n12803), .B2(n12907), .A(n12802), .ZN(P1_U2906) );
  INV_X1 U15992 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U15993 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12804) );
  OAI21_X1 U15994 ( .B1(n12805), .B2(n12907), .A(n12804), .ZN(P1_U2911) );
  INV_X1 U15995 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U15996 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12806) );
  OAI21_X1 U15997 ( .B1(n12807), .B2(n12907), .A(n12806), .ZN(P1_U2909) );
  INV_X1 U15998 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U15999 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12808) );
  OAI21_X1 U16000 ( .B1(n12809), .B2(n12907), .A(n12808), .ZN(P1_U2910) );
  INV_X1 U16001 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U16002 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12810) );
  OAI21_X1 U16003 ( .B1(n12811), .B2(n12907), .A(n12810), .ZN(P1_U2912) );
  OAI211_X1 U16004 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16479), .B(n19388), .ZN(n12816) );
  OAI21_X1 U16005 ( .B1(n12813), .B2(n12812), .A(n11393), .ZN(n20055) );
  AOI21_X1 U16006 ( .B1(n16474), .B2(n20055), .A(n12814), .ZN(n12815) );
  OAI211_X1 U16007 ( .C1(n19385), .C2(n20922), .A(n12816), .B(n12815), .ZN(
        n12819) );
  NOR2_X1 U16008 ( .A1(n12817), .A2(n16477), .ZN(n12818) );
  AOI211_X1 U16009 ( .C1(n12820), .C2(n19391), .A(n12819), .B(n12818), .ZN(
        n12821) );
  OAI21_X1 U16010 ( .B1(n15080), .B2(n19404), .A(n12821), .ZN(P2_U3045) );
  MUX2_X1 U16011 ( .A(n10769), .B(n12824), .S(n12766), .Z(n12825) );
  OAI21_X1 U16012 ( .B1(n20043), .B2(n15185), .A(n12825), .ZN(P2_U2885) );
  INV_X1 U16013 ( .A(n12826), .ZN(n12828) );
  NAND2_X1 U16014 ( .A1(n12828), .A2(n12827), .ZN(n12830) );
  NOR2_X1 U16015 ( .A1(n16438), .A2(n12766), .ZN(n12831) );
  AOI21_X1 U16016 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n12766), .A(n12831), .ZN(
        n12832) );
  OAI21_X1 U16017 ( .B1(n19672), .B2(n15185), .A(n12832), .ZN(P2_U2884) );
  OR2_X1 U16018 ( .A1(n12833), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12835) );
  AND2_X1 U16019 ( .A1(n12835), .A2(n12834), .ZN(n13465) );
  INV_X1 U16020 ( .A(n13465), .ZN(n12853) );
  NAND2_X1 U16021 ( .A1(n14403), .A2(n14408), .ZN(n12867) );
  NOR2_X1 U16022 ( .A1(n12863), .A2(n12836), .ZN(n13205) );
  INV_X1 U16023 ( .A(n13073), .ZN(n14351) );
  NAND4_X1 U16024 ( .A1(n12837), .A2(n13205), .A3(n14351), .A4(n11737), .ZN(
        n13068) );
  OR2_X1 U16025 ( .A1(n13068), .A2(n14410), .ZN(n12838) );
  NAND2_X1 U16026 ( .A1(n12867), .A2(n12838), .ZN(n12839) );
  NOR2_X2 U16027 ( .A1(n11737), .A2(n12842), .ZN(n14011) );
  NOR2_X1 U16028 ( .A1(n11797), .A2(n12842), .ZN(n13103) );
  INV_X1 U16029 ( .A(n13103), .ZN(n12846) );
  NAND2_X1 U16030 ( .A1(n14331), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12845) );
  NAND2_X1 U16031 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12844) );
  OAI211_X1 U16032 ( .C1(n12846), .C2(n11666), .A(n12845), .B(n12844), .ZN(
        n12847) );
  AOI21_X1 U16033 ( .B1(n12841), .B2(n14011), .A(n12847), .ZN(n12917) );
  NAND2_X1 U16034 ( .A1(n12848), .A2(n13671), .ZN(n12849) );
  NAND2_X1 U16035 ( .A1(n12849), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12851) );
  OR2_X1 U16036 ( .A1(n12851), .A2(n12917), .ZN(n12921) );
  INV_X1 U16037 ( .A(n12921), .ZN(n12850) );
  AOI21_X1 U16038 ( .B1(n12917), .B2(n12851), .A(n12850), .ZN(n12890) );
  INV_X1 U16039 ( .A(n12890), .ZN(n13472) );
  NAND2_X2 U16040 ( .A1(n20204), .A2(n13073), .ZN(n14624) );
  OAI222_X1 U16041 ( .A1(n12853), .A2(n20194), .B1(n12852), .B2(n20204), .C1(
        n13472), .C2(n14624), .ZN(P1_U2872) );
  OAI21_X1 U16042 ( .B1(n12855), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12854), .ZN(n12888) );
  NAND2_X1 U16043 ( .A1(n20177), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n12887) );
  INV_X1 U16044 ( .A(n12887), .ZN(n12857) );
  NOR2_X1 U16045 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12856), .ZN(
        n12990) );
  AOI211_X1 U16046 ( .C1(n16256), .C2(n13465), .A(n12857), .B(n12990), .ZN(
        n12859) );
  OAI21_X1 U16047 ( .B1(n14900), .B2(n12991), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12858) );
  OAI211_X1 U16048 ( .C1(n12888), .C2(n16259), .A(n12859), .B(n12858), .ZN(
        P1_U3031) );
  NAND4_X1 U16049 ( .A1(n12860), .A2(n20747), .A3(n12180), .A4(n15907), .ZN(
        n13067) );
  INV_X1 U16050 ( .A(n13067), .ZN(n12861) );
  NOR3_X1 U16051 ( .A1(n15930), .A2(n14408), .A3(n15929), .ZN(n15900) );
  OAI22_X1 U16052 ( .A1(n14948), .A2(n12862), .B1(n12861), .B2(n15900), .ZN(
        n12865) );
  OR2_X1 U16053 ( .A1(n13425), .A2(n12863), .ZN(n12864) );
  NAND4_X1 U16054 ( .A1(n12867), .A2(n12866), .A3(n12865), .A4(n12864), .ZN(
        n12870) );
  NAND2_X1 U16055 ( .A1(n12881), .A2(n13438), .ZN(n13207) );
  OR2_X1 U16056 ( .A1(n15881), .A2(n20094), .ZN(n12872) );
  NOR2_X1 U16057 ( .A1(n11886), .A2(n16271), .ZN(n13234) );
  NAND2_X1 U16058 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13234), .ZN(n12871) );
  AND2_X1 U16059 ( .A1(n12872), .A2(n12871), .ZN(n12875) );
  NAND2_X1 U16060 ( .A1(n11886), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n12873) );
  NAND2_X1 U16061 ( .A1(n12875), .A2(n12873), .ZN(n14966) );
  INV_X1 U16062 ( .A(n13343), .ZN(n13126) );
  NOR2_X1 U16063 ( .A1(n11921), .A2(n13126), .ZN(n12874) );
  XOR2_X1 U16064 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12874), .Z(
        n20172) );
  INV_X1 U16065 ( .A(n12875), .ZN(n12876) );
  NAND4_X1 U16066 ( .A1(n20172), .A2(n14949), .A3(n12171), .A4(n12876), .ZN(
        n12877) );
  OAI21_X1 U16067 ( .B1(n12878), .B2(n14966), .A(n12877), .ZN(P1_U3468) );
  NOR2_X1 U16068 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20661), .ZN(n20740) );
  NAND2_X1 U16069 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20740), .ZN(n16265) );
  INV_X1 U16070 ( .A(n16265), .ZN(n12879) );
  AND2_X2 U16071 ( .A1(n20548), .A2(n12879), .ZN(n16069) );
  OR2_X1 U16072 ( .A1(n12882), .A2(n20548), .ZN(n20746) );
  AND2_X1 U16073 ( .A1(n20746), .A2(n11886), .ZN(n12883) );
  INV_X1 U16074 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20453) );
  NAND2_X1 U16075 ( .A1(n20453), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12885) );
  NOR2_X1 U16076 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12842), .ZN(n20739) );
  INV_X1 U16077 ( .A(n20739), .ZN(n12884) );
  NAND2_X1 U16078 ( .A1(n12885), .A2(n12884), .ZN(n12910) );
  OAI21_X1 U16079 ( .B1(n16104), .B2(n12910), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12886) );
  OAI211_X1 U16080 ( .C1(n12888), .C2(n20100), .A(n12887), .B(n12886), .ZN(
        n12889) );
  AOI21_X1 U16081 ( .B1(n12890), .B2(n16069), .A(n12889), .ZN(n12891) );
  INV_X1 U16082 ( .A(n12891), .ZN(P1_U2999) );
  INV_X1 U16083 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U16084 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12892) );
  OAI21_X1 U16085 ( .B1(n12893), .B2(n12907), .A(n12892), .ZN(P1_U2917) );
  INV_X1 U16086 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U16087 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12894) );
  OAI21_X1 U16088 ( .B1(n12895), .B2(n12907), .A(n12894), .ZN(P1_U2920) );
  INV_X1 U16089 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U16090 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12896) );
  OAI21_X1 U16091 ( .B1(n12897), .B2(n12907), .A(n12896), .ZN(P1_U2915) );
  INV_X1 U16092 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16093 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12898) );
  OAI21_X1 U16094 ( .B1(n12899), .B2(n12907), .A(n12898), .ZN(P1_U2919) );
  INV_X1 U16095 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U16096 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12900) );
  OAI21_X1 U16097 ( .B1(n12901), .B2(n12907), .A(n12900), .ZN(P1_U2918) );
  INV_X1 U16098 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U16099 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12902) );
  OAI21_X1 U16100 ( .B1(n12903), .B2(n12907), .A(n12902), .ZN(P1_U2916) );
  INV_X1 U16101 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16102 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12904) );
  OAI21_X1 U16103 ( .B1(n12905), .B2(n12907), .A(n12904), .ZN(P1_U2913) );
  INV_X1 U16104 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16105 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12906) );
  OAI21_X1 U16106 ( .B1(n12908), .B2(n12907), .A(n12906), .ZN(P1_U2914) );
  XNOR2_X1 U16107 ( .A(n12909), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12999) );
  INV_X1 U16108 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U16109 ( .A1(n20177), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n12993) );
  OAI21_X1 U16110 ( .B1(n16120), .B2(n13446), .A(n12993), .ZN(n12925) );
  XNOR2_X2 U16111 ( .A(n12912), .B(n12911), .ZN(n13130) );
  NAND2_X1 U16112 ( .A1(n13130), .A2(n14011), .ZN(n12916) );
  INV_X1 U16113 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12913) );
  OAI22_X1 U16114 ( .A1(n14294), .A2(n12913), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13446), .ZN(n12914) );
  AOI21_X1 U16115 ( .B1(n13103), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12914), .ZN(n12915) );
  INV_X1 U16116 ( .A(n12917), .ZN(n12919) );
  NOR2_X1 U16117 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12918) );
  OR2_X1 U16118 ( .A1(n12919), .A2(n14303), .ZN(n12920) );
  NAND2_X1 U16119 ( .A1(n12921), .A2(n12920), .ZN(n12922) );
  NAND2_X1 U16120 ( .A1(n12923), .A2(n12922), .ZN(n13029) );
  OAI21_X1 U16121 ( .B1(n12923), .B2(n12922), .A(n13029), .ZN(n13427) );
  NOR2_X1 U16122 ( .A1(n13427), .A2(n14832), .ZN(n12924) );
  AOI211_X1 U16123 ( .C1(n16114), .C2(n13446), .A(n12925), .B(n12924), .ZN(
        n12926) );
  OAI21_X1 U16124 ( .B1(n12999), .B2(n20100), .A(n12926), .ZN(P1_U2998) );
  NAND2_X1 U16125 ( .A1(n12928), .A2(n12927), .ZN(n12931) );
  INV_X1 U16126 ( .A(n12929), .ZN(n12930) );
  AND2_X1 U16127 ( .A1(n12931), .A2(n12930), .ZN(n19399) );
  XNOR2_X1 U16128 ( .A(n20043), .B(n19399), .ZN(n12936) );
  INV_X1 U16129 ( .A(n20055), .ZN(n12932) );
  NAND2_X1 U16130 ( .A1(n20050), .A2(n12932), .ZN(n12933) );
  OAI21_X1 U16131 ( .B1(n20050), .B2(n12932), .A(n12933), .ZN(n19297) );
  NOR2_X1 U16132 ( .A1(n19297), .A2(n19298), .ZN(n19296) );
  INV_X1 U16133 ( .A(n12933), .ZN(n12934) );
  NOR2_X1 U16134 ( .A1(n19296), .A2(n12934), .ZN(n12935) );
  NOR2_X1 U16135 ( .A1(n12935), .A2(n12936), .ZN(n13179) );
  AOI21_X1 U16136 ( .B1(n12936), .B2(n12935), .A(n13179), .ZN(n12939) );
  INV_X1 U16137 ( .A(n19415), .ZN(n16347) );
  AOI22_X1 U16138 ( .A1(n19278), .A2(n16347), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19294), .ZN(n12938) );
  INV_X1 U16139 ( .A(n19399), .ZN(n20045) );
  NAND2_X1 U16140 ( .A1(n20045), .A2(n19295), .ZN(n12937) );
  OAI211_X1 U16141 ( .C1(n12939), .C2(n19299), .A(n12938), .B(n12937), .ZN(
        P2_U2917) );
  AND2_X1 U16142 ( .A1(n11818), .A2(n15929), .ZN(n12940) );
  INV_X2 U16143 ( .A(n12975), .ZN(n20259) );
  NAND2_X1 U16144 ( .A1(n14353), .A2(DATAI_2_), .ZN(n12942) );
  NAND2_X1 U16145 ( .A1(n14642), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12941) );
  AND2_X1 U16146 ( .A1(n12942), .A2(n12941), .ZN(n13157) );
  INV_X1 U16147 ( .A(n13157), .ZN(n14700) );
  NAND2_X1 U16148 ( .A1(n20244), .A2(n14700), .ZN(n13018) );
  AND2_X2 U16149 ( .A1(n12975), .A2(n11809), .ZN(n20254) );
  AOI22_X1 U16150 ( .A1(n20254), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U16151 ( .A1(n13018), .A2(n12943), .ZN(P1_U2954) );
  NAND2_X1 U16152 ( .A1(n14353), .A2(DATAI_4_), .ZN(n12945) );
  NAND2_X1 U16153 ( .A1(n14642), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12944) );
  AND2_X1 U16154 ( .A1(n12945), .A2(n12944), .ZN(n13677) );
  INV_X1 U16155 ( .A(n13677), .ZN(n14687) );
  NAND2_X1 U16156 ( .A1(n20244), .A2(n14687), .ZN(n13013) );
  AOI22_X1 U16157 ( .A1(n20254), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n12946) );
  NAND2_X1 U16158 ( .A1(n13013), .A2(n12946), .ZN(P1_U2956) );
  NAND2_X1 U16159 ( .A1(n14353), .A2(DATAI_3_), .ZN(n12948) );
  NAND2_X1 U16160 ( .A1(n14642), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12947) );
  AND2_X1 U16161 ( .A1(n12948), .A2(n12947), .ZN(n13143) );
  INV_X1 U16162 ( .A(n13143), .ZN(n14693) );
  NAND2_X1 U16163 ( .A1(n20244), .A2(n14693), .ZN(n13011) );
  AOI22_X1 U16164 ( .A1(n20254), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n12949) );
  NAND2_X1 U16165 ( .A1(n13011), .A2(n12949), .ZN(P1_U2955) );
  NAND2_X1 U16166 ( .A1(n14353), .A2(DATAI_7_), .ZN(n12951) );
  NAND2_X1 U16167 ( .A1(n14642), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12950) );
  AND2_X1 U16168 ( .A1(n12951), .A2(n12950), .ZN(n13526) );
  INV_X1 U16169 ( .A(n13526), .ZN(n14670) );
  NAND2_X1 U16170 ( .A1(n20244), .A2(n14670), .ZN(n13009) );
  AOI22_X1 U16171 ( .A1(n20254), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n12952) );
  NAND2_X1 U16172 ( .A1(n13009), .A2(n12952), .ZN(P1_U2959) );
  NAND2_X1 U16173 ( .A1(n14353), .A2(DATAI_5_), .ZN(n12954) );
  NAND2_X1 U16174 ( .A1(n14642), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12953) );
  AND2_X1 U16175 ( .A1(n12954), .A2(n12953), .ZN(n13259) );
  INV_X1 U16176 ( .A(n13259), .ZN(n14681) );
  NAND2_X1 U16177 ( .A1(n20244), .A2(n14681), .ZN(n13005) );
  AOI22_X1 U16178 ( .A1(n20254), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n12955) );
  NAND2_X1 U16179 ( .A1(n13005), .A2(n12955), .ZN(P1_U2957) );
  NAND2_X1 U16180 ( .A1(n14353), .A2(DATAI_6_), .ZN(n12957) );
  NAND2_X1 U16181 ( .A1(n14642), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12956) );
  AND2_X1 U16182 ( .A1(n12957), .A2(n12956), .ZN(n13670) );
  INV_X1 U16183 ( .A(n13670), .ZN(n14676) );
  NAND2_X1 U16184 ( .A1(n20244), .A2(n14676), .ZN(n13020) );
  AOI22_X1 U16185 ( .A1(n20254), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n12958) );
  NAND2_X1 U16186 ( .A1(n13020), .A2(n12958), .ZN(P1_U2958) );
  INV_X1 U16187 ( .A(n12841), .ZN(n13462) );
  AND3_X1 U16188 ( .A1(n12112), .A2(n12960), .A3(n12959), .ZN(n12961) );
  AND3_X1 U16189 ( .A1(n12962), .A2(n12961), .A3(n9907), .ZN(n14945) );
  OAI22_X1 U16190 ( .A1(n13462), .A2(n14945), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14944), .ZN(n15880) );
  INV_X1 U16191 ( .A(n14957), .ZN(n14962) );
  OAI22_X1 U16192 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20661), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14962), .ZN(n12963) );
  AOI21_X1 U16193 ( .B1(n15880), .B2(n14949), .A(n12963), .ZN(n12967) );
  INV_X1 U16194 ( .A(n14966), .ZN(n12966) );
  AND2_X1 U16195 ( .A1(n14948), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15879) );
  NAND2_X1 U16196 ( .A1(n15879), .A2(n14949), .ZN(n12965) );
  NAND2_X1 U16197 ( .A1(n12966), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12964) );
  OAI211_X1 U16198 ( .C1(n12967), .C2(n12966), .A(n12965), .B(n12964), .ZN(
        P1_U3474) );
  XNOR2_X1 U16199 ( .A(n12968), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12972) );
  OR2_X1 U16200 ( .A1(n12969), .A2(n12985), .ZN(n12970) );
  NAND2_X1 U16201 ( .A1(n13055), .A2(n12970), .ZN(n19169) );
  MUX2_X1 U16202 ( .A(n19168), .B(n19169), .S(n15159), .Z(n12971) );
  OAI21_X1 U16203 ( .B1(n12972), .B2(n15185), .A(n12971), .ZN(P2_U2880) );
  INV_X1 U16204 ( .A(n20254), .ZN(n13002) );
  INV_X1 U16205 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12978) );
  INV_X1 U16206 ( .A(n20244), .ZN(n12977) );
  INV_X1 U16207 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12973) );
  NOR2_X1 U16208 ( .A1(n14353), .A2(n12973), .ZN(n12974) );
  AOI21_X1 U16209 ( .B1(DATAI_15_), .B2(n14353), .A(n12974), .ZN(n14721) );
  INV_X1 U16210 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12976) );
  OAI222_X1 U16211 ( .A1(n13002), .A2(n12978), .B1(n12977), .B2(n14721), .C1(
        n12976), .C2(n12975), .ZN(P1_U2967) );
  OR2_X1 U16212 ( .A1(n12979), .A2(n13463), .ZN(n12980) );
  NAND2_X1 U16213 ( .A1(n13455), .A2(n12980), .ZN(n12995) );
  INV_X1 U16214 ( .A(n20204), .ZN(n14615) );
  AOI22_X1 U16215 ( .A1(n20199), .A2(n12995), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14615), .ZN(n12981) );
  OAI21_X1 U16216 ( .B1(n13427), .B2(n14624), .A(n12981), .ZN(P1_U2871) );
  NOR2_X1 U16217 ( .A1(n12982), .A2(n13669), .ZN(n12984) );
  INV_X1 U16218 ( .A(n12968), .ZN(n12983) );
  OAI211_X1 U16219 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n12984), .A(
        n12983), .B(n15149), .ZN(n12988) );
  AOI21_X1 U16220 ( .B1(n12986), .B2(n13779), .A(n12985), .ZN(n19184) );
  NAND2_X1 U16221 ( .A1(n19184), .A2(n15159), .ZN(n12987) );
  OAI211_X1 U16222 ( .C1(n15159), .C2(n12989), .A(n12988), .B(n12987), .ZN(
        P2_U2881) );
  OAI21_X1 U16223 ( .B1(n12991), .B2(n12990), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U16224 ( .A1(n12993), .A2(n12992), .ZN(n12994) );
  AOI21_X1 U16225 ( .B1(n16256), .B2(n12995), .A(n12994), .ZN(n12998) );
  OAI211_X1 U16226 ( .C1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n14900), .A(
        n14910), .B(n12996), .ZN(n12997) );
  OAI211_X1 U16227 ( .C1(n12999), .C2(n16259), .A(n12998), .B(n12997), .ZN(
        P1_U3030) );
  NAND2_X1 U16228 ( .A1(n14353), .A2(DATAI_1_), .ZN(n13001) );
  NAND2_X1 U16229 ( .A1(n14642), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13000) );
  AND2_X1 U16230 ( .A1(n13001), .A2(n13000), .ZN(n13131) );
  INV_X1 U16231 ( .A(n13131), .ZN(n14707) );
  NAND2_X1 U16232 ( .A1(n20244), .A2(n14707), .ZN(n13007) );
  AOI22_X1 U16233 ( .A1(n20254), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U16234 ( .A1(n13007), .A2(n13003), .ZN(P1_U2953) );
  AOI22_X1 U16235 ( .A1(n20254), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13004) );
  NAND2_X1 U16236 ( .A1(n13005), .A2(n13004), .ZN(P1_U2942) );
  AOI22_X1 U16237 ( .A1(n20254), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13006) );
  NAND2_X1 U16238 ( .A1(n13007), .A2(n13006), .ZN(P1_U2938) );
  AOI22_X1 U16239 ( .A1(n20254), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13008) );
  NAND2_X1 U16240 ( .A1(n13009), .A2(n13008), .ZN(P1_U2944) );
  AOI22_X1 U16241 ( .A1(n20254), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13010) );
  NAND2_X1 U16242 ( .A1(n13011), .A2(n13010), .ZN(P1_U2940) );
  AOI22_X1 U16243 ( .A1(n20254), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13012) );
  NAND2_X1 U16244 ( .A1(n13013), .A2(n13012), .ZN(P1_U2941) );
  NAND2_X1 U16245 ( .A1(n14353), .A2(DATAI_0_), .ZN(n13015) );
  NAND2_X1 U16246 ( .A1(n14642), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13014) );
  AND2_X1 U16247 ( .A1(n13015), .A2(n13014), .ZN(n13151) );
  INV_X1 U16248 ( .A(n13151), .ZN(n14714) );
  NAND2_X1 U16249 ( .A1(n20244), .A2(n14714), .ZN(n13022) );
  AOI22_X1 U16250 ( .A1(n20254), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U16251 ( .A1(n13022), .A2(n13016), .ZN(P1_U2937) );
  AOI22_X1 U16252 ( .A1(n20254), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U16253 ( .A1(n13018), .A2(n13017), .ZN(P1_U2939) );
  AOI22_X1 U16254 ( .A1(n20254), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16255 ( .A1(n13020), .A2(n13019), .ZN(P1_U2943) );
  AOI22_X1 U16256 ( .A1(n20254), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13021) );
  NAND2_X1 U16257 ( .A1(n13022), .A2(n13021), .ZN(P1_U2952) );
  INV_X1 U16258 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13024) );
  XNOR2_X1 U16259 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13694) );
  AOI21_X1 U16260 ( .B1(n14188), .B2(n13694), .A(n14330), .ZN(n13023) );
  OAI21_X1 U16261 ( .B1(n14294), .B2(n13024), .A(n13023), .ZN(n13025) );
  AOI21_X1 U16262 ( .B1(n13103), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13025), .ZN(n13026) );
  NAND2_X1 U16263 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  NAND2_X1 U16264 ( .A1(n14330), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13081) );
  NAND2_X1 U16265 ( .A1(n13028), .A2(n13081), .ZN(n13033) );
  INV_X1 U16266 ( .A(n13082), .ZN(n13032) );
  AOI21_X1 U16267 ( .B1(n13033), .B2(n13029), .A(n13032), .ZN(n13691) );
  INV_X1 U16268 ( .A(n13691), .ZN(n13078) );
  NAND2_X1 U16269 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  AND2_X1 U16270 ( .A1(n13095), .A2(n13036), .ZN(n13692) );
  AOI22_X1 U16271 ( .A1(n20199), .A2(n13692), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14615), .ZN(n13037) );
  OAI21_X1 U16272 ( .B1(n13078), .B2(n14624), .A(n13037), .ZN(P1_U2870) );
  XNOR2_X1 U16273 ( .A(n13039), .B(n13038), .ZN(n13053) );
  AOI22_X1 U16274 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20177), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13040) );
  OAI21_X1 U16275 ( .B1(n16111), .B2(n13694), .A(n13040), .ZN(n13041) );
  AOI21_X1 U16276 ( .B1(n13691), .B2(n16069), .A(n13041), .ZN(n13042) );
  OAI21_X1 U16277 ( .B1(n20100), .B2(n13053), .A(n13042), .ZN(P1_U2997) );
  NOR2_X1 U16278 ( .A1(n13046), .A2(n12996), .ZN(n13043) );
  OAI21_X1 U16279 ( .B1(n13901), .B2(n13043), .A(n14919), .ZN(n16208) );
  NOR2_X1 U16280 ( .A1(n20984), .A2(n12996), .ZN(n13044) );
  AOI21_X1 U16281 ( .B1(n13044), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13171), .ZN(n13050) );
  AOI21_X1 U16282 ( .B1(n20984), .B2(n13045), .A(n13901), .ZN(n14884) );
  NAND3_X1 U16283 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14884), .A3(
        n13046), .ZN(n13049) );
  INV_X1 U16284 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13566) );
  NOR2_X1 U16285 ( .A1(n9736), .A2(n13566), .ZN(n13047) );
  AOI21_X1 U16286 ( .B1(n16256), .B2(n13692), .A(n13047), .ZN(n13048) );
  OAI211_X1 U16287 ( .C1(n13050), .C2(n14920), .A(n13049), .B(n13048), .ZN(
        n13051) );
  AOI21_X1 U16288 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n16208), .A(
        n13051), .ZN(n13052) );
  OAI21_X1 U16289 ( .B1(n16259), .B2(n13053), .A(n13052), .ZN(P1_U3029) );
  AND2_X1 U16290 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  OR2_X1 U16291 ( .A1(n13062), .A2(n13056), .ZN(n19158) );
  OAI211_X1 U16292 ( .C1(n10218), .C2(n10226), .A(n15149), .B(n13057), .ZN(
        n13059) );
  NAND2_X1 U16293 ( .A1(n12766), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13058) );
  OAI211_X1 U16294 ( .C1(n19158), .C2(n12766), .A(n13059), .B(n13058), .ZN(
        P2_U2879) );
  XOR2_X1 U16295 ( .A(n13057), .B(n13117), .Z(n13066) );
  OR2_X1 U16296 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  AND2_X1 U16297 ( .A1(n13060), .A2(n13063), .ZN(n19145) );
  NOR2_X1 U16298 ( .A1(n15159), .A2(n11021), .ZN(n13064) );
  AOI21_X1 U16299 ( .B1(n19145), .B2(n15159), .A(n13064), .ZN(n13065) );
  OAI21_X1 U16300 ( .B1(n13066), .B2(n15185), .A(n13065), .ZN(P2_U2878) );
  OAI21_X1 U16301 ( .B1(n13068), .B2(n14411), .A(n13067), .ZN(n13069) );
  NAND2_X1 U16302 ( .A1(n11804), .A2(n13073), .ZN(n13072) );
  NAND2_X1 U16303 ( .A1(n13139), .A2(n13073), .ZN(n13074) );
  INV_X1 U16304 ( .A(n13075), .ZN(n13077) );
  INV_X1 U16305 ( .A(n14354), .ZN(n13076) );
  OAI222_X1 U16306 ( .A1(n9731), .A2(n13427), .B1(n13131), .B2(n14722), .C1(
        n16046), .C2(n12913), .ZN(P1_U2903) );
  INV_X1 U16307 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20230) );
  OAI222_X1 U16308 ( .A1(n9731), .A2(n13472), .B1(n13151), .B2(n14722), .C1(
        n16046), .C2(n20230), .ZN(P1_U2904) );
  OAI222_X1 U16309 ( .A1(n9731), .A2(n13078), .B1(n13157), .B2(n14722), .C1(
        n16046), .C2(n13024), .ZN(P1_U2902) );
  XNOR2_X1 U16310 ( .A(n13080), .B(n13079), .ZN(n13245) );
  INV_X1 U16311 ( .A(n14011), .ZN(n13971) );
  INV_X1 U16312 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13085) );
  OAI21_X1 U16313 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13083), .A(
        n13249), .ZN(n13529) );
  AOI22_X1 U16314 ( .A1(n14188), .A2(n13529), .B1(n14330), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13084) );
  OAI21_X1 U16315 ( .B1(n14294), .B2(n13085), .A(n13084), .ZN(n13086) );
  AOI21_X1 U16316 ( .B1(n13103), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13086), .ZN(n13087) );
  NOR2_X1 U16317 ( .A1(n13088), .A2(n13089), .ZN(n13090) );
  NOR2_X1 U16318 ( .A1(n13109), .A2(n13090), .ZN(n13527) );
  NAND2_X1 U16319 ( .A1(n20177), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13242) );
  NAND2_X1 U16320 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13091) );
  OAI211_X1 U16321 ( .C1(n16111), .C2(n13529), .A(n13242), .B(n13091), .ZN(
        n13092) );
  AOI21_X1 U16322 ( .B1(n13527), .B2(n16069), .A(n13092), .ZN(n13093) );
  OAI21_X1 U16323 ( .B1(n13245), .B2(n20100), .A(n13093), .ZN(P1_U2996) );
  INV_X1 U16324 ( .A(n13527), .ZN(n13098) );
  INV_X1 U16325 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13531) );
  AND2_X1 U16326 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  NOR2_X1 U16327 ( .A1(n13111), .A2(n13096), .ZN(n13535) );
  INV_X1 U16328 ( .A(n13535), .ZN(n13097) );
  OAI222_X1 U16329 ( .A1(n13098), .A2(n14624), .B1(n13531), .B2(n20204), .C1(
        n13097), .C2(n20194), .ZN(P1_U2869) );
  OAI222_X1 U16330 ( .A1(n9731), .A2(n13098), .B1(n13143), .B2(n14722), .C1(
        n16046), .C2(n13085), .ZN(P1_U2901) );
  NAND2_X1 U16331 ( .A1(n13099), .A2(n14011), .ZN(n13107) );
  INV_X1 U16332 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13100) );
  XNOR2_X1 U16333 ( .A(n13249), .B(n13100), .ZN(n20187) );
  INV_X1 U16334 ( .A(n20187), .ZN(n13105) );
  INV_X1 U16335 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13101) );
  OAI22_X1 U16336 ( .A1(n14294), .A2(n13101), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13100), .ZN(n13102) );
  AOI21_X1 U16337 ( .B1(n13103), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13102), .ZN(n13104) );
  MUX2_X1 U16338 ( .A(n13105), .B(n13104), .S(n14303), .Z(n13106) );
  NAND2_X1 U16339 ( .A1(n13107), .A2(n13106), .ZN(n13108) );
  NAND2_X1 U16340 ( .A1(n13109), .A2(n13108), .ZN(n13246) );
  OAI21_X1 U16341 ( .B1(n13109), .B2(n13108), .A(n13246), .ZN(n13190) );
  OAI222_X1 U16342 ( .A1(n9731), .A2(n13190), .B1(n13677), .B2(n14722), .C1(
        n16046), .C2(n13101), .ZN(P1_U2900) );
  OR2_X1 U16343 ( .A1(n13111), .A2(n13110), .ZN(n13112) );
  NAND2_X1 U16344 ( .A1(n16252), .A2(n13112), .ZN(n20174) );
  INV_X1 U16345 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13113) );
  OAI222_X1 U16346 ( .A1(n20174), .A2(n20194), .B1(n20204), .B2(n13113), .C1(
        n13190), .C2(n14624), .ZN(P1_U2868) );
  INV_X1 U16347 ( .A(n13060), .ZN(n13115) );
  OAI21_X1 U16348 ( .B1(n13115), .B2(n10229), .A(n13114), .ZN(n19132) );
  INV_X1 U16349 ( .A(n13116), .ZN(n13121) );
  INV_X1 U16350 ( .A(n13117), .ZN(n13119) );
  OAI21_X1 U16351 ( .B1(n13057), .B2(n13119), .A(n13118), .ZN(n13120) );
  NAND3_X1 U16352 ( .A1(n13121), .A2(n15149), .A3(n13120), .ZN(n13123) );
  NAND2_X1 U16353 ( .A1(n12766), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13122) );
  OAI211_X1 U16354 ( .C1(n19132), .C2(n12766), .A(n13123), .B(n13122), .ZN(
        P2_U2877) );
  NAND2_X1 U16355 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20598) );
  NOR2_X1 U16356 ( .A1(n20598), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13132) );
  NAND2_X1 U16357 ( .A1(n9769), .A2(n13124), .ZN(n20606) );
  NOR2_X1 U16358 ( .A1(n13125), .A2(n13126), .ZN(n20597) );
  INV_X1 U16359 ( .A(n13127), .ZN(n20450) );
  NOR3_X2 U16360 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20449), .A3(
        n20598), .ZN(n13719) );
  AOI21_X1 U16361 ( .B1(n20597), .B2(n20450), .A(n13719), .ZN(n13134) );
  OAI211_X1 U16362 ( .C1(n20606), .C2(n20453), .A(n20548), .B(n13134), .ZN(
        n13128) );
  OAI211_X1 U16363 ( .C1(n20548), .C2(n13132), .A(n20607), .B(n13128), .ZN(
        n13129) );
  INV_X1 U16364 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13138) );
  OR2_X1 U16365 ( .A1(n13130), .A2(n12848), .ZN(n20447) );
  NOR2_X2 U16366 ( .A1(n20606), .A2(n20447), .ZN(n13718) );
  NAND2_X1 U16367 ( .A1(n16069), .A2(n14642), .ZN(n13155) );
  NAND2_X1 U16368 ( .A1(n14353), .A2(n16069), .ZN(n13156) );
  AOI22_X1 U16369 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n13682), .B1(DATAI_17_), 
        .B2(n13681), .ZN(n20619) );
  INV_X1 U16370 ( .A(n20619), .ZN(n20563) );
  OR2_X1 U16371 ( .A1(n20606), .A2(n20394), .ZN(n20547) );
  AOI22_X1 U16372 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n13682), .B1(DATAI_25_), 
        .B2(n13681), .ZN(n20566) );
  INV_X1 U16373 ( .A(n20566), .ZN(n20616) );
  AOI22_X1 U16374 ( .A1(n13718), .A2(n20563), .B1(n20588), .B2(n20616), .ZN(
        n13137) );
  NOR2_X2 U16375 ( .A1(n13131), .A2(n13676), .ZN(n20615) );
  INV_X1 U16376 ( .A(n13132), .ZN(n13133) );
  OAI22_X1 U16377 ( .A1(n13134), .A2(n20601), .B1(n13133), .B2(n12842), .ZN(
        n13720) );
  NOR2_X2 U16378 ( .A1(n13680), .A2(n11809), .ZN(n20614) );
  AOI22_X1 U16379 ( .A1(n20615), .A2(n13720), .B1(n20614), .B2(n13719), .ZN(
        n13136) );
  OAI211_X1 U16380 ( .C1(n13724), .C2(n13138), .A(n13137), .B(n13136), .ZN(
        P1_U3138) );
  INV_X1 U16381 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U16382 ( .A1(DATAI_21_), .A2(n13681), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n13682), .ZN(n20643) );
  INV_X1 U16383 ( .A(n20643), .ZN(n20579) );
  AOI22_X1 U16384 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13682), .B1(DATAI_29_), 
        .B2(n13681), .ZN(n20582) );
  INV_X1 U16385 ( .A(n20582), .ZN(n20640) );
  AOI22_X1 U16386 ( .A1(n13718), .A2(n20579), .B1(n20588), .B2(n20640), .ZN(
        n13141) );
  NOR2_X2 U16387 ( .A1(n13259), .A2(n13676), .ZN(n20639) );
  NOR2_X2 U16388 ( .A1(n13680), .A2(n13139), .ZN(n20638) );
  AOI22_X1 U16389 ( .A1(n20639), .A2(n13720), .B1(n20638), .B2(n13719), .ZN(
        n13140) );
  OAI211_X1 U16390 ( .C1(n13724), .C2(n13142), .A(n13141), .B(n13140), .ZN(
        P1_U3142) );
  INV_X1 U16391 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U16392 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n13682), .B1(DATAI_19_), 
        .B2(n13681), .ZN(n20631) );
  INV_X1 U16393 ( .A(n20631), .ZN(n20571) );
  AOI22_X1 U16394 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13682), .B1(DATAI_27_), 
        .B2(n13681), .ZN(n20574) );
  INV_X1 U16395 ( .A(n20574), .ZN(n20628) );
  AOI22_X1 U16396 ( .A1(n13718), .A2(n20571), .B1(n20588), .B2(n20628), .ZN(
        n13146) );
  NOR2_X2 U16397 ( .A1(n13143), .A2(n13676), .ZN(n20627) );
  NOR2_X2 U16398 ( .A1(n13680), .A2(n13144), .ZN(n20626) );
  AOI22_X1 U16399 ( .A1(n20627), .A2(n13720), .B1(n20626), .B2(n13719), .ZN(
        n13145) );
  OAI211_X1 U16400 ( .C1(n13724), .C2(n13147), .A(n13146), .B(n13145), .ZN(
        P1_U3140) );
  INV_X1 U16401 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U16402 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n13682), .B1(DATAI_23_), 
        .B2(n13681), .ZN(n20660) );
  INV_X1 U16403 ( .A(n20660), .ZN(n20587) );
  AOI22_X1 U16404 ( .A1(DATAI_31_), .A2(n13681), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n13682), .ZN(n20594) );
  INV_X1 U16405 ( .A(n20594), .ZN(n20654) );
  AOI22_X1 U16406 ( .A1(n13718), .A2(n20587), .B1(n20588), .B2(n20654), .ZN(
        n13149) );
  NOR2_X2 U16407 ( .A1(n13526), .A2(n13676), .ZN(n20653) );
  NOR2_X2 U16408 ( .A1(n13680), .A2(n14351), .ZN(n20651) );
  AOI22_X1 U16409 ( .A1(n20653), .A2(n13720), .B1(n20651), .B2(n13719), .ZN(
        n13148) );
  OAI211_X1 U16410 ( .C1(n13724), .C2(n13150), .A(n13149), .B(n13148), .ZN(
        P1_U3144) );
  INV_X1 U16411 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U16412 ( .A1(DATAI_16_), .A2(n13681), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n13682), .ZN(n20613) );
  INV_X1 U16413 ( .A(n20613), .ZN(n20546) );
  AOI22_X1 U16414 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13682), .B1(DATAI_24_), 
        .B2(n13681), .ZN(n20562) );
  INV_X1 U16415 ( .A(n20562), .ZN(n20610) );
  AOI22_X1 U16416 ( .A1(n13718), .A2(n20546), .B1(n20588), .B2(n20610), .ZN(
        n13153) );
  NOR2_X2 U16417 ( .A1(n13151), .A2(n13676), .ZN(n20604) );
  NOR2_X2 U16418 ( .A1(n13680), .A2(n13449), .ZN(n20603) );
  AOI22_X1 U16419 ( .A1(n20604), .A2(n13720), .B1(n20603), .B2(n13719), .ZN(
        n13152) );
  OAI211_X1 U16420 ( .C1(n13724), .C2(n13154), .A(n13153), .B(n13152), .ZN(
        P1_U3137) );
  INV_X1 U16421 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13161) );
  INV_X1 U16422 ( .A(DATAI_18_), .ZN(n20954) );
  OAI22_X1 U16423 ( .A1(n20954), .A2(n13156), .B1(n14703), .B2(n13155), .ZN(
        n20567) );
  AOI22_X1 U16424 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n13682), .B1(DATAI_26_), 
        .B2(n13681), .ZN(n20570) );
  INV_X1 U16425 ( .A(n20570), .ZN(n20622) );
  AOI22_X1 U16426 ( .A1(n13718), .A2(n20567), .B1(n20588), .B2(n20622), .ZN(
        n13160) );
  NOR2_X2 U16427 ( .A1(n13157), .A2(n13676), .ZN(n20621) );
  NOR2_X2 U16428 ( .A1(n13680), .A2(n13158), .ZN(n20620) );
  AOI22_X1 U16429 ( .A1(n20621), .A2(n13720), .B1(n20620), .B2(n13719), .ZN(
        n13159) );
  OAI211_X1 U16430 ( .C1(n13724), .C2(n13161), .A(n13160), .B(n13159), .ZN(
        P1_U3139) );
  XNOR2_X1 U16431 ( .A(n13116), .B(n13199), .ZN(n13166) );
  NAND2_X1 U16432 ( .A1(n13114), .A2(n13162), .ZN(n13163) );
  AND2_X1 U16433 ( .A1(n13197), .A2(n13163), .ZN(n19121) );
  NOR2_X1 U16434 ( .A1(n15159), .A2(n19113), .ZN(n13164) );
  AOI21_X1 U16435 ( .B1(n19121), .B2(n15159), .A(n13164), .ZN(n13165) );
  OAI21_X1 U16436 ( .B1(n13166), .B2(n15185), .A(n13165), .ZN(P2_U2876) );
  XNOR2_X1 U16437 ( .A(n13168), .B(n13167), .ZN(n13195) );
  AOI21_X1 U16438 ( .B1(n14885), .B2(n13171), .A(n16208), .ZN(n13169) );
  INV_X1 U16439 ( .A(n13169), .ZN(n13240) );
  INV_X1 U16440 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20683) );
  NOR2_X1 U16441 ( .A1(n9736), .A2(n20683), .ZN(n13191) );
  NOR2_X1 U16442 ( .A1(n20174), .A2(n16220), .ZN(n13170) );
  AOI211_X1 U16443 ( .C1(n13240), .C2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13191), .B(n13170), .ZN(n13173) );
  NAND3_X1 U16444 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14884), .ZN(n14926) );
  OAI211_X1 U16445 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n16250), .B(n13825), .ZN(n13172) );
  OAI211_X1 U16446 ( .C1(n16259), .C2(n13195), .A(n13173), .B(n13172), .ZN(
        P1_U3027) );
  INV_X1 U16447 ( .A(n13174), .ZN(n13175) );
  NAND2_X1 U16448 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  OAI21_X1 U16449 ( .B1(n13178), .B2(n13177), .A(n12982), .ZN(n19216) );
  AOI21_X1 U16450 ( .B1(n19399), .B2(n20043), .A(n13179), .ZN(n19290) );
  OR2_X1 U16451 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  NAND2_X1 U16452 ( .A1(n13182), .A2(n13184), .ZN(n20038) );
  XNOR2_X1 U16453 ( .A(n19672), .B(n20038), .ZN(n19289) );
  NOR2_X1 U16454 ( .A1(n19290), .A2(n19289), .ZN(n19288) );
  INV_X1 U16455 ( .A(n19672), .ZN(n20034) );
  INV_X1 U16456 ( .A(n20038), .ZN(n19287) );
  NOR2_X1 U16457 ( .A1(n20034), .A2(n19287), .ZN(n13185) );
  XNOR2_X1 U16458 ( .A(n13184), .B(n13183), .ZN(n19212) );
  OAI21_X1 U16459 ( .B1(n19288), .B2(n13185), .A(n19212), .ZN(n19282) );
  XOR2_X1 U16460 ( .A(n19216), .B(n19282), .Z(n13189) );
  INV_X1 U16461 ( .A(n19212), .ZN(n13186) );
  AOI22_X1 U16462 ( .A1(n19295), .A2(n13186), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19294), .ZN(n13188) );
  INV_X1 U16463 ( .A(n15731), .ZN(n16342) );
  NAND2_X1 U16464 ( .A1(n19278), .A2(n16342), .ZN(n13187) );
  OAI211_X1 U16465 ( .C1(n13189), .C2(n19299), .A(n13188), .B(n13187), .ZN(
        P2_U2915) );
  INV_X1 U16466 ( .A(n13190), .ZN(n20183) );
  AOI21_X1 U16467 ( .B1(n16104), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13191), .ZN(n13192) );
  OAI21_X1 U16468 ( .B1(n16111), .B2(n20187), .A(n13192), .ZN(n13193) );
  AOI21_X1 U16469 ( .B1(n20183), .B2(n16069), .A(n13193), .ZN(n13194) );
  OAI21_X1 U16470 ( .B1(n13195), .B2(n20100), .A(n13194), .ZN(P1_U2995) );
  AND2_X1 U16471 ( .A1(n13197), .A2(n13196), .ZN(n13198) );
  OR2_X1 U16472 ( .A1(n13198), .A2(n13421), .ZN(n13325) );
  AND2_X1 U16473 ( .A1(n13116), .A2(n13199), .ZN(n13202) );
  OAI211_X1 U16474 ( .C1(n13202), .C2(n13201), .A(n15149), .B(n13200), .ZN(
        n13204) );
  NAND2_X1 U16475 ( .A1(n12766), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13203) );
  OAI211_X1 U16476 ( .C1(n13325), .C2(n12766), .A(n13204), .B(n13203), .ZN(
        P2_U2875) );
  NOR2_X1 U16477 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20661), .ZN(n13232) );
  INV_X1 U16478 ( .A(n13125), .ZN(n20270) );
  INV_X1 U16479 ( .A(n14945), .ZN(n13225) );
  NAND2_X1 U16480 ( .A1(n14945), .A2(n13205), .ZN(n13223) );
  XNOR2_X1 U16481 ( .A(n13206), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14953) );
  INV_X1 U16482 ( .A(n14403), .ZN(n13208) );
  NAND2_X1 U16483 ( .A1(n13208), .A2(n13207), .ZN(n13218) );
  XNOR2_X1 U16484 ( .A(n11892), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13209) );
  AOI22_X1 U16485 ( .A1(n13218), .A2(n14953), .B1(n14948), .B2(n13209), .ZN(
        n13210) );
  OAI21_X1 U16486 ( .B1(n13223), .B2(n14953), .A(n13210), .ZN(n13211) );
  AOI21_X1 U16487 ( .B1(n20270), .B2(n13225), .A(n13211), .ZN(n14960) );
  INV_X1 U16488 ( .A(n14960), .ZN(n13212) );
  MUX2_X1 U16489 ( .A(n13212), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15881), .Z(n15886) );
  AOI22_X1 U16490 ( .A1(n13232), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15886), .B2(n20661), .ZN(n13228) );
  INV_X1 U16491 ( .A(n13206), .ZN(n13214) );
  OAI21_X1 U16492 ( .B1(n13214), .B2(n13213), .A(n9985), .ZN(n13215) );
  NAND2_X1 U16493 ( .A1(n13215), .A2(n9751), .ZN(n14963) );
  MUX2_X1 U16494 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13220), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13216) );
  OAI21_X1 U16495 ( .B1(n13217), .B2(n13216), .A(n14948), .ZN(n13222) );
  MUX2_X1 U16496 ( .A(n13217), .B(n9985), .S(n13206), .Z(n13219) );
  OAI21_X1 U16497 ( .B1(n13220), .B2(n13219), .A(n13218), .ZN(n13221) );
  OAI211_X1 U16498 ( .C1(n13223), .C2(n14963), .A(n13222), .B(n13221), .ZN(
        n13224) );
  AOI21_X1 U16499 ( .B1(n20271), .B2(n13225), .A(n13224), .ZN(n14965) );
  INV_X1 U16500 ( .A(n14965), .ZN(n13226) );
  MUX2_X1 U16501 ( .A(n13226), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15881), .Z(n15890) );
  AOI22_X1 U16502 ( .A1(n13232), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20661), .B2(n15890), .ZN(n13227) );
  NOR2_X1 U16503 ( .A1(n13228), .A2(n13227), .ZN(n15896) );
  INV_X1 U16504 ( .A(n15896), .ZN(n13233) );
  AOI21_X1 U16505 ( .B1(n20172), .B2(n12171), .A(n15881), .ZN(n13230) );
  AOI211_X1 U16506 ( .C1(n15881), .C2(n12878), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n13230), .ZN(n13231) );
  AOI21_X1 U16507 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13232), .A(
        n13231), .ZN(n15898) );
  OAI21_X1 U16508 ( .B1(n13233), .B2(n13229), .A(n15898), .ZN(n13236) );
  OAI21_X1 U16509 ( .B1(n13236), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13234), .ZN(
        n13235) );
  NAND2_X1 U16510 ( .A1(n13235), .A2(n13676), .ZN(n20262) );
  NOR2_X1 U16511 ( .A1(n13236), .A2(n16271), .ZN(n15903) );
  NOR2_X1 U16512 ( .A1(n20661), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14942) );
  OAI22_X1 U16513 ( .A1(n12848), .A2(n20601), .B1(n13462), .B2(n14942), .ZN(
        n13237) );
  OAI21_X1 U16514 ( .B1(n15903), .B2(n13237), .A(n20262), .ZN(n13238) );
  OAI21_X1 U16515 ( .B1(n20262), .B2(n20449), .A(n13238), .ZN(P1_U3478) );
  AOI22_X1 U16516 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13240), .B1(
        n16250), .B2(n13239), .ZN(n13241) );
  NAND2_X1 U16517 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  AOI21_X1 U16518 ( .B1(n13535), .B2(n16256), .A(n13243), .ZN(n13244) );
  OAI21_X1 U16519 ( .B1(n13245), .B2(n16259), .A(n13244), .ZN(P1_U3028) );
  INV_X1 U16520 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13258) );
  INV_X1 U16521 ( .A(n13249), .ZN(n13247) );
  AOI21_X1 U16522 ( .B1(n13247), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13250) );
  OR2_X1 U16523 ( .A1(n13250), .A2(n13507), .ZN(n20168) );
  AOI22_X1 U16524 ( .A1(n20168), .A2(n14188), .B1(n14330), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13251) );
  OAI21_X1 U16525 ( .B1(n14294), .B2(n13258), .A(n13251), .ZN(n13252) );
  NAND2_X1 U16526 ( .A1(n13246), .A2(n13256), .ZN(n13257) );
  AND2_X1 U16527 ( .A1(n13514), .A2(n13257), .ZN(n20201) );
  INV_X1 U16528 ( .A(n20201), .ZN(n13260) );
  OAI222_X1 U16529 ( .A1(n13260), .A2(n9731), .B1(n13259), .B2(n14722), .C1(
        n13258), .C2(n16046), .ZN(P1_U2899) );
  INV_X1 U16530 ( .A(n20262), .ZN(n13268) );
  INV_X1 U16531 ( .A(n20512), .ZN(n20520) );
  MUX2_X1 U16532 ( .A(n20606), .B(n20423), .S(n13130), .Z(n13262) );
  NAND3_X1 U16533 ( .A1(n20520), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n13262), 
        .ZN(n13265) );
  AOI21_X1 U16534 ( .B1(n20268), .B2(n20453), .A(n20601), .ZN(n13264) );
  INV_X1 U16535 ( .A(n14942), .ZN(n13263) );
  AOI22_X1 U16536 ( .A1(n13265), .A2(n13264), .B1(n13263), .B2(n20271), .ZN(
        n13267) );
  NAND2_X1 U16537 ( .A1(n13268), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13266) );
  OAI21_X1 U16538 ( .B1(n13268), .B2(n13267), .A(n13266), .ZN(P1_U3475) );
  XNOR2_X1 U16539 ( .A(n13270), .B(n13269), .ZN(n13271) );
  XNOR2_X1 U16540 ( .A(n13272), .B(n13271), .ZN(n16442) );
  INV_X1 U16541 ( .A(n13273), .ZN(n13275) );
  MUX2_X1 U16542 ( .A(n13275), .B(n13274), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13277) );
  INV_X1 U16543 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19975) );
  AOI22_X1 U16544 ( .A1(n16474), .A2(n19287), .B1(n19180), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n13276) );
  OAI211_X1 U16545 ( .C1(n16438), .C2(n19404), .A(n13277), .B(n13276), .ZN(
        n13282) );
  OR2_X1 U16546 ( .A1(n13280), .A2(n13279), .ZN(n16436) );
  AND3_X1 U16547 ( .A1(n13278), .A2(n16436), .A3(n19391), .ZN(n13281) );
  AOI211_X1 U16548 ( .C1(n16442), .C2(n19395), .A(n13282), .B(n13281), .ZN(
        n13283) );
  INV_X1 U16549 ( .A(n13283), .ZN(P2_U3043) );
  NAND2_X1 U16550 ( .A1(n13130), .A2(n12848), .ZN(n20477) );
  NOR2_X2 U16551 ( .A1(n20606), .A2(n20477), .ZN(n20655) );
  OAI21_X1 U16552 ( .B1(n20655), .B2(n13718), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13286) );
  NAND2_X1 U16553 ( .A1(n20597), .A2(n11887), .ZN(n13285) );
  AOI21_X1 U16554 ( .B1(n13286), .B2(n13285), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n13288) );
  OR2_X1 U16555 ( .A1(n13290), .A2(n12842), .ZN(n20485) );
  INV_X1 U16556 ( .A(n20485), .ZN(n13287) );
  NAND2_X1 U16557 ( .A1(n20264), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20486) );
  NAND2_X1 U16558 ( .A1(n20486), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20481) );
  OAI211_X1 U16559 ( .C1(n13712), .C2(n13288), .A(n20553), .B(n20481), .ZN(
        n13289) );
  INV_X1 U16560 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U16561 ( .A1(n20655), .A2(n20587), .B1(n13718), .B2(n20654), .ZN(
        n13293) );
  NAND2_X1 U16562 ( .A1(n13290), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20557) );
  NAND3_X1 U16563 ( .A1(n20597), .A2(n11887), .A3(n20548), .ZN(n13291) );
  OAI21_X1 U16564 ( .B1(n20557), .B2(n20486), .A(n13291), .ZN(n13713) );
  AOI22_X1 U16565 ( .A1(n20653), .A2(n13713), .B1(n20651), .B2(n13712), .ZN(
        n13292) );
  OAI211_X1 U16566 ( .C1(n13717), .C2(n13294), .A(n13293), .B(n13292), .ZN(
        P1_U3152) );
  INV_X1 U16567 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16568 ( .A1(n20655), .A2(n20546), .B1(n13718), .B2(n20610), .ZN(
        n13296) );
  AOI22_X1 U16569 ( .A1(n20604), .A2(n13713), .B1(n20603), .B2(n13712), .ZN(
        n13295) );
  OAI211_X1 U16570 ( .C1(n13717), .C2(n13297), .A(n13296), .B(n13295), .ZN(
        P1_U3145) );
  INV_X1 U16571 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16572 ( .A1(n20655), .A2(n20579), .B1(n13718), .B2(n20640), .ZN(
        n13299) );
  AOI22_X1 U16573 ( .A1(n20639), .A2(n13713), .B1(n20638), .B2(n13712), .ZN(
        n13298) );
  OAI211_X1 U16574 ( .C1(n13717), .C2(n13300), .A(n13299), .B(n13298), .ZN(
        P1_U3150) );
  INV_X1 U16575 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13303) );
  AOI22_X1 U16576 ( .A1(n20655), .A2(n20563), .B1(n13718), .B2(n20616), .ZN(
        n13302) );
  AOI22_X1 U16577 ( .A1(n20615), .A2(n13713), .B1(n20614), .B2(n13712), .ZN(
        n13301) );
  OAI211_X1 U16578 ( .C1(n13717), .C2(n13303), .A(n13302), .B(n13301), .ZN(
        P1_U3146) );
  INV_X1 U16579 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U16580 ( .A1(n20655), .A2(n20567), .B1(n13718), .B2(n20622), .ZN(
        n13305) );
  AOI22_X1 U16581 ( .A1(n20621), .A2(n13713), .B1(n20620), .B2(n13712), .ZN(
        n13304) );
  OAI211_X1 U16582 ( .C1(n13717), .C2(n13306), .A(n13305), .B(n13304), .ZN(
        P1_U3147) );
  INV_X1 U16583 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U16584 ( .A1(n20655), .A2(n20571), .B1(n13718), .B2(n20628), .ZN(
        n13308) );
  AOI22_X1 U16585 ( .A1(n20627), .A2(n13713), .B1(n20626), .B2(n13712), .ZN(
        n13307) );
  OAI211_X1 U16586 ( .C1(n13717), .C2(n13309), .A(n13308), .B(n13307), .ZN(
        P1_U3148) );
  NOR2_X1 U16587 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13310), .ZN(n13637) );
  NOR2_X1 U16588 ( .A1(n13312), .A2(n13311), .ZN(n15614) );
  AOI21_X1 U16589 ( .B1(n13311), .B2(n13312), .A(n15614), .ZN(n15632) );
  INV_X1 U16590 ( .A(n15632), .ZN(n19263) );
  AOI21_X1 U16591 ( .B1(n19114), .B2(n13321), .A(n9840), .ZN(n19120) );
  AOI21_X1 U16592 ( .B1(n19139), .B2(n13319), .A(n13322), .ZN(n19144) );
  AOI21_X1 U16593 ( .B1(n15396), .B2(n13317), .A(n13320), .ZN(n19164) );
  AOI21_X1 U16594 ( .B1(n16432), .B2(n13315), .A(n13318), .ZN(n19191) );
  AOI21_X1 U16595 ( .B1(n16446), .B2(n13314), .A(n13316), .ZN(n16433) );
  OAI22_X1 U16596 ( .A1(n19309), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19240) );
  INV_X1 U16597 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15073) );
  OAI22_X1 U16598 ( .A1(n19309), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15073), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15072) );
  AND2_X1 U16599 ( .A1(n19240), .A2(n15072), .ZN(n15059) );
  OAI21_X1 U16600 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13314), .ZN(n15061) );
  NAND2_X1 U16601 ( .A1(n15059), .A2(n15061), .ZN(n15049) );
  NOR2_X1 U16602 ( .A1(n16433), .A2(n15049), .ZN(n19205) );
  OAI21_X1 U16603 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13316), .A(
        n13315), .ZN(n19207) );
  NAND2_X1 U16604 ( .A1(n19205), .A2(n19207), .ZN(n19189) );
  NOR2_X1 U16605 ( .A1(n19191), .A2(n19189), .ZN(n19181) );
  OAI21_X1 U16606 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13318), .A(
        n13317), .ZN(n19182) );
  NAND2_X1 U16607 ( .A1(n19181), .A2(n19182), .ZN(n19163) );
  NOR2_X1 U16608 ( .A1(n19164), .A2(n19163), .ZN(n19151) );
  OAI21_X1 U16609 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13320), .A(
        n13319), .ZN(n19152) );
  NAND2_X1 U16610 ( .A1(n19151), .A2(n19152), .ZN(n19142) );
  NOR2_X1 U16611 ( .A1(n19144), .A2(n19142), .ZN(n19125) );
  OAI21_X1 U16612 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13322), .A(
        n13321), .ZN(n19126) );
  NAND2_X1 U16613 ( .A1(n19125), .A2(n19126), .ZN(n19118) );
  NOR2_X1 U16614 ( .A1(n19120), .A2(n19118), .ZN(n14984) );
  NOR2_X1 U16615 ( .A1(n19206), .A2(n14984), .ZN(n13323) );
  OAI21_X1 U16616 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9840), .A(
        n14983), .ZN(n16400) );
  XNOR2_X1 U16617 ( .A(n13323), .B(n16400), .ZN(n13324) );
  NAND4_X1 U16618 ( .A1(n12754), .A2(n19309), .A3(n19770), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19955) );
  INV_X1 U16619 ( .A(n19955), .ZN(n19185) );
  NAND2_X1 U16620 ( .A1(n13324), .A2(n19185), .ZN(n13341) );
  INV_X1 U16621 ( .A(n13325), .ZN(n16397) );
  NAND2_X1 U16622 ( .A1(n20074), .A2(n10688), .ZN(n13327) );
  NAND2_X1 U16623 ( .A1(n19770), .A2(n20756), .ZN(n13329) );
  NAND2_X1 U16624 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13329), .ZN(n13326) );
  NOR2_X1 U16625 ( .A1(n13328), .A2(n19228), .ZN(n13339) );
  INV_X1 U16626 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15084) );
  NAND2_X1 U16627 ( .A1(n13329), .A2(n15084), .ZN(n13330) );
  AOI21_X1 U16628 ( .B1(n13331), .B2(n13330), .A(n13637), .ZN(n13332) );
  INV_X1 U16629 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13337) );
  OR4_X1 U16630 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), 
        .A3(n19309), .A4(n20037), .ZN(n13645) );
  NAND2_X1 U16631 ( .A1(n19955), .A2(n13645), .ZN(n13334) );
  OR2_X1 U16632 ( .A1(n19180), .A2(n13334), .ZN(n13335) );
  NAND2_X1 U16633 ( .A1(n19178), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19174) );
  AOI22_X1 U16634 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19223), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19236), .ZN(n13336) );
  OAI211_X1 U16635 ( .C1(n19197), .C2(n13337), .A(n13336), .B(n15581), .ZN(
        n13338) );
  AOI211_X1 U16636 ( .C1(n16397), .C2(n16282), .A(n13339), .B(n13338), .ZN(
        n13340) );
  OAI211_X1 U16637 ( .C1(n19213), .C2(n19263), .A(n13341), .B(n13340), .ZN(
        P2_U2843) );
  NAND2_X1 U16638 ( .A1(n13683), .A2(n20548), .ZN(n13342) );
  NAND2_X1 U16639 ( .A1(n20548), .A2(n20453), .ZN(n20549) );
  OAI21_X1 U16640 ( .B1(n20442), .B2(n13342), .A(n20549), .ZN(n13347) );
  OR2_X1 U16641 ( .A1(n13125), .A2(n13343), .ZN(n20393) );
  NOR2_X1 U16642 ( .A1(n20393), .A2(n20551), .ZN(n13345) );
  INV_X1 U16643 ( .A(n20557), .ZN(n13344) );
  INV_X1 U16644 ( .A(n20264), .ZN(n13399) );
  NOR2_X1 U16645 ( .A1(n13399), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20334) );
  AOI22_X1 U16646 ( .A1(n13347), .A2(n13345), .B1(n13344), .B2(n20334), .ZN(
        n13690) );
  INV_X1 U16647 ( .A(n20604), .ZN(n13352) );
  OR2_X1 U16648 ( .A1(n20599), .A2(n20419), .ZN(n13486) );
  NOR2_X1 U16649 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13486), .ZN(
        n13686) );
  INV_X1 U16650 ( .A(n13345), .ZN(n13346) );
  NOR2_X1 U16651 ( .A1(n20334), .A2(n12842), .ZN(n20330) );
  AOI21_X1 U16652 ( .B1(n13347), .B2(n13346), .A(n20330), .ZN(n13348) );
  OAI211_X1 U16653 ( .C1(n13686), .C2(n20554), .A(n20553), .B(n13348), .ZN(
        n13678) );
  NAND2_X1 U16654 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13351) );
  INV_X1 U16655 ( .A(n20442), .ZN(n13684) );
  OAI22_X1 U16656 ( .A1(n13684), .A2(n20562), .B1(n20613), .B2(n13683), .ZN(
        n13349) );
  AOI21_X1 U16657 ( .B1(n13686), .B2(n20603), .A(n13349), .ZN(n13350) );
  OAI211_X1 U16658 ( .C1(n13690), .C2(n13352), .A(n13351), .B(n13350), .ZN(
        P1_U3081) );
  INV_X1 U16659 ( .A(n20627), .ZN(n13356) );
  NAND2_X1 U16660 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13355) );
  OAI22_X1 U16661 ( .A1(n13684), .A2(n20574), .B1(n20631), .B2(n13683), .ZN(
        n13353) );
  AOI21_X1 U16662 ( .B1(n13686), .B2(n20626), .A(n13353), .ZN(n13354) );
  OAI211_X1 U16663 ( .C1(n13690), .C2(n13356), .A(n13355), .B(n13354), .ZN(
        P1_U3084) );
  INV_X1 U16664 ( .A(n20621), .ZN(n13360) );
  NAND2_X1 U16665 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13359) );
  INV_X1 U16666 ( .A(n20567), .ZN(n20625) );
  OAI22_X1 U16667 ( .A1(n13684), .A2(n20570), .B1(n13683), .B2(n20625), .ZN(
        n13357) );
  AOI21_X1 U16668 ( .B1(n13686), .B2(n20620), .A(n13357), .ZN(n13358) );
  OAI211_X1 U16669 ( .C1(n13690), .C2(n13360), .A(n13359), .B(n13358), .ZN(
        P1_U3083) );
  INV_X1 U16670 ( .A(n20615), .ZN(n13364) );
  NAND2_X1 U16671 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13363) );
  OAI22_X1 U16672 ( .A1(n13684), .A2(n20566), .B1(n20619), .B2(n13683), .ZN(
        n13361) );
  AOI21_X1 U16673 ( .B1(n13686), .B2(n20614), .A(n13361), .ZN(n13362) );
  OAI211_X1 U16674 ( .C1(n13690), .C2(n13364), .A(n13363), .B(n13362), .ZN(
        P1_U3082) );
  INV_X1 U16675 ( .A(n20639), .ZN(n13368) );
  NAND2_X1 U16676 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13367) );
  OAI22_X1 U16677 ( .A1(n13684), .A2(n20582), .B1(n20643), .B2(n13683), .ZN(
        n13365) );
  AOI21_X1 U16678 ( .B1(n13686), .B2(n20638), .A(n13365), .ZN(n13366) );
  OAI211_X1 U16679 ( .C1(n13690), .C2(n13368), .A(n13367), .B(n13366), .ZN(
        P1_U3086) );
  INV_X1 U16680 ( .A(n20653), .ZN(n13372) );
  NAND2_X1 U16681 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13371) );
  OAI22_X1 U16682 ( .A1(n13684), .A2(n20594), .B1(n20660), .B2(n13683), .ZN(
        n13369) );
  AOI21_X1 U16683 ( .B1(n13686), .B2(n20651), .A(n13369), .ZN(n13370) );
  OAI211_X1 U16684 ( .C1(n13690), .C2(n13372), .A(n13371), .B(n13370), .ZN(
        P1_U3088) );
  XNOR2_X1 U16685 ( .A(n13374), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13375) );
  XNOR2_X1 U16686 ( .A(n13373), .B(n13375), .ZN(n13392) );
  NAND3_X1 U16687 ( .A1(n13376), .A2(n13384), .A3(n16441), .ZN(n13383) );
  INV_X1 U16688 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19976) );
  OAI22_X1 U16689 ( .A1(n19976), .A2(n19210), .B1(n16424), .B2(n19207), .ZN(
        n13381) );
  AOI21_X1 U16690 ( .B1(n13379), .B2(n13378), .A(n13777), .ZN(n19217) );
  INV_X1 U16691 ( .A(n19217), .ZN(n14376) );
  NOR2_X1 U16692 ( .A1(n14376), .A2(n16439), .ZN(n13380) );
  AOI211_X1 U16693 ( .C1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n16409), .A(
        n13381), .B(n13380), .ZN(n13382) );
  OAI211_X1 U16694 ( .C1(n13392), .C2(n16427), .A(n13383), .B(n13382), .ZN(
        P2_U3010) );
  NAND3_X1 U16695 ( .A1(n13376), .A2(n13384), .A3(n19395), .ZN(n13391) );
  NOR2_X1 U16696 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13782), .ZN(
        n13386) );
  NOR2_X1 U16697 ( .A1(n19976), .A2(n19210), .ZN(n13385) );
  AOI211_X1 U16698 ( .C1(n13387), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13386), .B(n13385), .ZN(n13388) );
  OAI21_X1 U16699 ( .B1(n19400), .B2(n19212), .A(n13388), .ZN(n13389) );
  AOI21_X1 U16700 ( .B1(n19217), .B2(n16475), .A(n13389), .ZN(n13390) );
  OAI211_X1 U16701 ( .C1(n13392), .C2(n15702), .A(n13391), .B(n13390), .ZN(
        P2_U3042) );
  NAND2_X1 U16702 ( .A1(n20272), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20514) );
  NAND2_X1 U16703 ( .A1(n13393), .A2(n20557), .ZN(n20329) );
  INV_X1 U16704 ( .A(n20329), .ZN(n20480) );
  INV_X1 U16705 ( .A(n20394), .ZN(n13394) );
  NOR2_X2 U16706 ( .A1(n20423), .A2(n20510), .ZN(n13757) );
  OAI21_X1 U16707 ( .B1(n20473), .B2(n13757), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13396) );
  AND2_X1 U16708 ( .A1(n20271), .A2(n13125), .ZN(n20515) );
  AOI21_X1 U16709 ( .B1(n20515), .B2(n20551), .A(n10216), .ZN(n13400) );
  NAND2_X1 U16710 ( .A1(n13396), .A2(n13400), .ZN(n13397) );
  OAI211_X1 U16711 ( .C1(n10216), .C2(n20554), .A(n20480), .B(n13397), .ZN(
        n13398) );
  INV_X1 U16712 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16713 ( .A1(n20473), .A2(n20587), .B1(n13757), .B2(n20654), .ZN(
        n13402) );
  NAND2_X1 U16714 ( .A1(n13399), .A2(n20265), .ZN(n20556) );
  OAI22_X1 U16715 ( .A1(n13400), .A2(n20601), .B1(n20485), .B2(n20556), .ZN(
        n13725) );
  AOI22_X1 U16716 ( .A1(n20653), .A2(n13725), .B1(n20651), .B2(n10216), .ZN(
        n13401) );
  OAI211_X1 U16717 ( .C1(n13729), .C2(n13403), .A(n13402), .B(n13401), .ZN(
        P1_U3104) );
  INV_X1 U16718 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U16719 ( .A1(n20473), .A2(n20563), .B1(n13757), .B2(n20616), .ZN(
        n13405) );
  AOI22_X1 U16720 ( .A1(n20615), .A2(n13725), .B1(n20614), .B2(n10216), .ZN(
        n13404) );
  OAI211_X1 U16721 ( .C1(n13729), .C2(n13406), .A(n13405), .B(n13404), .ZN(
        P1_U3098) );
  INV_X1 U16722 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U16723 ( .A1(n20473), .A2(n20546), .B1(n13757), .B2(n20610), .ZN(
        n13408) );
  AOI22_X1 U16724 ( .A1(n20604), .A2(n13725), .B1(n20603), .B2(n10216), .ZN(
        n13407) );
  OAI211_X1 U16725 ( .C1(n13729), .C2(n13409), .A(n13408), .B(n13407), .ZN(
        P1_U3097) );
  INV_X1 U16726 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U16727 ( .A1(n20473), .A2(n20579), .B1(n13757), .B2(n20640), .ZN(
        n13411) );
  AOI22_X1 U16728 ( .A1(n20639), .A2(n13725), .B1(n20638), .B2(n10216), .ZN(
        n13410) );
  OAI211_X1 U16729 ( .C1(n13729), .C2(n13412), .A(n13411), .B(n13410), .ZN(
        P1_U3102) );
  INV_X1 U16730 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U16731 ( .A1(n20473), .A2(n20567), .B1(n13757), .B2(n20622), .ZN(
        n13414) );
  AOI22_X1 U16732 ( .A1(n20621), .A2(n13725), .B1(n20620), .B2(n10216), .ZN(
        n13413) );
  OAI211_X1 U16733 ( .C1(n13729), .C2(n13415), .A(n13414), .B(n13413), .ZN(
        P1_U3099) );
  INV_X1 U16734 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U16735 ( .A1(n20473), .A2(n20571), .B1(n13757), .B2(n20628), .ZN(
        n13417) );
  AOI22_X1 U16736 ( .A1(n20627), .A2(n13725), .B1(n20626), .B2(n10216), .ZN(
        n13416) );
  OAI211_X1 U16737 ( .C1(n13729), .C2(n13418), .A(n13417), .B(n13416), .ZN(
        P1_U3100) );
  XNOR2_X1 U16738 ( .A(n13200), .B(n13474), .ZN(n13424) );
  NOR2_X1 U16739 ( .A1(n13421), .A2(n13420), .ZN(n13422) );
  OR2_X1 U16740 ( .A1(n13419), .A2(n13422), .ZN(n16389) );
  MUX2_X1 U16741 ( .A(n16389), .B(n11293), .S(n12766), .Z(n13423) );
  OAI21_X1 U16742 ( .B1(n13424), .B2(n15185), .A(n13423), .ZN(P2_U2874) );
  INV_X1 U16743 ( .A(n13425), .ZN(n13426) );
  NAND2_X1 U16744 ( .A1(n20745), .A2(n13426), .ZN(n20169) );
  INV_X1 U16745 ( .A(n13427), .ZN(n13440) );
  NOR3_X1 U16746 ( .A1(n20554), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16268) );
  INV_X1 U16747 ( .A(n16268), .ZN(n15910) );
  NOR2_X1 U16748 ( .A1(n15910), .A2(n11886), .ZN(n13430) );
  AND2_X1 U16749 ( .A1(n14188), .A2(n20740), .ZN(n13428) );
  OR2_X1 U16750 ( .A1(n20177), .A2(n13428), .ZN(n13429) );
  INV_X1 U16751 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14816) );
  INV_X1 U16752 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15971) );
  INV_X1 U16753 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13433) );
  INV_X1 U16754 ( .A(n14232), .ZN(n13434) );
  INV_X1 U16755 ( .A(n14276), .ZN(n13435) );
  INV_X1 U16756 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20999) );
  NAND2_X1 U16757 ( .A1(n20745), .A2(n13438), .ZN(n13439) );
  NAND2_X1 U16758 ( .A1(n20141), .A2(n13439), .ZN(n20182) );
  NAND2_X1 U16759 ( .A1(n13440), .A2(n20182), .ZN(n13461) );
  OAI21_X1 U16760 ( .B1(n13449), .B2(P1_EBX_REG_31__SCAN_IN), .A(n11818), .ZN(
        n13443) );
  NAND2_X1 U16761 ( .A1(n20747), .A2(n20453), .ZN(n13452) );
  INV_X1 U16762 ( .A(n13452), .ZN(n13441) );
  OAI21_X1 U16763 ( .B1(n12180), .B2(n13442), .A(n13441), .ZN(n13450) );
  AND2_X1 U16764 ( .A1(n13443), .A2(n13450), .ZN(n13444) );
  NAND2_X1 U16765 ( .A1(n20745), .A2(n13444), .ZN(n20136) );
  NOR2_X1 U16766 ( .A1(n14379), .A2(n20661), .ZN(n13445) );
  INV_X1 U16767 ( .A(n15994), .ZN(n15942) );
  AOI22_X1 U16768 ( .A1(n20126), .A2(n13446), .B1(n15942), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13448) );
  NAND2_X1 U16769 ( .A1(n20178), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13447) );
  OAI211_X1 U16770 ( .C1(n20136), .C2(n12182), .A(n13448), .B(n13447), .ZN(
        n13459) );
  NOR2_X1 U16771 ( .A1(n13450), .A2(n13449), .ZN(n13451) );
  INV_X1 U16772 ( .A(n20745), .ZN(n13454) );
  NAND2_X1 U16773 ( .A1(n13452), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13453) );
  NOR2_X1 U16774 ( .A1(n13454), .A2(n13453), .ZN(n13464) );
  INV_X1 U16775 ( .A(n13455), .ZN(n13456) );
  NAND2_X1 U16776 ( .A1(n13464), .A2(n13456), .ZN(n13457) );
  OAI21_X1 U16777 ( .B1(n20152), .B2(P1_REIP_REG_1__SCAN_IN), .A(n13457), .ZN(
        n13458) );
  NOR2_X1 U16778 ( .A1(n13459), .A2(n13458), .ZN(n13460) );
  OAI211_X1 U16779 ( .C1(n20169), .C2(n20551), .A(n13461), .B(n13460), .ZN(
        P1_U2839) );
  INV_X1 U16780 ( .A(n20182), .ZN(n13471) );
  NAND2_X1 U16781 ( .A1(n20152), .A2(n15994), .ZN(n15996) );
  NOR2_X1 U16782 ( .A1(n13462), .A2(n20169), .ZN(n13469) );
  NAND2_X1 U16783 ( .A1(n20159), .A2(n13465), .ZN(n13467) );
  OAI21_X1 U16784 ( .B1(n20178), .B2(n20126), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13466) );
  OAI211_X1 U16785 ( .C1(n20136), .C2(n12852), .A(n13467), .B(n13466), .ZN(
        n13468) );
  AOI211_X1 U16786 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n15996), .A(n13469), .B(
        n13468), .ZN(n13470) );
  OAI21_X1 U16787 ( .B1(n13472), .B2(n13471), .A(n13470), .ZN(P1_U2840) );
  OAI21_X1 U16788 ( .B1(n13200), .B2(n13474), .A(n13473), .ZN(n13476) );
  NAND3_X1 U16789 ( .A1(n13476), .A2(n15149), .A3(n13475), .ZN(n13480) );
  OR2_X1 U16790 ( .A1(n13419), .A2(n13477), .ZN(n13478) );
  AND2_X1 U16791 ( .A1(n13731), .A2(n13478), .ZN(n19097) );
  NAND2_X1 U16792 ( .A1(n19097), .A2(n15159), .ZN(n13479) );
  OAI211_X1 U16793 ( .C1(n15159), .C2(n13481), .A(n13480), .B(n13479), .ZN(
        P2_U2873) );
  INV_X1 U16794 ( .A(n20423), .ZN(n13483) );
  OR2_X1 U16795 ( .A1(n13130), .A2(n20601), .ZN(n13482) );
  NAND2_X1 U16796 ( .A1(n13482), .A2(n20549), .ZN(n20519) );
  INV_X1 U16797 ( .A(n20519), .ZN(n14940) );
  OAI21_X1 U16798 ( .B1(n20393), .B2(n20513), .A(n13488), .ZN(n13485) );
  AOI211_X1 U16799 ( .C1(n13483), .C2(n14940), .A(n20601), .B(n13485), .ZN(
        n13484) );
  INV_X1 U16800 ( .A(n20607), .ZN(n20364) );
  AOI211_X2 U16801 ( .C1(n20601), .C2(n13486), .A(n13484), .B(n20364), .ZN(
        n13764) );
  INV_X1 U16802 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13491) );
  AOI22_X1 U16803 ( .A1(n13758), .A2(n20610), .B1(n13757), .B2(n20546), .ZN(
        n13490) );
  INV_X1 U16804 ( .A(n13485), .ZN(n13487) );
  OAI22_X1 U16805 ( .A1(n13487), .A2(n20601), .B1(n13486), .B2(n12842), .ZN(
        n13760) );
  INV_X1 U16806 ( .A(n13488), .ZN(n13759) );
  AOI22_X1 U16807 ( .A1(n20604), .A2(n13760), .B1(n13759), .B2(n20603), .ZN(
        n13489) );
  OAI211_X1 U16808 ( .C1(n13764), .C2(n13491), .A(n13490), .B(n13489), .ZN(
        P1_U3089) );
  INV_X1 U16809 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13494) );
  AOI22_X1 U16810 ( .A1(n13758), .A2(n20622), .B1(n13757), .B2(n20567), .ZN(
        n13493) );
  AOI22_X1 U16811 ( .A1(n20621), .A2(n13760), .B1(n13759), .B2(n20620), .ZN(
        n13492) );
  OAI211_X1 U16812 ( .C1(n13764), .C2(n13494), .A(n13493), .B(n13492), .ZN(
        P1_U3091) );
  INV_X1 U16813 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U16814 ( .A1(n13758), .A2(n20628), .B1(n13757), .B2(n20571), .ZN(
        n13496) );
  AOI22_X1 U16815 ( .A1(n20627), .A2(n13760), .B1(n13759), .B2(n20626), .ZN(
        n13495) );
  OAI211_X1 U16816 ( .C1(n13764), .C2(n13497), .A(n13496), .B(n13495), .ZN(
        P1_U3092) );
  INV_X1 U16817 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U16818 ( .A1(n13758), .A2(n20616), .B1(n13757), .B2(n20563), .ZN(
        n13499) );
  AOI22_X1 U16819 ( .A1(n20615), .A2(n13760), .B1(n13759), .B2(n20614), .ZN(
        n13498) );
  OAI211_X1 U16820 ( .C1(n13764), .C2(n13500), .A(n13499), .B(n13498), .ZN(
        P1_U3090) );
  INV_X1 U16821 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U16822 ( .A1(n13758), .A2(n20640), .B1(n13757), .B2(n20579), .ZN(
        n13502) );
  AOI22_X1 U16823 ( .A1(n20639), .A2(n13760), .B1(n13759), .B2(n20638), .ZN(
        n13501) );
  OAI211_X1 U16824 ( .C1(n13764), .C2(n13503), .A(n13502), .B(n13501), .ZN(
        P1_U3094) );
  INV_X1 U16825 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U16826 ( .A1(n13758), .A2(n20654), .B1(n13757), .B2(n20587), .ZN(
        n13505) );
  AOI22_X1 U16827 ( .A1(n20653), .A2(n13760), .B1(n13759), .B2(n20651), .ZN(
        n13504) );
  OAI211_X1 U16828 ( .C1(n13764), .C2(n13506), .A(n13505), .B(n13504), .ZN(
        P1_U3096) );
  INV_X1 U16829 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13511) );
  NOR2_X1 U16830 ( .A1(n13507), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13508) );
  OR2_X1 U16831 ( .A1(n13516), .A2(n13508), .ZN(n20158) );
  INV_X1 U16832 ( .A(n14330), .ZN(n14051) );
  INV_X1 U16833 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20148) );
  NOR2_X1 U16834 ( .A1(n14051), .A2(n20148), .ZN(n13509) );
  AOI21_X1 U16835 ( .B1(n20158), .B2(n14188), .A(n13509), .ZN(n13510) );
  OAI21_X1 U16836 ( .B1(n14294), .B2(n13511), .A(n13510), .ZN(n13512) );
  NAND2_X1 U16837 ( .A1(n13515), .A2(n14011), .ZN(n13521) );
  INV_X1 U16838 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13525) );
  NOR2_X1 U16839 ( .A1(n13516), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13517) );
  OR2_X1 U16840 ( .A1(n13551), .A2(n13517), .ZN(n20145) );
  AOI22_X1 U16841 ( .A1(n20145), .A2(n14188), .B1(n14330), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13518) );
  OAI21_X1 U16842 ( .B1(n14294), .B2(n13525), .A(n13518), .ZN(n13519) );
  INV_X1 U16843 ( .A(n13519), .ZN(n13520) );
  NAND2_X1 U16844 ( .A1(n13521), .A2(n13520), .ZN(n13523) );
  NOR2_X1 U16845 ( .A1(n13522), .A2(n13523), .ZN(n13524) );
  OR2_X1 U16846 ( .A1(n13556), .A2(n13524), .ZN(n20195) );
  OAI222_X1 U16847 ( .A1(n20195), .A2(n9731), .B1(n13526), .B2(n14722), .C1(
        n13525), .C2(n16046), .ZN(P1_U2897) );
  INV_X1 U16848 ( .A(n20271), .ZN(n13540) );
  NAND2_X1 U16849 ( .A1(n13527), .A2(n20182), .ZN(n13539) );
  INV_X1 U16850 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20116) );
  NOR2_X1 U16851 ( .A1(n20116), .A2(n13566), .ZN(n13528) );
  OAI21_X1 U16852 ( .B1(n20152), .B2(n13528), .A(n15994), .ZN(n13700) );
  INV_X1 U16853 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20685) );
  NAND3_X1 U16854 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(n20685), .ZN(n13534) );
  INV_X1 U16855 ( .A(n13529), .ZN(n13530) );
  AOI22_X1 U16856 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n13530), .ZN(n13533) );
  OR2_X1 U16857 ( .A1(n20136), .A2(n13531), .ZN(n13532) );
  OAI211_X1 U16858 ( .C1(n13534), .C2(n20152), .A(n13533), .B(n13532), .ZN(
        n13537) );
  AND2_X1 U16859 ( .A1(n20159), .A2(n13535), .ZN(n13536) );
  AOI211_X1 U16860 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n13700), .A(n13537), .B(
        n13536), .ZN(n13538) );
  OAI211_X1 U16861 ( .C1(n13540), .C2(n20169), .A(n13539), .B(n13538), .ZN(
        P1_U2837) );
  AOI22_X1 U16862 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13544) );
  AOI22_X1 U16863 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13543) );
  AOI22_X1 U16864 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13542) );
  BUF_X1 U16865 ( .A(n11701), .Z(n14239) );
  AOI22_X1 U16866 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13541) );
  NAND4_X1 U16867 ( .A1(n13544), .A2(n13543), .A3(n13542), .A4(n13541), .ZN(
        n13550) );
  AOI22_X1 U16868 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13548) );
  AOI22_X1 U16869 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13547) );
  AOI22_X1 U16870 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13546) );
  AOI22_X1 U16871 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13545) );
  NAND4_X1 U16872 ( .A1(n13548), .A2(n13547), .A3(n13546), .A4(n13545), .ZN(
        n13549) );
  OAI21_X1 U16873 ( .B1(n13550), .B2(n13549), .A(n14011), .ZN(n13555) );
  XNOR2_X1 U16874 ( .A(n13551), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13817) );
  NAND2_X1 U16875 ( .A1(n13817), .A2(n12918), .ZN(n13554) );
  NAND2_X1 U16876 ( .A1(n14331), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U16877 ( .A1(n14330), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13552) );
  NAND4_X1 U16878 ( .A1(n13555), .A2(n13554), .A3(n13553), .A4(n13552), .ZN(
        n13557) );
  OR2_X1 U16879 ( .A1(n13556), .A2(n13557), .ZN(n13558) );
  NAND2_X1 U16880 ( .A1(n13808), .A2(n13558), .ZN(n13821) );
  INV_X1 U16881 ( .A(DATAI_8_), .ZN(n13560) );
  NAND2_X1 U16882 ( .A1(n14642), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13559) );
  OAI21_X1 U16883 ( .B1(n14642), .B2(n13560), .A(n13559), .ZN(n20231) );
  AOI22_X1 U16884 ( .A1(n16043), .A2(n20231), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14724), .ZN(n13561) );
  OAI21_X1 U16885 ( .B1(n13821), .B2(n9731), .A(n13561), .ZN(P1_U2896) );
  AND2_X1 U16886 ( .A1(n13514), .A2(n13562), .ZN(n13563) );
  NOR2_X1 U16887 ( .A1(n13522), .A2(n13563), .ZN(n20155) );
  INV_X1 U16888 ( .A(n20155), .ZN(n13565) );
  OAI222_X1 U16889 ( .A1(n9731), .A2(n13565), .B1(n13670), .B2(n14722), .C1(
        n16046), .C2(n13511), .ZN(P1_U2898) );
  INV_X1 U16890 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13564) );
  XNOR2_X1 U16891 ( .A(n10063), .B(n16230), .ZN(n16240) );
  OAI222_X1 U16892 ( .A1(n14624), .A2(n13565), .B1(n13564), .B2(n20204), .C1(
        n20194), .C2(n16240), .ZN(P1_U2866) );
  INV_X1 U16893 ( .A(n13817), .ZN(n13578) );
  NOR4_X1 U16894 ( .A1(n20683), .A2(n20685), .A3(n20116), .A4(n13566), .ZN(
        n13567) );
  NAND3_X1 U16895 ( .A1(n13567), .A2(P1_REIP_REG_6__SCAN_IN), .A3(
        P1_REIP_REG_5__SCAN_IN), .ZN(n13872) );
  NOR2_X1 U16896 ( .A1(n20152), .A2(n13872), .ZN(n20133) );
  NAND2_X1 U16897 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20133), .ZN(n13576) );
  INV_X1 U16898 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U16899 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .ZN(n20119) );
  OR2_X1 U16900 ( .A1(n20152), .A2(n13567), .ZN(n13568) );
  NAND2_X1 U16901 ( .A1(n13568), .A2(n15994), .ZN(n20181) );
  INV_X1 U16902 ( .A(n20181), .ZN(n13571) );
  AND2_X1 U16903 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n13569) );
  OR2_X1 U16904 ( .A1(n20152), .A2(n13569), .ZN(n13570) );
  NAND2_X1 U16905 ( .A1(n13571), .A2(n13570), .ZN(n20150) );
  AOI21_X1 U16906 ( .B1(n15996), .B2(n20119), .A(n20150), .ZN(n20131) );
  OAI21_X1 U16907 ( .B1(n16231), .B2(n13572), .A(n16217), .ZN(n13823) );
  INV_X1 U16908 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21038) );
  OAI22_X1 U16909 ( .A1(n13823), .A2(n20175), .B1(n21038), .B2(n20136), .ZN(
        n13573) );
  AOI211_X1 U16910 ( .C1(n20178), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20177), .B(n13573), .ZN(n13574) );
  OAI221_X1 U16911 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n13576), .C1(n13575), 
        .C2(n20131), .A(n13574), .ZN(n13577) );
  AOI21_X1 U16912 ( .B1(n20126), .B2(n13578), .A(n13577), .ZN(n13579) );
  OAI21_X1 U16913 ( .B1(n20141), .B2(n13821), .A(n13579), .ZN(P1_U2832) );
  INV_X1 U16914 ( .A(n13600), .ZN(n13623) );
  AND2_X1 U16915 ( .A1(n13607), .A2(n13581), .ZN(n13595) );
  NOR2_X1 U16916 ( .A1(n9742), .A2(n15720), .ZN(n13597) );
  INV_X1 U16917 ( .A(n13620), .ZN(n13619) );
  INV_X1 U16918 ( .A(n11161), .ZN(n13582) );
  OAI22_X1 U16919 ( .A1(n13595), .A2(n13597), .B1(n13619), .B2(n13582), .ZN(
        n13588) );
  INV_X1 U16920 ( .A(n13597), .ZN(n13586) );
  NAND2_X1 U16921 ( .A1(n10697), .A2(n13583), .ZN(n13585) );
  NAND2_X1 U16922 ( .A1(n13585), .A2(n13584), .ZN(n13591) );
  OAI211_X1 U16923 ( .C1(n11161), .C2(n13619), .A(n13586), .B(n13591), .ZN(
        n13587) );
  MUX2_X1 U16924 ( .A(n13588), .B(n13587), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13589) );
  AOI211_X1 U16925 ( .C1(n13580), .C2(n13623), .A(n10820), .B(n13589), .ZN(
        n15723) );
  MUX2_X1 U16926 ( .A(n13590), .B(n15723), .S(n13601), .Z(n13635) );
  INV_X1 U16927 ( .A(n13591), .ZN(n13594) );
  NOR3_X1 U16928 ( .A1(n13619), .A2(n13592), .A3(n11161), .ZN(n13593) );
  AOI21_X1 U16929 ( .B1(n13594), .B2(n13586), .A(n13593), .ZN(n13599) );
  INV_X1 U16930 ( .A(n13595), .ZN(n13596) );
  OAI21_X1 U16931 ( .B1(n10786), .B2(n13597), .A(n13596), .ZN(n13598) );
  OAI211_X1 U16932 ( .C1(n10769), .C2(n13600), .A(n13599), .B(n13598), .ZN(
        n15719) );
  INV_X1 U16933 ( .A(n13601), .ZN(n13626) );
  NAND2_X1 U16934 ( .A1(n13626), .A2(n13602), .ZN(n13603) );
  OAI21_X1 U16935 ( .B1(n15719), .B2(n13626), .A(n13603), .ZN(n13634) );
  AOI22_X1 U16936 ( .A1(n13643), .A2(n13605), .B1(n11366), .B2(n13604), .ZN(
        n13606) );
  OAI21_X1 U16937 ( .B1(n13643), .B2(n13607), .A(n13606), .ZN(n20066) );
  NOR2_X1 U16938 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n13613) );
  AOI21_X1 U16939 ( .B1(n11564), .B2(n20756), .A(n13608), .ZN(n13609) );
  NAND3_X1 U16940 ( .A1(n11366), .A2(n13610), .A3(n13609), .ZN(n18999) );
  INV_X1 U16941 ( .A(n13611), .ZN(n13612) );
  OAI211_X1 U16942 ( .C1(n13613), .C2(n18999), .A(n13612), .B(n20068), .ZN(
        n13614) );
  AOI211_X1 U16943 ( .C1(n13626), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20066), .B(n13614), .ZN(n13633) );
  NOR2_X1 U16944 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13634), .ZN(
        n13630) );
  NAND2_X1 U16945 ( .A1(n9774), .A2(n13623), .ZN(n13618) );
  INV_X1 U16946 ( .A(n13615), .ZN(n13616) );
  OR2_X1 U16947 ( .A1(n13616), .A2(n11364), .ZN(n13621) );
  OAI21_X1 U16948 ( .B1(n10788), .B2(n10794), .A(n13621), .ZN(n13617) );
  OAI211_X1 U16949 ( .C1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n13619), .A(
        n13618), .B(n13617), .ZN(n15711) );
  INV_X1 U16950 ( .A(n15711), .ZN(n13624) );
  MUX2_X1 U16951 ( .A(n13621), .B(n13620), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13622) );
  AOI21_X1 U16952 ( .B1(n19231), .B2(n13623), .A(n13622), .ZN(n15704) );
  AOI22_X1 U16953 ( .A1(n13624), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n15704), .ZN(n13625) );
  AOI21_X1 U16954 ( .B1(n10880), .B2(n15711), .A(n13625), .ZN(n13627) );
  NOR2_X1 U16955 ( .A1(n13627), .A2(n13626), .ZN(n13628) );
  OAI21_X1 U16956 ( .B1(n13630), .B2(n20047), .A(n13628), .ZN(n13629) );
  AOI222_X1 U16957 ( .A1(n13635), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n13635), .B2(n13629), .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n13629), .ZN(n13631) );
  OAI221_X1 U16958 ( .B1(n13631), .B2(n13630), .C1(n13631), .C2(n20047), .A(
        n15937), .ZN(n13632) );
  OAI211_X1 U16959 ( .C1(n13635), .C2(n13634), .A(n13633), .B(n13632), .ZN(
        n13651) );
  INV_X1 U16960 ( .A(n20756), .ZN(n19952) );
  NOR2_X1 U16961 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19309), .ZN(n19953) );
  NAND2_X1 U16962 ( .A1(n19952), .A2(n19953), .ZN(n15932) );
  OAI21_X1 U16963 ( .B1(n13636), .B2(n16486), .A(n15932), .ZN(n13650) );
  INV_X1 U16964 ( .A(n13637), .ZN(n13638) );
  OR2_X1 U16965 ( .A1(n13639), .A2(n13638), .ZN(n13641) );
  OAI21_X1 U16966 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n13651), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13640) );
  NAND2_X1 U16967 ( .A1(n13641), .A2(n13640), .ZN(n13647) );
  INV_X1 U16968 ( .A(n20072), .ZN(n13655) );
  AND2_X1 U16969 ( .A1(n13655), .A2(n13648), .ZN(n13642) );
  NOR2_X1 U16970 ( .A1(n13647), .A2(n13642), .ZN(n19957) );
  INV_X1 U16971 ( .A(n19957), .ZN(n16487) );
  OAI21_X1 U16972 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n19309), .ZN(n20080) );
  OAI21_X1 U16973 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n15714), .A(n20080), 
        .ZN(n13644) );
  OAI21_X1 U16974 ( .B1(n16487), .B2(n20756), .A(n13644), .ZN(n13646) );
  OAI211_X1 U16975 ( .C1(n13648), .C2(n13647), .A(n13646), .B(n13645), .ZN(
        n13649) );
  AOI211_X1 U16976 ( .C1(n13651), .C2(n19304), .A(n13650), .B(n13649), .ZN(
        n13652) );
  INV_X1 U16977 ( .A(n13652), .ZN(P2_U3176) );
  OAI222_X1 U16978 ( .A1(n13821), .A2(n14624), .B1(n20204), .B2(n21038), .C1(
        n13823), .C2(n20194), .ZN(P1_U2864) );
  NOR2_X2 U16979 ( .A1(n19737), .A2(n19893), .ZN(n19927) );
  NOR2_X2 U16980 ( .A1(n19673), .A2(n19579), .ZN(n19465) );
  OAI21_X1 U16981 ( .B1(n19927), .B2(n19465), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13653) );
  NAND2_X1 U16982 ( .A1(n13653), .A2(n20029), .ZN(n13666) );
  INV_X1 U16983 ( .A(n13666), .ZN(n13657) );
  NAND2_X1 U16984 ( .A1(n12315), .A2(n20047), .ZN(n19501) );
  OR2_X1 U16985 ( .A1(n19501), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19443) );
  NOR2_X1 U16986 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19443), .ZN(
        n19432) );
  INV_X1 U16987 ( .A(n19432), .ZN(n13660) );
  AND2_X1 U16988 ( .A1(n19882), .A2(n13660), .ZN(n13665) );
  INV_X1 U16989 ( .A(n20080), .ZN(n13654) );
  AOI211_X1 U16990 ( .C1(n13663), .C2(n20037), .A(n20029), .B(n19432), .ZN(
        n13656) );
  INV_X1 U16991 ( .A(n19931), .ZN(n19832) );
  AOI22_X1 U16992 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19435), .ZN(n19598) );
  INV_X1 U16993 ( .A(n19465), .ZN(n13661) );
  NAND2_X1 U16994 ( .A1(n13659), .A2(n19430), .ZN(n19458) );
  OAI22_X1 U16995 ( .A1(n19598), .A2(n13661), .B1(n13660), .B2(n19458), .ZN(
        n13662) );
  AOI21_X1 U16996 ( .B1(n19927), .B2(n19832), .A(n13662), .ZN(n13668) );
  OAI21_X1 U16997 ( .B1(n13663), .B2(n19432), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13664) );
  NOR2_X2 U16998 ( .A1(n19277), .A2(n9715), .ZN(n19925) );
  NAND2_X1 U16999 ( .A1(n19436), .A2(n19925), .ZN(n13667) );
  OAI211_X1 U17000 ( .C1(n19439), .C2(n13669), .A(n13668), .B(n13667), .ZN(
        P2_U3053) );
  NOR2_X2 U17001 ( .A1(n13670), .A2(n13676), .ZN(n20645) );
  INV_X1 U17002 ( .A(n20645), .ZN(n13675) );
  NAND2_X1 U17003 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13674) );
  AOI22_X1 U17004 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13682), .B1(DATAI_30_), 
        .B2(n13681), .ZN(n20586) );
  AOI22_X1 U17005 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13682), .B1(DATAI_22_), 
        .B2(n13681), .ZN(n20649) );
  OAI22_X1 U17006 ( .A1(n13684), .A2(n20586), .B1(n20649), .B2(n13683), .ZN(
        n13672) );
  AOI21_X1 U17007 ( .B1(n13686), .B2(n20644), .A(n13672), .ZN(n13673) );
  OAI211_X1 U17008 ( .C1(n13690), .C2(n13675), .A(n13674), .B(n13673), .ZN(
        P1_U3087) );
  NOR2_X2 U17009 ( .A1(n13677), .A2(n13676), .ZN(n20633) );
  INV_X1 U17010 ( .A(n20633), .ZN(n13689) );
  NAND2_X1 U17011 ( .A1(n13678), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13688) );
  NOR2_X2 U17012 ( .A1(n13680), .A2(n13679), .ZN(n20632) );
  AOI22_X1 U17013 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13682), .B1(DATAI_28_), 
        .B2(n13681), .ZN(n20578) );
  AOI22_X1 U17014 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n13682), .B1(DATAI_20_), 
        .B2(n13681), .ZN(n20637) );
  OAI22_X1 U17015 ( .A1(n13684), .A2(n20578), .B1(n20637), .B2(n13683), .ZN(
        n13685) );
  AOI21_X1 U17016 ( .B1(n13686), .B2(n20632), .A(n13685), .ZN(n13687) );
  OAI211_X1 U17017 ( .C1(n13690), .C2(n13689), .A(n13688), .B(n13687), .ZN(
        P1_U3085) );
  NAND2_X1 U17018 ( .A1(n13691), .A2(n20182), .ZN(n13702) );
  OAI21_X1 U17019 ( .B1(n20152), .B2(n20116), .A(n13566), .ZN(n13699) );
  INV_X1 U17020 ( .A(n13692), .ZN(n13697) );
  INV_X1 U17021 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13693) );
  OAI22_X1 U17022 ( .A1(n13694), .A2(n20186), .B1(n20162), .B2(n13693), .ZN(
        n13695) );
  AOI21_X1 U17023 ( .B1(n20170), .B2(P1_EBX_REG_2__SCAN_IN), .A(n13695), .ZN(
        n13696) );
  OAI21_X1 U17024 ( .B1(n20175), .B2(n13697), .A(n13696), .ZN(n13698) );
  AOI21_X1 U17025 ( .B1(n13700), .B2(n13699), .A(n13698), .ZN(n13701) );
  OAI211_X1 U17026 ( .C1(n20169), .C2(n13125), .A(n13702), .B(n13701), .ZN(
        P1_U2838) );
  INV_X1 U17027 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13705) );
  INV_X1 U17028 ( .A(n20649), .ZN(n20583) );
  INV_X1 U17029 ( .A(n20586), .ZN(n20646) );
  AOI22_X1 U17030 ( .A1(n20655), .A2(n20583), .B1(n13718), .B2(n20646), .ZN(
        n13704) );
  AOI22_X1 U17031 ( .A1(n20645), .A2(n13713), .B1(n20644), .B2(n13712), .ZN(
        n13703) );
  OAI211_X1 U17032 ( .C1(n13717), .C2(n13705), .A(n13704), .B(n13703), .ZN(
        P1_U3151) );
  INV_X1 U17033 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13708) );
  AOI22_X1 U17034 ( .A1(n13718), .A2(n20583), .B1(n20588), .B2(n20646), .ZN(
        n13707) );
  AOI22_X1 U17035 ( .A1(n20645), .A2(n13720), .B1(n20644), .B2(n13719), .ZN(
        n13706) );
  OAI211_X1 U17036 ( .C1(n13724), .C2(n13708), .A(n13707), .B(n13706), .ZN(
        P1_U3143) );
  INV_X1 U17037 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U17038 ( .A1(n20473), .A2(n20583), .B1(n13757), .B2(n20646), .ZN(
        n13710) );
  AOI22_X1 U17039 ( .A1(n20645), .A2(n13725), .B1(n20644), .B2(n10216), .ZN(
        n13709) );
  OAI211_X1 U17040 ( .C1(n13729), .C2(n13711), .A(n13710), .B(n13709), .ZN(
        P1_U3103) );
  INV_X1 U17041 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13716) );
  INV_X1 U17042 ( .A(n20637), .ZN(n20575) );
  INV_X1 U17043 ( .A(n20578), .ZN(n20634) );
  AOI22_X1 U17044 ( .A1(n20655), .A2(n20575), .B1(n13718), .B2(n20634), .ZN(
        n13715) );
  AOI22_X1 U17045 ( .A1(n20633), .A2(n13713), .B1(n20632), .B2(n13712), .ZN(
        n13714) );
  OAI211_X1 U17046 ( .C1(n13717), .C2(n13716), .A(n13715), .B(n13714), .ZN(
        P1_U3149) );
  INV_X1 U17047 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U17048 ( .A1(n13718), .A2(n20575), .B1(n20588), .B2(n20634), .ZN(
        n13722) );
  AOI22_X1 U17049 ( .A1(n20633), .A2(n13720), .B1(n20632), .B2(n13719), .ZN(
        n13721) );
  OAI211_X1 U17050 ( .C1(n13724), .C2(n13723), .A(n13722), .B(n13721), .ZN(
        P1_U3141) );
  INV_X1 U17051 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13728) );
  AOI22_X1 U17052 ( .A1(n20473), .A2(n20575), .B1(n13757), .B2(n20634), .ZN(
        n13727) );
  AOI22_X1 U17053 ( .A1(n20633), .A2(n13725), .B1(n20632), .B2(n10216), .ZN(
        n13726) );
  OAI211_X1 U17054 ( .C1(n13729), .C2(n13728), .A(n13727), .B(n13726), .ZN(
        P1_U3101) );
  XNOR2_X1 U17055 ( .A(n13475), .B(n13730), .ZN(n13736) );
  INV_X1 U17056 ( .A(n13731), .ZN(n13734) );
  INV_X1 U17057 ( .A(n13732), .ZN(n13733) );
  OAI21_X1 U17058 ( .B1(n13734), .B2(n13733), .A(n15181), .ZN(n19085) );
  MUX2_X1 U17059 ( .A(n11072), .B(n19085), .S(n15159), .Z(n13735) );
  OAI21_X1 U17060 ( .B1(n13736), .B2(n15185), .A(n13735), .ZN(P2_U2872) );
  NAND3_X1 U17061 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n12315), .A3(
        n10880), .ZN(n19556) );
  NOR2_X1 U17062 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19556), .ZN(
        n19544) );
  INV_X1 U17063 ( .A(n19544), .ZN(n13748) );
  NAND2_X1 U17064 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13748), .ZN(n13737) );
  OR2_X1 U17065 ( .A1(n13738), .A2(n13737), .ZN(n13745) );
  OAI21_X1 U17066 ( .B1(n19546), .B2(n19564), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13741) );
  INV_X1 U17067 ( .A(n13739), .ZN(n13740) );
  NOR2_X1 U17068 ( .A1(n13740), .A2(n19707), .ZN(n19778) );
  NAND2_X1 U17069 ( .A1(n19778), .A2(n12315), .ZN(n13743) );
  AOI22_X1 U17070 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13748), .B1(n13741), 
        .B2(n13743), .ZN(n13742) );
  NAND3_X1 U17071 ( .A1(n13745), .A2(n13742), .A3(n19889), .ZN(n19547) );
  INV_X1 U17072 ( .A(n19547), .ZN(n13753) );
  INV_X1 U17073 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13752) );
  OAI21_X1 U17074 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13743), .A(n12754), 
        .ZN(n13744) );
  AND2_X1 U17075 ( .A1(n13745), .A2(n13744), .ZN(n19545) );
  NOR2_X2 U17076 ( .A1(n19244), .A2(n9715), .ZN(n19887) );
  INV_X1 U17077 ( .A(n19886), .ZN(n13749) );
  AOI22_X1 U17078 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19435), .ZN(n19749) );
  INV_X1 U17079 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18316) );
  INV_X1 U17080 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16565) );
  AOI22_X1 U17081 ( .A1(n19564), .A2(n19896), .B1(n19546), .B2(n19820), .ZN(
        n13747) );
  OAI21_X1 U17082 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n13750) );
  AOI21_X1 U17083 ( .B1(n19545), .B2(n19887), .A(n13750), .ZN(n13751) );
  OAI21_X1 U17084 ( .B1(n13753), .B2(n13752), .A(n13751), .ZN(P2_U3080) );
  INV_X1 U17085 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13756) );
  AOI22_X1 U17086 ( .A1(n13758), .A2(n20646), .B1(n13757), .B2(n20583), .ZN(
        n13755) );
  AOI22_X1 U17087 ( .A1(n20645), .A2(n13760), .B1(n13759), .B2(n20644), .ZN(
        n13754) );
  OAI211_X1 U17088 ( .C1(n13764), .C2(n13756), .A(n13755), .B(n13754), .ZN(
        P1_U3095) );
  INV_X1 U17089 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U17090 ( .A1(n13758), .A2(n20634), .B1(n13757), .B2(n20575), .ZN(
        n13762) );
  AOI22_X1 U17091 ( .A1(n20633), .A2(n13760), .B1(n13759), .B2(n20632), .ZN(
        n13761) );
  OAI211_X1 U17092 ( .C1(n13764), .C2(n13763), .A(n13762), .B(n13761), .ZN(
        P1_U3093) );
  OAI21_X1 U17093 ( .B1(n13767), .B2(n13766), .A(n13765), .ZN(n16426) );
  INV_X1 U17094 ( .A(n13769), .ZN(n13773) );
  OAI21_X1 U17095 ( .B1(n13773), .B2(n9720), .A(n13771), .ZN(n13772) );
  OAI21_X1 U17096 ( .B1(n13768), .B2(n13773), .A(n13772), .ZN(n16428) );
  INV_X1 U17097 ( .A(n16428), .ZN(n13791) );
  OAI21_X1 U17098 ( .B1(n13776), .B2(n13775), .A(n13774), .ZN(n19285) );
  OR2_X1 U17099 ( .A1(n13778), .A2(n13777), .ZN(n13780) );
  NAND2_X1 U17100 ( .A1(n13780), .A2(n13779), .ZN(n19199) );
  INV_X1 U17101 ( .A(n19199), .ZN(n13788) );
  INV_X1 U17102 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19978) );
  NOR2_X1 U17103 ( .A1(n19978), .A2(n19210), .ZN(n13787) );
  OAI21_X1 U17104 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n13781), .ZN(n13783) );
  OAI22_X1 U17105 ( .A1(n13785), .A2(n13784), .B1(n13783), .B2(n13782), .ZN(
        n13786) );
  AOI211_X1 U17106 ( .C1(n16475), .C2(n13788), .A(n13787), .B(n13786), .ZN(
        n13789) );
  OAI21_X1 U17107 ( .B1(n19285), .B2(n19400), .A(n13789), .ZN(n13790) );
  AOI21_X1 U17108 ( .B1(n13791), .B2(n19391), .A(n13790), .ZN(n13792) );
  OAI21_X1 U17109 ( .B1(n16477), .B2(n16426), .A(n13792), .ZN(P2_U3041) );
  XOR2_X1 U17110 ( .A(n20122), .B(n13793), .Z(n20125) );
  AOI22_X1 U17111 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13797) );
  AOI22_X1 U17112 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9761), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13796) );
  AOI22_X1 U17113 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13795) );
  AOI22_X1 U17114 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13794) );
  NAND4_X1 U17115 ( .A1(n13797), .A2(n13796), .A3(n13795), .A4(n13794), .ZN(
        n13803) );
  AOI22_X1 U17116 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13801) );
  AOI22_X1 U17117 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U17118 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13799) );
  AOI22_X1 U17119 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13798) );
  NAND4_X1 U17120 ( .A1(n13801), .A2(n13800), .A3(n13799), .A4(n13798), .ZN(
        n13802) );
  OR2_X1 U17121 ( .A1(n13803), .A2(n13802), .ZN(n13804) );
  AOI22_X1 U17122 ( .A1(n14011), .A2(n13804), .B1(n14330), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U17123 ( .A1(n14331), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13805) );
  OAI211_X1 U17124 ( .C1(n20125), .C2(n14303), .A(n13806), .B(n13805), .ZN(
        n13807) );
  INV_X1 U17125 ( .A(n13807), .ZN(n13809) );
  NAND2_X1 U17126 ( .A1(n13808), .A2(n13809), .ZN(n13810) );
  NAND2_X1 U17127 ( .A1(n9839), .A2(n13810), .ZN(n20189) );
  INV_X1 U17128 ( .A(DATAI_9_), .ZN(n13812) );
  NAND2_X1 U17129 ( .A1(n14642), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13811) );
  OAI21_X1 U17130 ( .B1(n14642), .B2(n13812), .A(n13811), .ZN(n20233) );
  AOI22_X1 U17131 ( .A1(n16043), .A2(n20233), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14724), .ZN(n13813) );
  OAI21_X1 U17132 ( .B1(n20189), .B2(n9731), .A(n13813), .ZN(P1_U2895) );
  XNOR2_X1 U17133 ( .A(n13814), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13815) );
  XNOR2_X1 U17134 ( .A(n13816), .B(n13815), .ZN(n13822) );
  NAND2_X1 U17135 ( .A1(n13822), .A2(n16116), .ZN(n13820) );
  NOR2_X1 U17136 ( .A1(n9736), .A2(n13575), .ZN(n13831) );
  NOR2_X1 U17137 ( .A1(n16111), .A2(n13817), .ZN(n13818) );
  AOI211_X1 U17138 ( .C1(n16104), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13831), .B(n13818), .ZN(n13819) );
  OAI211_X1 U17139 ( .C1(n14832), .C2(n13821), .A(n13820), .B(n13819), .ZN(
        P1_U2991) );
  INV_X1 U17140 ( .A(n13822), .ZN(n13834) );
  INV_X1 U17141 ( .A(n13823), .ZN(n13832) );
  OR2_X1 U17142 ( .A1(n13825), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16248) );
  INV_X1 U17143 ( .A(n13901), .ZN(n14923) );
  NOR2_X1 U17144 ( .A1(n16204), .A2(n14920), .ZN(n13824) );
  AOI211_X1 U17145 ( .C1(n14923), .C2(n13825), .A(n13824), .B(n16208), .ZN(
        n16263) );
  OAI21_X1 U17146 ( .B1(n14926), .B2(n16248), .A(n16263), .ZN(n16242) );
  AOI21_X1 U17147 ( .B1(n13827), .B2(n14910), .A(n16242), .ZN(n16238) );
  INV_X1 U17148 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13829) );
  INV_X1 U17149 ( .A(n16250), .ZN(n13826) );
  NOR3_X1 U17150 ( .A1(n14918), .A2(n13827), .A3(n13826), .ZN(n16234) );
  INV_X1 U17151 ( .A(n16234), .ZN(n16212) );
  OAI21_X1 U17152 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16213), .ZN(n13828) );
  OAI22_X1 U17153 ( .A1(n16238), .A2(n13829), .B1(n16212), .B2(n13828), .ZN(
        n13830) );
  AOI211_X1 U17154 ( .C1(n16256), .C2(n13832), .A(n13831), .B(n13830), .ZN(
        n13833) );
  OAI21_X1 U17155 ( .B1(n16259), .B2(n13834), .A(n13833), .ZN(P1_U3023) );
  NAND2_X1 U17156 ( .A1(n13835), .A2(n13836), .ZN(n15164) );
  OAI21_X1 U17157 ( .B1(n13835), .B2(n13836), .A(n15164), .ZN(n15177) );
  OAI21_X1 U17158 ( .B1(n13837), .B2(n13838), .A(n15557), .ZN(n13839) );
  INV_X1 U17159 ( .A(n13839), .ZN(n19065) );
  NOR2_X2 U17160 ( .A1(n13841), .A2(n15187), .ZN(n19247) );
  INV_X1 U17161 ( .A(n19247), .ZN(n15254) );
  INV_X1 U17162 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14710) );
  NOR2_X2 U17163 ( .A1(n13841), .A2(n13840), .ZN(n19248) );
  INV_X1 U17164 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19342) );
  OAI22_X1 U17165 ( .A1(n15250), .A2(n19410), .B1(n19275), .B2(n19342), .ZN(
        n13842) );
  AOI21_X1 U17166 ( .B1(n19248), .B2(BUF2_REG_17__SCAN_IN), .A(n13842), .ZN(
        n13843) );
  OAI21_X1 U17167 ( .B1(n15254), .B2(n14710), .A(n13843), .ZN(n13844) );
  AOI21_X1 U17168 ( .B1(n19065), .B2(n19295), .A(n13844), .ZN(n13845) );
  OAI21_X1 U17169 ( .B1(n19299), .B2(n15177), .A(n13845), .ZN(P2_U2902) );
  XNOR2_X1 U17170 ( .A(n13846), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14841) );
  AOI22_X1 U17171 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U17172 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13849) );
  AOI22_X1 U17173 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13848) );
  AOI22_X1 U17174 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13847) );
  NAND4_X1 U17175 ( .A1(n13850), .A2(n13849), .A3(n13848), .A4(n13847), .ZN(
        n13856) );
  AOI22_X1 U17176 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U17177 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U17178 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13852) );
  AOI22_X1 U17179 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13851) );
  NAND4_X1 U17180 ( .A1(n13854), .A2(n13853), .A3(n13852), .A4(n13851), .ZN(
        n13855) );
  NOR2_X1 U17181 ( .A1(n13856), .A2(n13855), .ZN(n13859) );
  NAND2_X1 U17182 ( .A1(n14331), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13858) );
  NAND2_X1 U17183 ( .A1(n14330), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13857) );
  OAI211_X1 U17184 ( .C1(n13971), .C2(n13859), .A(n13858), .B(n13857), .ZN(
        n13860) );
  AOI21_X1 U17185 ( .B1(n14841), .B2(n12918), .A(n13860), .ZN(n13862) );
  AOI21_X1 U17186 ( .B1(n13862), .B2(n9839), .A(n13921), .ZN(n14843) );
  INV_X1 U17187 ( .A(n14624), .ZN(n20200) );
  NAND2_X1 U17188 ( .A1(n16219), .A2(n13863), .ZN(n13864) );
  NAND2_X1 U17189 ( .A1(n13981), .A2(n13864), .ZN(n16209) );
  OAI22_X1 U17190 ( .A1(n16209), .A2(n20194), .B1(n13870), .B2(n20204), .ZN(
        n13865) );
  AOI21_X1 U17191 ( .B1(n14843), .B2(n20200), .A(n13865), .ZN(n13866) );
  INV_X1 U17192 ( .A(n13866), .ZN(P1_U2862) );
  INV_X1 U17193 ( .A(n14843), .ZN(n13878) );
  INV_X1 U17194 ( .A(DATAI_10_), .ZN(n13868) );
  NAND2_X1 U17195 ( .A1(n14642), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13867) );
  OAI21_X1 U17196 ( .B1(n14642), .B2(n13868), .A(n13867), .ZN(n20235) );
  AOI22_X1 U17197 ( .A1(n16043), .A2(n20235), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14724), .ZN(n13869) );
  OAI21_X1 U17198 ( .B1(n13878), .B2(n9731), .A(n13869), .ZN(P1_U2894) );
  NAND3_X1 U17199 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .A3(P1_REIP_REG_7__SCAN_IN), .ZN(n13871) );
  NOR2_X1 U17200 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n13871), .ZN(n13876) );
  OAI22_X1 U17201 ( .A1(n13870), .A2(n20136), .B1(n20186), .B2(n14841), .ZN(
        n13875) );
  INV_X1 U17202 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20835) );
  NOR3_X1 U17203 ( .A1(n20835), .A2(n13872), .A3(n13871), .ZN(n16026) );
  OAI21_X1 U17204 ( .B1(n20152), .B2(n16026), .A(n15994), .ZN(n16037) );
  AOI22_X1 U17205 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20178), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n16037), .ZN(n13873) );
  OAI211_X1 U17206 ( .C1(n16209), .C2(n20175), .A(n13873), .B(n9736), .ZN(
        n13874) );
  AOI211_X1 U17207 ( .C1(n20133), .C2(n13876), .A(n13875), .B(n13874), .ZN(
        n13877) );
  OAI21_X1 U17208 ( .B1(n13878), .B2(n20141), .A(n13877), .ZN(P1_U2830) );
  XNOR2_X1 U17209 ( .A(n16090), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13879) );
  XNOR2_X1 U17210 ( .A(n13880), .B(n13879), .ZN(n16224) );
  NAND2_X1 U17211 ( .A1(n16224), .A2(n16116), .ZN(n13883) );
  NAND2_X1 U17212 ( .A1(n20177), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16221) );
  OAI21_X1 U17213 ( .B1(n16120), .B2(n20122), .A(n16221), .ZN(n13881) );
  AOI21_X1 U17214 ( .B1(n16114), .B2(n20125), .A(n13881), .ZN(n13882) );
  OAI211_X1 U17215 ( .C1(n14832), .C2(n20189), .A(n13883), .B(n13882), .ZN(
        P1_U2990) );
  INV_X1 U17216 ( .A(n13884), .ZN(n15163) );
  NAND2_X1 U17217 ( .A1(n15166), .A2(n13885), .ZN(n15148) );
  OAI21_X1 U17218 ( .B1(n15166), .B2(n13885), .A(n15148), .ZN(n15162) );
  XOR2_X1 U17219 ( .A(n13886), .B(n15559), .Z(n19040) );
  NAND2_X1 U17220 ( .A1(n19040), .A2(n19295), .ZN(n13890) );
  INV_X1 U17221 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19337) );
  OAI22_X1 U17222 ( .A1(n15250), .A2(n19422), .B1(n19275), .B2(n19337), .ZN(
        n13888) );
  INV_X1 U17223 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14696) );
  NOR2_X1 U17224 ( .A1(n15254), .A2(n14696), .ZN(n13887) );
  AOI211_X1 U17225 ( .C1(n19248), .C2(BUF2_REG_19__SCAN_IN), .A(n13888), .B(
        n13887), .ZN(n13889) );
  OAI211_X1 U17226 ( .C1(n19299), .C2(n15162), .A(n13890), .B(n13889), .ZN(
        P2_U2900) );
  NAND2_X1 U17227 ( .A1(n14834), .A2(n16076), .ZN(n13895) );
  INV_X1 U17228 ( .A(n13892), .ZN(n13893) );
  AOI21_X1 U17229 ( .B1(n13895), .B2(n13894), .A(n13893), .ZN(n13897) );
  MUX2_X1 U17230 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n12227), .S(
        n16090), .Z(n13896) );
  XNOR2_X1 U17231 ( .A(n13897), .B(n13896), .ZN(n13996) );
  NAND2_X1 U17232 ( .A1(n14541), .A2(n13898), .ZN(n13899) );
  NAND2_X1 U17233 ( .A1(n14612), .A2(n13899), .ZN(n16018) );
  INV_X1 U17234 ( .A(n14899), .ZN(n13903) );
  OAI21_X1 U17235 ( .B1(n13901), .B2(n13900), .A(n14919), .ZN(n14908) );
  AOI21_X1 U17236 ( .B1(n14885), .B2(n13902), .A(n14908), .ZN(n16196) );
  OAI21_X1 U17237 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13903), .A(
        n16196), .ZN(n13904) );
  NAND2_X1 U17238 ( .A1(n13904), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13905) );
  NAND2_X1 U17239 ( .A1(n20177), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n13992) );
  OAI211_X1 U17240 ( .C1(n16220), .C2(n16018), .A(n13905), .B(n13992), .ZN(
        n13906) );
  AOI21_X1 U17241 ( .B1(n12227), .B2(n16140), .A(n13906), .ZN(n13907) );
  OAI21_X1 U17242 ( .B1(n13996), .B2(n16259), .A(n13907), .ZN(P1_U3017) );
  INV_X1 U17243 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13986) );
  OAI21_X1 U17244 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13908), .A(
        n13948), .ZN(n16097) );
  AOI22_X1 U17245 ( .A1(n14188), .A2(n16097), .B1(n14330), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13909) );
  OAI21_X1 U17246 ( .B1(n14294), .B2(n13986), .A(n13909), .ZN(n13979) );
  AOI22_X1 U17247 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14221), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17248 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U17249 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U17250 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13910) );
  NAND4_X1 U17251 ( .A1(n13913), .A2(n13912), .A3(n13911), .A4(n13910), .ZN(
        n13919) );
  AOI22_X1 U17252 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U17253 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U17254 ( .A1(n14308), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U17255 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13914) );
  NAND4_X1 U17256 ( .A1(n13917), .A2(n13916), .A3(n13915), .A4(n13914), .ZN(
        n13918) );
  OR2_X1 U17257 ( .A1(n13919), .A2(n13918), .ZN(n13920) );
  AND2_X1 U17258 ( .A1(n14011), .A2(n13920), .ZN(n14534) );
  NAND2_X1 U17259 ( .A1(n13921), .A2(n14534), .ZN(n13922) );
  XOR2_X1 U17260 ( .A(n14548), .B(n13923), .Z(n14828) );
  AOI22_X1 U17261 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U17262 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U17263 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U17264 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13924) );
  NAND4_X1 U17265 ( .A1(n13927), .A2(n13926), .A3(n13925), .A4(n13924), .ZN(
        n13933) );
  AOI22_X1 U17266 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14126), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U17267 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14239), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U17268 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U17269 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13928) );
  NAND4_X1 U17270 ( .A1(n13931), .A2(n13930), .A3(n13929), .A4(n13928), .ZN(
        n13932) );
  OR2_X1 U17271 ( .A1(n13933), .A2(n13932), .ZN(n13934) );
  AOI22_X1 U17272 ( .A1(n14011), .A2(n13934), .B1(n14330), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13936) );
  NAND2_X1 U17273 ( .A1(n14331), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13935) );
  OAI211_X1 U17274 ( .C1(n14828), .C2(n14303), .A(n13936), .B(n13935), .ZN(
        n14537) );
  INV_X1 U17275 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17276 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U17277 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11845), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17278 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13938) );
  AOI22_X1 U17279 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13937) );
  NAND4_X1 U17280 ( .A1(n13940), .A2(n13939), .A3(n13938), .A4(n13937), .ZN(
        n13946) );
  AOI22_X1 U17281 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14006), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U17282 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U17283 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U17284 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13941) );
  NAND4_X1 U17285 ( .A1(n13944), .A2(n13943), .A3(n13942), .A4(n13941), .ZN(
        n13945) );
  OR2_X1 U17286 ( .A1(n13946), .A2(n13945), .ZN(n13947) );
  NAND2_X1 U17287 ( .A1(n14011), .A2(n13947), .ZN(n13951) );
  XOR2_X1 U17288 ( .A(n16028), .B(n13948), .Z(n16086) );
  INV_X1 U17289 ( .A(n16086), .ZN(n13949) );
  AOI22_X1 U17290 ( .A1(n14330), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n14188), .B2(n13949), .ZN(n13950) );
  OAI211_X1 U17291 ( .C1(n13952), .C2(n14294), .A(n13951), .B(n13950), .ZN(
        n14536) );
  AND2_X1 U17292 ( .A1(n14537), .A2(n14536), .ZN(n13953) );
  NAND2_X1 U17293 ( .A1(n13955), .A2(n21042), .ZN(n13957) );
  INV_X1 U17294 ( .A(n14014), .ZN(n13956) );
  NAND2_X1 U17295 ( .A1(n13957), .A2(n13956), .ZN(n13991) );
  AOI22_X1 U17296 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U17297 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13960) );
  AOI22_X1 U17298 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13959) );
  AOI22_X1 U17299 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13958) );
  NAND4_X1 U17300 ( .A1(n13961), .A2(n13960), .A3(n13959), .A4(n13958), .ZN(
        n13967) );
  AOI22_X1 U17301 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13965) );
  AOI22_X1 U17302 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14239), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U17303 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U17304 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13962) );
  NAND4_X1 U17305 ( .A1(n13965), .A2(n13964), .A3(n13963), .A4(n13962), .ZN(
        n13966) );
  NOR2_X1 U17306 ( .A1(n13967), .A2(n13966), .ZN(n13970) );
  NAND2_X1 U17307 ( .A1(n14331), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13969) );
  NAND2_X1 U17308 ( .A1(n14330), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13968) );
  OAI211_X1 U17309 ( .C1(n13971), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        n13972) );
  AOI21_X1 U17310 ( .B1(n13991), .B2(n14188), .A(n13972), .ZN(n14019) );
  OR2_X1 U17311 ( .A1(n14021), .A2(n14019), .ZN(n14609) );
  NAND2_X1 U17312 ( .A1(n14021), .A2(n14019), .ZN(n13973) );
  INV_X1 U17313 ( .A(n16021), .ZN(n13977) );
  INV_X1 U17314 ( .A(DATAI_14_), .ZN(n13975) );
  NAND2_X1 U17315 ( .A1(n14642), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13974) );
  OAI21_X1 U17316 ( .B1(n14642), .B2(n13975), .A(n13974), .ZN(n20243) );
  AOI22_X1 U17317 ( .A1(n16043), .A2(n20243), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14724), .ZN(n13976) );
  OAI21_X1 U17318 ( .B1(n13977), .B2(n9731), .A(n13976), .ZN(P1_U2890) );
  OR2_X1 U17319 ( .A1(n13921), .A2(n13979), .ZN(n13980) );
  AND2_X1 U17320 ( .A1(n13978), .A2(n13980), .ZN(n14535) );
  XOR2_X1 U17321 ( .A(n14534), .B(n14535), .Z(n16094) );
  INV_X1 U17322 ( .A(n16094), .ZN(n13988) );
  AOI21_X1 U17323 ( .B1(n13982), .B2(n13981), .A(n14621), .ZN(n16197) );
  AOI22_X1 U17324 ( .A1(n16197), .A2(n20199), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14615), .ZN(n13983) );
  OAI21_X1 U17325 ( .B1(n13988), .B2(n14624), .A(n13983), .ZN(P1_U2861) );
  INV_X1 U17326 ( .A(DATAI_11_), .ZN(n13985) );
  NAND2_X1 U17327 ( .A1(n14642), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13984) );
  OAI21_X1 U17328 ( .B1(n14642), .B2(n13985), .A(n13984), .ZN(n20237) );
  INV_X1 U17329 ( .A(n20237), .ZN(n13987) );
  OAI222_X1 U17330 ( .A1(n13988), .A2(n9731), .B1(n13987), .B2(n14722), .C1(
        n13986), .C2(n16046), .ZN(P1_U2893) );
  OAI22_X1 U17331 ( .A1(n16018), .A2(n20194), .B1(n16017), .B2(n20204), .ZN(
        n13989) );
  AOI21_X1 U17332 ( .B1(n16021), .B2(n20200), .A(n13989), .ZN(n13990) );
  INV_X1 U17333 ( .A(n13990), .ZN(P1_U2858) );
  INV_X1 U17334 ( .A(n13991), .ZN(n16020) );
  NAND2_X1 U17335 ( .A1(n16114), .A2(n16020), .ZN(n13993) );
  OAI211_X1 U17336 ( .C1(n16120), .C2(n21042), .A(n13993), .B(n13992), .ZN(
        n13994) );
  AOI21_X1 U17337 ( .B1(n16021), .B2(n16069), .A(n13994), .ZN(n13995) );
  OAI21_X1 U17338 ( .B1(n13996), .B2(n20100), .A(n13995), .ZN(P1_U2985) );
  INV_X1 U17339 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18777) );
  NAND3_X1 U17340 ( .A1(n17334), .A2(n15854), .A3(n18777), .ZN(n18308) );
  NOR2_X1 U17341 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18308), .ZN(n13998) );
  NAND3_X1 U17342 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18926)
         );
  NAND2_X1 U17343 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18307) );
  NAND2_X1 U17344 ( .A1(n18937), .A2(n18986), .ZN(n18973) );
  NAND2_X1 U17345 ( .A1(n18777), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18829) );
  AOI21_X1 U17346 ( .B1(n18307), .B2(n18973), .A(n18952), .ZN(n13997) );
  INV_X1 U17347 ( .A(n13997), .ZN(n18317) );
  OAI21_X1 U17348 ( .B1(n13998), .B2(n18926), .A(n18367), .ZN(n18314) );
  INV_X1 U17349 ( .A(n18314), .ZN(n13999) );
  INV_X1 U17350 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16668) );
  NOR2_X1 U17351 ( .A1(n18937), .A2(n16668), .ZN(n17968) );
  NAND2_X1 U17352 ( .A1(n21062), .A2(n18307), .ZN(n18976) );
  NOR2_X1 U17353 ( .A1(n17968), .A2(n18976), .ZN(n15841) );
  AOI21_X1 U17354 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15841), .ZN(n15842) );
  NOR2_X1 U17355 ( .A1(n13999), .A2(n15842), .ZN(n14001) );
  NAND3_X1 U17356 ( .A1(n18986), .A2(n21062), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18672) );
  INV_X1 U17357 ( .A(n18672), .ZN(n15843) );
  NOR2_X1 U17358 ( .A1(n21062), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18366) );
  OR2_X1 U17359 ( .A1(n18366), .A2(n13999), .ZN(n15840) );
  OR2_X1 U17360 ( .A1(n15843), .A2(n15840), .ZN(n14000) );
  MUX2_X1 U17361 ( .A(n14001), .B(n14000), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI22_X1 U17362 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14005) );
  AOI22_X1 U17363 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14004) );
  AOI22_X1 U17364 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14003) );
  AOI22_X1 U17365 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14002) );
  NAND4_X1 U17366 ( .A1(n14005), .A2(n14004), .A3(n14003), .A4(n14002), .ZN(
        n14013) );
  AOI22_X1 U17367 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U17368 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U17369 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14008) );
  AOI22_X1 U17370 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14007) );
  NAND4_X1 U17371 ( .A1(n14010), .A2(n14009), .A3(n14008), .A4(n14007), .ZN(
        n14012) );
  OAI21_X1 U17372 ( .B1(n14013), .B2(n14012), .A(n14011), .ZN(n14018) );
  XOR2_X1 U17373 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n14014), .Z(
        n16081) );
  INV_X1 U17374 ( .A(n16081), .ZN(n14015) );
  AOI22_X1 U17375 ( .A1(n14330), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n14188), .B2(n14015), .ZN(n14017) );
  NAND2_X1 U17376 ( .A1(n14331), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n14016) );
  INV_X1 U17377 ( .A(n14944), .ZN(n14022) );
  AOI22_X1 U17378 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14027) );
  AOI22_X1 U17379 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U17380 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14025) );
  AOI22_X1 U17381 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14024) );
  NAND4_X1 U17382 ( .A1(n14027), .A2(n14026), .A3(n14025), .A4(n14024), .ZN(
        n14033) );
  AOI22_X1 U17383 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U17384 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17385 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14029) );
  AOI22_X1 U17386 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14028) );
  NAND4_X1 U17387 ( .A1(n14031), .A2(n14030), .A3(n14029), .A4(n14028), .ZN(
        n14032) );
  NOR2_X1 U17388 ( .A1(n14033), .A2(n14032), .ZN(n14036) );
  AOI21_X1 U17389 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14816), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14034) );
  AOI21_X1 U17390 ( .B1(n14331), .B2(P1_EAX_REG_16__SCAN_IN), .A(n14034), .ZN(
        n14035) );
  OAI21_X1 U17391 ( .B1(n14297), .B2(n14036), .A(n14035), .ZN(n14039) );
  XNOR2_X1 U17392 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B(n14037), .ZN(
        n16005) );
  NAND2_X1 U17393 ( .A1(n16005), .A2(n12918), .ZN(n14038) );
  NAND2_X1 U17394 ( .A1(n14039), .A2(n14038), .ZN(n14602) );
  XOR2_X1 U17395 ( .A(n14525), .B(n14040), .Z(n16068) );
  AOI22_X1 U17396 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U17397 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14043) );
  AOI22_X1 U17398 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14042) );
  AOI22_X1 U17399 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14041) );
  NAND4_X1 U17400 ( .A1(n14044), .A2(n14043), .A3(n14042), .A4(n14041), .ZN(
        n14050) );
  AOI22_X1 U17401 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14048) );
  AOI22_X1 U17402 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14047) );
  AOI22_X1 U17403 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U17404 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14045) );
  NAND4_X1 U17405 ( .A1(n14048), .A2(n14047), .A3(n14046), .A4(n14045), .ZN(
        n14049) );
  OR2_X1 U17406 ( .A1(n14050), .A2(n14049), .ZN(n14053) );
  OAI22_X1 U17407 ( .A1(n14294), .A2(n12899), .B1(n14051), .B2(n14525), .ZN(
        n14052) );
  AOI21_X1 U17408 ( .B1(n14324), .B2(n14053), .A(n14052), .ZN(n14054) );
  OAI21_X1 U17409 ( .B1(n16068), .B2(n14303), .A(n14054), .ZN(n14519) );
  XNOR2_X1 U17410 ( .A(n14055), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15987) );
  AOI22_X1 U17411 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14221), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U17412 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U17413 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14056), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14058) );
  AOI22_X1 U17414 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14057) );
  NAND4_X1 U17415 ( .A1(n14060), .A2(n14059), .A3(n14058), .A4(n14057), .ZN(
        n14066) );
  AOI22_X1 U17416 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U17417 ( .A1(n14308), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U17418 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U17419 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14061) );
  NAND4_X1 U17420 ( .A1(n14064), .A2(n14063), .A3(n14062), .A4(n14061), .ZN(
        n14065) );
  OAI21_X1 U17421 ( .B1(n14066), .B2(n14065), .A(n14324), .ZN(n14070) );
  INV_X1 U17422 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14067) );
  OAI22_X1 U17423 ( .A1(n14294), .A2(n12901), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14067), .ZN(n14068) );
  INV_X1 U17424 ( .A(n14068), .ZN(n14069) );
  AOI21_X1 U17425 ( .B1(n14070), .B2(n14069), .A(n14188), .ZN(n14071) );
  AOI21_X1 U17426 ( .B1(n15987), .B2(n14188), .A(n14071), .ZN(n14593) );
  AOI22_X1 U17427 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14126), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14075) );
  AOI22_X1 U17428 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14074) );
  AOI22_X1 U17429 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14073) );
  AOI22_X1 U17430 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14072) );
  NAND4_X1 U17431 ( .A1(n14075), .A2(n14074), .A3(n14073), .A4(n14072), .ZN(
        n14081) );
  AOI22_X1 U17432 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14079) );
  AOI22_X1 U17433 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17434 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U17435 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14076) );
  NAND4_X1 U17436 ( .A1(n14079), .A2(n14078), .A3(n14077), .A4(n14076), .ZN(
        n14080) );
  NOR2_X1 U17437 ( .A1(n14081), .A2(n14080), .ZN(n14084) );
  OAI21_X1 U17438 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20453), .A(
        n12842), .ZN(n14083) );
  NAND2_X1 U17439 ( .A1(n14331), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n14082) );
  OAI211_X1 U17440 ( .C1(n14297), .C2(n14084), .A(n14083), .B(n14082), .ZN(
        n14087) );
  OAI21_X1 U17441 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n14085), .A(
        n14102), .ZN(n16062) );
  OR2_X1 U17442 ( .A1(n14303), .A2(n16062), .ZN(n14086) );
  NAND2_X1 U17443 ( .A1(n14087), .A2(n14086), .ZN(n14588) );
  AOI22_X1 U17444 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17445 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n14126), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U17446 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14221), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U17447 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14089) );
  NAND4_X1 U17448 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14098) );
  AOI22_X1 U17449 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n14006), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U17450 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11845), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17451 ( .A1(n11833), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U17452 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n14192), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14093) );
  NAND4_X1 U17453 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        n14097) );
  NOR2_X1 U17454 ( .A1(n14098), .A2(n14097), .ZN(n14101) );
  OAI21_X1 U17455 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15971), .A(n14303), 
        .ZN(n14099) );
  AOI21_X1 U17456 ( .B1(n14331), .B2(P1_EAX_REG_20__SCAN_IN), .A(n14099), .ZN(
        n14100) );
  OAI21_X1 U17457 ( .B1(n14297), .B2(n14101), .A(n14100), .ZN(n14104) );
  XNOR2_X1 U17458 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n14102), .ZN(
        n16052) );
  NAND2_X1 U17459 ( .A1(n14188), .A2(n16052), .ZN(n14103) );
  AOI22_X1 U17460 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14221), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U17461 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17462 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U17463 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14106) );
  NAND4_X1 U17464 ( .A1(n14109), .A2(n14108), .A3(n14107), .A4(n14106), .ZN(
        n14115) );
  AOI22_X1 U17465 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17466 ( .A1(n14308), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U17467 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U17468 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14110) );
  NAND4_X1 U17469 ( .A1(n14113), .A2(n14112), .A3(n14111), .A4(n14110), .ZN(
        n14114) );
  NOR2_X1 U17470 ( .A1(n14115), .A2(n14114), .ZN(n14118) );
  OAI21_X1 U17471 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20453), .A(
        n12842), .ZN(n14117) );
  NAND2_X1 U17472 ( .A1(n14331), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n14116) );
  OAI211_X1 U17473 ( .C1(n14297), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        n14121) );
  OAI21_X1 U17474 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n14119), .A(
        n14136), .ZN(n16051) );
  OR2_X1 U17475 ( .A1(n14303), .A2(n16051), .ZN(n14120) );
  NAND2_X1 U17476 ( .A1(n14571), .A2(n14572), .ZN(n14562) );
  INV_X2 U17477 ( .A(n14562), .ZN(n14141) );
  AOI22_X1 U17478 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17479 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14124) );
  AOI22_X1 U17480 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14239), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U17481 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14122) );
  NAND4_X1 U17482 ( .A1(n14125), .A2(n14124), .A3(n14123), .A4(n14122), .ZN(
        n14132) );
  AOI22_X1 U17483 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14130) );
  AOI22_X1 U17484 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14129) );
  AOI22_X1 U17485 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14128) );
  AOI22_X1 U17486 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14127) );
  NAND4_X1 U17487 ( .A1(n14130), .A2(n14129), .A3(n14128), .A4(n14127), .ZN(
        n14131) );
  NOR2_X1 U17488 ( .A1(n14132), .A2(n14131), .ZN(n14135) );
  INV_X1 U17489 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20900) );
  AOI21_X1 U17490 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20900), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14133) );
  AOI21_X1 U17491 ( .B1(n14331), .B2(P1_EAX_REG_22__SCAN_IN), .A(n14133), .ZN(
        n14134) );
  OAI21_X1 U17492 ( .B1(n14297), .B2(n14135), .A(n14134), .ZN(n14139) );
  NAND2_X1 U17493 ( .A1(n20900), .A2(n14136), .ZN(n14137) );
  AND2_X1 U17494 ( .A1(n14137), .A2(n14167), .ZN(n15944) );
  NAND2_X1 U17495 ( .A1(n15944), .A2(n12918), .ZN(n14138) );
  NAND2_X1 U17496 ( .A1(n14139), .A2(n14138), .ZN(n14563) );
  AOI22_X1 U17497 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14105), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U17498 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U17499 ( .A1(n14192), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17500 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14142) );
  NAND4_X1 U17501 ( .A1(n14145), .A2(n14144), .A3(n14143), .A4(n14142), .ZN(
        n14151) );
  AOI22_X1 U17502 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U17503 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9759), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17504 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17505 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14146) );
  NAND4_X1 U17506 ( .A1(n14149), .A2(n14148), .A3(n14147), .A4(n14146), .ZN(
        n14150) );
  NOR2_X1 U17507 ( .A1(n14151), .A2(n14150), .ZN(n14171) );
  AOI22_X1 U17508 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14221), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U17509 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U17510 ( .A1(n14314), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17511 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11846), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14152) );
  NAND4_X1 U17512 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14161) );
  AOI22_X1 U17513 ( .A1(n9758), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U17514 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U17515 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14157) );
  AOI22_X1 U17516 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14156) );
  NAND4_X1 U17517 ( .A1(n14159), .A2(n14158), .A3(n14157), .A4(n14156), .ZN(
        n14160) );
  NOR2_X1 U17518 ( .A1(n14161), .A2(n14160), .ZN(n14172) );
  XNOR2_X1 U17519 ( .A(n14171), .B(n14172), .ZN(n14165) );
  NAND2_X1 U17520 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14162) );
  OAI211_X1 U17521 ( .C1(n14294), .C2(n12905), .A(n14303), .B(n14162), .ZN(
        n14163) );
  INV_X1 U17522 ( .A(n14163), .ZN(n14164) );
  OAI21_X1 U17523 ( .B1(n14297), .B2(n14165), .A(n14164), .ZN(n14170) );
  INV_X1 U17524 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14166) );
  NAND2_X1 U17525 ( .A1(n14167), .A2(n14166), .ZN(n14168) );
  AND2_X1 U17526 ( .A1(n14187), .A2(n14168), .ZN(n14792) );
  NAND2_X1 U17527 ( .A1(n14792), .A2(n12918), .ZN(n14169) );
  NAND2_X1 U17528 ( .A1(n14170), .A2(n14169), .ZN(n14503) );
  NOR2_X1 U17529 ( .A1(n14172), .A2(n14171), .ZN(n14204) );
  AOI22_X1 U17530 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14176) );
  AOI22_X1 U17531 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U17532 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U17533 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14173) );
  NAND4_X1 U17534 ( .A1(n14176), .A2(n14175), .A3(n14174), .A4(n14173), .ZN(
        n14182) );
  AOI22_X1 U17535 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14180) );
  AOI22_X1 U17536 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U17537 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14178) );
  AOI22_X1 U17538 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14177) );
  NAND4_X1 U17539 ( .A1(n14180), .A2(n14179), .A3(n14178), .A4(n14177), .ZN(
        n14181) );
  OR2_X1 U17540 ( .A1(n14182), .A2(n14181), .ZN(n14203) );
  INV_X1 U17541 ( .A(n14203), .ZN(n14183) );
  XNOR2_X1 U17542 ( .A(n14204), .B(n14183), .ZN(n14184) );
  NAND2_X1 U17543 ( .A1(n14184), .A2(n14324), .ZN(n14191) );
  NAND2_X1 U17544 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14185) );
  OAI211_X1 U17545 ( .C1(n14294), .C2(n12811), .A(n14303), .B(n14185), .ZN(
        n14186) );
  INV_X1 U17546 ( .A(n14186), .ZN(n14190) );
  XNOR2_X1 U17547 ( .A(n14187), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14784) );
  AOI21_X1 U17548 ( .B1(n14191), .B2(n14190), .A(n14189), .ZN(n14492) );
  AOI22_X1 U17549 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U17550 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14195) );
  AOI22_X1 U17551 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U17552 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14193) );
  NAND4_X1 U17553 ( .A1(n14196), .A2(n14195), .A3(n14194), .A4(n14193), .ZN(
        n14202) );
  AOI22_X1 U17554 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14200) );
  AOI22_X1 U17555 ( .A1(n14239), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14199) );
  AOI22_X1 U17556 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14198) );
  AOI22_X1 U17557 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14023), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14197) );
  NAND4_X1 U17558 ( .A1(n14200), .A2(n14199), .A3(n14198), .A4(n14197), .ZN(
        n14201) );
  NOR2_X1 U17559 ( .A1(n14202), .A2(n14201), .ZN(n14216) );
  NAND2_X1 U17560 ( .A1(n14204), .A2(n14203), .ZN(n14215) );
  XNOR2_X1 U17561 ( .A(n14216), .B(n14215), .ZN(n14208) );
  NAND2_X1 U17562 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14205) );
  OAI211_X1 U17563 ( .C1(n14294), .C2(n12805), .A(n14303), .B(n14205), .ZN(
        n14206) );
  INV_X1 U17564 ( .A(n14206), .ZN(n14207) );
  OAI21_X1 U17565 ( .B1(n14208), .B2(n14297), .A(n14207), .ZN(n14214) );
  INV_X1 U17566 ( .A(n14209), .ZN(n14211) );
  INV_X1 U17567 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14210) );
  NAND2_X1 U17568 ( .A1(n14211), .A2(n14210), .ZN(n14212) );
  NAND2_X1 U17569 ( .A1(n14232), .A2(n14212), .ZN(n14777) );
  NOR2_X1 U17570 ( .A1(n14216), .A2(n14215), .ZN(n14247) );
  AOI22_X1 U17571 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14220) );
  AOI22_X1 U17572 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14219) );
  AOI22_X1 U17573 ( .A1(n14126), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14218) );
  AOI22_X1 U17574 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14217) );
  NAND4_X1 U17575 ( .A1(n14220), .A2(n14219), .A3(n14218), .A4(n14217), .ZN(
        n14227) );
  AOI22_X1 U17576 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9767), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14225) );
  AOI22_X1 U17577 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14224) );
  AOI22_X1 U17578 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14223) );
  AOI22_X1 U17579 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14222) );
  NAND4_X1 U17580 ( .A1(n14225), .A2(n14224), .A3(n14223), .A4(n14222), .ZN(
        n14226) );
  OR2_X1 U17581 ( .A1(n14227), .A2(n14226), .ZN(n14246) );
  XNOR2_X1 U17582 ( .A(n14247), .B(n14246), .ZN(n14231) );
  NAND2_X1 U17583 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14228) );
  OAI211_X1 U17584 ( .C1(n14294), .C2(n12809), .A(n14303), .B(n14228), .ZN(
        n14229) );
  INV_X1 U17585 ( .A(n14229), .ZN(n14230) );
  OAI21_X1 U17586 ( .B1(n14231), .B2(n14297), .A(n14230), .ZN(n14234) );
  XNOR2_X1 U17587 ( .A(n14232), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14468) );
  NAND2_X1 U17588 ( .A1(n14468), .A2(n12918), .ZN(n14233) );
  NAND2_X1 U17589 ( .A1(n14234), .A2(n14233), .ZN(n14467) );
  AOI22_X1 U17590 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n14006), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U17591 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U17592 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U17593 ( .A1(n14314), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14235) );
  NAND4_X1 U17594 ( .A1(n14238), .A2(n14237), .A3(n14236), .A4(n14235), .ZN(
        n14245) );
  AOI22_X1 U17595 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11845), .B1(
        n9760), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14243) );
  AOI22_X1 U17596 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14239), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U17597 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n14221), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U17598 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14240) );
  NAND4_X1 U17599 ( .A1(n14243), .A2(n14242), .A3(n14241), .A4(n14240), .ZN(
        n14244) );
  NOR2_X1 U17600 ( .A1(n14245), .A2(n14244), .ZN(n14260) );
  NAND2_X1 U17601 ( .A1(n14247), .A2(n14246), .ZN(n14259) );
  XNOR2_X1 U17602 ( .A(n14260), .B(n14259), .ZN(n14251) );
  NAND2_X1 U17603 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14248) );
  OAI211_X1 U17604 ( .C1(n14294), .C2(n12807), .A(n14303), .B(n14248), .ZN(
        n14249) );
  INV_X1 U17605 ( .A(n14249), .ZN(n14250) );
  OAI21_X1 U17606 ( .B1(n14251), .B2(n14297), .A(n14250), .ZN(n14257) );
  INV_X1 U17607 ( .A(n14252), .ZN(n14254) );
  INV_X1 U17608 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U17609 ( .A1(n14254), .A2(n14253), .ZN(n14255) );
  NAND2_X1 U17610 ( .A1(n14276), .A2(n14255), .ZN(n14761) );
  NAND2_X1 U17611 ( .A1(n14257), .A2(n14256), .ZN(n14453) );
  NOR2_X1 U17612 ( .A1(n14260), .A2(n14259), .ZN(n14292) );
  AOI22_X1 U17613 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11777), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14264) );
  AOI22_X1 U17614 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14263) );
  AOI22_X1 U17615 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14262) );
  AOI22_X1 U17616 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14261) );
  NAND4_X1 U17617 ( .A1(n14264), .A2(n14263), .A3(n14262), .A4(n14261), .ZN(
        n14271) );
  AOI22_X1 U17618 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9768), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14269) );
  AOI22_X1 U17619 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14268) );
  AOI22_X1 U17620 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14267) );
  AOI22_X1 U17621 ( .A1(n11833), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14266) );
  NAND4_X1 U17622 ( .A1(n14269), .A2(n14268), .A3(n14267), .A4(n14266), .ZN(
        n14270) );
  OR2_X1 U17623 ( .A1(n14271), .A2(n14270), .ZN(n14291) );
  XNOR2_X1 U17624 ( .A(n14292), .B(n14291), .ZN(n14275) );
  NAND2_X1 U17625 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14272) );
  OAI211_X1 U17626 ( .C1(n14294), .C2(n12801), .A(n14303), .B(n14272), .ZN(
        n14273) );
  INV_X1 U17627 ( .A(n14273), .ZN(n14274) );
  OAI21_X1 U17628 ( .B1(n14275), .B2(n14297), .A(n14274), .ZN(n14278) );
  XNOR2_X1 U17629 ( .A(n14276), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14747) );
  NAND2_X1 U17630 ( .A1(n14747), .A2(n12918), .ZN(n14277) );
  NAND2_X1 U17631 ( .A1(n14278), .A2(n14277), .ZN(n14440) );
  AOI22_X1 U17632 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14126), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U17633 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U17634 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14280) );
  AOI22_X1 U17635 ( .A1(n9768), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14279) );
  NAND4_X1 U17636 ( .A1(n14282), .A2(n14281), .A3(n14280), .A4(n14279), .ZN(
        n14290) );
  AOI22_X1 U17637 ( .A1(n14283), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14288) );
  AOI22_X1 U17638 ( .A1(n14284), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14287) );
  AOI22_X1 U17639 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14286) );
  AOI22_X1 U17640 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14285) );
  NAND4_X1 U17641 ( .A1(n14288), .A2(n14287), .A3(n14286), .A4(n14285), .ZN(
        n14289) );
  NOR2_X1 U17642 ( .A1(n14290), .A2(n14289), .ZN(n14307) );
  NAND2_X1 U17643 ( .A1(n14292), .A2(n14291), .ZN(n14306) );
  XNOR2_X1 U17644 ( .A(n14307), .B(n14306), .ZN(n14298) );
  NAND2_X1 U17645 ( .A1(n12842), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14293) );
  OAI211_X1 U17646 ( .C1(n14294), .C2(n12799), .A(n14303), .B(n14293), .ZN(
        n14295) );
  INV_X1 U17647 ( .A(n14295), .ZN(n14296) );
  OAI21_X1 U17648 ( .B1(n14298), .B2(n14297), .A(n14296), .ZN(n14305) );
  INV_X1 U17649 ( .A(n14299), .ZN(n14301) );
  INV_X1 U17650 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14300) );
  NAND2_X1 U17651 ( .A1(n14301), .A2(n14300), .ZN(n14302) );
  NAND2_X1 U17652 ( .A1(n14327), .A2(n14302), .ZN(n14736) );
  NOR2_X1 U17653 ( .A1(n14307), .A2(n14306), .ZN(n14323) );
  AOI22_X1 U17654 ( .A1(n14006), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14126), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U17655 ( .A1(n11845), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14308), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U17656 ( .A1(n9767), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U17657 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11703), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14309) );
  NAND4_X1 U17658 ( .A1(n14312), .A2(n14311), .A3(n14310), .A4(n14309), .ZN(
        n14321) );
  AOI22_X1 U17659 ( .A1(n14105), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14284), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U17660 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14192), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U17661 ( .A1(n9761), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14313), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U17662 ( .A1(n14221), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14314), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14316) );
  NAND4_X1 U17663 ( .A1(n14319), .A2(n14318), .A3(n14317), .A4(n14316), .ZN(
        n14320) );
  NOR2_X1 U17664 ( .A1(n14321), .A2(n14320), .ZN(n14322) );
  XNOR2_X1 U17665 ( .A(n14323), .B(n14322), .ZN(n14325) );
  NAND2_X1 U17666 ( .A1(n14325), .A2(n14324), .ZN(n14329) );
  NOR2_X1 U17667 ( .A1(n20999), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14326) );
  AOI211_X1 U17668 ( .C1(n14331), .C2(P1_EAX_REG_30__SCAN_IN), .A(n14326), .B(
        n12918), .ZN(n14328) );
  XNOR2_X1 U17669 ( .A(n14327), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14727) );
  AOI22_X1 U17670 ( .A1(n14329), .A2(n14328), .B1(n14727), .B2(n12918), .ZN(
        n14414) );
  AOI22_X1 U17671 ( .A1(n14331), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n14330), .ZN(n14332) );
  NAND2_X1 U17672 ( .A1(n14384), .A2(n20154), .ZN(n14350) );
  INV_X1 U17673 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20719) );
  INV_X1 U17674 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14418) );
  NOR2_X1 U17675 ( .A1(n20719), .A2(n14418), .ZN(n14345) );
  INV_X1 U17676 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15951) );
  INV_X1 U17677 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14520) );
  INV_X1 U17678 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20697) );
  NAND3_X1 U17679 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n16026), .ZN(n14542) );
  NOR2_X1 U17680 ( .A1(n20697), .A2(n14542), .ZN(n16015) );
  NAND2_X1 U17681 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16015), .ZN(n15992) );
  NAND2_X1 U17682 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15997) );
  NOR3_X1 U17683 ( .A1(n14520), .A2(n15992), .A3(n15997), .ZN(n15963) );
  NAND4_X1 U17684 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15963), .A3(
        P1_REIP_REG_18__SCAN_IN), .A4(P1_REIP_REG_19__SCAN_IN), .ZN(n15957) );
  NOR2_X1 U17685 ( .A1(n15951), .A2(n15957), .ZN(n15943) );
  NAND2_X1 U17686 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15943), .ZN(n14508) );
  INV_X1 U17687 ( .A(n14508), .ZN(n14335) );
  AND2_X1 U17688 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14335), .ZN(n14494) );
  OR2_X1 U17689 ( .A1(n20152), .A2(n14494), .ZN(n14336) );
  NAND2_X1 U17690 ( .A1(n14336), .A2(n15994), .ZN(n14516) );
  NOR2_X1 U17691 ( .A1(n20152), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14337) );
  NOR2_X1 U17692 ( .A1(n14516), .A2(n14337), .ZN(n14483) );
  AND2_X1 U17693 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14341) );
  OR2_X1 U17694 ( .A1(n20152), .A2(n14341), .ZN(n14338) );
  AND2_X1 U17695 ( .A1(n14483), .A2(n14338), .ZN(n14472) );
  NAND2_X1 U17696 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14343) );
  NAND2_X1 U17697 ( .A1(n15996), .A2(n14343), .ZN(n14339) );
  AND2_X1 U17698 ( .A1(n14472), .A2(n14339), .ZN(n14446) );
  OAI21_X1 U17699 ( .B1(n14345), .B2(n20152), .A(n14446), .ZN(n14419) );
  INV_X1 U17700 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14552) );
  INV_X1 U17701 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14382) );
  OAI22_X1 U17702 ( .A1(n14552), .A2(n20136), .B1(n20162), .B2(n14382), .ZN(
        n14348) );
  NAND2_X1 U17703 ( .A1(n14494), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14340) );
  OR2_X1 U17704 ( .A1(n20152), .A2(n14340), .ZN(n14487) );
  INV_X1 U17705 ( .A(n14341), .ZN(n14342) );
  NOR2_X1 U17706 ( .A1(n14487), .A2(n14342), .ZN(n14459) );
  INV_X1 U17707 ( .A(n14343), .ZN(n14344) );
  NAND2_X1 U17708 ( .A1(n14459), .A2(n14344), .ZN(n14434) );
  INV_X1 U17709 ( .A(n14345), .ZN(n14346) );
  NOR3_X1 U17710 ( .A1(n14434), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14346), 
        .ZN(n14347) );
  AOI211_X1 U17711 ( .C1(n14419), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14348), 
        .B(n14347), .ZN(n14349) );
  OAI211_X1 U17712 ( .C1(n14553), .C2(n20175), .A(n14350), .B(n14349), .ZN(
        P1_U2809) );
  INV_X1 U17713 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n14357) );
  AND2_X1 U17714 ( .A1(n16046), .A2(n14351), .ZN(n14352) );
  AOI22_X1 U17715 ( .A1(n14713), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14724), .ZN(n14355) );
  OAI211_X1 U17716 ( .C1(n14717), .C2(n14357), .A(n14356), .B(n14355), .ZN(
        P1_U2873) );
  NAND2_X1 U17717 ( .A1(n14358), .A2(n19391), .ZN(n14372) );
  INV_X1 U17718 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n16276) );
  NAND2_X1 U17719 ( .A1(n11525), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14360) );
  NAND2_X1 U17720 ( .A1(n11554), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n14359) );
  OAI211_X1 U17721 ( .C1(n14361), .C2(n16276), .A(n14360), .B(n14359), .ZN(
        n14362) );
  NAND2_X1 U17722 ( .A1(n19241), .A2(n16474), .ZN(n14369) );
  AND2_X1 U17723 ( .A1(n16479), .A2(n14370), .ZN(n14364) );
  OAI21_X1 U17724 ( .B1(n14365), .B2(n14364), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14367) );
  AND2_X1 U17725 ( .A1(n14367), .A2(n14366), .ZN(n14368) );
  XOR2_X1 U17726 ( .A(n12982), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14375)
         );
  MUX2_X1 U17727 ( .A(n19198), .B(n19199), .S(n15159), .Z(n14374) );
  OAI21_X1 U17728 ( .B1(n14375), .B2(n15185), .A(n14374), .ZN(P2_U2882) );
  MUX2_X1 U17729 ( .A(n14377), .B(n14376), .S(n15159), .Z(n14378) );
  OAI21_X1 U17730 ( .B1(n19216), .B2(n15185), .A(n14378), .ZN(P2_U2883) );
  NAND2_X1 U17731 ( .A1(n16114), .A2(n14379), .ZN(n14381) );
  OAI211_X1 U17732 ( .C1(n14382), .C2(n16120), .A(n14381), .B(n14380), .ZN(
        n14383) );
  OAI21_X1 U17733 ( .B1(n14386), .B2(n20100), .A(n14385), .ZN(P1_U2968) );
  INV_X1 U17734 ( .A(n14387), .ZN(n14388) );
  XNOR2_X1 U17735 ( .A(n14389), .B(n14388), .ZN(n19396) );
  NOR2_X1 U17736 ( .A1(n16424), .A2(n15061), .ZN(n14396) );
  INV_X1 U17737 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14394) );
  AOI21_X1 U17738 ( .B1(n14392), .B2(n14391), .A(n14390), .ZN(n19392) );
  AOI22_X1 U17739 ( .A1(n19392), .A2(n16435), .B1(P2_REIP_REG_2__SCAN_IN), 
        .B2(n19180), .ZN(n14393) );
  OAI21_X1 U17740 ( .B1(n14394), .B2(n16445), .A(n14393), .ZN(n14395) );
  AOI211_X1 U17741 ( .C1(n19396), .C2(n16441), .A(n14396), .B(n14395), .ZN(
        n14397) );
  OAI21_X1 U17742 ( .B1(n10769), .B2(n16439), .A(n14397), .ZN(P2_U3012) );
  NAND2_X1 U17743 ( .A1(n14398), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14400)
         );
  NAND3_X1 U17744 ( .A1(n14400), .A2(n14399), .A3(n20097), .ZN(P1_U2801) );
  AOI21_X1 U17745 ( .B1(n14401), .B2(n12173), .A(n15907), .ZN(n14402) );
  INV_X1 U17746 ( .A(n14402), .ZN(n14405) );
  NAND2_X1 U17747 ( .A1(n14403), .A2(n15907), .ZN(n14404) );
  OAI211_X1 U17748 ( .C1(n14406), .C2(n12166), .A(n14405), .B(n14404), .ZN(
        n15893) );
  INV_X1 U17749 ( .A(n14407), .ZN(n14409) );
  AOI22_X1 U17750 ( .A1(n14409), .A2(n12173), .B1(n14408), .B2(n14411), .ZN(
        n20093) );
  NAND3_X1 U17751 ( .A1(n14411), .A2(n15930), .A3(n14410), .ZN(n14412) );
  NAND2_X1 U17752 ( .A1(n14412), .A2(n20747), .ZN(n20743) );
  NAND2_X1 U17753 ( .A1(n20093), .A2(n20743), .ZN(n15891) );
  AND2_X1 U17754 ( .A1(n15891), .A2(n14413), .ZN(n20102) );
  MUX2_X1 U17755 ( .A(P1_MORE_REG_SCAN_IN), .B(n15893), .S(n20102), .Z(
        P1_U3484) );
  INV_X1 U17756 ( .A(n14730), .ZN(n14631) );
  OAI22_X1 U17757 ( .A1(n14426), .A2(n12179), .B1(n14415), .B2(n14441), .ZN(
        n14417) );
  XNOR2_X1 U17758 ( .A(n14417), .B(n14416), .ZN(n14848) );
  INV_X1 U17759 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14555) );
  NOR2_X1 U17760 ( .A1(n14434), .A2(n14418), .ZN(n14420) );
  OAI21_X1 U17761 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14420), .A(n14419), 
        .ZN(n14422) );
  AOI22_X1 U17762 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n14727), .ZN(n14421) );
  OAI211_X1 U17763 ( .C1(n20136), .C2(n14555), .A(n14422), .B(n14421), .ZN(
        n14423) );
  AOI21_X1 U17764 ( .B1(n14848), .B2(n20159), .A(n14423), .ZN(n14424) );
  OAI21_X1 U17765 ( .B1(n14631), .B2(n20141), .A(n14424), .ZN(P1_U2810) );
  AND2_X1 U17766 ( .A1(n14441), .A2(n14425), .ZN(n14427) );
  INV_X1 U17767 ( .A(n14428), .ZN(n14430) );
  NAND2_X1 U17768 ( .A1(n14738), .A2(n20154), .ZN(n14438) );
  INV_X1 U17769 ( .A(n14446), .ZN(n14436) );
  INV_X1 U17770 ( .A(n14736), .ZN(n14431) );
  AOI22_X1 U17771 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n14431), .ZN(n14433) );
  OR2_X1 U17772 ( .A1(n20136), .A2(n14556), .ZN(n14432) );
  OAI211_X1 U17773 ( .C1(n14434), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14433), 
        .B(n14432), .ZN(n14435) );
  AOI21_X1 U17774 ( .B1(n14436), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14435), 
        .ZN(n14437) );
  OAI211_X1 U17775 ( .C1(n20175), .C2(n14855), .A(n14438), .B(n14437), .ZN(
        P1_U2811) );
  AOI21_X1 U17776 ( .B1(n14440), .B2(n14439), .A(n14428), .ZN(n14751) );
  INV_X1 U17777 ( .A(n14751), .ZN(n14647) );
  AOI21_X1 U17778 ( .B1(n14442), .B2(n9788), .A(n10068), .ZN(n14867) );
  AOI21_X1 U17779 ( .B1(n14459), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14445) );
  AOI22_X1 U17780 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n14747), .ZN(n14444) );
  NAND2_X1 U17781 ( .A1(n20170), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14443) );
  OAI211_X1 U17782 ( .C1(n14446), .C2(n14445), .A(n14444), .B(n14443), .ZN(
        n14447) );
  AOI21_X1 U17783 ( .B1(n14867), .B2(n20159), .A(n14447), .ZN(n14448) );
  OAI21_X1 U17784 ( .B1(n14647), .B2(n20141), .A(n14448), .ZN(P1_U2812) );
  OR2_X1 U17785 ( .A1(n14464), .A2(n14449), .ZN(n14450) );
  NAND2_X1 U17786 ( .A1(n9788), .A2(n14450), .ZN(n14878) );
  INV_X1 U17787 ( .A(n14439), .ZN(n14452) );
  AOI21_X1 U17788 ( .B1(n14453), .B2(n14466), .A(n14452), .ZN(n14763) );
  NAND2_X1 U17789 ( .A1(n14763), .A2(n20154), .ZN(n14461) );
  INV_X1 U17790 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14458) );
  INV_X1 U17791 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n20840) );
  INV_X1 U17792 ( .A(n14761), .ZN(n14454) );
  AOI22_X1 U17793 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n14454), .ZN(n14455) );
  OAI21_X1 U17794 ( .B1(n20136), .B2(n20840), .A(n14455), .ZN(n14457) );
  NOR2_X1 U17795 ( .A1(n14472), .A2(n14458), .ZN(n14456) );
  AOI211_X1 U17796 ( .C1(n14459), .C2(n14458), .A(n14457), .B(n14456), .ZN(
        n14460) );
  OAI211_X1 U17797 ( .C1(n20175), .C2(n14878), .A(n14461), .B(n14460), .ZN(
        P1_U2813) );
  NOR2_X1 U17798 ( .A1(n14478), .A2(n14462), .ZN(n14463) );
  OR2_X1 U17799 ( .A1(n14464), .A2(n14463), .ZN(n16121) );
  AOI21_X1 U17800 ( .B1(n14467), .B2(n14465), .A(n14451), .ZN(n14770) );
  NAND2_X1 U17801 ( .A1(n14770), .A2(n20154), .ZN(n14476) );
  INV_X1 U17802 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14469) );
  INV_X1 U17803 ( .A(n14468), .ZN(n14768) );
  OAI22_X1 U17804 ( .A1(n14469), .A2(n20162), .B1(n20186), .B2(n14768), .ZN(
        n14474) );
  INV_X1 U17805 ( .A(n14487), .ZN(n14470) );
  AOI21_X1 U17806 ( .B1(n14470), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_26__SCAN_IN), .ZN(n14471) );
  NOR2_X1 U17807 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  AOI211_X1 U17808 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20170), .A(n14474), .B(
        n14473), .ZN(n14475) );
  OAI211_X1 U17809 ( .C1(n20175), .C2(n16121), .A(n14476), .B(n14475), .ZN(
        P1_U2814) );
  AND2_X1 U17810 ( .A1(n14498), .A2(n14477), .ZN(n14479) );
  OR2_X1 U17811 ( .A1(n14479), .A2(n14478), .ZN(n16131) );
  OAI21_X1 U17812 ( .B1(n14480), .B2(n14482), .A(n14465), .ZN(n14664) );
  INV_X1 U17813 ( .A(n14664), .ZN(n14779) );
  NAND2_X1 U17814 ( .A1(n14779), .A2(n20154), .ZN(n14491) );
  INV_X1 U17815 ( .A(n14483), .ZN(n14489) );
  INV_X1 U17816 ( .A(n14777), .ZN(n14484) );
  AOI22_X1 U17817 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n14484), .ZN(n14486) );
  INV_X1 U17818 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14559) );
  OR2_X1 U17819 ( .A1(n20136), .A2(n14559), .ZN(n14485) );
  OAI211_X1 U17820 ( .C1(n14487), .C2(P1_REIP_REG_25__SCAN_IN), .A(n14486), 
        .B(n14485), .ZN(n14488) );
  AOI21_X1 U17821 ( .B1(n14489), .B2(P1_REIP_REG_25__SCAN_IN), .A(n14488), 
        .ZN(n14490) );
  OAI211_X1 U17822 ( .C1(n20175), .C2(n16131), .A(n14491), .B(n14490), .ZN(
        P1_U2815) );
  AOI21_X1 U17823 ( .B1(n10142), .B2(n9779), .A(n14480), .ZN(n14788) );
  INV_X1 U17824 ( .A(n14788), .ZN(n14669) );
  INV_X1 U17825 ( .A(n20152), .ZN(n16016) );
  INV_X1 U17826 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14493) );
  NAND3_X1 U17827 ( .A1(n16016), .A2(n14494), .A3(n14493), .ZN(n14496) );
  AOI22_X1 U17828 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n14784), .ZN(n14495) );
  OAI211_X1 U17829 ( .C1(n12255), .C2(n20136), .A(n14496), .B(n14495), .ZN(
        n14497) );
  AOI21_X1 U17830 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14516), .A(n14497), 
        .ZN(n14502) );
  INV_X1 U17831 ( .A(n14498), .ZN(n14499) );
  AOI21_X1 U17832 ( .B1(n14500), .B2(n14512), .A(n14499), .ZN(n14890) );
  NAND2_X1 U17833 ( .A1(n14890), .A2(n20159), .ZN(n14501) );
  OAI211_X1 U17834 ( .C1(n14669), .C2(n20141), .A(n14502), .B(n14501), .ZN(
        P1_U2816) );
  INV_X1 U17835 ( .A(n14503), .ZN(n14506) );
  INV_X1 U17836 ( .A(n14504), .ZN(n14505) );
  INV_X1 U17837 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14507) );
  OAI21_X1 U17838 ( .B1(n20152), .B2(n14508), .A(n14507), .ZN(n14515) );
  INV_X1 U17839 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14561) );
  AOI22_X1 U17840 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n14792), .ZN(n14509) );
  OAI21_X1 U17841 ( .B1(n20136), .B2(n14561), .A(n14509), .ZN(n14514) );
  NAND2_X1 U17842 ( .A1(n14567), .A2(n14510), .ZN(n14511) );
  NAND2_X1 U17843 ( .A1(n14512), .A2(n14511), .ZN(n16142) );
  NOR2_X1 U17844 ( .A1(n16142), .A2(n20175), .ZN(n14513) );
  AOI211_X1 U17845 ( .C1(n14516), .C2(n14515), .A(n14514), .B(n14513), .ZN(
        n14517) );
  OAI21_X1 U17846 ( .B1(n14791), .B2(n20141), .A(n14517), .ZN(P1_U2817) );
  OAI21_X1 U17847 ( .B1(n14518), .B2(n14519), .A(n9817), .ZN(n14706) );
  NOR2_X1 U17848 ( .A1(n20152), .A2(n15992), .ZN(n16008) );
  INV_X1 U17849 ( .A(n16008), .ZN(n14521) );
  OAI21_X1 U17850 ( .B1(n15997), .B2(n14521), .A(n14520), .ZN(n14531) );
  OAI21_X1 U17851 ( .B1(n20152), .B2(n15963), .A(n15994), .ZN(n15986) );
  INV_X1 U17852 ( .A(n14605), .ZN(n14524) );
  INV_X1 U17853 ( .A(n14522), .ZN(n14523) );
  OAI21_X1 U17854 ( .B1(n14524), .B2(n14523), .A(n9816), .ZN(n16176) );
  OAI21_X1 U17855 ( .B1(n20162), .B2(n14525), .A(n9736), .ZN(n14528) );
  INV_X1 U17856 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14526) );
  NOR2_X1 U17857 ( .A1(n20136), .A2(n14526), .ZN(n14527) );
  AOI211_X1 U17858 ( .C1(n16068), .C2(n20126), .A(n14528), .B(n14527), .ZN(
        n14529) );
  OAI21_X1 U17859 ( .B1(n16176), .B2(n20175), .A(n14529), .ZN(n14530) );
  AOI21_X1 U17860 ( .B1(n14531), .B2(n15986), .A(n14530), .ZN(n14532) );
  OAI21_X1 U17861 ( .B1(n14706), .B2(n20141), .A(n14532), .ZN(P1_U2823) );
  INV_X1 U17862 ( .A(n13978), .ZN(n14533) );
  AOI21_X1 U17863 ( .B1(n14535), .B2(n14534), .A(n14533), .ZN(n14619) );
  INV_X1 U17864 ( .A(n14536), .ZN(n14618) );
  NOR2_X1 U17865 ( .A1(n14619), .A2(n14618), .ZN(n14617) );
  OAI21_X1 U17866 ( .B1(n14617), .B2(n14537), .A(n14021), .ZN(n14831) );
  OR2_X1 U17867 ( .A1(n14538), .A2(n14539), .ZN(n14540) );
  AND2_X1 U17868 ( .A1(n14541), .A2(n14540), .ZN(n16191) );
  INV_X1 U17869 ( .A(n14542), .ZN(n14544) );
  NAND2_X1 U17870 ( .A1(n15994), .A2(n14544), .ZN(n14543) );
  NAND2_X1 U17871 ( .A1(n15996), .A2(n14543), .ZN(n16035) );
  AOI22_X1 U17872 ( .A1(n20170), .A2(P1_EBX_REG_13__SCAN_IN), .B1(n20126), 
        .B2(n14828), .ZN(n14547) );
  NAND2_X1 U17873 ( .A1(n20697), .A2(n14544), .ZN(n14545) );
  OR2_X1 U17874 ( .A1(n20152), .A2(n14545), .ZN(n14546) );
  OAI211_X1 U17875 ( .C1(n16035), .C2(n20697), .A(n14547), .B(n14546), .ZN(
        n14550) );
  OAI21_X1 U17876 ( .B1(n20162), .B2(n14548), .A(n9736), .ZN(n14549) );
  AOI211_X1 U17877 ( .C1(n16191), .C2(n20159), .A(n14550), .B(n14549), .ZN(
        n14551) );
  OAI21_X1 U17878 ( .B1(n14831), .B2(n20141), .A(n14551), .ZN(P1_U2827) );
  OAI22_X1 U17879 ( .A1(n14553), .A2(n20194), .B1(n20204), .B2(n14552), .ZN(
        P1_U2841) );
  INV_X1 U17880 ( .A(n14848), .ZN(n14554) );
  OAI222_X1 U17881 ( .A1(n14624), .A2(n14631), .B1(n14555), .B2(n20204), .C1(
        n14554), .C2(n20194), .ZN(P1_U2842) );
  INV_X1 U17882 ( .A(n14738), .ZN(n14639) );
  OAI222_X1 U17883 ( .A1(n14624), .A2(n14639), .B1(n14556), .B2(n20204), .C1(
        n14855), .C2(n20194), .ZN(P1_U2843) );
  AOI22_X1 U17884 ( .A1(n14867), .A2(n20199), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14615), .ZN(n14557) );
  OAI21_X1 U17885 ( .B1(n14647), .B2(n14624), .A(n14557), .ZN(P1_U2844) );
  INV_X1 U17886 ( .A(n14763), .ZN(n14653) );
  OAI222_X1 U17887 ( .A1(n14624), .A2(n14653), .B1(n20840), .B2(n20204), .C1(
        n14878), .C2(n20194), .ZN(P1_U2845) );
  INV_X1 U17888 ( .A(n14770), .ZN(n14659) );
  OAI222_X1 U17889 ( .A1(n14624), .A2(n14659), .B1(n14558), .B2(n20204), .C1(
        n16121), .C2(n20194), .ZN(P1_U2846) );
  OAI222_X1 U17890 ( .A1(n14624), .A2(n14664), .B1(n14559), .B2(n20204), .C1(
        n16131), .C2(n20194), .ZN(P1_U2847) );
  AOI22_X1 U17891 ( .A1(n14890), .A2(n20199), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14615), .ZN(n14560) );
  OAI21_X1 U17892 ( .B1(n14669), .B2(n14624), .A(n14560), .ZN(P1_U2848) );
  OAI222_X1 U17893 ( .A1(n14791), .A2(n14624), .B1(n14561), .B2(n20204), .C1(
        n16142), .C2(n20194), .ZN(P1_U2849) );
  NAND2_X1 U17894 ( .A1(n14562), .A2(n14563), .ZN(n14564) );
  AND2_X1 U17895 ( .A1(n14504), .A2(n14564), .ZN(n15949) );
  OR2_X1 U17896 ( .A1(n9846), .A2(n14565), .ZN(n14566) );
  NAND2_X1 U17897 ( .A1(n14567), .A2(n14566), .ZN(n16149) );
  OAI22_X1 U17898 ( .A1(n16149), .A2(n20194), .B1(n14568), .B2(n20204), .ZN(
        n14569) );
  INV_X1 U17899 ( .A(n14569), .ZN(n14570) );
  OAI21_X1 U17900 ( .B1(n14805), .B2(n14624), .A(n14570), .ZN(P1_U2850) );
  OR2_X1 U17901 ( .A1(n14571), .A2(n14572), .ZN(n14573) );
  AND2_X1 U17902 ( .A1(n14562), .A2(n14573), .ZN(n16048) );
  INV_X1 U17903 ( .A(n16048), .ZN(n14686) );
  INV_X1 U17904 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14576) );
  AND2_X1 U17905 ( .A1(n14585), .A2(n14574), .ZN(n14575) );
  OR2_X1 U17906 ( .A1(n9846), .A2(n14575), .ZN(n15959) );
  OAI222_X1 U17907 ( .A1(n14686), .A2(n14624), .B1(n14576), .B2(n20204), .C1(
        n15959), .C2(n20194), .ZN(P1_U2851) );
  INV_X1 U17908 ( .A(n14577), .ZN(n14581) );
  INV_X1 U17909 ( .A(n14579), .ZN(n14580) );
  AOI21_X1 U17910 ( .B1(n14581), .B2(n14580), .A(n14571), .ZN(n16053) );
  INV_X1 U17911 ( .A(n16053), .ZN(n14692) );
  INV_X1 U17912 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14586) );
  INV_X1 U17913 ( .A(n14591), .ZN(n14583) );
  NAND2_X1 U17914 ( .A1(n14583), .A2(n10061), .ZN(n14584) );
  NAND2_X1 U17915 ( .A1(n14585), .A2(n14584), .ZN(n15965) );
  OAI222_X1 U17916 ( .A1(n14692), .A2(n14624), .B1(n14586), .B2(n20204), .C1(
        n15965), .C2(n20194), .ZN(P1_U2852) );
  AOI21_X1 U17917 ( .B1(n14588), .B2(n14595), .A(n14579), .ZN(n16059) );
  INV_X1 U17918 ( .A(n16059), .ZN(n14699) );
  AND2_X1 U17919 ( .A1(n14598), .A2(n14589), .ZN(n14590) );
  NOR2_X1 U17920 ( .A1(n14591), .A2(n14590), .ZN(n16157) );
  AOI22_X1 U17921 ( .A1(n16157), .A2(n20199), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14615), .ZN(n14592) );
  OAI21_X1 U17922 ( .B1(n14699), .B2(n14624), .A(n14592), .ZN(P1_U2853) );
  NAND2_X1 U17923 ( .A1(n9817), .A2(n14593), .ZN(n14594) );
  AND2_X1 U17924 ( .A1(n14595), .A2(n14594), .ZN(n15989) );
  NAND2_X1 U17925 ( .A1(n9816), .A2(n14596), .ZN(n14597) );
  NAND2_X1 U17926 ( .A1(n14598), .A2(n14597), .ZN(n16168) );
  OAI22_X1 U17927 ( .A1(n16168), .A2(n20194), .B1(n15983), .B2(n20204), .ZN(
        n14599) );
  AOI21_X1 U17928 ( .B1(n15989), .B2(n20200), .A(n14599), .ZN(n14600) );
  INV_X1 U17929 ( .A(n14600), .ZN(P1_U2854) );
  OAI222_X1 U17930 ( .A1(n16176), .A2(n20194), .B1(n14526), .B2(n20204), .C1(
        n14706), .C2(n14624), .ZN(P1_U2855) );
  INV_X1 U17931 ( .A(n14601), .ZN(n14608) );
  AOI21_X1 U17932 ( .B1(n14602), .B2(n14608), .A(n14518), .ZN(n16000) );
  OR2_X1 U17933 ( .A1(n14611), .A2(n14603), .ZN(n14604) );
  NAND2_X1 U17934 ( .A1(n14605), .A2(n14604), .ZN(n16001) );
  OAI22_X1 U17935 ( .A1(n16001), .A2(n20194), .B1(n15999), .B2(n20204), .ZN(
        n14606) );
  AOI21_X1 U17936 ( .B1(n16000), .B2(n20200), .A(n14606), .ZN(n14607) );
  INV_X1 U17937 ( .A(n14607), .ZN(P1_U2856) );
  AOI21_X1 U17938 ( .B1(n14610), .B2(n14609), .A(n14601), .ZN(n16082) );
  INV_X1 U17939 ( .A(n16082), .ZN(n14723) );
  AOI21_X1 U17940 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(n16183) );
  AOI22_X1 U17941 ( .A1(n16183), .A2(n20199), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14615), .ZN(n14614) );
  OAI21_X1 U17942 ( .B1(n14723), .B2(n14624), .A(n14614), .ZN(P1_U2857) );
  AOI22_X1 U17943 ( .A1(n16191), .A2(n20199), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14615), .ZN(n14616) );
  OAI21_X1 U17944 ( .B1(n14831), .B2(n14624), .A(n14616), .ZN(P1_U2859) );
  AOI21_X1 U17945 ( .B1(n14619), .B2(n14618), .A(n14617), .ZN(n16085) );
  INV_X1 U17946 ( .A(n16085), .ZN(n14625) );
  INV_X1 U17947 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14623) );
  NOR2_X1 U17948 ( .A1(n14621), .A2(n14620), .ZN(n14622) );
  OR2_X1 U17949 ( .A1(n14538), .A2(n14622), .ZN(n16029) );
  OAI222_X1 U17950 ( .A1(n14625), .A2(n14624), .B1(n14623), .B2(n20204), .C1(
        n16029), .C2(n20194), .ZN(P1_U2860) );
  INV_X1 U17951 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U17952 ( .A1(n14713), .A2(DATAI_30_), .ZN(n14627) );
  AOI22_X1 U17953 ( .A1(n13075), .A2(n20243), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n14724), .ZN(n14626) );
  OAI211_X1 U17954 ( .C1(n14717), .C2(n14628), .A(n14627), .B(n14626), .ZN(
        n14629) );
  INV_X1 U17955 ( .A(n14629), .ZN(n14630) );
  OAI21_X1 U17956 ( .B1(n14631), .B2(n9731), .A(n14630), .ZN(P1_U2874) );
  INV_X1 U17957 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14636) );
  NAND2_X1 U17958 ( .A1(n14713), .A2(DATAI_29_), .ZN(n14635) );
  INV_X1 U17959 ( .A(DATAI_13_), .ZN(n14633) );
  NAND2_X1 U17960 ( .A1(n14642), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14632) );
  OAI21_X1 U17961 ( .B1(n14642), .B2(n14633), .A(n14632), .ZN(n20241) );
  AOI22_X1 U17962 ( .A1(n13075), .A2(n20241), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n14724), .ZN(n14634) );
  OAI211_X1 U17963 ( .C1(n14717), .C2(n14636), .A(n14635), .B(n14634), .ZN(
        n14637) );
  INV_X1 U17964 ( .A(n14637), .ZN(n14638) );
  OAI21_X1 U17965 ( .B1(n14639), .B2(n9731), .A(n14638), .ZN(P1_U2875) );
  NAND2_X1 U17966 ( .A1(n14713), .A2(DATAI_28_), .ZN(n14644) );
  INV_X1 U17967 ( .A(DATAI_12_), .ZN(n14641) );
  NAND2_X1 U17968 ( .A1(n14642), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14640) );
  OAI21_X1 U17969 ( .B1(n14642), .B2(n14641), .A(n14640), .ZN(n20239) );
  AOI22_X1 U17970 ( .A1(n13075), .A2(n20239), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n14724), .ZN(n14643) );
  OAI211_X1 U17971 ( .C1(n14717), .C2(n16559), .A(n14644), .B(n14643), .ZN(
        n14645) );
  INV_X1 U17972 ( .A(n14645), .ZN(n14646) );
  OAI21_X1 U17973 ( .B1(n14647), .B2(n9731), .A(n14646), .ZN(P1_U2876) );
  INV_X1 U17974 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14650) );
  NAND2_X1 U17975 ( .A1(n14713), .A2(DATAI_27_), .ZN(n14649) );
  AOI22_X1 U17976 ( .A1(n13075), .A2(n20237), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14724), .ZN(n14648) );
  OAI211_X1 U17977 ( .C1(n14717), .C2(n14650), .A(n14649), .B(n14648), .ZN(
        n14651) );
  INV_X1 U17978 ( .A(n14651), .ZN(n14652) );
  OAI21_X1 U17979 ( .B1(n14653), .B2(n9731), .A(n14652), .ZN(P1_U2877) );
  INV_X1 U17980 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n14656) );
  NAND2_X1 U17981 ( .A1(n14713), .A2(DATAI_26_), .ZN(n14655) );
  AOI22_X1 U17982 ( .A1(n13075), .A2(n20235), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n14724), .ZN(n14654) );
  OAI211_X1 U17983 ( .C1(n14656), .C2(n14717), .A(n14655), .B(n14654), .ZN(
        n14657) );
  INV_X1 U17984 ( .A(n14657), .ZN(n14658) );
  OAI21_X1 U17985 ( .B1(n14659), .B2(n9731), .A(n14658), .ZN(P1_U2878) );
  NAND2_X1 U17986 ( .A1(n14713), .A2(DATAI_25_), .ZN(n14661) );
  AOI22_X1 U17987 ( .A1(n13075), .A2(n20233), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n14724), .ZN(n14660) );
  OAI211_X1 U17988 ( .C1(n16563), .C2(n14717), .A(n14661), .B(n14660), .ZN(
        n14662) );
  INV_X1 U17989 ( .A(n14662), .ZN(n14663) );
  OAI21_X1 U17990 ( .B1(n14664), .B2(n9731), .A(n14663), .ZN(P1_U2879) );
  NAND2_X1 U17991 ( .A1(n14713), .A2(DATAI_24_), .ZN(n14666) );
  AOI22_X1 U17992 ( .A1(n13075), .A2(n20231), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n14724), .ZN(n14665) );
  OAI211_X1 U17993 ( .C1(n16565), .C2(n14717), .A(n14666), .B(n14665), .ZN(
        n14667) );
  INV_X1 U17994 ( .A(n14667), .ZN(n14668) );
  OAI21_X1 U17995 ( .B1(n14669), .B2(n9731), .A(n14668), .ZN(P1_U2880) );
  INV_X1 U17996 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14673) );
  NAND2_X1 U17997 ( .A1(n14713), .A2(DATAI_23_), .ZN(n14672) );
  AOI22_X1 U17998 ( .A1(n13075), .A2(n14670), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14724), .ZN(n14671) );
  OAI211_X1 U17999 ( .C1(n14673), .C2(n14717), .A(n14672), .B(n14671), .ZN(
        n14674) );
  INV_X1 U18000 ( .A(n14674), .ZN(n14675) );
  OAI21_X1 U18001 ( .B1(n14791), .B2(n9731), .A(n14675), .ZN(P1_U2881) );
  NAND2_X1 U18002 ( .A1(n14713), .A2(DATAI_22_), .ZN(n14678) );
  AOI22_X1 U18003 ( .A1(n13075), .A2(n14676), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n14724), .ZN(n14677) );
  OAI211_X1 U18004 ( .C1(n16568), .C2(n14717), .A(n14678), .B(n14677), .ZN(
        n14679) );
  INV_X1 U18005 ( .A(n14679), .ZN(n14680) );
  OAI21_X1 U18006 ( .B1(n14805), .B2(n9731), .A(n14680), .ZN(P1_U2882) );
  INV_X1 U18007 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15253) );
  NAND2_X1 U18008 ( .A1(n14713), .A2(DATAI_21_), .ZN(n14683) );
  AOI22_X1 U18009 ( .A1(n13075), .A2(n14681), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n14724), .ZN(n14682) );
  OAI211_X1 U18010 ( .C1(n15253), .C2(n14717), .A(n14683), .B(n14682), .ZN(
        n14684) );
  INV_X1 U18011 ( .A(n14684), .ZN(n14685) );
  OAI21_X1 U18012 ( .B1(n14686), .B2(n9731), .A(n14685), .ZN(P1_U2883) );
  NAND2_X1 U18013 ( .A1(n14713), .A2(DATAI_20_), .ZN(n14689) );
  AOI22_X1 U18014 ( .A1(n13075), .A2(n14687), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14724), .ZN(n14688) );
  OAI211_X1 U18015 ( .C1(n16571), .C2(n14717), .A(n14689), .B(n14688), .ZN(
        n14690) );
  INV_X1 U18016 ( .A(n14690), .ZN(n14691) );
  OAI21_X1 U18017 ( .B1(n14692), .B2(n9731), .A(n14691), .ZN(P1_U2884) );
  NAND2_X1 U18018 ( .A1(n14713), .A2(DATAI_19_), .ZN(n14695) );
  AOI22_X1 U18019 ( .A1(n13075), .A2(n14693), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n14724), .ZN(n14694) );
  OAI211_X1 U18020 ( .C1(n14696), .C2(n14717), .A(n14695), .B(n14694), .ZN(
        n14697) );
  INV_X1 U18021 ( .A(n14697), .ZN(n14698) );
  OAI21_X1 U18022 ( .B1(n14699), .B2(n9731), .A(n14698), .ZN(P1_U2885) );
  INV_X1 U18023 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14703) );
  NAND2_X1 U18024 ( .A1(n14713), .A2(DATAI_18_), .ZN(n14702) );
  AOI22_X1 U18025 ( .A1(n13075), .A2(n14700), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n14724), .ZN(n14701) );
  OAI211_X1 U18026 ( .C1(n14703), .C2(n14717), .A(n14702), .B(n14701), .ZN(
        n14704) );
  AOI21_X1 U18027 ( .B1(n15989), .B2(n16044), .A(n14704), .ZN(n14705) );
  INV_X1 U18028 ( .A(n14705), .ZN(P1_U2886) );
  INV_X1 U18029 ( .A(n14706), .ZN(n16070) );
  NAND2_X1 U18030 ( .A1(n14713), .A2(DATAI_17_), .ZN(n14709) );
  AOI22_X1 U18031 ( .A1(n13075), .A2(n14707), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n14724), .ZN(n14708) );
  OAI211_X1 U18032 ( .C1(n14710), .C2(n14717), .A(n14709), .B(n14708), .ZN(
        n14711) );
  AOI21_X1 U18033 ( .B1(n16070), .B2(n16044), .A(n14711), .ZN(n14712) );
  INV_X1 U18034 ( .A(n14712), .ZN(P1_U2887) );
  INV_X1 U18035 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14718) );
  NAND2_X1 U18036 ( .A1(n14713), .A2(DATAI_16_), .ZN(n14716) );
  AOI22_X1 U18037 ( .A1(n13075), .A2(n14714), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n14724), .ZN(n14715) );
  OAI211_X1 U18038 ( .C1(n14718), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        n14719) );
  AOI21_X1 U18039 ( .B1(n16000), .B2(n16044), .A(n14719), .ZN(n14720) );
  INV_X1 U18040 ( .A(n14720), .ZN(P1_U2888) );
  OAI222_X1 U18041 ( .A1(n9731), .A2(n14723), .B1(n14722), .B2(n14721), .C1(
        n16046), .C2(n12978), .ZN(P1_U2889) );
  AOI22_X1 U18042 ( .A1(n16043), .A2(n20241), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14724), .ZN(n14725) );
  OAI21_X1 U18043 ( .B1(n14831), .B2(n9731), .A(n14725), .ZN(P1_U2891) );
  AOI21_X1 U18044 ( .B1(n14726), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9834), .ZN(n14853) );
  NAND2_X1 U18045 ( .A1(n16114), .A2(n14727), .ZN(n14728) );
  NAND2_X1 U18046 ( .A1(n20177), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14846) );
  OAI211_X1 U18047 ( .C1(n16120), .C2(n20999), .A(n14728), .B(n14846), .ZN(
        n14729) );
  AOI21_X1 U18048 ( .B1(n14730), .B2(n16069), .A(n14729), .ZN(n14731) );
  OAI21_X1 U18049 ( .B1(n14853), .B2(n20100), .A(n14731), .ZN(P1_U2969) );
  MUX2_X1 U18050 ( .A(n14733), .B(n14732), .S(n16090), .Z(n14734) );
  XNOR2_X1 U18051 ( .A(n14734), .B(n14856), .ZN(n14862) );
  NAND2_X1 U18052 ( .A1(n20177), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14854) );
  NAND2_X1 U18053 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14735) );
  OAI211_X1 U18054 ( .C1(n16111), .C2(n14736), .A(n14854), .B(n14735), .ZN(
        n14737) );
  AOI21_X1 U18055 ( .B1(n14738), .B2(n16069), .A(n14737), .ZN(n14739) );
  OAI21_X1 U18056 ( .B1(n20100), .B2(n14862), .A(n14739), .ZN(P1_U2970) );
  NAND2_X1 U18057 ( .A1(n14741), .A2(n14894), .ZN(n14773) );
  NAND2_X1 U18058 ( .A1(n14741), .A2(n14740), .ZN(n14756) );
  AND2_X1 U18059 ( .A1(n14753), .A2(n14765), .ZN(n14742) );
  NAND2_X1 U18060 ( .A1(n16090), .A2(n14765), .ZN(n14743) );
  NOR2_X1 U18061 ( .A1(n14744), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14745) );
  AOI211_X1 U18062 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14894), .A(
        n14758), .B(n14745), .ZN(n14746) );
  XNOR2_X1 U18063 ( .A(n14746), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14873) );
  INV_X1 U18064 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14749) );
  NAND2_X1 U18065 ( .A1(n16114), .A2(n14747), .ZN(n14748) );
  NAND2_X1 U18066 ( .A1(n20177), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14868) );
  OAI211_X1 U18067 ( .C1(n16120), .C2(n14749), .A(n14748), .B(n14868), .ZN(
        n14750) );
  AOI21_X1 U18068 ( .B1(n14751), .B2(n16069), .A(n14750), .ZN(n14752) );
  OAI21_X1 U18069 ( .B1(n20100), .B2(n14873), .A(n14752), .ZN(P1_U2971) );
  INV_X1 U18070 ( .A(n14753), .ZN(n14754) );
  OR2_X1 U18071 ( .A1(n16090), .A2(n14754), .ZN(n14755) );
  NAND2_X1 U18072 ( .A1(n14756), .A2(n14755), .ZN(n14757) );
  OR2_X1 U18073 ( .A1(n14758), .A2(n14766), .ZN(n14759) );
  INV_X1 U18074 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14874) );
  XNOR2_X1 U18075 ( .A(n14759), .B(n14874), .ZN(n14882) );
  NAND2_X1 U18076 ( .A1(n20177), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14877) );
  NAND2_X1 U18077 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14760) );
  OAI211_X1 U18078 ( .C1(n16111), .C2(n14761), .A(n14877), .B(n14760), .ZN(
        n14762) );
  AOI21_X1 U18079 ( .B1(n14763), .B2(n16069), .A(n14762), .ZN(n14764) );
  OAI21_X1 U18080 ( .B1(n20100), .B2(n14882), .A(n14764), .ZN(P1_U2972) );
  AOI22_X1 U18081 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20177), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n14767) );
  OAI21_X1 U18082 ( .B1(n16111), .B2(n14768), .A(n14767), .ZN(n14769) );
  AOI21_X1 U18083 ( .B1(n14770), .B2(n16069), .A(n14769), .ZN(n14771) );
  OAI21_X1 U18084 ( .B1(n20100), .B2(n16122), .A(n14771), .ZN(P1_U2973) );
  INV_X1 U18085 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16148) );
  AND2_X1 U18086 ( .A1(n14772), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14782) );
  MUX2_X1 U18087 ( .A(n14894), .B(n14782), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n14774) );
  OAI211_X1 U18088 ( .C1(n16148), .C2(n16090), .A(n14774), .B(n14773), .ZN(
        n14775) );
  XNOR2_X1 U18089 ( .A(n14775), .B(n16136), .ZN(n16130) );
  AOI22_X1 U18090 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20177), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n14776) );
  OAI21_X1 U18091 ( .B1(n16111), .B2(n14777), .A(n14776), .ZN(n14778) );
  AOI21_X1 U18092 ( .B1(n14779), .B2(n16069), .A(n14778), .ZN(n14780) );
  OAI21_X1 U18093 ( .B1(n20100), .B2(n16130), .A(n14780), .ZN(P1_U2974) );
  NOR2_X1 U18094 ( .A1(n14782), .A2(n14741), .ZN(n14781) );
  MUX2_X1 U18095 ( .A(n14782), .B(n14781), .S(n14894), .Z(n14783) );
  XNOR2_X1 U18096 ( .A(n14783), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14892) );
  INV_X1 U18097 ( .A(n14784), .ZN(n14786) );
  AOI22_X1 U18098 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20177), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n14785) );
  OAI21_X1 U18099 ( .B1(n16111), .B2(n14786), .A(n14785), .ZN(n14787) );
  AOI21_X1 U18100 ( .B1(n14788), .B2(n16069), .A(n14787), .ZN(n14789) );
  OAI21_X1 U18101 ( .B1(n20100), .B2(n14892), .A(n14789), .ZN(P1_U2975) );
  XNOR2_X1 U18102 ( .A(n16090), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14790) );
  XNOR2_X1 U18103 ( .A(n14741), .B(n14790), .ZN(n16141) );
  INV_X1 U18104 ( .A(n14791), .ZN(n14796) );
  INV_X1 U18105 ( .A(n14792), .ZN(n14794) );
  AOI22_X1 U18106 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20177), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14793) );
  OAI21_X1 U18107 ( .B1(n16111), .B2(n14794), .A(n14793), .ZN(n14795) );
  AOI21_X1 U18108 ( .B1(n14796), .B2(n16069), .A(n14795), .ZN(n14797) );
  OAI21_X1 U18109 ( .B1(n16141), .B2(n20100), .A(n14797), .ZN(P1_U2976) );
  INV_X1 U18110 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14798) );
  OAI22_X1 U18111 ( .A1(n16120), .A2(n20900), .B1(n9736), .B2(n14798), .ZN(
        n14799) );
  AOI21_X1 U18112 ( .B1(n15944), .B2(n16114), .A(n14799), .ZN(n14804) );
  NAND2_X1 U18113 ( .A1(n14801), .A2(n14800), .ZN(n14802) );
  XOR2_X1 U18114 ( .A(n12249), .B(n14802), .Z(n16152) );
  NAND2_X1 U18115 ( .A1(n16152), .A2(n16116), .ZN(n14803) );
  OAI211_X1 U18116 ( .C1(n14805), .C2(n14832), .A(n14804), .B(n14803), .ZN(
        P1_U2977) );
  OAI21_X1 U18117 ( .B1(n14806), .B2(n14808), .A(n14807), .ZN(n16169) );
  AOI22_X1 U18118 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20177), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14809) );
  OAI21_X1 U18119 ( .B1(n15987), .B2(n16111), .A(n14809), .ZN(n14810) );
  AOI21_X1 U18120 ( .B1(n15989), .B2(n16069), .A(n14810), .ZN(n14811) );
  OAI21_X1 U18121 ( .B1(n20100), .B2(n16169), .A(n14811), .ZN(P1_U2981) );
  OR2_X1 U18122 ( .A1(n14834), .A2(n14812), .ZN(n16078) );
  AOI21_X1 U18123 ( .B1(n16078), .B2(n16063), .A(n16073), .ZN(n14813) );
  XOR2_X1 U18124 ( .A(n14814), .B(n14813), .Z(n14917) );
  NAND2_X1 U18125 ( .A1(n16000), .A2(n16069), .ZN(n14819) );
  INV_X1 U18126 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14815) );
  OAI22_X1 U18127 ( .A1(n16120), .A2(n14816), .B1(n9736), .B2(n14815), .ZN(
        n14817) );
  AOI21_X1 U18128 ( .B1(n16114), .B2(n16005), .A(n14817), .ZN(n14818) );
  OAI211_X1 U18129 ( .C1(n14917), .C2(n20100), .A(n14819), .B(n14818), .ZN(
        P1_U2983) );
  INV_X1 U18130 ( .A(n14820), .ZN(n14821) );
  AOI22_X1 U18131 ( .A1(n12073), .A2(n14822), .B1(n14894), .B2(n14821), .ZN(
        n14930) );
  INV_X1 U18132 ( .A(n14824), .ZN(n14823) );
  AOI21_X1 U18133 ( .B1(n14894), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14823), .ZN(n14929) );
  NAND2_X1 U18134 ( .A1(n14930), .A2(n14929), .ZN(n14928) );
  NAND2_X1 U18135 ( .A1(n14928), .A2(n14824), .ZN(n14825) );
  XOR2_X1 U18136 ( .A(n14826), .B(n14825), .Z(n16192) );
  NAND2_X1 U18137 ( .A1(n16192), .A2(n16116), .ZN(n14830) );
  OAI22_X1 U18138 ( .A1(n16120), .A2(n14548), .B1(n9736), .B2(n20697), .ZN(
        n14827) );
  AOI21_X1 U18139 ( .B1(n16114), .B2(n14828), .A(n14827), .ZN(n14829) );
  OAI211_X1 U18140 ( .C1(n14832), .C2(n14831), .A(n14830), .B(n14829), .ZN(
        P1_U2986) );
  NAND2_X1 U18141 ( .A1(n14833), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14836) );
  XNOR2_X1 U18142 ( .A(n14834), .B(n14837), .ZN(n14835) );
  MUX2_X1 U18143 ( .A(n14836), .B(n14835), .S(n16090), .Z(n14839) );
  INV_X1 U18144 ( .A(n14833), .ZN(n14838) );
  NAND3_X1 U18145 ( .A1(n14838), .A2(n14894), .A3(n14837), .ZN(n16091) );
  NAND2_X1 U18146 ( .A1(n14839), .A2(n16091), .ZN(n16211) );
  INV_X1 U18147 ( .A(n16211), .ZN(n14845) );
  AOI22_X1 U18148 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20177), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14840) );
  OAI21_X1 U18149 ( .B1(n16111), .B2(n14841), .A(n14840), .ZN(n14842) );
  AOI21_X1 U18150 ( .B1(n14843), .B2(n16069), .A(n14842), .ZN(n14844) );
  OAI21_X1 U18151 ( .B1(n14845), .B2(n20100), .A(n14844), .ZN(P1_U2989) );
  INV_X1 U18152 ( .A(n14846), .ZN(n14847) );
  AOI21_X1 U18153 ( .B1(n14848), .B2(n16256), .A(n14847), .ZN(n14852) );
  OAI21_X1 U18154 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14850), .A(
        n14849), .ZN(n14851) );
  OAI211_X1 U18155 ( .C1(n14853), .C2(n16259), .A(n14852), .B(n14851), .ZN(
        P1_U3001) );
  INV_X1 U18156 ( .A(n14866), .ZN(n14875) );
  NOR2_X1 U18157 ( .A1(n14863), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14860) );
  OAI21_X1 U18158 ( .B1(n14855), .B2(n16220), .A(n14854), .ZN(n14859) );
  NOR2_X1 U18159 ( .A1(n14857), .A2(n14856), .ZN(n14858) );
  AOI211_X1 U18160 ( .C1(n14875), .C2(n14860), .A(n14859), .B(n14858), .ZN(
        n14861) );
  OAI21_X1 U18161 ( .B1(n14862), .B2(n16259), .A(n14861), .ZN(P1_U3002) );
  INV_X1 U18162 ( .A(n14863), .ZN(n14865) );
  NOR3_X1 U18163 ( .A1(n14866), .A2(n14865), .A3(n14864), .ZN(n14871) );
  INV_X1 U18164 ( .A(n14867), .ZN(n14869) );
  OAI21_X1 U18165 ( .B1(n14869), .B2(n16220), .A(n14868), .ZN(n14870) );
  AOI211_X1 U18166 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n14880), .A(
        n14871), .B(n14870), .ZN(n14872) );
  OAI21_X1 U18167 ( .B1(n14873), .B2(n16259), .A(n14872), .ZN(P1_U3003) );
  NAND2_X1 U18168 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  OAI211_X1 U18169 ( .C1(n14878), .C2(n16220), .A(n14877), .B(n14876), .ZN(
        n14879) );
  AOI21_X1 U18170 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14880), .A(
        n14879), .ZN(n14881) );
  OAI21_X1 U18171 ( .B1(n14882), .B2(n16259), .A(n14881), .ZN(P1_U3004) );
  OAI22_X1 U18172 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14883), .B1(
        n14493), .B2(n9736), .ZN(n14889) );
  OAI21_X1 U18173 ( .B1(n14885), .B2(n14884), .A(n16148), .ZN(n14887) );
  AOI21_X1 U18174 ( .B1(n14887), .B2(n16147), .A(n14886), .ZN(n14888) );
  AOI211_X1 U18175 ( .C1(n14890), .C2(n16256), .A(n14889), .B(n14888), .ZN(
        n14891) );
  OAI21_X1 U18176 ( .B1(n14892), .B2(n16259), .A(n14891), .ZN(P1_U3007) );
  NAND2_X1 U18177 ( .A1(n16090), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14893) );
  NOR2_X1 U18178 ( .A1(n14807), .A2(n14893), .ZN(n15914) );
  INV_X1 U18179 ( .A(n15914), .ZN(n14896) );
  NAND2_X1 U18180 ( .A1(n14895), .A2(n14894), .ZN(n15916) );
  NAND2_X1 U18181 ( .A1(n14896), .A2(n15916), .ZN(n14897) );
  XNOR2_X1 U18182 ( .A(n14897), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16056) );
  AOI221_X1 U18183 ( .B1(n14900), .B2(n16160), .C1(n14899), .C2(n16160), .A(
        n9883), .ZN(n14901) );
  OAI22_X1 U18184 ( .A1(n16056), .A2(n16259), .B1(n14902), .B2(n14901), .ZN(
        n14906) );
  NOR4_X1 U18185 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16189), .A3(
        n16160), .A4(n16159), .ZN(n14905) );
  INV_X1 U18186 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14903) );
  OAI22_X1 U18187 ( .A1(n15965), .A2(n16220), .B1(n9736), .B2(n14903), .ZN(
        n14904) );
  OR3_X1 U18188 ( .A1(n14906), .A2(n14905), .A3(n14904), .ZN(P1_U3011) );
  NAND2_X1 U18189 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16140), .ZN(
        n16174) );
  NOR2_X1 U18190 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16174), .ZN(
        n16184) );
  AOI21_X1 U18191 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14907), .A(
        n14920), .ZN(n14909) );
  AOI211_X1 U18192 ( .C1(n12227), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        n16165) );
  INV_X1 U18193 ( .A(n16165), .ZN(n16185) );
  OAI21_X1 U18194 ( .B1(n16184), .B2(n16185), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14911) );
  INV_X1 U18195 ( .A(n14911), .ZN(n14915) );
  NOR3_X1 U18196 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14912), .A3(
        n16174), .ZN(n14914) );
  OAI22_X1 U18197 ( .A1(n16001), .A2(n16220), .B1(n14815), .B2(n9736), .ZN(
        n14913) );
  NOR3_X1 U18198 ( .A1(n14915), .A2(n14914), .A3(n14913), .ZN(n14916) );
  OAI21_X1 U18199 ( .B1(n14917), .B2(n16259), .A(n14916), .ZN(P1_U3015) );
  NOR3_X1 U18200 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14918), .A3(
        n14924), .ZN(n16198) );
  INV_X1 U18201 ( .A(n16198), .ZN(n14925) );
  OAI221_X1 U18202 ( .B1(n14920), .B2(n16204), .C1(n14920), .C2(n14927), .A(
        n14919), .ZN(n14921) );
  AOI221_X1 U18203 ( .B1(n14924), .B2(n14923), .C1(n14922), .C2(n14923), .A(
        n14921), .ZN(n16203) );
  OAI21_X1 U18204 ( .B1(n14926), .B2(n14925), .A(n16203), .ZN(n14934) );
  NAND3_X1 U18205 ( .A1(n14927), .A2(n16239), .A3(n16250), .ZN(n14932) );
  OAI21_X1 U18206 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(n14931) );
  INV_X1 U18207 ( .A(n14931), .ZN(n16089) );
  OAI22_X1 U18208 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14932), .B1(
        n16089), .B2(n16259), .ZN(n14933) );
  AOI21_X1 U18209 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14934), .A(
        n14933), .ZN(n14936) );
  NAND2_X1 U18210 ( .A1(n16241), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14935) );
  OAI211_X1 U18211 ( .C1(n16220), .C2(n16029), .A(n14936), .B(n14935), .ZN(
        P1_U3019) );
  OAI21_X1 U18212 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13130), .A(n20519), 
        .ZN(n14937) );
  OAI21_X1 U18213 ( .B1(n14942), .B2(n20551), .A(n14937), .ZN(n14938) );
  MUX2_X1 U18214 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14938), .S(
        n20262), .Z(P1_U3477) );
  AND2_X1 U18215 ( .A1(n20548), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14939) );
  NAND2_X1 U18216 ( .A1(n13130), .A2(n14939), .ZN(n20605) );
  MUX2_X1 U18217 ( .A(n20605), .B(n14940), .S(n9769), .Z(n14941) );
  OAI21_X1 U18218 ( .B1(n14942), .B2(n13125), .A(n14941), .ZN(n14943) );
  MUX2_X1 U18219 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14943), .S(
        n20262), .Z(P1_U3476) );
  NOR3_X1 U18220 ( .A1(n14944), .A2(n13229), .A3(n13206), .ZN(n14947) );
  NOR2_X1 U18221 ( .A1(n20551), .A2(n14945), .ZN(n14946) );
  AOI211_X1 U18222 ( .C1(n14948), .C2(n11892), .A(n14947), .B(n14946), .ZN(
        n15882) );
  INV_X1 U18223 ( .A(n14949), .ZN(n14964) );
  OAI22_X1 U18224 ( .A1(n12087), .A2(n12996), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14954) );
  NOR2_X1 U18225 ( .A1(n20661), .A2(n20984), .ZN(n14956) );
  NOR3_X1 U18226 ( .A1(n13229), .A2(n13206), .A3(n14962), .ZN(n14950) );
  AOI21_X1 U18227 ( .B1(n14954), .B2(n14956), .A(n14950), .ZN(n14951) );
  OAI21_X1 U18228 ( .B1(n15882), .B2(n14964), .A(n14951), .ZN(n14952) );
  MUX2_X1 U18229 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14952), .S(
        n14966), .Z(P1_U3473) );
  INV_X1 U18230 ( .A(n14953), .ZN(n14958) );
  INV_X1 U18231 ( .A(n14954), .ZN(n14955) );
  AOI22_X1 U18232 ( .A1(n14958), .A2(n14957), .B1(n14956), .B2(n14955), .ZN(
        n14959) );
  OAI21_X1 U18233 ( .B1(n14960), .B2(n14964), .A(n14959), .ZN(n14961) );
  MUX2_X1 U18234 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14961), .S(
        n14966), .Z(P1_U3472) );
  OAI22_X1 U18235 ( .A1(n14965), .A2(n14964), .B1(n14963), .B2(n14962), .ZN(
        n14967) );
  MUX2_X1 U18236 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14967), .S(
        n14966), .Z(P1_U3469) );
  OR2_X1 U18237 ( .A1(n14969), .A2(n14968), .ZN(n14971) );
  NAND2_X1 U18238 ( .A1(n14975), .A2(n16306), .ZN(n14972) );
  AND2_X1 U18239 ( .A1(n14973), .A2(n14972), .ZN(n15280) );
  INV_X1 U18240 ( .A(n15280), .ZN(n16315) );
  OR2_X1 U18241 ( .A1(n9864), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14974) );
  NAND2_X1 U18242 ( .A1(n14975), .A2(n14974), .ZN(n15291) );
  AND2_X1 U18243 ( .A1(n14977), .A2(n15029), .ZN(n14976) );
  OR2_X1 U18244 ( .A1(n14976), .A2(n9864), .ZN(n15300) );
  OAI21_X1 U18245 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n14978), .A(
        n14977), .ZN(n16327) );
  AOI21_X1 U18246 ( .B1(n16362), .B2(n14979), .A(n14978), .ZN(n16354) );
  INV_X1 U18247 ( .A(n16354), .ZN(n16337) );
  OAI21_X1 U18248 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14980), .A(
        n14979), .ZN(n15869) );
  NAND2_X1 U18249 ( .A1(n15337), .A2(n14991), .ZN(n14982) );
  INV_X1 U18250 ( .A(n14980), .ZN(n14981) );
  AND2_X1 U18251 ( .A1(n14982), .A2(n14981), .ZN(n15339) );
  AOI21_X1 U18252 ( .B1(n14989), .B2(n15358), .A(n9863), .ZN(n19035) );
  AOI21_X1 U18253 ( .B1(n15369), .B2(n14987), .A(n14990), .ZN(n15368) );
  AOI21_X1 U18254 ( .B1(n19090), .B2(n14985), .A(n14988), .ZN(n19084) );
  AOI21_X1 U18255 ( .B1(n19102), .B2(n14983), .A(n14986), .ZN(n19108) );
  NAND2_X1 U18256 ( .A1(n14984), .A2(n16400), .ZN(n19106) );
  NOR2_X1 U18257 ( .A1(n19108), .A2(n19106), .ZN(n19091) );
  OAI21_X1 U18258 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14986), .A(
        n14985), .ZN(n19092) );
  NAND2_X1 U18259 ( .A1(n19091), .A2(n19092), .ZN(n19082) );
  NOR2_X1 U18260 ( .A1(n19084), .A2(n19082), .ZN(n19069) );
  OAI21_X1 U18261 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14988), .A(
        n14987), .ZN(n19070) );
  NAND2_X1 U18262 ( .A1(n19069), .A2(n19070), .ZN(n19057) );
  NOR2_X1 U18263 ( .A1(n15368), .A2(n19057), .ZN(n19044) );
  OAI21_X1 U18264 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14990), .A(
        n14989), .ZN(n19045) );
  NAND2_X1 U18265 ( .A1(n19044), .A2(n19045), .ZN(n19033) );
  NOR2_X1 U18266 ( .A1(n19035), .A2(n19033), .ZN(n19028) );
  OAI21_X1 U18267 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9863), .A(
        n14991), .ZN(n19027) );
  NAND2_X1 U18268 ( .A1(n19028), .A2(n19027), .ZN(n15037) );
  OAI21_X1 U18269 ( .B1(n15339), .B2(n15037), .A(n19190), .ZN(n15868) );
  NAND2_X1 U18270 ( .A1(n15869), .A2(n15868), .ZN(n15867) );
  NAND2_X1 U18271 ( .A1(n19190), .A2(n15867), .ZN(n16336) );
  NAND2_X1 U18272 ( .A1(n16337), .A2(n16336), .ZN(n16335) );
  NAND2_X1 U18273 ( .A1(n19190), .A2(n16335), .ZN(n16326) );
  NAND2_X1 U18274 ( .A1(n16327), .A2(n16326), .ZN(n16325) );
  NAND2_X1 U18275 ( .A1(n19190), .A2(n16325), .ZN(n15025) );
  NAND2_X1 U18276 ( .A1(n15300), .A2(n15025), .ZN(n15024) );
  NAND2_X1 U18277 ( .A1(n19190), .A2(n15024), .ZN(n15014) );
  NAND2_X1 U18278 ( .A1(n15291), .A2(n15014), .ZN(n15013) );
  NAND2_X1 U18279 ( .A1(n19190), .A2(n15013), .ZN(n16314) );
  NAND2_X1 U18280 ( .A1(n16315), .A2(n16314), .ZN(n16313) );
  NAND2_X1 U18281 ( .A1(n19190), .A2(n16313), .ZN(n16300) );
  NAND2_X1 U18282 ( .A1(n16301), .A2(n16300), .ZN(n16299) );
  NAND2_X1 U18283 ( .A1(n19190), .A2(n16299), .ZN(n14994) );
  NOR2_X1 U18284 ( .A1(n14992), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14993) );
  OR2_X1 U18285 ( .A1(n15259), .A2(n14993), .ZN(n15273) );
  NAND2_X1 U18286 ( .A1(n15273), .A2(n14994), .ZN(n16273) );
  OAI211_X1 U18287 ( .C1(n14994), .C2(n15273), .A(n19185), .B(n16273), .ZN(
        n15003) );
  OAI21_X1 U18288 ( .B1(n15203), .B2(n14996), .A(n14995), .ZN(n15414) );
  INV_X1 U18289 ( .A(n15414), .ZN(n15197) );
  INV_X1 U18290 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14998) );
  AOI22_X1 U18291 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19223), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19222), .ZN(n14997) );
  OAI21_X1 U18292 ( .B1(n14998), .B2(n19174), .A(n14997), .ZN(n15001) );
  NOR2_X1 U18293 ( .A1(n14999), .A2(n19228), .ZN(n15000) );
  AOI211_X1 U18294 ( .C1(n15197), .C2(n19224), .A(n15001), .B(n15000), .ZN(
        n15002) );
  OAI211_X1 U18295 ( .C1(n15090), .C2(n19200), .A(n15003), .B(n15002), .ZN(
        P2_U2826) );
  INV_X1 U18296 ( .A(n15100), .ZN(n15004) );
  AOI21_X1 U18297 ( .B1(n15005), .B2(n15023), .A(n15004), .ZN(n15447) );
  NAND2_X1 U18298 ( .A1(n15007), .A2(n15006), .ZN(n15008) );
  AND2_X1 U18299 ( .A1(n15210), .A2(n15008), .ZN(n15449) );
  INV_X1 U18300 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20937) );
  OAI22_X1 U18301 ( .A1(n20937), .A2(n19178), .B1(n15009), .B2(n19197), .ZN(
        n15010) );
  INV_X1 U18302 ( .A(n15010), .ZN(n15011) );
  OAI21_X1 U18303 ( .B1(n19174), .B2(n10094), .A(n15011), .ZN(n15012) );
  AOI21_X1 U18304 ( .B1(n15449), .B2(n19224), .A(n15012), .ZN(n15016) );
  OAI211_X1 U18305 ( .C1(n15291), .C2(n15014), .A(n19185), .B(n15013), .ZN(
        n15015) );
  OAI211_X1 U18306 ( .C1(n15017), .C2(n19228), .A(n15016), .B(n15015), .ZN(
        n15018) );
  AOI21_X1 U18307 ( .B1(n15447), .B2(n16282), .A(n15018), .ZN(n15019) );
  INV_X1 U18308 ( .A(n15019), .ZN(P2_U2829) );
  OR2_X1 U18309 ( .A1(n15020), .A2(n15021), .ZN(n15022) );
  AND2_X1 U18310 ( .A1(n15023), .A2(n15022), .ZN(n15468) );
  INV_X1 U18311 ( .A(n15468), .ZN(n15033) );
  OAI211_X1 U18312 ( .C1(n15025), .C2(n15300), .A(n19185), .B(n15024), .ZN(
        n15032) );
  XOR2_X1 U18313 ( .A(n15026), .B(n15230), .Z(n15460) );
  NAND2_X1 U18314 ( .A1(n15460), .A2(n19224), .ZN(n15028) );
  AOI22_X1 U18315 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19223), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19222), .ZN(n15027) );
  OAI211_X1 U18316 ( .C1(n19174), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        n15030) );
  AOI21_X1 U18317 ( .B1(n9819), .B2(n19194), .A(n15030), .ZN(n15031) );
  OAI211_X1 U18318 ( .C1(n19200), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        P2_U2830) );
  OAI21_X1 U18319 ( .B1(n15034), .B2(n15036), .A(n15035), .ZN(n15517) );
  AND2_X1 U18320 ( .A1(n19190), .A2(n15037), .ZN(n19026) );
  OAI21_X1 U18321 ( .B1(n15339), .B2(n19026), .A(n19185), .ZN(n15038) );
  AOI21_X1 U18322 ( .B1(n19026), .B2(n15339), .A(n15038), .ZN(n15047) );
  OR2_X1 U18323 ( .A1(n15152), .A2(n15040), .ZN(n15041) );
  NAND2_X1 U18324 ( .A1(n15039), .A2(n15041), .ZN(n15509) );
  INV_X1 U18325 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15144) );
  OAI22_X1 U18326 ( .A1(n21000), .A2(n19178), .B1(n15144), .B2(n19197), .ZN(
        n15042) );
  AOI21_X1 U18327 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19236), .A(
        n15042), .ZN(n15045) );
  NAND2_X1 U18328 ( .A1(n15043), .A2(n19194), .ZN(n15044) );
  OAI211_X1 U18329 ( .C1(n15509), .C2(n19200), .A(n15045), .B(n15044), .ZN(
        n15046) );
  NOR2_X1 U18330 ( .A1(n15047), .A2(n15046), .ZN(n15048) );
  OAI21_X1 U18331 ( .B1(n15517), .B2(n19213), .A(n15048), .ZN(P2_U2834) );
  NAND2_X1 U18332 ( .A1(n19190), .A2(n15049), .ZN(n15050) );
  XNOR2_X1 U18333 ( .A(n16433), .B(n15050), .ZN(n15051) );
  NAND2_X1 U18334 ( .A1(n15051), .A2(n19185), .ZN(n15058) );
  NOR2_X1 U18335 ( .A1(n19178), .A2(n19975), .ZN(n15053) );
  OAI22_X1 U18336 ( .A1(n19213), .A2(n20038), .B1(n19174), .B2(n16446), .ZN(
        n15052) );
  AOI211_X1 U18337 ( .C1(n19222), .C2(P2_EBX_REG_3__SCAN_IN), .A(n15053), .B(
        n15052), .ZN(n15054) );
  OAI21_X1 U18338 ( .B1(n15055), .B2(n19228), .A(n15054), .ZN(n15056) );
  AOI21_X1 U18339 ( .B1(n13580), .B2(n16282), .A(n15056), .ZN(n15057) );
  OAI211_X1 U18340 ( .C1(n19233), .C2(n19672), .A(n15058), .B(n15057), .ZN(
        P2_U2852) );
  INV_X1 U18341 ( .A(n15061), .ZN(n15062) );
  NOR2_X1 U18342 ( .A1(n19206), .A2(n15059), .ZN(n15071) );
  INV_X1 U18343 ( .A(n15071), .ZN(n15060) );
  AOI221_X1 U18344 ( .B1(n15062), .B2(n15071), .C1(n15061), .C2(n15060), .A(
        n19955), .ZN(n15063) );
  INV_X1 U18345 ( .A(n15063), .ZN(n15070) );
  AOI22_X1 U18346 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19223), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n19222), .ZN(n15065) );
  NAND2_X1 U18347 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19236), .ZN(
        n15064) );
  OAI211_X1 U18348 ( .C1(n19228), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15068) );
  NOR2_X1 U18349 ( .A1(n19399), .A2(n19213), .ZN(n15067) );
  OAI211_X1 U18350 ( .C1(n20043), .C2(n19233), .A(n15070), .B(n15069), .ZN(
        P2_U2853) );
  OAI21_X1 U18351 ( .B1(n19240), .B2(n15072), .A(n15071), .ZN(n15707) );
  INV_X1 U18352 ( .A(n19233), .ZN(n19218) );
  AOI22_X1 U18353 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19223), .B1(
        P2_EBX_REG_1__SCAN_IN), .B2(n19222), .ZN(n15075) );
  NOR2_X1 U18354 ( .A1(n19190), .A2(n19955), .ZN(n19235) );
  NAND2_X1 U18355 ( .A1(n19235), .A2(n15073), .ZN(n15074) );
  OAI211_X1 U18356 ( .C1(n15073), .C2(n19174), .A(n15075), .B(n15074), .ZN(
        n15076) );
  AOI21_X1 U18357 ( .B1(n19194), .B2(n15077), .A(n15076), .ZN(n15079) );
  NAND2_X1 U18358 ( .A1(n20055), .A2(n19224), .ZN(n15078) );
  OAI211_X1 U18359 ( .C1(n15080), .C2(n19200), .A(n15079), .B(n15078), .ZN(
        n15081) );
  AOI21_X1 U18360 ( .B1(n20053), .B2(n19218), .A(n15081), .ZN(n15082) );
  OAI21_X1 U18361 ( .B1(n15707), .B2(n19955), .A(n15082), .ZN(P2_U2854) );
  NAND2_X1 U18362 ( .A1(n16274), .A2(n15159), .ZN(n15083) );
  OAI21_X1 U18363 ( .B1(n15159), .B2(n15084), .A(n15083), .ZN(P2_U2856) );
  OR2_X1 U18364 ( .A1(n15086), .A2(n15085), .ZN(n15195) );
  NAND3_X1 U18365 ( .A1(n15195), .A2(n15087), .A3(n15149), .ZN(n15089) );
  NAND2_X1 U18366 ( .A1(n12766), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15088) );
  OAI211_X1 U18367 ( .C1(n15090), .C2(n12766), .A(n15089), .B(n15088), .ZN(
        P2_U2858) );
  NOR2_X1 U18368 ( .A1(n9745), .A2(n15091), .ZN(n15093) );
  XNOR2_X1 U18369 ( .A(n15093), .B(n15092), .ZN(n15208) );
  NOR2_X1 U18370 ( .A1(n16297), .A2(n12766), .ZN(n15094) );
  AOI21_X1 U18371 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n12766), .A(n15094), .ZN(
        n15095) );
  OAI21_X1 U18372 ( .B1(n15208), .B2(n15185), .A(n15095), .ZN(P2_U2859) );
  OAI21_X1 U18373 ( .B1(n15096), .B2(n15098), .A(n15097), .ZN(n15216) );
  NAND2_X1 U18374 ( .A1(n15100), .A2(n15099), .ZN(n15101) );
  NAND2_X1 U18375 ( .A1(n15102), .A2(n15101), .ZN(n15432) );
  NOR2_X1 U18376 ( .A1(n15432), .A2(n12766), .ZN(n15103) );
  AOI21_X1 U18377 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n12766), .A(n15103), .ZN(
        n15104) );
  OAI21_X1 U18378 ( .B1(n15216), .B2(n15185), .A(n15104), .ZN(P2_U2860) );
  INV_X1 U18379 ( .A(n15447), .ZN(n15110) );
  AOI21_X1 U18380 ( .B1(n15107), .B2(n15106), .A(n15105), .ZN(n15217) );
  NAND2_X1 U18381 ( .A1(n15217), .A2(n15149), .ZN(n15109) );
  NAND2_X1 U18382 ( .A1(n12766), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15108) );
  OAI211_X1 U18383 ( .C1(n15110), .C2(n12766), .A(n15109), .B(n15108), .ZN(
        P2_U2861) );
  OAI21_X1 U18384 ( .B1(n15113), .B2(n15112), .A(n15111), .ZN(n15226) );
  NOR2_X1 U18385 ( .A1(n15159), .A2(n15114), .ZN(n15115) );
  AOI21_X1 U18386 ( .B1(n15468), .B2(n15159), .A(n15115), .ZN(n15116) );
  OAI21_X1 U18387 ( .B1(n15226), .B2(n15185), .A(n15116), .ZN(P2_U2862) );
  AOI21_X1 U18388 ( .B1(n9847), .B2(n15117), .A(n9746), .ZN(n15118) );
  XOR2_X1 U18389 ( .A(n15119), .B(n15118), .Z(n15235) );
  NOR2_X1 U18390 ( .A1(n15124), .A2(n15120), .ZN(n15121) );
  OR2_X1 U18391 ( .A1(n15020), .A2(n15121), .ZN(n16319) );
  MUX2_X1 U18392 ( .A(n16319), .B(n11115), .S(n12766), .Z(n15122) );
  OAI21_X1 U18393 ( .B1(n15235), .B2(n15185), .A(n15122), .ZN(P2_U2863) );
  AND2_X1 U18394 ( .A1(n15133), .A2(n15123), .ZN(n15125) );
  OR2_X1 U18395 ( .A1(n15125), .A2(n15124), .ZN(n16357) );
  AOI21_X1 U18396 ( .B1(n15128), .B2(n15127), .A(n15126), .ZN(n15236) );
  NAND2_X1 U18397 ( .A1(n15236), .A2(n15149), .ZN(n15130) );
  NAND2_X1 U18398 ( .A1(n12766), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15129) );
  OAI211_X1 U18399 ( .C1(n16357), .C2(n12766), .A(n15130), .B(n15129), .ZN(
        P2_U2864) );
  NAND2_X1 U18400 ( .A1(n15039), .A2(n15131), .ZN(n15132) );
  NAND2_X1 U18401 ( .A1(n15133), .A2(n15132), .ZN(n15874) );
  AOI21_X1 U18402 ( .B1(n15134), .B2(n15140), .A(n12455), .ZN(n15248) );
  NAND2_X1 U18403 ( .A1(n15248), .A2(n15149), .ZN(n15136) );
  NAND2_X1 U18404 ( .A1(n12766), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15135) );
  OAI211_X1 U18405 ( .C1(n15874), .C2(n12766), .A(n15136), .B(n15135), .ZN(
        P2_U2865) );
  NAND2_X1 U18406 ( .A1(n15138), .A2(n15137), .ZN(n15139) );
  AND2_X1 U18407 ( .A1(n15140), .A2(n15139), .ZN(n15256) );
  NAND2_X1 U18408 ( .A1(n15256), .A2(n15149), .ZN(n15143) );
  INV_X1 U18409 ( .A(n15509), .ZN(n15141) );
  NAND2_X1 U18410 ( .A1(n15141), .A2(n15159), .ZN(n15142) );
  OAI211_X1 U18411 ( .C1(n15159), .C2(n15144), .A(n15143), .B(n15142), .ZN(
        P2_U2866) );
  INV_X1 U18412 ( .A(n15145), .ZN(n15147) );
  AOI21_X1 U18413 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(n16343) );
  NAND2_X1 U18414 ( .A1(n16343), .A2(n15149), .ZN(n15154) );
  AND2_X1 U18415 ( .A1(n15156), .A2(n15150), .ZN(n15151) );
  NOR2_X1 U18416 ( .A1(n15152), .A2(n15151), .ZN(n19025) );
  NAND2_X1 U18417 ( .A1(n19025), .A2(n15159), .ZN(n15153) );
  OAI211_X1 U18418 ( .C1(n15159), .C2(n11049), .A(n15154), .B(n15153), .ZN(
        P2_U2867) );
  NAND2_X1 U18419 ( .A1(n12766), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15161) );
  INV_X1 U18420 ( .A(n15156), .ZN(n15157) );
  AOI21_X1 U18421 ( .B1(n15158), .B2(n15155), .A(n15157), .ZN(n19039) );
  NAND2_X1 U18422 ( .A1(n19039), .A2(n15159), .ZN(n15160) );
  OAI211_X1 U18423 ( .C1(n15162), .C2(n15185), .A(n15161), .B(n15160), .ZN(
        P2_U2868) );
  AND2_X1 U18424 ( .A1(n15164), .A2(n15163), .ZN(n15165) );
  OR2_X1 U18425 ( .A1(n15166), .A2(n15165), .ZN(n16348) );
  OR2_X1 U18426 ( .A1(n15171), .A2(n15167), .ZN(n15168) );
  AND2_X1 U18427 ( .A1(n15168), .A2(n15155), .ZN(n16366) );
  INV_X1 U18428 ( .A(n16366), .ZN(n19051) );
  MUX2_X1 U18429 ( .A(n19051), .B(n15169), .S(n12766), .Z(n15170) );
  OAI21_X1 U18430 ( .B1(n16348), .B2(n15185), .A(n15170), .ZN(P2_U2869) );
  INV_X1 U18431 ( .A(n15171), .ZN(n15174) );
  NAND2_X1 U18432 ( .A1(n15183), .A2(n15172), .ZN(n15173) );
  NAND2_X1 U18433 ( .A1(n15174), .A2(n15173), .ZN(n19063) );
  NOR2_X1 U18434 ( .A1(n19063), .A2(n12766), .ZN(n15175) );
  AOI21_X1 U18435 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n12766), .A(n15175), .ZN(
        n15176) );
  OAI21_X1 U18436 ( .B1(n15177), .B2(n15185), .A(n15176), .ZN(P2_U2870) );
  NOR2_X1 U18437 ( .A1(n9801), .A2(n15178), .ZN(n15179) );
  OR2_X1 U18438 ( .A1(n13835), .A2(n15179), .ZN(n19249) );
  NAND2_X1 U18439 ( .A1(n15181), .A2(n15180), .ZN(n15182) );
  NAND2_X1 U18440 ( .A1(n15183), .A2(n15182), .ZN(n15582) );
  MUX2_X1 U18441 ( .A(n15582), .B(n11062), .S(n12766), .Z(n15184) );
  OAI21_X1 U18442 ( .B1(n19249), .B2(n15185), .A(n15184), .ZN(P2_U2871) );
  AOI22_X1 U18443 ( .A1(n19248), .A2(BUF2_REG_30__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n15191) );
  NAND2_X1 U18444 ( .A1(n15187), .A2(BUF2_REG_14__SCAN_IN), .ZN(n15189) );
  INV_X1 U18445 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n15186) );
  OR2_X1 U18446 ( .A1(n15187), .A2(n15186), .ZN(n15188) );
  NAND2_X1 U18447 ( .A1(n15189), .A2(n15188), .ZN(n19377) );
  AOI22_X1 U18448 ( .A1(n19246), .A2(n19377), .B1(n19294), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n15190) );
  OAI211_X1 U18449 ( .C1(n16285), .C2(n16349), .A(n15191), .B(n15190), .ZN(
        n15192) );
  AOI21_X1 U18450 ( .B1(n15193), .B2(n19280), .A(n15192), .ZN(n15194) );
  INV_X1 U18451 ( .A(n15194), .ZN(P2_U2889) );
  NAND3_X1 U18452 ( .A1(n15195), .A2(n15087), .A3(n19280), .ZN(n15200) );
  OAI22_X1 U18453 ( .A1(n15250), .A2(n19260), .B1(n19275), .B2(n20903), .ZN(
        n15196) );
  AOI21_X1 U18454 ( .B1(n19295), .B2(n15197), .A(n15196), .ZN(n15199) );
  AOI22_X1 U18455 ( .A1(n19248), .A2(BUF2_REG_29__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15198) );
  NAND3_X1 U18456 ( .A1(n15200), .A2(n15199), .A3(n15198), .ZN(P2_U2890) );
  NOR2_X1 U18457 ( .A1(n15211), .A2(n15201), .ZN(n15202) );
  INV_X1 U18458 ( .A(n16296), .ZN(n15205) );
  OAI22_X1 U18459 ( .A1(n15250), .A2(n19262), .B1(n19275), .B2(n19320), .ZN(
        n15204) );
  AOI21_X1 U18460 ( .B1(n15205), .B2(n19295), .A(n15204), .ZN(n15207) );
  AOI22_X1 U18461 ( .A1(n19248), .A2(BUF2_REG_28__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15206) );
  OAI211_X1 U18462 ( .C1(n15208), .C2(n19299), .A(n15207), .B(n15206), .ZN(
        P2_U2891) );
  AND2_X1 U18463 ( .A1(n15210), .A2(n15209), .ZN(n15212) );
  OR2_X1 U18464 ( .A1(n15212), .A2(n15211), .ZN(n16318) );
  INV_X1 U18465 ( .A(n16318), .ZN(n15435) );
  OAI22_X1 U18466 ( .A1(n15250), .A2(n19264), .B1(n19275), .B2(n19322), .ZN(
        n15213) );
  AOI21_X1 U18467 ( .B1(n15435), .B2(n19295), .A(n15213), .ZN(n15215) );
  AOI22_X1 U18468 ( .A1(n19248), .A2(BUF2_REG_27__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15214) );
  OAI211_X1 U18469 ( .C1(n15216), .C2(n19299), .A(n15215), .B(n15214), .ZN(
        P2_U2892) );
  NAND2_X1 U18470 ( .A1(n15217), .A2(n19280), .ZN(n15221) );
  AOI22_X1 U18471 ( .A1(n19246), .A2(n19266), .B1(n19294), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15220) );
  AOI22_X1 U18472 ( .A1(n19248), .A2(BUF2_REG_26__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15219) );
  NAND2_X1 U18473 ( .A1(n19295), .A2(n15449), .ZN(n15218) );
  NAND4_X1 U18474 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        P2_U2893) );
  INV_X1 U18475 ( .A(n19269), .ZN(n15222) );
  OAI22_X1 U18476 ( .A1(n15250), .A2(n15222), .B1(n19275), .B2(n19326), .ZN(
        n15223) );
  AOI21_X1 U18477 ( .B1(n19295), .B2(n15460), .A(n15223), .ZN(n15225) );
  AOI22_X1 U18478 ( .A1(n19248), .A2(BUF2_REG_25__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15224) );
  OAI211_X1 U18479 ( .C1(n15226), .C2(n19299), .A(n15225), .B(n15224), .ZN(
        P2_U2894) );
  NOR2_X1 U18480 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  OR2_X1 U18481 ( .A1(n15230), .A2(n15229), .ZN(n16330) );
  INV_X1 U18482 ( .A(n16330), .ZN(n15232) );
  INV_X1 U18483 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19328) );
  OAI22_X1 U18484 ( .A1(n15250), .A2(n19272), .B1(n19275), .B2(n19328), .ZN(
        n15231) );
  AOI21_X1 U18485 ( .B1(n19295), .B2(n15232), .A(n15231), .ZN(n15234) );
  AOI22_X1 U18486 ( .A1(n19248), .A2(BUF2_REG_24__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15233) );
  OAI211_X1 U18487 ( .C1(n15235), .C2(n19299), .A(n15234), .B(n15233), .ZN(
        P2_U2895) );
  NAND2_X1 U18488 ( .A1(n15236), .A2(n19280), .ZN(n15242) );
  INV_X1 U18489 ( .A(n19433), .ZN(n15237) );
  AOI22_X1 U18490 ( .A1(n19246), .A2(n15237), .B1(n19294), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15241) );
  AOI22_X1 U18491 ( .A1(n19248), .A2(BUF2_REG_23__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15240) );
  XNOR2_X1 U18492 ( .A(n15238), .B(n9845), .ZN(n16332) );
  NAND2_X1 U18493 ( .A1(n19295), .A2(n16332), .ZN(n15239) );
  NAND4_X1 U18494 ( .A1(n15242), .A2(n15241), .A3(n15240), .A4(n15239), .ZN(
        P2_U2896) );
  XNOR2_X1 U18495 ( .A(n15243), .B(n15035), .ZN(n15878) );
  AOI22_X1 U18496 ( .A1(n19248), .A2(BUF2_REG_22__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15246) );
  INV_X1 U18497 ( .A(n19426), .ZN(n15244) );
  AOI22_X1 U18498 ( .A1(n19246), .A2(n15244), .B1(n19294), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15245) );
  OAI211_X1 U18499 ( .C1(n16349), .C2(n15878), .A(n15246), .B(n15245), .ZN(
        n15247) );
  AOI21_X1 U18500 ( .B1(n15248), .B2(n19280), .A(n15247), .ZN(n15249) );
  INV_X1 U18501 ( .A(n15249), .ZN(P2_U2897) );
  OAI22_X1 U18502 ( .A1(n15250), .A2(n19277), .B1(n19275), .B2(n20873), .ZN(
        n15251) );
  AOI21_X1 U18503 ( .B1(n19248), .B2(BUF2_REG_21__SCAN_IN), .A(n15251), .ZN(
        n15252) );
  OAI21_X1 U18504 ( .B1(n15254), .B2(n15253), .A(n15252), .ZN(n15255) );
  AOI21_X1 U18505 ( .B1(n15256), .B2(n19280), .A(n15255), .ZN(n15257) );
  OAI21_X1 U18506 ( .B1(n15517), .B2(n16349), .A(n15257), .ZN(P2_U2898) );
  NAND2_X1 U18507 ( .A1(n15258), .A2(n16435), .ZN(n15264) );
  XNOR2_X1 U18508 ( .A(n15259), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16290) );
  NAND2_X1 U18509 ( .A1(n16409), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15260) );
  OAI211_X1 U18510 ( .C1(n16290), .C2(n16424), .A(n15261), .B(n15260), .ZN(
        n15262) );
  AOI21_X1 U18511 ( .B1(n16287), .B2(n16421), .A(n15262), .ZN(n15263) );
  OAI211_X1 U18512 ( .C1(n15265), .C2(n16425), .A(n15264), .B(n15263), .ZN(
        P2_U2984) );
  NAND2_X1 U18513 ( .A1(n15267), .A2(n15266), .ZN(n15269) );
  XOR2_X1 U18514 ( .A(n15269), .B(n15268), .Z(n15422) );
  AOI21_X1 U18515 ( .B1(n15271), .B2(n11653), .A(n15270), .ZN(n15410) );
  NAND2_X1 U18516 ( .A1(n15410), .A2(n16435), .ZN(n15276) );
  NAND2_X1 U18517 ( .A1(n19180), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15413) );
  NAND2_X1 U18518 ( .A1(n16409), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15272) );
  OAI211_X1 U18519 ( .C1(n15273), .C2(n16424), .A(n15413), .B(n15272), .ZN(
        n15274) );
  AOI21_X1 U18520 ( .B1(n15416), .B2(n16421), .A(n15274), .ZN(n15275) );
  OAI211_X1 U18521 ( .C1(n15422), .C2(n16425), .A(n15276), .B(n15275), .ZN(
        P2_U2985) );
  XNOR2_X1 U18522 ( .A(n15277), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15445) );
  AOI21_X1 U18523 ( .B1(n15437), .B2(n15278), .A(n11652), .ZN(n15443) );
  NAND2_X1 U18524 ( .A1(n19180), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15433) );
  OAI21_X1 U18525 ( .B1(n16445), .B2(n16306), .A(n15433), .ZN(n15279) );
  AOI21_X1 U18526 ( .B1(n15280), .B2(n16434), .A(n15279), .ZN(n15281) );
  OAI21_X1 U18527 ( .B1(n15432), .B2(n16439), .A(n15281), .ZN(n15282) );
  AOI21_X1 U18528 ( .B1(n15443), .B2(n16435), .A(n15282), .ZN(n15283) );
  OAI21_X1 U18529 ( .B1(n15445), .B2(n16425), .A(n15283), .ZN(P2_U2987) );
  NOR2_X1 U18530 ( .A1(n15309), .A2(n15463), .ZN(n15298) );
  OAI21_X1 U18531 ( .B1(n15298), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15278), .ZN(n15457) );
  INV_X1 U18532 ( .A(n15285), .ZN(n15286) );
  OAI21_X1 U18533 ( .B1(n15286), .B2(n15296), .A(n15294), .ZN(n15288) );
  XNOR2_X1 U18534 ( .A(n15288), .B(n15287), .ZN(n15455) );
  NAND2_X1 U18535 ( .A1(n15447), .A2(n16421), .ZN(n15290) );
  NOR2_X1 U18536 ( .A1(n19210), .A2(n20937), .ZN(n15448) );
  AOI21_X1 U18537 ( .B1(n16409), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15448), .ZN(n15289) );
  OAI211_X1 U18538 ( .C1(n16424), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        n15292) );
  AOI21_X1 U18539 ( .B1(n15455), .B2(n16441), .A(n15292), .ZN(n15293) );
  OAI21_X1 U18540 ( .B1(n15457), .B2(n16427), .A(n15293), .ZN(P2_U2988) );
  INV_X1 U18541 ( .A(n15294), .ZN(n15295) );
  NOR2_X1 U18542 ( .A1(n15296), .A2(n15295), .ZN(n15297) );
  XNOR2_X1 U18543 ( .A(n15285), .B(n15297), .ZN(n15471) );
  INV_X1 U18544 ( .A(n15298), .ZN(n15459) );
  NAND2_X1 U18545 ( .A1(n15309), .A2(n15463), .ZN(n15458) );
  NAND3_X1 U18546 ( .A1(n15459), .A2(n16435), .A3(n15458), .ZN(n15303) );
  NAND2_X1 U18547 ( .A1(n19180), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U18548 ( .A1(n16409), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15299) );
  OAI211_X1 U18549 ( .C1(n15300), .C2(n16424), .A(n15462), .B(n15299), .ZN(
        n15301) );
  AOI21_X1 U18550 ( .B1(n15468), .B2(n16421), .A(n15301), .ZN(n15302) );
  OAI211_X1 U18551 ( .C1(n16425), .C2(n15471), .A(n15303), .B(n15302), .ZN(
        P2_U2989) );
  NOR2_X1 U18552 ( .A1(n15306), .A2(n11121), .ZN(n15307) );
  XNOR2_X1 U18553 ( .A(n9719), .B(n15307), .ZN(n15482) );
  AOI21_X1 U18554 ( .B1(n15474), .B2(n15308), .A(n15284), .ZN(n15472) );
  NAND2_X1 U18555 ( .A1(n15472), .A2(n16435), .ZN(n15313) );
  OAI22_X1 U18556 ( .A1(n11542), .A2(n19210), .B1(n16424), .B2(n16327), .ZN(
        n15311) );
  NOR2_X1 U18557 ( .A1(n16319), .A2(n16439), .ZN(n15310) );
  AOI211_X1 U18558 ( .C1(n16409), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15311), .B(n15310), .ZN(n15312) );
  OAI211_X1 U18559 ( .C1(n15482), .C2(n16425), .A(n15313), .B(n15312), .ZN(
        P2_U2990) );
  INV_X1 U18560 ( .A(n15314), .ZN(n15315) );
  OAI21_X1 U18561 ( .B1(n15315), .B2(n15514), .A(n15487), .ZN(n15317) );
  NAND2_X1 U18562 ( .A1(n15317), .A2(n15484), .ZN(n15508) );
  NAND2_X1 U18563 ( .A1(n15320), .A2(n15319), .ZN(n15321) );
  XNOR2_X1 U18564 ( .A(n15318), .B(n15321), .ZN(n15505) );
  INV_X1 U18565 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20005) );
  OAI22_X1 U18566 ( .A1(n20005), .A2(n19210), .B1(n16424), .B2(n15869), .ZN(
        n15322) );
  AOI21_X1 U18567 ( .B1(n16409), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15322), .ZN(n15323) );
  OAI21_X1 U18568 ( .B1(n15874), .B2(n16439), .A(n15323), .ZN(n15324) );
  AOI21_X1 U18569 ( .B1(n15505), .B2(n16441), .A(n15324), .ZN(n15325) );
  OAI21_X1 U18570 ( .B1(n15508), .B2(n16427), .A(n15325), .ZN(P2_U2992) );
  OAI21_X1 U18571 ( .B1(n15624), .B2(n9938), .A(n10228), .ZN(n15328) );
  INV_X1 U18572 ( .A(n15329), .ZN(n15375) );
  NAND2_X1 U18573 ( .A1(n15332), .A2(n15331), .ZN(n15364) );
  NAND2_X1 U18574 ( .A1(n15552), .A2(n15549), .ZN(n15351) );
  NAND2_X1 U18575 ( .A1(n15334), .A2(n15333), .ZN(n15345) );
  XNOR2_X1 U18576 ( .A(n15335), .B(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15336) );
  XOR2_X1 U18577 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15314), .Z(
        n15519) );
  NAND2_X1 U18578 ( .A1(n19180), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15510) );
  OAI21_X1 U18579 ( .B1(n16445), .B2(n15337), .A(n15510), .ZN(n15338) );
  AOI21_X1 U18580 ( .B1(n16434), .B2(n15339), .A(n15338), .ZN(n15340) );
  OAI21_X1 U18581 ( .B1(n15509), .B2(n16439), .A(n15340), .ZN(n15341) );
  AOI21_X1 U18582 ( .B1(n15519), .B2(n16435), .A(n15341), .ZN(n15342) );
  OAI21_X1 U18583 ( .B1(n15521), .B2(n16425), .A(n15342), .ZN(P2_U2993) );
  NOR2_X1 U18584 ( .A1(n15343), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15344) );
  OR2_X1 U18585 ( .A1(n15314), .A2(n15344), .ZN(n15537) );
  NAND2_X1 U18586 ( .A1(n15346), .A2(n15345), .ZN(n15522) );
  NAND3_X1 U18587 ( .A1(n15523), .A2(n15522), .A3(n16441), .ZN(n15350) );
  NOR2_X1 U18588 ( .A1(n19210), .A2(n20002), .ZN(n15531) );
  AOI21_X1 U18589 ( .B1(n16409), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15531), .ZN(n15347) );
  OAI21_X1 U18590 ( .B1(n16424), .B2(n19027), .A(n15347), .ZN(n15348) );
  AOI21_X1 U18591 ( .B1(n19025), .B2(n16421), .A(n15348), .ZN(n15349) );
  OAI211_X1 U18592 ( .C1(n16427), .C2(n15537), .A(n15350), .B(n15349), .ZN(
        P2_U2994) );
  NAND2_X1 U18593 ( .A1(n15351), .A2(n15550), .ZN(n15356) );
  INV_X1 U18594 ( .A(n15352), .ZN(n15354) );
  NAND2_X1 U18595 ( .A1(n15354), .A2(n15353), .ZN(n15355) );
  XNOR2_X1 U18596 ( .A(n15356), .B(n15355), .ZN(n15548) );
  NAND2_X1 U18597 ( .A1(n19035), .A2(n16434), .ZN(n15357) );
  NAND2_X1 U18598 ( .A1(n19180), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15538) );
  OAI211_X1 U18599 ( .C1(n16445), .C2(n15358), .A(n15357), .B(n15538), .ZN(
        n15361) );
  INV_X1 U18600 ( .A(n15359), .ZN(n15555) );
  NOR2_X1 U18601 ( .A1(n15359), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15544) );
  NOR3_X1 U18602 ( .A1(n15544), .A2(n15343), .A3(n16427), .ZN(n15360) );
  AOI211_X1 U18603 ( .C1(n16421), .C2(n19039), .A(n15361), .B(n15360), .ZN(
        n15362) );
  OAI21_X1 U18604 ( .B1(n15548), .B2(n16425), .A(n15362), .ZN(P2_U2995) );
  XOR2_X1 U18605 ( .A(n15364), .B(n15363), .Z(n15578) );
  INV_X1 U18606 ( .A(n15569), .ZN(n15377) );
  INV_X1 U18607 ( .A(n15365), .ZN(n15366) );
  AOI211_X1 U18608 ( .C1(n15377), .C2(n15367), .A(n15366), .B(n16427), .ZN(
        n15373) );
  NAND2_X1 U18609 ( .A1(n19180), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15572) );
  INV_X1 U18610 ( .A(n15572), .ZN(n15372) );
  NOR2_X1 U18611 ( .A1(n19063), .A2(n16439), .ZN(n15371) );
  INV_X1 U18612 ( .A(n15368), .ZN(n19059) );
  OAI22_X1 U18613 ( .A1(n15369), .A2(n16445), .B1(n16424), .B2(n19059), .ZN(
        n15370) );
  NOR4_X1 U18614 ( .A1(n15373), .A2(n15372), .A3(n15371), .A4(n15370), .ZN(
        n15374) );
  OAI21_X1 U18615 ( .B1(n15578), .B2(n16425), .A(n15374), .ZN(P2_U2997) );
  XNOR2_X1 U18616 ( .A(n15376), .B(n15375), .ZN(n15583) );
  INV_X1 U18617 ( .A(n15591), .ZN(n15378) );
  OAI211_X1 U18618 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15378), .A(
        n15377), .B(n16435), .ZN(n15382) );
  INV_X1 U18619 ( .A(n15582), .ZN(n19076) );
  AOI22_X1 U18620 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n19180), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16409), .ZN(n15379) );
  OAI21_X1 U18621 ( .B1(n16424), .B2(n19070), .A(n15379), .ZN(n15380) );
  AOI21_X1 U18622 ( .B1(n19076), .B2(n16421), .A(n15380), .ZN(n15381) );
  OAI211_X1 U18623 ( .C1(n15583), .C2(n16425), .A(n15382), .B(n15381), .ZN(
        P2_U2998) );
  OAI21_X1 U18624 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n9781), .A(
        n9925), .ZN(n15665) );
  NAND2_X1 U18625 ( .A1(n15385), .A2(n15384), .ZN(n15389) );
  INV_X1 U18626 ( .A(n15386), .ZN(n15669) );
  NOR2_X1 U18627 ( .A1(n15387), .A2(n15669), .ZN(n15388) );
  XOR2_X1 U18628 ( .A(n15389), .B(n15388), .Z(n15663) );
  INV_X1 U18629 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20870) );
  OAI22_X1 U18630 ( .A1(n20870), .A2(n15581), .B1(n16424), .B2(n19126), .ZN(
        n15391) );
  OAI22_X1 U18631 ( .A1(n19132), .A2(n16439), .B1(n10097), .B2(n16445), .ZN(
        n15390) );
  AOI211_X1 U18632 ( .C1(n15663), .C2(n16441), .A(n15391), .B(n15390), .ZN(
        n15392) );
  OAI21_X1 U18633 ( .B1(n15665), .B2(n16427), .A(n15392), .ZN(P2_U3004) );
  XNOR2_X1 U18634 ( .A(n15393), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15692) );
  NAND2_X1 U18635 ( .A1(n16414), .A2(n16416), .ZN(n15395) );
  XNOR2_X1 U18636 ( .A(n15394), .B(n15395), .ZN(n15690) );
  OAI22_X1 U18637 ( .A1(n15396), .A2(n16445), .B1(n19982), .B2(n15581), .ZN(
        n15399) );
  INV_X1 U18638 ( .A(n19164), .ZN(n15397) );
  OAI22_X1 U18639 ( .A1(n16439), .A2(n19169), .B1(n16424), .B2(n15397), .ZN(
        n15398) );
  AOI211_X1 U18640 ( .C1(n15690), .C2(n16441), .A(n15399), .B(n15398), .ZN(
        n15400) );
  OAI21_X1 U18641 ( .B1(n15692), .B2(n16427), .A(n15400), .ZN(P2_U3007) );
  XNOR2_X1 U18642 ( .A(n15401), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15703) );
  OAI21_X1 U18643 ( .B1(n15404), .B2(n15403), .A(n15402), .ZN(n15405) );
  INV_X1 U18644 ( .A(n15405), .ZN(n15700) );
  OAI22_X1 U18645 ( .A1(n19980), .A2(n15581), .B1(n16424), .B2(n19182), .ZN(
        n15408) );
  INV_X1 U18646 ( .A(n19184), .ZN(n15406) );
  OAI22_X1 U18647 ( .A1(n16439), .A2(n15406), .B1(n16445), .B2(n10101), .ZN(
        n15407) );
  AOI211_X1 U18648 ( .C1(n15700), .C2(n16441), .A(n15408), .B(n15407), .ZN(
        n15409) );
  OAI21_X1 U18649 ( .B1(n15703), .B2(n16427), .A(n15409), .ZN(P2_U3008) );
  NAND2_X1 U18650 ( .A1(n15410), .A2(n19391), .ZN(n15421) );
  INV_X1 U18651 ( .A(n15441), .ZN(n15411) );
  NAND2_X1 U18652 ( .A1(n10214), .A2(n15411), .ZN(n15412) );
  OAI211_X1 U18653 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15571), .A(
        n15412), .B(n15438), .ZN(n15428) );
  OAI21_X1 U18654 ( .B1(n19400), .B2(n15414), .A(n15413), .ZN(n15415) );
  AOI21_X1 U18655 ( .B1(n15416), .B2(n16475), .A(n15415), .ZN(n15417) );
  OAI21_X1 U18656 ( .B1(n15418), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15417), .ZN(n15419) );
  AOI21_X1 U18657 ( .B1(n15428), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15419), .ZN(n15420) );
  OAI211_X1 U18658 ( .C1(n15422), .C2(n16477), .A(n15421), .B(n15420), .ZN(
        P2_U3017) );
  NAND2_X1 U18659 ( .A1(n15423), .A2(n19395), .ZN(n15430) );
  OAI21_X1 U18660 ( .B1(n15441), .B2(n15437), .A(n10214), .ZN(n15427) );
  NOR2_X1 U18661 ( .A1(n16297), .A2(n19404), .ZN(n15426) );
  OAI21_X1 U18662 ( .B1(n19400), .B2(n16296), .A(n15424), .ZN(n15425) );
  OAI211_X1 U18663 ( .C1(n15702), .C2(n15431), .A(n15430), .B(n15429), .ZN(
        P2_U3018) );
  INV_X1 U18664 ( .A(n15432), .ZN(n16312) );
  INV_X1 U18665 ( .A(n15433), .ZN(n15434) );
  AOI21_X1 U18666 ( .B1(n16474), .B2(n15435), .A(n15434), .ZN(n15436) );
  OAI21_X1 U18667 ( .B1(n15438), .B2(n15437), .A(n15436), .ZN(n15439) );
  AOI21_X1 U18668 ( .B1(n16312), .B2(n16475), .A(n15439), .ZN(n15440) );
  OAI21_X1 U18669 ( .B1(n15441), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15440), .ZN(n15442) );
  AOI21_X1 U18670 ( .B1(n15443), .B2(n19391), .A(n15442), .ZN(n15444) );
  OAI21_X1 U18671 ( .B1(n15445), .B2(n16477), .A(n15444), .ZN(P2_U3019) );
  AOI211_X1 U18672 ( .C1(n15463), .C2(n15452), .A(n11251), .B(n15465), .ZN(
        n15454) );
  NAND2_X1 U18673 ( .A1(n15447), .A2(n16475), .ZN(n15451) );
  AOI21_X1 U18674 ( .B1(n16474), .B2(n15449), .A(n15448), .ZN(n15450) );
  OAI211_X1 U18675 ( .C1(n15464), .C2(n15452), .A(n15451), .B(n15450), .ZN(
        n15453) );
  AOI211_X1 U18676 ( .C1(n15455), .C2(n19395), .A(n15454), .B(n15453), .ZN(
        n15456) );
  OAI21_X1 U18677 ( .B1(n15457), .B2(n15702), .A(n15456), .ZN(P2_U3020) );
  NAND3_X1 U18678 ( .A1(n15459), .A2(n19391), .A3(n15458), .ZN(n15470) );
  NAND2_X1 U18679 ( .A1(n16474), .A2(n15460), .ZN(n15461) );
  OAI211_X1 U18680 ( .C1(n15464), .C2(n15463), .A(n15462), .B(n15461), .ZN(
        n15467) );
  NOR2_X1 U18681 ( .A1(n15465), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15466) );
  AOI211_X1 U18682 ( .C1(n15468), .C2(n16475), .A(n15467), .B(n15466), .ZN(
        n15469) );
  OAI211_X1 U18683 ( .C1(n15471), .C2(n16477), .A(n15470), .B(n15469), .ZN(
        P2_U3021) );
  NAND2_X1 U18684 ( .A1(n15472), .A2(n19391), .ZN(n15481) );
  AND2_X1 U18685 ( .A1(n15473), .A2(n15515), .ZN(n15475) );
  AOI22_X1 U18686 ( .A1(n19180), .A2(P2_REIP_REG_24__SCAN_IN), .B1(n15475), 
        .B2(n15474), .ZN(n15476) );
  OAI21_X1 U18687 ( .B1(n19400), .B2(n16330), .A(n15476), .ZN(n15478) );
  NOR2_X1 U18688 ( .A1(n16319), .A2(n19404), .ZN(n15477) );
  AOI211_X1 U18689 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n15479), .A(
        n15478), .B(n15477), .ZN(n15480) );
  OAI211_X1 U18690 ( .C1(n15482), .C2(n16477), .A(n15481), .B(n15480), .ZN(
        P2_U3022) );
  INV_X1 U18691 ( .A(n15308), .ZN(n15483) );
  INV_X1 U18692 ( .A(n16359), .ZN(n15497) );
  NAND2_X1 U18693 ( .A1(n15515), .A2(n15514), .ZN(n15485) );
  NAND2_X1 U18694 ( .A1(n15511), .A2(n15485), .ZN(n15504) );
  NAND2_X1 U18695 ( .A1(n15515), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15501) );
  AOI221_X1 U18696 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C1(n15487), .C2(n15486), .A(
        n15501), .ZN(n15489) );
  NOR2_X1 U18697 ( .A1(n19210), .A2(n21070), .ZN(n15488) );
  AOI211_X1 U18698 ( .C1(n16474), .C2(n16332), .A(n15489), .B(n15488), .ZN(
        n15490) );
  OAI21_X1 U18699 ( .B1(n16357), .B2(n19404), .A(n15490), .ZN(n15491) );
  AOI21_X1 U18700 ( .B1(n15504), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15491), .ZN(n15496) );
  OR2_X1 U18701 ( .A1(n15493), .A2(n15492), .ZN(n16355) );
  NAND3_X1 U18702 ( .A1(n16355), .A2(n19395), .A3(n15494), .ZN(n15495) );
  OAI211_X1 U18703 ( .C1(n15497), .C2(n15702), .A(n15496), .B(n15495), .ZN(
        P2_U3023) );
  INV_X1 U18704 ( .A(n15878), .ZN(n15499) );
  NOR2_X1 U18705 ( .A1(n20005), .A2(n19210), .ZN(n15498) );
  AOI21_X1 U18706 ( .B1(n16474), .B2(n15499), .A(n15498), .ZN(n15500) );
  OAI21_X1 U18707 ( .B1(n15874), .B2(n19404), .A(n15500), .ZN(n15503) );
  NOR2_X1 U18708 ( .A1(n15501), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15502) );
  AOI211_X1 U18709 ( .C1(n15504), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15503), .B(n15502), .ZN(n15507) );
  NAND2_X1 U18710 ( .A1(n15505), .A2(n19395), .ZN(n15506) );
  OAI211_X1 U18711 ( .C1(n15508), .C2(n15702), .A(n15507), .B(n15506), .ZN(
        P2_U3024) );
  NOR2_X1 U18712 ( .A1(n15509), .A2(n19404), .ZN(n15513) );
  OAI21_X1 U18713 ( .B1(n15511), .B2(n15514), .A(n15510), .ZN(n15512) );
  AOI211_X1 U18714 ( .C1(n15515), .C2(n15514), .A(n15513), .B(n15512), .ZN(
        n15516) );
  OAI21_X1 U18715 ( .B1(n15517), .B2(n19400), .A(n15516), .ZN(n15518) );
  AOI21_X1 U18716 ( .B1(n15519), .B2(n19391), .A(n15518), .ZN(n15520) );
  OAI21_X1 U18717 ( .B1(n15521), .B2(n16477), .A(n15520), .ZN(P2_U3025) );
  NAND3_X1 U18718 ( .A1(n15523), .A2(n15522), .A3(n19395), .ZN(n15536) );
  NOR2_X1 U18719 ( .A1(n15525), .A2(n15524), .ZN(n15526) );
  XNOR2_X1 U18720 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15533) );
  INV_X1 U18721 ( .A(n15646), .ZN(n15568) );
  AOI21_X1 U18722 ( .B1(n15528), .B2(n16479), .A(n15527), .ZN(n15560) );
  NOR3_X1 U18723 ( .A1(n15568), .A2(n15560), .A3(n15529), .ZN(n15530) );
  AOI211_X1 U18724 ( .C1(n19025), .C2(n16475), .A(n15531), .B(n15530), .ZN(
        n15532) );
  OAI21_X1 U18725 ( .B1(n15543), .B2(n15533), .A(n15532), .ZN(n15534) );
  AOI21_X1 U18726 ( .B1(n10220), .B2(n16474), .A(n15534), .ZN(n15535) );
  OAI211_X1 U18727 ( .C1(n15537), .C2(n15702), .A(n15536), .B(n15535), .ZN(
        P2_U3026) );
  INV_X1 U18728 ( .A(n15538), .ZN(n15541) );
  NOR3_X1 U18729 ( .A1(n15568), .A2(n15560), .A3(n15539), .ZN(n15540) );
  AOI211_X1 U18730 ( .C1(n19039), .C2(n16475), .A(n15541), .B(n15540), .ZN(
        n15542) );
  OAI21_X1 U18731 ( .B1(n15543), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15542), .ZN(n15546) );
  NOR3_X1 U18732 ( .A1(n15544), .A2(n15343), .A3(n15702), .ZN(n15545) );
  AOI211_X1 U18733 ( .C1(n16474), .C2(n19040), .A(n15546), .B(n15545), .ZN(
        n15547) );
  OAI21_X1 U18734 ( .B1(n15548), .B2(n16477), .A(n15547), .ZN(P2_U3027) );
  NAND2_X1 U18735 ( .A1(n15550), .A2(n15549), .ZN(n15551) );
  XNOR2_X1 U18736 ( .A(n15552), .B(n15551), .ZN(n16364) );
  NAND2_X1 U18737 ( .A1(n15365), .A2(n15553), .ZN(n15554) );
  NAND2_X1 U18738 ( .A1(n15555), .A2(n15554), .ZN(n16363) );
  INV_X1 U18739 ( .A(n16363), .ZN(n15566) );
  NAND2_X1 U18740 ( .A1(n15557), .A2(n15556), .ZN(n15558) );
  NAND2_X1 U18741 ( .A1(n15559), .A2(n15558), .ZN(n19052) );
  INV_X1 U18742 ( .A(n15560), .ZN(n15561) );
  OAI21_X1 U18743 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15562), .A(
        n15561), .ZN(n15564) );
  AOI22_X1 U18744 ( .A1(n16366), .A2(n16475), .B1(P2_REIP_REG_18__SCAN_IN), 
        .B2(n19180), .ZN(n15563) );
  OAI211_X1 U18745 ( .C1(n19052), .C2(n19400), .A(n15564), .B(n15563), .ZN(
        n15565) );
  AOI21_X1 U18746 ( .B1(n15566), .B2(n19391), .A(n15565), .ZN(n15567) );
  OAI21_X1 U18747 ( .B1(n16364), .B2(n16477), .A(n15567), .ZN(P2_U3028) );
  AOI21_X1 U18748 ( .B1(n15630), .B2(n9808), .A(n15568), .ZN(n15604) );
  AOI21_X1 U18749 ( .B1(n15702), .B2(n19387), .A(n15569), .ZN(n15570) );
  OAI21_X1 U18750 ( .B1(n19063), .B2(n19404), .A(n15572), .ZN(n15576) );
  INV_X1 U18751 ( .A(n16452), .ZN(n15573) );
  AOI22_X1 U18752 ( .A1(n16375), .A2(n19391), .B1(n9808), .B2(n15573), .ZN(
        n15586) );
  NOR3_X1 U18753 ( .A1(n15586), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15574), .ZN(n15575) );
  AOI211_X1 U18754 ( .C1(n16474), .C2(n19065), .A(n15576), .B(n15575), .ZN(
        n15577) );
  AND2_X1 U18755 ( .A1(n15596), .A2(n15579), .ZN(n15580) );
  NOR2_X1 U18756 ( .A1(n13837), .A2(n15580), .ZN(n19251) );
  INV_X1 U18757 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19997) );
  OAI22_X1 U18758 ( .A1(n15582), .A2(n19404), .B1(n19997), .B2(n15581), .ZN(
        n15585) );
  NOR2_X1 U18759 ( .A1(n15583), .A2(n16477), .ZN(n15584) );
  AOI211_X1 U18760 ( .C1(n16474), .C2(n19251), .A(n15585), .B(n15584), .ZN(
        n15588) );
  OR3_X1 U18761 ( .A1(n15586), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15601), .ZN(n15587) );
  OAI211_X1 U18762 ( .C1(n15590), .C2(n15589), .A(n15588), .B(n15587), .ZN(
        P2_U3030) );
  NAND2_X1 U18763 ( .A1(n15593), .A2(n15592), .ZN(n15594) );
  XNOR2_X1 U18764 ( .A(n15595), .B(n15594), .ZN(n16372) );
  OAI21_X1 U18765 ( .B1(n16447), .B2(n15597), .A(n15596), .ZN(n19256) );
  NOR2_X1 U18766 ( .A1(n15598), .A2(n16452), .ZN(n15600) );
  INV_X1 U18767 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19995) );
  NOR2_X1 U18768 ( .A1(n19995), .A2(n19210), .ZN(n15599) );
  AOI21_X1 U18769 ( .B1(n15601), .B2(n15600), .A(n15599), .ZN(n15602) );
  OAI21_X1 U18770 ( .B1(n19085), .B2(n19404), .A(n15602), .ZN(n15603) );
  AOI21_X1 U18771 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15604), .A(
        n15603), .ZN(n15605) );
  OAI21_X1 U18772 ( .B1(n19256), .B2(n19400), .A(n15605), .ZN(n15606) );
  AOI21_X1 U18773 ( .B1(n16372), .B2(n19395), .A(n15606), .ZN(n15607) );
  OAI21_X1 U18774 ( .B1(n16369), .B2(n15702), .A(n15607), .ZN(P2_U3031) );
  OAI21_X1 U18775 ( .B1(n15621), .B2(n20891), .A(n11290), .ZN(n15608) );
  NAND2_X1 U18776 ( .A1(n16376), .A2(n15608), .ZN(n16388) );
  NAND2_X1 U18777 ( .A1(n15610), .A2(n15609), .ZN(n15612) );
  XOR2_X1 U18778 ( .A(n15612), .B(n15611), .Z(n16390) );
  OAI21_X1 U18779 ( .B1(n15614), .B2(n15613), .A(n16449), .ZN(n19261) );
  OR2_X1 U18780 ( .A1(n16452), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15633) );
  NAND2_X1 U18781 ( .A1(n15633), .A2(n15630), .ZN(n16456) );
  NAND2_X1 U18782 ( .A1(n16456), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15618) );
  NOR2_X1 U18783 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16452), .ZN(
        n16457) );
  INV_X1 U18784 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19992) );
  NOR2_X1 U18785 ( .A1(n19992), .A2(n19210), .ZN(n15616) );
  NOR2_X1 U18786 ( .A1(n16389), .A2(n19404), .ZN(n15615) );
  AOI211_X1 U18787 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16457), .A(
        n15616), .B(n15615), .ZN(n15617) );
  OAI211_X1 U18788 ( .C1(n19261), .C2(n19400), .A(n15618), .B(n15617), .ZN(
        n15619) );
  AOI21_X1 U18789 ( .B1(n16390), .B2(n19395), .A(n15619), .ZN(n15620) );
  OAI21_X1 U18790 ( .B1(n16388), .B2(n15702), .A(n15620), .ZN(P2_U3033) );
  XNOR2_X1 U18791 ( .A(n15621), .B(n20891), .ZN(n16395) );
  INV_X1 U18792 ( .A(n15622), .ZN(n15623) );
  NAND2_X1 U18793 ( .A1(n15624), .A2(n15623), .ZN(n15627) );
  NOR2_X1 U18794 ( .A1(n9938), .A2(n15625), .ZN(n15626) );
  XNOR2_X1 U18795 ( .A(n15627), .B(n15626), .ZN(n16394) );
  NAND2_X1 U18796 ( .A1(n16397), .A2(n16475), .ZN(n15629) );
  NAND2_X1 U18797 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n11600), .ZN(n15628) );
  OAI211_X1 U18798 ( .C1(n20891), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        n15631) );
  AOI21_X1 U18799 ( .B1(n15632), .B2(n16474), .A(n15631), .ZN(n15634) );
  OAI211_X1 U18800 ( .C1(n16394), .C2(n16477), .A(n15634), .B(n15633), .ZN(
        n15635) );
  INV_X1 U18801 ( .A(n15635), .ZN(n15636) );
  OAI21_X1 U18802 ( .B1(n16395), .B2(n15702), .A(n15636), .ZN(P2_U3034) );
  AOI21_X1 U18803 ( .B1(n15638), .B2(n9925), .A(n15637), .ZN(n16401) );
  INV_X1 U18804 ( .A(n16401), .ZN(n15654) );
  NAND2_X1 U18805 ( .A1(n15640), .A2(n15639), .ZN(n15643) );
  NAND2_X1 U18806 ( .A1(n10215), .A2(n15641), .ZN(n15642) );
  XNOR2_X1 U18807 ( .A(n15643), .B(n15642), .ZN(n16402) );
  INV_X1 U18808 ( .A(n15644), .ZN(n15658) );
  AOI211_X1 U18809 ( .C1(n15657), .C2(n15638), .A(n15645), .B(n15658), .ZN(
        n15652) );
  NAND2_X1 U18810 ( .A1(n15676), .A2(n15646), .ZN(n15656) );
  OAI21_X1 U18811 ( .B1(n9795), .B2(n15647), .A(n13311), .ZN(n19265) );
  INV_X1 U18812 ( .A(n19265), .ZN(n15648) );
  NAND2_X1 U18813 ( .A1(n15648), .A2(n16474), .ZN(n15650) );
  AOI22_X1 U18814 ( .A1(n19121), .A2(n16475), .B1(P2_REIP_REG_11__SCAN_IN), 
        .B2(n19180), .ZN(n15649) );
  OAI211_X1 U18815 ( .C1(n15638), .C2(n15656), .A(n15650), .B(n15649), .ZN(
        n15651) );
  AOI211_X1 U18816 ( .C1(n16402), .C2(n19395), .A(n15652), .B(n15651), .ZN(
        n15653) );
  OAI21_X1 U18817 ( .B1(n15654), .B2(n15702), .A(n15653), .ZN(P2_U3035) );
  NAND2_X1 U18818 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n11600), .ZN(n15655) );
  OAI221_X1 U18819 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15658), 
        .C1(n15657), .C2(n15656), .A(n15655), .ZN(n15662) );
  AOI21_X1 U18820 ( .B1(n15659), .B2(n15660), .A(n9795), .ZN(n19134) );
  INV_X1 U18821 ( .A(n19134), .ZN(n19268) );
  OAI22_X1 U18822 ( .A1(n19268), .A2(n19400), .B1(n19404), .B2(n19132), .ZN(
        n15661) );
  AOI211_X1 U18823 ( .C1(n15663), .C2(n19395), .A(n15662), .B(n15661), .ZN(
        n15664) );
  OAI21_X1 U18824 ( .B1(n15665), .B2(n15702), .A(n15664), .ZN(P2_U3036) );
  INV_X1 U18825 ( .A(n9716), .ZN(n15668) );
  AOI21_X1 U18826 ( .B1(n15668), .B2(n15667), .A(n9781), .ZN(n16406) );
  INV_X1 U18827 ( .A(n16406), .ZN(n15682) );
  NOR2_X1 U18828 ( .A1(n15670), .A2(n15669), .ZN(n15671) );
  XNOR2_X1 U18829 ( .A(n15672), .B(n15671), .ZN(n16405) );
  OAI21_X1 U18830 ( .B1(n15673), .B2(n15674), .A(n15659), .ZN(n19271) );
  NAND2_X1 U18831 ( .A1(n15667), .A2(n15675), .ZN(n15677) );
  NAND2_X1 U18832 ( .A1(n15677), .A2(n15676), .ZN(n15679) );
  AOI22_X1 U18833 ( .A1(n16475), .A2(n19145), .B1(P2_REIP_REG_9__SCAN_IN), 
        .B2(n19180), .ZN(n15678) );
  OAI211_X1 U18834 ( .C1(n19271), .C2(n19400), .A(n15679), .B(n15678), .ZN(
        n15680) );
  AOI21_X1 U18835 ( .B1(n16405), .B2(n19395), .A(n15680), .ZN(n15681) );
  OAI21_X1 U18836 ( .B1(n15682), .B2(n15702), .A(n15681), .ZN(P2_U3037) );
  NOR2_X1 U18837 ( .A1(n19982), .A2(n19210), .ZN(n15683) );
  AOI221_X1 U18838 ( .B1(n16469), .B2(n11253), .C1(n16464), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15683), .ZN(n15684) );
  INV_X1 U18839 ( .A(n15684), .ZN(n15689) );
  OR2_X1 U18840 ( .A1(n15686), .A2(n15685), .ZN(n15687) );
  NAND2_X1 U18841 ( .A1(n15687), .A2(n16462), .ZN(n19274) );
  OAI22_X1 U18842 ( .A1(n19274), .A2(n19400), .B1(n19404), .B2(n19169), .ZN(
        n15688) );
  AOI211_X1 U18843 ( .C1(n15690), .C2(n19395), .A(n15689), .B(n15688), .ZN(
        n15691) );
  OAI21_X1 U18844 ( .B1(n15692), .B2(n15702), .A(n15691), .ZN(P2_U3039) );
  XNOR2_X1 U18845 ( .A(n15694), .B(n15693), .ZN(n19276) );
  AOI22_X1 U18846 ( .A1(n16475), .A2(n19184), .B1(n19180), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15697) );
  NAND2_X1 U18847 ( .A1(n15695), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15696) );
  OAI211_X1 U18848 ( .C1(n19276), .C2(n19400), .A(n15697), .B(n15696), .ZN(
        n15698) );
  AOI211_X1 U18849 ( .C1(n15700), .C2(n19395), .A(n15699), .B(n15698), .ZN(
        n15701) );
  OAI21_X1 U18850 ( .B1(n15703), .B2(n15702), .A(n15701), .ZN(P2_U3040) );
  INV_X1 U18851 ( .A(n15714), .ZN(n15724) );
  OAI22_X1 U18852 ( .A1(n19190), .A2(n20916), .B1(n19240), .B2(n19206), .ZN(
        n15708) );
  INV_X1 U18853 ( .A(n15718), .ZN(n20031) );
  OAI222_X1 U18854 ( .A1(n15724), .A2(n15705), .B1(n19950), .B2(n15708), .C1(
        n20031), .C2(n15704), .ZN(n15706) );
  MUX2_X1 U18855 ( .A(n15706), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15725), .Z(P2_U3601) );
  OAI21_X1 U18856 ( .B1(n19190), .B2(n20922), .A(n15707), .ZN(n15717) );
  INV_X1 U18857 ( .A(n15717), .ZN(n15710) );
  INV_X1 U18858 ( .A(n15708), .ZN(n15709) );
  NOR2_X1 U18859 ( .A1(n15709), .A2(n19950), .ZN(n15716) );
  AOI222_X1 U18860 ( .A1(n15711), .A2(n15718), .B1(n20053), .B2(n15714), .C1(
        n15710), .C2(n15716), .ZN(n15713) );
  NAND2_X1 U18861 ( .A1(n15725), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15712) );
  OAI21_X1 U18862 ( .B1(n15713), .B2(n15725), .A(n15712), .ZN(P2_U3600) );
  AOI222_X1 U18863 ( .A1(n15719), .A2(n15718), .B1(n15717), .B2(n15716), .C1(
        n15715), .C2(n15714), .ZN(n15722) );
  NAND2_X1 U18864 ( .A1(n15725), .A2(n15720), .ZN(n15721) );
  OAI21_X1 U18865 ( .B1(n15722), .B2(n15725), .A(n15721), .ZN(P2_U3599) );
  OAI22_X1 U18866 ( .A1(n19672), .A2(n15724), .B1(n15723), .B2(n20031), .ZN(
        n15726) );
  MUX2_X1 U18867 ( .A(n15726), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15725), .Z(P2_U3596) );
  INV_X1 U18868 ( .A(n19436), .ZN(n15738) );
  INV_X1 U18869 ( .A(n19887), .ZN(n15730) );
  INV_X1 U18870 ( .A(n19439), .ZN(n15735) );
  INV_X1 U18871 ( .A(n19927), .ZN(n19947) );
  AOI22_X1 U18872 ( .A1(n19896), .A2(n19465), .B1(n19432), .B2(n19886), .ZN(
        n15727) );
  OAI21_X1 U18873 ( .B1(n19899), .B2(n19947), .A(n15727), .ZN(n15728) );
  AOI21_X1 U18874 ( .B1(n15735), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n15728), .ZN(n15729) );
  OAI21_X1 U18875 ( .B1(n15738), .B2(n15730), .A(n15729), .ZN(P2_U3048) );
  NOR2_X2 U18876 ( .A1(n15731), .A2(n9715), .ZN(n19919) );
  INV_X1 U18877 ( .A(n19919), .ZN(n15737) );
  INV_X1 U18878 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n20975) );
  INV_X1 U18879 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16559) );
  AOI22_X1 U18880 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19435), .ZN(n19870) );
  INV_X1 U18881 ( .A(n19870), .ZN(n19920) );
  NOR2_X2 U18882 ( .A1(n15732), .A2(n19414), .ZN(n19918) );
  AOI22_X1 U18883 ( .A1(n19920), .A2(n19465), .B1(n19432), .B2(n19918), .ZN(
        n15733) );
  OAI21_X1 U18884 ( .B1(n19923), .B2(n19947), .A(n15733), .ZN(n15734) );
  AOI21_X1 U18885 ( .B1(n15735), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n15734), .ZN(n15736) );
  OAI21_X1 U18886 ( .B1(n15738), .B2(n15737), .A(n15736), .ZN(P2_U3052) );
  INV_X1 U18887 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16757) );
  INV_X1 U18888 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16788) );
  INV_X1 U18889 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17152) );
  INV_X1 U18890 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17154) );
  INV_X1 U18891 ( .A(n18768), .ZN(n15740) );
  INV_X1 U18892 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17218) );
  INV_X1 U18893 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16856) );
  INV_X1 U18894 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17267) );
  INV_X1 U18895 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17249) );
  INV_X1 U18896 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20977) );
  NAND2_X1 U18897 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17028) );
  NOR2_X1 U18898 ( .A1(n20977), .A2(n17028), .ZN(n17350) );
  NAND3_X1 U18899 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17350), .ZN(n17352) );
  NAND4_X1 U18900 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n15744) );
  NOR4_X1 U18901 ( .A1(n17267), .A2(n17249), .A3(n17352), .A4(n15744), .ZN(
        n15745) );
  NAND3_X1 U18902 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n15745), .ZN(n15837) );
  NAND2_X1 U18903 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .ZN(n17216) );
  NOR4_X1 U18904 ( .A1(n17218), .A2(n16856), .A3(n15837), .A4(n17216), .ZN(
        n17198) );
  NAND2_X1 U18905 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17198), .ZN(n17197) );
  NOR2_X1 U18906 ( .A1(n17365), .A2(n17197), .ZN(n17182) );
  NAND2_X1 U18907 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17182), .ZN(n17181) );
  NAND2_X1 U18908 ( .A1(n18361), .A2(n17169), .ZN(n17151) );
  NAND2_X1 U18909 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17136), .ZN(n17122) );
  NOR2_X1 U18910 ( .A1(n16788), .A2(n17122), .ZN(n17103) );
  NAND2_X1 U18911 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17103), .ZN(n17097) );
  NAND2_X1 U18912 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17096), .ZN(n17087) );
  INV_X1 U18913 ( .A(n17087), .ZN(n17092) );
  NAND2_X1 U18914 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17092), .ZN(n15824) );
  AND2_X1 U18915 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17049) );
  NOR2_X1 U18916 ( .A1(n17456), .A2(n17365), .ZN(n17349) );
  INV_X1 U18917 ( .A(n17349), .ZN(n17368) );
  NOR2_X2 U18918 ( .A1(n17365), .A2(n18361), .ZN(n17366) );
  NAND2_X1 U18919 ( .A1(n17355), .A2(n17087), .ZN(n15746) );
  OAI21_X1 U18920 ( .B1(n17049), .B2(n17368), .A(n15746), .ZN(n17082) );
  AOI22_X1 U18921 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15747) );
  OAI21_X1 U18922 ( .B1(n15789), .B2(n20925), .A(n15747), .ZN(n15756) );
  AOI22_X1 U18923 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15754) );
  OAI22_X1 U18924 ( .A1(n17300), .A2(n17123), .B1(n17263), .B2(n15826), .ZN(
        n15752) );
  AOI22_X1 U18925 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15750) );
  AOI22_X1 U18926 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15749) );
  AOI22_X1 U18927 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15748) );
  NAND3_X1 U18928 ( .A1(n15750), .A2(n15749), .A3(n15748), .ZN(n15751) );
  AOI211_X1 U18929 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15752), .B(n15751), .ZN(n15753) );
  OAI211_X1 U18930 ( .C1(n9771), .C2(n20824), .A(n15754), .B(n15753), .ZN(
        n15755) );
  AOI211_X1 U18931 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15756), .B(n15755), .ZN(n15822) );
  AOI22_X1 U18932 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15757) );
  OAI21_X1 U18933 ( .B1(n10288), .B2(n17157), .A(n15757), .ZN(n15766) );
  AOI22_X1 U18934 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15764) );
  OAI22_X1 U18935 ( .A1(n17275), .A2(n18656), .B1(n17334), .B2(n17283), .ZN(
        n15762) );
  AOI22_X1 U18936 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15760) );
  AOI22_X1 U18937 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15759) );
  AOI22_X1 U18938 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15758) );
  NAND3_X1 U18939 ( .A1(n15760), .A2(n15759), .A3(n15758), .ZN(n15761) );
  AOI211_X1 U18940 ( .C1(n17290), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n15762), .B(n15761), .ZN(n15763) );
  OAI211_X1 U18941 ( .C1(n9814), .C2(n17274), .A(n15764), .B(n15763), .ZN(
        n15765) );
  AOI211_X1 U18942 ( .C1(n10331), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n15766), .B(n15765), .ZN(n17089) );
  AOI22_X1 U18943 ( .A1(n17237), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15767) );
  OAI21_X1 U18944 ( .B1(n10253), .B2(n17186), .A(n15767), .ZN(n15776) );
  AOI22_X1 U18945 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15774) );
  AOI22_X1 U18946 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15768) );
  OAI21_X1 U18947 ( .B1(n17263), .B2(n17316), .A(n15768), .ZN(n15772) );
  AOI22_X1 U18948 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15770) );
  AOI22_X1 U18949 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15769) );
  OAI211_X1 U18950 ( .C1(n17275), .C2(n18650), .A(n15770), .B(n15769), .ZN(
        n15771) );
  AOI211_X1 U18951 ( .C1(n17202), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n15772), .B(n15771), .ZN(n15773) );
  OAI211_X1 U18952 ( .C1(n17204), .C2(n21085), .A(n15774), .B(n15773), .ZN(
        n15775) );
  AOI211_X1 U18953 ( .C1(n9734), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n15776), .B(n15775), .ZN(n17099) );
  AOI22_X1 U18954 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U18955 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10329), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U18956 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15777) );
  OAI211_X1 U18957 ( .C1(n17187), .C2(n17203), .A(n15778), .B(n15777), .ZN(
        n15784) );
  AOI22_X1 U18958 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U18959 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15781) );
  AOI22_X1 U18960 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15780) );
  NAND2_X1 U18961 ( .A1(n17313), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15779) );
  NAND4_X1 U18962 ( .A1(n15782), .A2(n15781), .A3(n15780), .A4(n15779), .ZN(
        n15783) );
  AOI211_X1 U18963 ( .C1(n17202), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n15784), .B(n15783), .ZN(n15785) );
  OAI211_X1 U18964 ( .C1(n17263), .C2(n15787), .A(n15786), .B(n15785), .ZN(
        n17105) );
  AOI22_X1 U18965 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10327), .B1(
        n10286), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15798) );
  AOI22_X1 U18966 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17290), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17326), .ZN(n15788) );
  OAI21_X1 U18967 ( .B1(n15789), .B2(n18765), .A(n15788), .ZN(n15796) );
  OAI22_X1 U18968 ( .A1(n9814), .A2(n18593), .B1(n17334), .B2(n18365), .ZN(
        n15790) );
  AOI21_X1 U18969 ( .B1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n15818), .A(
        n15790), .ZN(n15794) );
  AOI22_X1 U18970 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17237), .ZN(n15793) );
  AOI22_X1 U18971 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17306), .ZN(n15792) );
  AOI22_X1 U18972 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17202), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n10289), .ZN(n15791) );
  NAND4_X1 U18973 ( .A1(n15794), .A2(n15793), .A3(n15792), .A4(n15791), .ZN(
        n15795) );
  AOI211_X1 U18974 ( .C1(n9726), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n15796), .B(n15795), .ZN(n15797) );
  OAI211_X1 U18975 ( .C1(n18670), .C2(n10288), .A(n15798), .B(n15797), .ZN(
        n17106) );
  NAND2_X1 U18976 ( .A1(n17105), .A2(n17106), .ZN(n17104) );
  NOR2_X1 U18977 ( .A1(n17099), .A2(n17104), .ZN(n17098) );
  INV_X1 U18978 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15809) );
  AOI22_X1 U18979 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15808) );
  AOI22_X1 U18980 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15800) );
  AOI22_X1 U18981 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15799) );
  OAI211_X1 U18982 ( .C1(n10404), .C2(n17171), .A(n15800), .B(n15799), .ZN(
        n15806) );
  AOI22_X1 U18983 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15804) );
  AOI22_X1 U18984 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15803) );
  AOI22_X1 U18985 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15802) );
  NAND2_X1 U18986 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n15801) );
  NAND4_X1 U18987 ( .A1(n15804), .A2(n15803), .A3(n15802), .A4(n15801), .ZN(
        n15805) );
  AOI211_X1 U18988 ( .C1(n10286), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n15806), .B(n15805), .ZN(n15807) );
  OAI211_X1 U18989 ( .C1(n17263), .C2(n15809), .A(n15808), .B(n15807), .ZN(
        n17094) );
  NAND2_X1 U18990 ( .A1(n17098), .A2(n17094), .ZN(n17093) );
  NOR2_X1 U18991 ( .A1(n17089), .A2(n17093), .ZN(n17088) );
  AOI22_X1 U18992 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15821) );
  AOI22_X1 U18993 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15820) );
  OAI22_X1 U18994 ( .A1(n17263), .A2(n15810), .B1(n17325), .B2(n18739), .ZN(
        n15817) );
  OAI22_X1 U18995 ( .A1(n17275), .A2(n18659), .B1(n17334), .B2(n17141), .ZN(
        n15811) );
  AOI21_X1 U18996 ( .B1(n9734), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n15811), .ZN(n15815) );
  AOI22_X1 U18997 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15814) );
  AOI22_X1 U18998 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15813) );
  AOI22_X1 U18999 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15812) );
  NAND4_X1 U19000 ( .A1(n15815), .A2(n15814), .A3(n15813), .A4(n15812), .ZN(
        n15816) );
  AOI211_X1 U19001 ( .C1(n15818), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n15817), .B(n15816), .ZN(n15819) );
  NAND3_X1 U19002 ( .A1(n15821), .A2(n15820), .A3(n15819), .ZN(n17085) );
  NAND2_X1 U19003 ( .A1(n17088), .A2(n17085), .ZN(n17084) );
  NOR2_X1 U19004 ( .A1(n15822), .A2(n17084), .ZN(n17079) );
  AOI21_X1 U19005 ( .B1(n15822), .B2(n17084), .A(n17079), .ZN(n17387) );
  AOI22_X1 U19006 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17082), .B1(n17387), 
        .B2(n17366), .ZN(n15823) );
  OAI21_X1 U19007 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n15824), .A(n15823), .ZN(
        P3_U2675) );
  AOI22_X1 U19008 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15825) );
  OAI21_X1 U19009 ( .B1(n10288), .B2(n20824), .A(n15825), .ZN(n15836) );
  INV_X1 U19010 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15834) );
  AOI22_X1 U19011 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15833) );
  OAI22_X1 U19012 ( .A1(n9814), .A2(n15826), .B1(n10404), .B2(n20925), .ZN(
        n15831) );
  AOI22_X1 U19013 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15829) );
  AOI22_X1 U19014 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15828) );
  AOI22_X1 U19015 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15827) );
  NAND3_X1 U19016 ( .A1(n15829), .A2(n15828), .A3(n15827), .ZN(n15830) );
  AOI211_X1 U19017 ( .C1(n10327), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n15831), .B(n15830), .ZN(n15832) );
  OAI211_X1 U19018 ( .C1(n17204), .C2(n15834), .A(n15833), .B(n15832), .ZN(
        n15835) );
  AOI211_X1 U19019 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n15836), .B(n15835), .ZN(n17467) );
  INV_X1 U19020 ( .A(n15837), .ZN(n15838) );
  NAND2_X1 U19021 ( .A1(n17362), .A2(n15838), .ZN(n17215) );
  AND2_X1 U19022 ( .A1(n17355), .A2(n17215), .ZN(n17246) );
  NOR2_X1 U19023 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17368), .ZN(n17247) );
  AOI22_X1 U19024 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17246), .B1(n15838), 
        .B2(n17247), .ZN(n15839) );
  OAI21_X1 U19025 ( .B1(n17467), .B2(n17355), .A(n15839), .ZN(P3_U2690) );
  NAND2_X1 U19026 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18474) );
  AOI221_X1 U19027 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18474), .C1(n15841), 
        .C2(n18474), .A(n15840), .ZN(n18313) );
  NOR2_X1 U19028 ( .A1(n15842), .A2(n18809), .ZN(n15844) );
  OAI21_X1 U19029 ( .B1(n15844), .B2(n15843), .A(n18314), .ZN(n18311) );
  AOI22_X1 U19030 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18313), .B1(
        n18311), .B2(n18814), .ZN(P3_U2865) );
  INV_X1 U19031 ( .A(n18979), .ZN(n18971) );
  NOR2_X1 U19032 ( .A1(n16489), .A2(n18971), .ZN(n15849) );
  INV_X1 U19033 ( .A(n15845), .ZN(n15846) );
  NAND2_X1 U19034 ( .A1(n18324), .A2(n17580), .ZN(n18826) );
  AOI21_X1 U19035 ( .B1(n15849), .B2(n17522), .A(n15847), .ZN(n15851) );
  NAND3_X1 U19036 ( .A1(n15852), .A2(n15851), .A3(n15940), .ZN(n18802) );
  NOR2_X1 U19037 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21062), .ZN(n18318) );
  INV_X1 U19038 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18309) );
  NOR2_X1 U19039 ( .A1(n18309), .A2(n18926), .ZN(n15853) );
  INV_X1 U19040 ( .A(n18957), .ZN(n18955) );
  AOI21_X1 U19041 ( .B1(n15854), .B2(n18777), .A(n18789), .ZN(n18824) );
  NAND3_X1 U19042 ( .A1(n18955), .A2(n18987), .A3(n18824), .ZN(n15855) );
  OAI21_X1 U19043 ( .B1(n18955), .B2(n18777), .A(n15855), .ZN(P3_U3284) );
  INV_X1 U19044 ( .A(n16541), .ZN(n15859) );
  NAND2_X1 U19045 ( .A1(n15856), .A2(n17637), .ZN(n16542) );
  OAI21_X1 U19046 ( .B1(n18305), .B2(n16542), .A(n15857), .ZN(n15858) );
  AOI21_X1 U19047 ( .B1(n15859), .B2(n18212), .A(n15858), .ZN(n15924) );
  INV_X1 U19048 ( .A(n18199), .ZN(n18235) );
  NOR2_X1 U19049 ( .A1(n18778), .A2(n18780), .ZN(n18186) );
  INV_X1 U19050 ( .A(n18186), .ZN(n18193) );
  AOI21_X1 U19051 ( .B1(n18009), .B2(n18193), .A(n15860), .ZN(n16544) );
  AOI22_X1 U19052 ( .A1(n18287), .A2(n16505), .B1(n18212), .B2(n16525), .ZN(
        n15927) );
  OAI21_X1 U19053 ( .B1(n18235), .B2(n16544), .A(n15927), .ZN(n15861) );
  AOI21_X1 U19054 ( .B1(n18292), .B2(n17638), .A(n15861), .ZN(n15866) );
  NAND2_X1 U19055 ( .A1(n15863), .A2(n15862), .ZN(n15864) );
  XOR2_X1 U19056 ( .A(n15864), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16531) );
  AOI22_X1 U19057 ( .A1(n18301), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18203), 
        .B2(n16531), .ZN(n15865) );
  OAI221_X1 U19058 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15924), 
        .C1(n16528), .C2(n15866), .A(n15865), .ZN(P3_U2833) );
  OAI211_X1 U19059 ( .C1(n15869), .C2(n15868), .A(n19185), .B(n15867), .ZN(
        n15871) );
  AOI22_X1 U19060 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19236), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19222), .ZN(n15870) );
  NAND2_X1 U19061 ( .A1(n15871), .A2(n15870), .ZN(n15872) );
  AOI21_X1 U19062 ( .B1(n19223), .B2(P2_REIP_REG_22__SCAN_IN), .A(n15872), 
        .ZN(n15877) );
  OAI22_X1 U19063 ( .A1(n15874), .A2(n19200), .B1(n15873), .B2(n19228), .ZN(
        n15875) );
  INV_X1 U19064 ( .A(n15875), .ZN(n15876) );
  OAI211_X1 U19065 ( .C1(n15878), .C2(n19213), .A(n15877), .B(n15876), .ZN(
        P2_U2833) );
  NOR3_X1 U19066 ( .A1(n15880), .A2(n15879), .A3(n20449), .ZN(n15885) );
  OAI22_X1 U19067 ( .A1(n15882), .A2(n15881), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15885), .ZN(n15883) );
  INV_X1 U19068 ( .A(n15883), .ZN(n15884) );
  AOI21_X1 U19069 ( .B1(n15885), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15884), .ZN(n15887) );
  OAI222_X1 U19070 ( .A1(n20272), .A2(n15887), .B1(n20272), .B2(n15886), .C1(
        n15887), .C2(n15886), .ZN(n15888) );
  INV_X1 U19071 ( .A(n15888), .ZN(n15889) );
  AOI222_X1 U19072 ( .A1(n20273), .A2(n15890), .B1(n20273), .B2(n15889), .C1(
        n15890), .C2(n15889), .ZN(n15899) );
  INV_X1 U19073 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15892) );
  INV_X1 U19074 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20101) );
  AOI21_X1 U19075 ( .B1(n15892), .B2(n20101), .A(n15891), .ZN(n15894) );
  NOR4_X1 U19076 ( .A1(n15896), .A2(n15895), .A3(n15894), .A4(n15893), .ZN(
        n15897) );
  OAI211_X1 U19077 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15899), .A(
        n15898), .B(n15897), .ZN(n15904) );
  NAND3_X1 U19078 ( .A1(n15901), .A2(n15900), .A3(n20453), .ZN(n15902) );
  OAI221_X1 U19079 ( .B1(n15905), .B2(n20739), .C1(n15905), .C2(n15929), .A(
        n15902), .ZN(n16266) );
  AOI221_X1 U19080 ( .B1(n11886), .B2(n20661), .C1(n15904), .C2(n20661), .A(
        n16266), .ZN(n15906) );
  NOR2_X1 U19081 ( .A1(n15906), .A2(n11886), .ZN(n16272) );
  OAI21_X1 U19082 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20747), .A(n16272), 
        .ZN(n16270) );
  AOI211_X1 U19083 ( .C1(n15905), .C2(n15904), .A(n15903), .B(n16270), .ZN(
        n15911) );
  AOI21_X1 U19084 ( .B1(n15907), .B2(n16268), .A(n15906), .ZN(n15908) );
  INV_X1 U19085 ( .A(n15908), .ZN(n15909) );
  AOI22_X1 U19086 ( .A1(n15911), .A2(n15910), .B1(n11886), .B2(n15909), .ZN(
        P1_U3161) );
  NAND2_X1 U19087 ( .A1(n16206), .A2(n15912), .ZN(n16150) );
  NAND2_X1 U19088 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15913) );
  NOR3_X1 U19089 ( .A1(n16189), .A2(n16159), .A3(n15913), .ZN(n16154) );
  AOI22_X1 U19090 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16241), .B1(n16154), 
        .B2(n15917), .ZN(n15921) );
  NAND2_X1 U19091 ( .A1(n15914), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15915) );
  OAI21_X1 U19092 ( .B1(n15916), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15915), .ZN(n15918) );
  XNOR2_X1 U19093 ( .A(n15918), .B(n15917), .ZN(n16047) );
  INV_X1 U19094 ( .A(n15959), .ZN(n15919) );
  AOI22_X1 U19095 ( .A1(n16047), .A2(n16244), .B1(n16256), .B2(n15919), .ZN(
        n15920) );
  OAI211_X1 U19096 ( .C1(n15917), .C2(n16150), .A(n15921), .B(n15920), .ZN(
        P1_U3010) );
  INV_X1 U19097 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18916) );
  NOR2_X1 U19098 ( .A1(n18199), .A2(n18916), .ZN(n16508) );
  NOR3_X1 U19099 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15924), .A3(
        n16528), .ZN(n15925) );
  OAI221_X1 U19100 ( .B1(n16518), .B2(n15928), .C1(n16518), .C2(n15927), .A(
        n15926), .ZN(P3_U2832) );
  INV_X1 U19101 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20680) );
  INV_X1 U19102 ( .A(HOLD), .ZN(n20852) );
  NOR2_X1 U19103 ( .A1(n20680), .A2(n20852), .ZN(n20667) );
  AOI22_X1 U19104 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15931) );
  NAND2_X1 U19105 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15929), .ZN(n20678) );
  OAI211_X1 U19106 ( .C1(n20667), .C2(n15931), .A(n15930), .B(n20678), .ZN(
        P1_U3195) );
  NAND2_X1 U19107 ( .A1(n15932), .A2(n16486), .ZN(n15933) );
  AOI211_X1 U19108 ( .C1(n15935), .C2(n19770), .A(n15934), .B(n15933), .ZN(
        P2_U3178) );
  OAI221_X1 U19109 ( .B1(n19001), .B2(n16486), .C1(n15936), .C2(n16486), .A(
        n9715), .ZN(n20062) );
  NOR2_X1 U19110 ( .A1(n15937), .A2(n20062), .ZN(P2_U3047) );
  OAI22_X4 U19111 ( .A1(n18832), .A2(n15940), .B1(n15939), .B2(n15938), .ZN(
        n17369) );
  NAND2_X1 U19112 ( .A1(n18361), .A2(n17369), .ZN(n17515) );
  INV_X1 U19113 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17578) );
  NAND2_X2 U19114 ( .A1(n17456), .A2(n17369), .ZN(n17506) );
  AOI22_X1 U19115 ( .A1(n17514), .A2(BUF2_REG_0__SCAN_IN), .B1(n17513), .B2(
        n17993), .ZN(n15941) );
  OAI221_X1 U19116 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17515), .C1(n17578), 
        .C2(n17369), .A(n15941), .ZN(P3_U2735) );
  OR2_X1 U19117 ( .A1(n20152), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15956) );
  OAI21_X1 U19118 ( .B1(n15942), .B2(n15957), .A(n15996), .ZN(n15966) );
  AOI21_X1 U19119 ( .B1(n15956), .B2(n15966), .A(n14798), .ZN(n15948) );
  NAND3_X1 U19120 ( .A1(n16016), .A2(n14798), .A3(n15943), .ZN(n15946) );
  AOI22_X1 U19121 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20178), .B1(
        n20126), .B2(n15944), .ZN(n15945) );
  OAI211_X1 U19122 ( .C1(n14568), .C2(n20136), .A(n15946), .B(n15945), .ZN(
        n15947) );
  AOI211_X1 U19123 ( .C1(n15949), .C2(n20154), .A(n15948), .B(n15947), .ZN(
        n15950) );
  OAI21_X1 U19124 ( .B1(n20175), .B2(n16149), .A(n15950), .ZN(P1_U2818) );
  NOR2_X1 U19125 ( .A1(n15951), .A2(n15966), .ZN(n15954) );
  INV_X1 U19126 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15952) );
  NOR2_X1 U19127 ( .A1(n20162), .A2(n15952), .ZN(n15953) );
  AOI211_X1 U19128 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n20170), .A(n15954), .B(
        n15953), .ZN(n15955) );
  OAI21_X1 U19129 ( .B1(n15957), .B2(n15956), .A(n15955), .ZN(n15958) );
  INV_X1 U19130 ( .A(n15958), .ZN(n15962) );
  NOR2_X1 U19131 ( .A1(n15959), .A2(n20175), .ZN(n15960) );
  AOI21_X1 U19132 ( .B1(n16048), .B2(n20154), .A(n15960), .ZN(n15961) );
  OAI211_X1 U19133 ( .C1(n16051), .C2(n20186), .A(n15962), .B(n15961), .ZN(
        P1_U2819) );
  AOI22_X1 U19134 ( .A1(n20170), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n20126), 
        .B2(n16052), .ZN(n15970) );
  INV_X1 U19135 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21063) );
  INV_X1 U19136 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20705) );
  NOR2_X1 U19137 ( .A1(n21063), .A2(n20705), .ZN(n15972) );
  INV_X1 U19138 ( .A(n15963), .ZN(n15964) );
  NOR2_X1 U19139 ( .A1(n20152), .A2(n15964), .ZN(n15985) );
  AOI21_X1 U19140 ( .B1(n15972), .B2(n15985), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15967) );
  OAI22_X1 U19141 ( .A1(n15967), .A2(n15966), .B1(n15965), .B2(n20175), .ZN(
        n15968) );
  AOI21_X1 U19142 ( .B1(n16053), .B2(n20154), .A(n15968), .ZN(n15969) );
  OAI211_X1 U19143 ( .C1(n15971), .C2(n20162), .A(n15970), .B(n15969), .ZN(
        P1_U2820) );
  AOI21_X1 U19144 ( .B1(n21063), .B2(n20705), .A(n15972), .ZN(n15973) );
  AOI22_X1 U19145 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n15986), .B1(n15985), 
        .B2(n15973), .ZN(n15974) );
  INV_X1 U19146 ( .A(n15974), .ZN(n15979) );
  INV_X1 U19147 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15977) );
  INV_X1 U19148 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15975) );
  OR2_X1 U19149 ( .A1(n20136), .A2(n15975), .ZN(n15976) );
  OAI211_X1 U19150 ( .C1(n15977), .C2(n20162), .A(n15976), .B(n9736), .ZN(
        n15978) );
  NOR2_X1 U19151 ( .A1(n15979), .A2(n15978), .ZN(n15981) );
  AOI22_X1 U19152 ( .A1(n16059), .A2(n20154), .B1(n20159), .B2(n16157), .ZN(
        n15980) );
  OAI211_X1 U19153 ( .C1(n16062), .C2(n20186), .A(n15981), .B(n15980), .ZN(
        P1_U2821) );
  AOI21_X1 U19154 ( .B1(n20178), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20177), .ZN(n15982) );
  OAI21_X1 U19155 ( .B1(n15983), .B2(n20136), .A(n15982), .ZN(n15984) );
  AOI221_X1 U19156 ( .B1(n15986), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n15985), 
        .C2(n21063), .A(n15984), .ZN(n15991) );
  NOR2_X1 U19157 ( .A1(n15987), .A2(n20186), .ZN(n15988) );
  AOI21_X1 U19158 ( .B1(n15989), .B2(n20154), .A(n15988), .ZN(n15990) );
  OAI211_X1 U19159 ( .C1(n20175), .C2(n16168), .A(n15991), .B(n15990), .ZN(
        P1_U2822) );
  INV_X1 U19160 ( .A(n15992), .ZN(n15993) );
  NAND2_X1 U19161 ( .A1(n15994), .A2(n15993), .ZN(n15995) );
  NAND2_X1 U19162 ( .A1(n15996), .A2(n15995), .ZN(n16024) );
  OAI211_X1 U19163 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n16008), .B(n15997), .ZN(n15998) );
  OAI211_X1 U19164 ( .C1(n15999), .C2(n20136), .A(n15998), .B(n9736), .ZN(
        n16004) );
  INV_X1 U19165 ( .A(n16000), .ZN(n16002) );
  OAI22_X1 U19166 ( .A1(n16002), .A2(n20141), .B1(n20175), .B2(n16001), .ZN(
        n16003) );
  AOI211_X1 U19167 ( .C1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n20178), .A(
        n16004), .B(n16003), .ZN(n16007) );
  NAND2_X1 U19168 ( .A1(n16005), .A2(n20126), .ZN(n16006) );
  OAI211_X1 U19169 ( .C1(n14815), .C2(n16024), .A(n16007), .B(n16006), .ZN(
        P1_U2824) );
  INV_X1 U19170 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20699) );
  AOI22_X1 U19171 ( .A1(n16081), .A2(n20126), .B1(n16008), .B2(n20699), .ZN(
        n16014) );
  INV_X1 U19172 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16009) );
  OAI21_X1 U19173 ( .B1(n20162), .B2(n16009), .A(n9736), .ZN(n16011) );
  NOR2_X1 U19174 ( .A1(n16024), .A2(n20699), .ZN(n16010) );
  AOI211_X1 U19175 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n20170), .A(n16011), .B(
        n16010), .ZN(n16013) );
  AOI22_X1 U19176 ( .A1(n16082), .A2(n20154), .B1(n20159), .B2(n16183), .ZN(
        n16012) );
  NAND3_X1 U19177 ( .A1(n16014), .A2(n16013), .A3(n16012), .ZN(P1_U2825) );
  AOI21_X1 U19178 ( .B1(n16016), .B2(n16015), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n16025) );
  OAI22_X1 U19179 ( .A1(n16018), .A2(n20175), .B1(n16017), .B2(n20136), .ZN(
        n16019) );
  AOI211_X1 U19180 ( .C1(n20178), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20177), .B(n16019), .ZN(n16023) );
  AOI22_X1 U19181 ( .A1(n16021), .A2(n20154), .B1(n16020), .B2(n20126), .ZN(
        n16022) );
  OAI211_X1 U19182 ( .C1(n16025), .C2(n16024), .A(n16023), .B(n16022), .ZN(
        P1_U2826) );
  INV_X1 U19183 ( .A(n16026), .ZN(n16027) );
  NOR2_X1 U19184 ( .A1(n20152), .A2(n16027), .ZN(n16036) );
  AOI21_X1 U19185 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16036), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16034) );
  OAI21_X1 U19186 ( .B1(n20162), .B2(n16028), .A(n9736), .ZN(n16031) );
  NOR2_X1 U19187 ( .A1(n16029), .A2(n20175), .ZN(n16030) );
  AOI211_X1 U19188 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n20170), .A(n16031), .B(
        n16030), .ZN(n16033) );
  AOI22_X1 U19189 ( .A1(n16086), .A2(n20126), .B1(n20154), .B2(n16085), .ZN(
        n16032) );
  OAI211_X1 U19190 ( .C1(n16035), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        P1_U2828) );
  INV_X1 U19191 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20694) );
  AOI22_X1 U19192 ( .A1(n20159), .A2(n16197), .B1(n16036), .B2(n20694), .ZN(
        n16042) );
  INV_X1 U19193 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16039) );
  AOI22_X1 U19194 ( .A1(n16037), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20170), 
        .B2(P1_EBX_REG_11__SCAN_IN), .ZN(n16038) );
  OAI211_X1 U19195 ( .C1(n20162), .C2(n16039), .A(n16038), .B(n9736), .ZN(
        n16040) );
  AOI21_X1 U19196 ( .B1(n20154), .B2(n16094), .A(n16040), .ZN(n16041) );
  OAI211_X1 U19197 ( .C1(n16097), .C2(n20186), .A(n16042), .B(n16041), .ZN(
        P1_U2829) );
  AOI22_X1 U19198 ( .A1(n16085), .A2(n16044), .B1(n20239), .B2(n16043), .ZN(
        n16045) );
  OAI21_X1 U19199 ( .B1(n16046), .B2(n13952), .A(n16045), .ZN(P1_U2892) );
  AOI22_X1 U19200 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16050) );
  AOI22_X1 U19201 ( .A1(n16048), .A2(n16069), .B1(n16116), .B2(n16047), .ZN(
        n16049) );
  OAI211_X1 U19202 ( .C1(n16111), .C2(n16051), .A(n16050), .B(n16049), .ZN(
        P1_U2978) );
  AOI22_X1 U19203 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n16055) );
  AOI22_X1 U19204 ( .A1(n16053), .A2(n16069), .B1(n16114), .B2(n16052), .ZN(
        n16054) );
  OAI211_X1 U19205 ( .C1(n16056), .C2(n20100), .A(n16055), .B(n16054), .ZN(
        P1_U2979) );
  AOI22_X1 U19206 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16061) );
  NOR2_X1 U19207 ( .A1(n16090), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16057) );
  MUX2_X1 U19208 ( .A(n16090), .B(n16057), .S(n14807), .Z(n16058) );
  XNOR2_X1 U19209 ( .A(n16058), .B(n16160), .ZN(n16158) );
  AOI22_X1 U19210 ( .A1(n16059), .A2(n16069), .B1(n16116), .B2(n16158), .ZN(
        n16060) );
  OAI211_X1 U19211 ( .C1(n16111), .C2(n16062), .A(n16061), .B(n16060), .ZN(
        P1_U2980) );
  NOR2_X1 U19212 ( .A1(n16090), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16066) );
  NAND2_X1 U19213 ( .A1(n16064), .A2(n16063), .ZN(n16065) );
  MUX2_X1 U19214 ( .A(n16066), .B(n16090), .S(n16065), .Z(n16067) );
  XNOR2_X1 U19215 ( .A(n16067), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16182) );
  AOI22_X1 U19216 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16072) );
  AOI22_X1 U19217 ( .A1(n16070), .A2(n16069), .B1(n16114), .B2(n16068), .ZN(
        n16071) );
  OAI211_X1 U19218 ( .C1(n20100), .C2(n16182), .A(n16072), .B(n16071), .ZN(
        P1_U2982) );
  INV_X1 U19219 ( .A(n16073), .ZN(n16075) );
  NAND2_X1 U19220 ( .A1(n16075), .A2(n16074), .ZN(n16080) );
  NAND3_X1 U19221 ( .A1(n16078), .A2(n16077), .A3(n16076), .ZN(n16079) );
  XOR2_X1 U19222 ( .A(n16080), .B(n16079), .Z(n16188) );
  AOI22_X1 U19223 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16084) );
  AOI22_X1 U19224 ( .A1(n16082), .A2(n16069), .B1(n16081), .B2(n16114), .ZN(
        n16083) );
  OAI211_X1 U19225 ( .C1(n16188), .C2(n20100), .A(n16084), .B(n16083), .ZN(
        P1_U2984) );
  AOI22_X1 U19226 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16088) );
  AOI22_X1 U19227 ( .A1(n16114), .A2(n16086), .B1(n16069), .B2(n16085), .ZN(
        n16087) );
  OAI211_X1 U19228 ( .C1(n16089), .C2(n20100), .A(n16088), .B(n16087), .ZN(
        P1_U2987) );
  AOI22_X1 U19229 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16096) );
  NAND3_X1 U19230 ( .A1(n12073), .A2(n16090), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16092) );
  NAND2_X1 U19231 ( .A1(n16092), .A2(n16091), .ZN(n16093) );
  XOR2_X1 U19232 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16093), .Z(
        n16199) );
  AOI22_X1 U19233 ( .A1(n16116), .A2(n16199), .B1(n16069), .B2(n16094), .ZN(
        n16095) );
  OAI211_X1 U19234 ( .C1(n16111), .C2(n16097), .A(n16096), .B(n16095), .ZN(
        P1_U2988) );
  AOI22_X1 U19235 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16103) );
  XNOR2_X1 U19236 ( .A(n16098), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16099) );
  XNOR2_X1 U19237 ( .A(n16100), .B(n16099), .ZN(n16233) );
  INV_X1 U19238 ( .A(n20195), .ZN(n16101) );
  AOI22_X1 U19239 ( .A1(n16233), .A2(n16116), .B1(n16069), .B2(n16101), .ZN(
        n16102) );
  OAI211_X1 U19240 ( .C1(n16111), .C2(n20145), .A(n16103), .B(n16102), .ZN(
        P1_U2992) );
  AOI22_X1 U19241 ( .A1(n16104), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16241), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16110) );
  NAND2_X1 U19242 ( .A1(n16106), .A2(n16105), .ZN(n16107) );
  XNOR2_X1 U19243 ( .A(n16108), .B(n16107), .ZN(n16243) );
  AOI22_X1 U19244 ( .A1(n16243), .A2(n16116), .B1(n16069), .B2(n20155), .ZN(
        n16109) );
  OAI211_X1 U19245 ( .C1(n16111), .C2(n20158), .A(n16110), .B(n16109), .ZN(
        P1_U2993) );
  INV_X1 U19246 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20161) );
  XNOR2_X1 U19247 ( .A(n16113), .B(n16112), .ZN(n16260) );
  INV_X1 U19248 ( .A(n16260), .ZN(n16117) );
  INV_X1 U19249 ( .A(n20168), .ZN(n16115) );
  AOI222_X1 U19250 ( .A1(n16117), .A2(n16116), .B1(n16115), .B2(n16114), .C1(
        n16069), .C2(n20201), .ZN(n16119) );
  AND2_X1 U19251 ( .A1(n20177), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16255) );
  INV_X1 U19252 ( .A(n16255), .ZN(n16118) );
  OAI211_X1 U19253 ( .C1(n20161), .C2(n16120), .A(n16119), .B(n16118), .ZN(
        P1_U2994) );
  OAI21_X1 U19254 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16129), .ZN(n16127) );
  INV_X1 U19255 ( .A(n16137), .ZN(n16124) );
  INV_X1 U19256 ( .A(n16121), .ZN(n16123) );
  AOI222_X1 U19257 ( .A1(n16124), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .B1(n16256), .B2(n16123), .C1(n16244), .C2(n9739), .ZN(n16126) );
  NAND2_X1 U19258 ( .A1(n16241), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16125) );
  OAI211_X1 U19259 ( .C1(n16128), .C2(n16127), .A(n16126), .B(n16125), .ZN(
        P1_U3005) );
  AOI22_X1 U19260 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n16241), .B1(n16129), 
        .B2(n16136), .ZN(n16135) );
  INV_X1 U19261 ( .A(n16130), .ZN(n16133) );
  INV_X1 U19262 ( .A(n16131), .ZN(n16132) );
  AOI22_X1 U19263 ( .A1(n16133), .A2(n16244), .B1(n16256), .B2(n16132), .ZN(
        n16134) );
  OAI211_X1 U19264 ( .C1(n16137), .C2(n16136), .A(n16135), .B(n16134), .ZN(
        P1_U3006) );
  AND2_X1 U19265 ( .A1(n16138), .A2(n16148), .ZN(n16139) );
  AOI22_X1 U19266 ( .A1(n16241), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n16140), 
        .B2(n16139), .ZN(n16146) );
  INV_X1 U19267 ( .A(n16141), .ZN(n16144) );
  INV_X1 U19268 ( .A(n16142), .ZN(n16143) );
  AOI22_X1 U19269 ( .A1(n16144), .A2(n16244), .B1(n16256), .B2(n16143), .ZN(
        n16145) );
  OAI211_X1 U19270 ( .C1(n16148), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        P1_U3008) );
  OAI22_X1 U19271 ( .A1(n16150), .A2(n12249), .B1(n16220), .B2(n16149), .ZN(
        n16151) );
  AOI21_X1 U19272 ( .B1(n16244), .B2(n16152), .A(n16151), .ZN(n16156) );
  OAI211_X1 U19273 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(n16154), .B(n16153), .ZN(
        n16155) );
  OAI211_X1 U19274 ( .C1(n14798), .C2(n9736), .A(n16156), .B(n16155), .ZN(
        P1_U3009) );
  AOI22_X1 U19275 ( .A1(n16158), .A2(n16244), .B1(n16256), .B2(n16157), .ZN(
        n16163) );
  NOR2_X1 U19276 ( .A1(n16189), .A2(n16159), .ZN(n16161) );
  AOI22_X1 U19277 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n9883), .B1(
        n16161), .B2(n16160), .ZN(n16162) );
  OAI211_X1 U19278 ( .C1(n20705), .C2(n9736), .A(n16163), .B(n16162), .ZN(
        P1_U3012) );
  NAND2_X1 U19279 ( .A1(n16166), .A2(n16164), .ZN(n16173) );
  OAI21_X1 U19280 ( .B1(n16167), .B2(n16166), .A(n16165), .ZN(n16178) );
  OAI22_X1 U19281 ( .A1(n16169), .A2(n16259), .B1(n16220), .B2(n16168), .ZN(
        n16170) );
  AOI21_X1 U19282 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16178), .A(
        n16170), .ZN(n16172) );
  NAND2_X1 U19283 ( .A1(n16241), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16171) );
  OAI211_X1 U19284 ( .C1(n16174), .C2(n16173), .A(n16172), .B(n16171), .ZN(
        P1_U3013) );
  NAND2_X1 U19285 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16175) );
  OAI21_X1 U19286 ( .B1(n16175), .B2(n16174), .A(n12078), .ZN(n16179) );
  INV_X1 U19287 ( .A(n16176), .ZN(n16177) );
  AOI22_X1 U19288 ( .A1(n16179), .A2(n16178), .B1(n16256), .B2(n16177), .ZN(
        n16181) );
  NAND2_X1 U19289 ( .A1(n16241), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16180) );
  OAI211_X1 U19290 ( .C1(n16182), .C2(n16259), .A(n16181), .B(n16180), .ZN(
        P1_U3014) );
  AOI22_X1 U19291 ( .A1(n16183), .A2(n16256), .B1(n16241), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n16187) );
  AOI21_X1 U19292 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16185), .A(
        n16184), .ZN(n16186) );
  OAI211_X1 U19293 ( .C1(n16188), .C2(n16259), .A(n16187), .B(n16186), .ZN(
        P1_U3016) );
  OAI22_X1 U19294 ( .A1(n20697), .A2(n9736), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16189), .ZN(n16190) );
  INV_X1 U19295 ( .A(n16190), .ZN(n16194) );
  AOI22_X1 U19296 ( .A1(n16192), .A2(n16244), .B1(n16256), .B2(n16191), .ZN(
        n16193) );
  OAI211_X1 U19297 ( .C1(n16196), .C2(n16195), .A(n16194), .B(n16193), .ZN(
        P1_U3018) );
  AOI22_X1 U19298 ( .A1(n16197), .A2(n16256), .B1(n16241), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16201) );
  AOI22_X1 U19299 ( .A1(n16244), .A2(n16199), .B1(n16198), .B2(n16250), .ZN(
        n16200) );
  OAI211_X1 U19300 ( .C1(n16203), .C2(n16202), .A(n16201), .B(n16200), .ZN(
        P1_U3020) );
  NAND2_X1 U19301 ( .A1(n16205), .A2(n16204), .ZN(n16207) );
  OAI21_X1 U19302 ( .B1(n16208), .B2(n16207), .A(n16206), .ZN(n16227) );
  OAI22_X1 U19303 ( .A1(n16209), .A2(n16220), .B1(n20835), .B2(n9736), .ZN(
        n16210) );
  AOI21_X1 U19304 ( .B1(n16244), .B2(n16211), .A(n16210), .ZN(n16215) );
  NOR2_X1 U19305 ( .A1(n16213), .A2(n16212), .ZN(n16223) );
  OAI221_X1 U19306 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14837), .C2(n16228), .A(
        n16223), .ZN(n16214) );
  OAI211_X1 U19307 ( .C1(n14837), .C2(n16227), .A(n16215), .B(n16214), .ZN(
        P1_U3021) );
  NAND2_X1 U19308 ( .A1(n16217), .A2(n16216), .ZN(n16218) );
  NAND2_X1 U19309 ( .A1(n16219), .A2(n16218), .ZN(n20188) );
  OR2_X1 U19310 ( .A1(n20188), .A2(n16220), .ZN(n16222) );
  AND2_X1 U19311 ( .A1(n16222), .A2(n16221), .ZN(n16226) );
  AOI22_X1 U19312 ( .A1(n16224), .A2(n16244), .B1(n16223), .B2(n16228), .ZN(
        n16225) );
  OAI211_X1 U19313 ( .C1(n16228), .C2(n16227), .A(n16226), .B(n16225), .ZN(
        P1_U3022) );
  INV_X1 U19314 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16237) );
  AOI21_X1 U19315 ( .B1(n10063), .B2(n16230), .A(n16229), .ZN(n16232) );
  OR2_X1 U19316 ( .A1(n16232), .A2(n16231), .ZN(n20193) );
  INV_X1 U19317 ( .A(n20193), .ZN(n20134) );
  AOI22_X1 U19318 ( .A1(n20134), .A2(n16256), .B1(n16241), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16236) );
  AOI22_X1 U19319 ( .A1(n16234), .A2(n16237), .B1(n16244), .B2(n16233), .ZN(
        n16235) );
  OAI211_X1 U19320 ( .C1(n16238), .C2(n16237), .A(n16236), .B(n16235), .ZN(
        P1_U3024) );
  NAND2_X1 U19321 ( .A1(n16239), .A2(n16250), .ZN(n16247) );
  INV_X1 U19322 ( .A(n16240), .ZN(n20146) );
  AOI22_X1 U19323 ( .A1(n20146), .A2(n16256), .B1(n16241), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16246) );
  AOI22_X1 U19324 ( .A1(n16244), .A2(n16243), .B1(n16242), .B2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16245) );
  OAI211_X1 U19325 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16247), .A(
        n16246), .B(n16245), .ZN(P1_U3025) );
  INV_X1 U19326 ( .A(n16248), .ZN(n16249) );
  NAND2_X1 U19327 ( .A1(n16250), .A2(n16249), .ZN(n16258) );
  NAND2_X1 U19328 ( .A1(n16252), .A2(n16251), .ZN(n16253) );
  AND2_X1 U19329 ( .A1(n16254), .A2(n16253), .ZN(n20198) );
  AOI21_X1 U19330 ( .B1(n20198), .B2(n16256), .A(n16255), .ZN(n16257) );
  OAI211_X1 U19331 ( .C1(n16260), .C2(n16259), .A(n16258), .B(n16257), .ZN(
        n16261) );
  INV_X1 U19332 ( .A(n16261), .ZN(n16262) );
  OAI21_X1 U19333 ( .B1(n16263), .B2(n12040), .A(n16262), .ZN(P1_U3026) );
  NAND4_X1 U19334 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n12842), .A4(n20747), .ZN(n16264) );
  AND2_X1 U19335 ( .A1(n16265), .A2(n16264), .ZN(n20662) );
  INV_X1 U19336 ( .A(n16266), .ZN(n16267) );
  AOI21_X1 U19337 ( .B1(n20662), .B2(n16271), .A(n16267), .ZN(n16269) );
  AOI211_X1 U19338 ( .C1(n20661), .C2(n16270), .A(n16269), .B(n16268), .ZN(
        P1_U3162) );
  OAI22_X1 U19339 ( .A1(n16272), .A2(n20554), .B1(n11886), .B2(n16271), .ZN(
        P1_U3466) );
  NAND2_X1 U19340 ( .A1(n19185), .A2(n19190), .ZN(n19239) );
  NAND2_X1 U19341 ( .A1(n19190), .A2(n16273), .ZN(n16289) );
  NAND2_X1 U19342 ( .A1(n16290), .A2(n16289), .ZN(n16288) );
  AOI22_X1 U19343 ( .A1(n19222), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19236), .ZN(n16275) );
  OAI21_X1 U19344 ( .B1(n16276), .B2(n19178), .A(n16275), .ZN(n16277) );
  AOI21_X1 U19345 ( .B1(n16278), .B2(n19194), .A(n16277), .ZN(n16279) );
  OAI21_X1 U19346 ( .B1(n19239), .B2(n16288), .A(n16283), .ZN(P2_U2824) );
  AOI22_X1 U19347 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19222), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19223), .ZN(n16294) );
  AOI22_X1 U19348 ( .A1(n16284), .A2(n19194), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19236), .ZN(n16293) );
  INV_X1 U19349 ( .A(n16285), .ZN(n16286) );
  AOI22_X1 U19350 ( .A1(n16287), .A2(n16282), .B1(n19224), .B2(n16286), .ZN(
        n16292) );
  OAI211_X1 U19351 ( .C1(n16290), .C2(n16289), .A(n19185), .B(n16288), .ZN(
        n16291) );
  NAND4_X1 U19352 ( .A1(n16294), .A2(n16293), .A3(n16292), .A4(n16291), .ZN(
        P2_U2825) );
  AOI22_X1 U19353 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19223), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19222), .ZN(n16305) );
  AOI22_X1 U19354 ( .A1(n16295), .A2(n19194), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19236), .ZN(n16304) );
  OAI22_X1 U19355 ( .A1(n16297), .A2(n19200), .B1(n16296), .B2(n19213), .ZN(
        n16298) );
  INV_X1 U19356 ( .A(n16298), .ZN(n16303) );
  OAI211_X1 U19357 ( .C1(n16301), .C2(n16300), .A(n19185), .B(n16299), .ZN(
        n16302) );
  NAND4_X1 U19358 ( .A1(n16305), .A2(n16304), .A3(n16303), .A4(n16302), .ZN(
        P2_U2827) );
  OAI22_X1 U19359 ( .A1(n19197), .A2(n16307), .B1(n19174), .B2(n16306), .ZN(
        n16308) );
  AOI21_X1 U19360 ( .B1(P2_REIP_REG_27__SCAN_IN), .B2(n19223), .A(n16308), 
        .ZN(n16309) );
  OAI21_X1 U19361 ( .B1(n16310), .B2(n19228), .A(n16309), .ZN(n16311) );
  AOI21_X1 U19362 ( .B1(n16312), .B2(n16282), .A(n16311), .ZN(n16317) );
  OAI211_X1 U19363 ( .C1(n16315), .C2(n16314), .A(n19185), .B(n16313), .ZN(
        n16316) );
  OAI211_X1 U19364 ( .C1(n19213), .C2(n16318), .A(n16317), .B(n16316), .ZN(
        P2_U2828) );
  INV_X1 U19365 ( .A(n16319), .ZN(n16324) );
  OAI22_X1 U19366 ( .A1(n19197), .A2(n11115), .B1(n19174), .B2(n10093), .ZN(
        n16320) );
  AOI21_X1 U19367 ( .B1(n19223), .B2(P2_REIP_REG_24__SCAN_IN), .A(n16320), 
        .ZN(n16321) );
  OAI21_X1 U19368 ( .B1(n16322), .B2(n19228), .A(n16321), .ZN(n16323) );
  AOI21_X1 U19369 ( .B1(n16324), .B2(n16282), .A(n16323), .ZN(n16329) );
  OAI211_X1 U19370 ( .C1(n16327), .C2(n16326), .A(n19185), .B(n16325), .ZN(
        n16328) );
  OAI211_X1 U19371 ( .C1(n19213), .C2(n16330), .A(n16329), .B(n16328), .ZN(
        P2_U2831) );
  AOI22_X1 U19372 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19223), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19222), .ZN(n16341) );
  AOI22_X1 U19373 ( .A1(n16331), .A2(n19194), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19236), .ZN(n16340) );
  INV_X1 U19374 ( .A(n16332), .ZN(n16333) );
  OAI22_X1 U19375 ( .A1(n16357), .A2(n19200), .B1(n16333), .B2(n19213), .ZN(
        n16334) );
  INV_X1 U19376 ( .A(n16334), .ZN(n16339) );
  OAI211_X1 U19377 ( .C1(n16337), .C2(n16336), .A(n19185), .B(n16335), .ZN(
        n16338) );
  NAND4_X1 U19378 ( .A1(n16341), .A2(n16340), .A3(n16339), .A4(n16338), .ZN(
        P2_U2832) );
  AOI22_X1 U19379 ( .A1(n19246), .A2(n16342), .B1(n19294), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16346) );
  AOI22_X1 U19380 ( .A1(n19248), .A2(BUF2_REG_20__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16345) );
  AOI22_X1 U19381 ( .A1(n10220), .A2(n19295), .B1(n19280), .B2(n16343), .ZN(
        n16344) );
  NAND3_X1 U19382 ( .A1(n16346), .A2(n16345), .A3(n16344), .ZN(P2_U2899) );
  AOI22_X1 U19383 ( .A1(n19246), .A2(n16347), .B1(n19294), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16353) );
  AOI22_X1 U19384 ( .A1(n19248), .A2(BUF2_REG_18__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16352) );
  OAI22_X1 U19385 ( .A1(n16349), .A2(n19052), .B1(n16348), .B2(n19299), .ZN(
        n16350) );
  INV_X1 U19386 ( .A(n16350), .ZN(n16351) );
  NAND3_X1 U19387 ( .A1(n16353), .A2(n16352), .A3(n16351), .ZN(P2_U2901) );
  AOI22_X1 U19388 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n11600), .B1(n16434), 
        .B2(n16354), .ZN(n16361) );
  NAND3_X1 U19389 ( .A1(n16355), .A2(n15494), .A3(n16441), .ZN(n16356) );
  OAI21_X1 U19390 ( .B1(n16439), .B2(n16357), .A(n16356), .ZN(n16358) );
  AOI21_X1 U19391 ( .B1(n16359), .B2(n16435), .A(n16358), .ZN(n16360) );
  OAI211_X1 U19392 ( .C1(n16362), .C2(n16445), .A(n16361), .B(n16360), .ZN(
        P2_U2991) );
  AOI22_X1 U19393 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16409), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19180), .ZN(n16368) );
  OAI22_X1 U19394 ( .A1(n16364), .A2(n16425), .B1(n16427), .B2(n16363), .ZN(
        n16365) );
  AOI21_X1 U19395 ( .B1(n16421), .B2(n16366), .A(n16365), .ZN(n16367) );
  OAI211_X1 U19396 ( .C1(n16424), .C2(n19045), .A(n16368), .B(n16367), .ZN(
        P2_U2996) );
  AOI22_X1 U19397 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n11600), .B1(n16434), 
        .B2(n19084), .ZN(n16374) );
  INV_X1 U19398 ( .A(n19085), .ZN(n16371) );
  INV_X1 U19399 ( .A(n16369), .ZN(n16370) );
  AOI222_X1 U19400 ( .A1(n16372), .A2(n16441), .B1(n16421), .B2(n16371), .C1(
        n16435), .C2(n16370), .ZN(n16373) );
  OAI211_X1 U19401 ( .C1(n19090), .C2(n16445), .A(n16374), .B(n16373), .ZN(
        P2_U2999) );
  AOI22_X1 U19402 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19180), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16409), .ZN(n16387) );
  AOI21_X1 U19403 ( .B1(n16377), .B2(n16376), .A(n16375), .ZN(n16455) );
  INV_X1 U19404 ( .A(n16378), .ZN(n16383) );
  AOI21_X1 U19405 ( .B1(n16380), .B2(n16382), .A(n16379), .ZN(n16381) );
  AOI21_X1 U19406 ( .B1(n16383), .B2(n16382), .A(n16381), .ZN(n16454) );
  AOI22_X1 U19407 ( .A1(n16455), .A2(n16435), .B1(n16441), .B2(n16454), .ZN(
        n16384) );
  INV_X1 U19408 ( .A(n16384), .ZN(n16385) );
  AOI21_X1 U19409 ( .B1(n16421), .B2(n19097), .A(n16385), .ZN(n16386) );
  OAI211_X1 U19410 ( .C1(n16424), .C2(n19092), .A(n16387), .B(n16386), .ZN(
        P2_U3000) );
  AOI22_X1 U19411 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n11600), .B1(n16434), 
        .B2(n19108), .ZN(n16393) );
  INV_X1 U19412 ( .A(n16388), .ZN(n16391) );
  INV_X1 U19413 ( .A(n16389), .ZN(n19109) );
  AOI222_X1 U19414 ( .A1(n16391), .A2(n16435), .B1(n16441), .B2(n16390), .C1(
        n16421), .C2(n19109), .ZN(n16392) );
  OAI211_X1 U19415 ( .C1(n19102), .C2(n16445), .A(n16393), .B(n16392), .ZN(
        P2_U3001) );
  AOI22_X1 U19416 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n11600), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16409), .ZN(n16399) );
  OAI22_X1 U19417 ( .A1(n16395), .A2(n16427), .B1(n16394), .B2(n16425), .ZN(
        n16396) );
  AOI21_X1 U19418 ( .B1(n16421), .B2(n16397), .A(n16396), .ZN(n16398) );
  OAI211_X1 U19419 ( .C1(n16424), .C2(n16400), .A(n16399), .B(n16398), .ZN(
        P2_U3002) );
  AOI22_X1 U19420 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n11600), .B1(n16434), 
        .B2(n19120), .ZN(n16404) );
  AOI222_X1 U19421 ( .A1(n16402), .A2(n16441), .B1(n16421), .B2(n19121), .C1(
        n16435), .C2(n16401), .ZN(n16403) );
  OAI211_X1 U19422 ( .C1(n19114), .C2(n16445), .A(n16404), .B(n16403), .ZN(
        P2_U3003) );
  AOI22_X1 U19423 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n11600), .B1(n16434), 
        .B2(n19144), .ZN(n16408) );
  AOI222_X1 U19424 ( .A1(n16406), .A2(n16435), .B1(n16441), .B2(n16405), .C1(
        n16421), .C2(n19145), .ZN(n16407) );
  OAI211_X1 U19425 ( .C1(n19139), .C2(n16445), .A(n16408), .B(n16407), .ZN(
        P2_U3005) );
  AOI22_X1 U19426 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n11600), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16409), .ZN(n16423) );
  INV_X1 U19427 ( .A(n19158), .ZN(n16466) );
  XOR2_X1 U19428 ( .A(n16410), .B(n16411), .Z(n16467) );
  NAND2_X1 U19429 ( .A1(n16413), .A2(n16412), .ZN(n16418) );
  INV_X1 U19430 ( .A(n16414), .ZN(n16415) );
  AOI21_X1 U19431 ( .B1(n15394), .B2(n16416), .A(n16415), .ZN(n16417) );
  XOR2_X1 U19432 ( .A(n16418), .B(n16417), .Z(n16465) );
  AOI22_X1 U19433 ( .A1(n16467), .A2(n16435), .B1(n16441), .B2(n16465), .ZN(
        n16419) );
  INV_X1 U19434 ( .A(n16419), .ZN(n16420) );
  AOI21_X1 U19435 ( .B1(n16421), .B2(n16466), .A(n16420), .ZN(n16422) );
  OAI211_X1 U19436 ( .C1(n16424), .C2(n19152), .A(n16423), .B(n16422), .ZN(
        P2_U3006) );
  AOI22_X1 U19437 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n11600), .B1(n16434), 
        .B2(n19191), .ZN(n16431) );
  OAI222_X1 U19438 ( .A1(n19199), .A2(n16439), .B1(n16428), .B2(n16427), .C1(
        n16426), .C2(n16425), .ZN(n16429) );
  INV_X1 U19439 ( .A(n16429), .ZN(n16430) );
  OAI211_X1 U19440 ( .C1(n16432), .C2(n16445), .A(n16431), .B(n16430), .ZN(
        P2_U3009) );
  AOI22_X1 U19441 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n11600), .B1(n16434), 
        .B2(n16433), .ZN(n16444) );
  NAND3_X1 U19442 ( .A1(n16436), .A2(n13278), .A3(n16435), .ZN(n16437) );
  OAI21_X1 U19443 ( .B1(n16439), .B2(n16438), .A(n16437), .ZN(n16440) );
  AOI21_X1 U19444 ( .B1(n16442), .B2(n16441), .A(n16440), .ZN(n16443) );
  OAI211_X1 U19445 ( .C1(n16446), .C2(n16445), .A(n16444), .B(n16443), .ZN(
        P2_U3011) );
  AOI21_X1 U19446 ( .B1(n16449), .B2(n16448), .A(n16447), .ZN(n19257) );
  INV_X1 U19447 ( .A(n16450), .ZN(n16451) );
  NOR3_X1 U19448 ( .A1(n16452), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16451), .ZN(n16453) );
  AOI21_X1 U19449 ( .B1(n16474), .B2(n19257), .A(n16453), .ZN(n16461) );
  AOI222_X1 U19450 ( .A1(n16455), .A2(n19391), .B1(n19395), .B2(n16454), .C1(
        n16475), .C2(n19097), .ZN(n16460) );
  NAND2_X1 U19451 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19180), .ZN(n16459) );
  OAI21_X1 U19452 ( .B1(n16457), .B2(n16456), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16458) );
  NAND4_X1 U19453 ( .A1(n16461), .A2(n16460), .A3(n16459), .A4(n16458), .ZN(
        P2_U3032) );
  AOI21_X1 U19454 ( .B1(n16463), .B2(n16462), .A(n15673), .ZN(n19157) );
  AOI22_X1 U19455 ( .A1(n16474), .A2(n19157), .B1(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16464), .ZN(n16473) );
  AOI222_X1 U19456 ( .A1(n16467), .A2(n19391), .B1(n16475), .B2(n16466), .C1(
        n16465), .C2(n19395), .ZN(n16472) );
  NAND2_X1 U19457 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19180), .ZN(n16471) );
  OAI211_X1 U19458 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16469), .B(n16468), .ZN(n16470) );
  NAND4_X1 U19459 ( .A1(n16473), .A2(n16472), .A3(n16471), .A4(n16470), .ZN(
        P2_U3038) );
  AOI22_X1 U19460 ( .A1(n19231), .A2(n16475), .B1(n16474), .B2(n19225), .ZN(
        n16483) );
  OR2_X1 U19461 ( .A1(n16477), .A2(n16476), .ZN(n16482) );
  NAND2_X1 U19462 ( .A1(n19391), .A2(n16478), .ZN(n16481) );
  NAND2_X1 U19463 ( .A1(n16479), .A2(n20916), .ZN(n16480) );
  AND4_X1 U19464 ( .A1(n16483), .A2(n16482), .A3(n16481), .A4(n16480), .ZN(
        n16485) );
  OAI211_X1 U19465 ( .C1(n19385), .C2(n20916), .A(n16485), .B(n16484), .ZN(
        P2_U3046) );
  OAI221_X1 U19466 ( .B1(n20037), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n20037), 
        .C2(n16487), .A(n16486), .ZN(P2_U3593) );
  NOR2_X1 U19467 ( .A1(n16489), .A2(n16488), .ZN(n18772) );
  INV_X1 U19468 ( .A(n17843), .ZN(n17803) );
  INV_X1 U19469 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20970) );
  INV_X1 U19470 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21028) );
  NAND2_X1 U19471 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17967) );
  NOR2_X1 U19472 ( .A1(n17909), .A2(n16937), .ZN(n16925) );
  INV_X1 U19473 ( .A(n16925), .ZN(n17902) );
  NOR2_X1 U19474 ( .A1(n17901), .A2(n17902), .ZN(n16490) );
  NAND4_X1 U19475 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(n16490), .ZN(n17828) );
  NAND2_X1 U19476 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17830) );
  INV_X1 U19477 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17772) );
  INV_X1 U19478 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17702) );
  NAND2_X1 U19479 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17674) );
  INV_X1 U19480 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17661) );
  INV_X1 U19481 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17634) );
  INV_X1 U19482 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16707) );
  NAND3_X1 U19483 ( .A1(n17673), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17660) );
  NOR2_X1 U19484 ( .A1(n17661), .A2(n17660), .ZN(n17633) );
  NAND3_X1 U19485 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n17633), .ZN(n16535) );
  NOR2_X1 U19486 ( .A1(n16707), .A2(n16535), .ZN(n16491) );
  NAND2_X1 U19487 ( .A1(n18974), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17995) );
  NOR2_X2 U19488 ( .A1(n18367), .A2(n18672), .ZN(n18704) );
  AOI21_X1 U19489 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17738), .A(
        n18704), .ZN(n17829) );
  INV_X1 U19490 ( .A(n17829), .ZN(n17785) );
  NAND2_X1 U19491 ( .A1(n16491), .A2(n17785), .ZN(n16513) );
  XNOR2_X1 U19492 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16493) );
  NAND2_X1 U19493 ( .A1(n16707), .A2(n17738), .ZN(n16521) );
  INV_X1 U19494 ( .A(n16521), .ZN(n16492) );
  OR2_X1 U19495 ( .A1(n18358), .A2(n16491), .ZN(n16534) );
  OAI211_X1 U19496 ( .C1(n16677), .C2(n17995), .A(n17996), .B(n16534), .ZN(
        n16524) );
  NOR2_X1 U19497 ( .A1(n16492), .A2(n16524), .ZN(n16511) );
  OAI22_X1 U19498 ( .A1(n16513), .A2(n16493), .B1(n16511), .B2(n20970), .ZN(
        n16494) );
  AOI211_X1 U19499 ( .C1(n17803), .C2(n16879), .A(n16495), .B(n16494), .ZN(
        n16501) );
  INV_X1 U19500 ( .A(n16496), .ZN(n16497) );
  OAI211_X1 U19501 ( .C1(n18000), .C2(n16502), .A(n16501), .B(n16500), .ZN(
        P3_U2799) );
  NAND3_X1 U19502 ( .A1(n16504), .A2(n16503), .A3(n17779), .ZN(n16519) );
  AOI22_X1 U19503 ( .A1(n17900), .A2(n16525), .B1(n9775), .B2(n16505), .ZN(
        n16517) );
  INV_X1 U19504 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16512) );
  OAI21_X1 U19505 ( .B1(n16507), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16506), .ZN(n16699) );
  INV_X1 U19506 ( .A(n16699), .ZN(n16509) );
  AOI21_X1 U19507 ( .B1(n16509), .B2(n17803), .A(n16508), .ZN(n16510) );
  OAI221_X1 U19508 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16513), .C1(
        n16512), .C2(n16511), .A(n16510), .ZN(n16514) );
  AOI21_X1 U19509 ( .B1(n17888), .B2(n16515), .A(n16514), .ZN(n16516) );
  OAI221_X1 U19510 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16519), 
        .C1(n16518), .C2(n16517), .A(n16516), .ZN(P3_U2800) );
  INV_X1 U19511 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18912) );
  NOR2_X1 U19512 ( .A1(n18199), .A2(n18912), .ZN(n16523) );
  OAI21_X1 U19513 ( .B1(n16677), .B2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16520), .ZN(n16711) );
  AOI21_X1 U19514 ( .B1(n17843), .B2(n16521), .A(n16711), .ZN(n16522) );
  AOI211_X1 U19515 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16524), .A(
        n16523), .B(n16522), .ZN(n16533) );
  NAND2_X1 U19516 ( .A1(n17900), .A2(n16525), .ZN(n16526) );
  AOI21_X1 U19517 ( .B1(n16541), .B2(n16528), .A(n16526), .ZN(n16530) );
  AOI211_X1 U19518 ( .C1(n16528), .C2(n16542), .A(n16527), .B(n18000), .ZN(
        n16529) );
  AOI211_X1 U19519 ( .C1(n17888), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        n16532) );
  OAI211_X1 U19520 ( .C1(n16535), .C2(n16534), .A(n16533), .B(n16532), .ZN(
        P3_U2801) );
  NOR2_X1 U19521 ( .A1(n16536), .A2(n18773), .ZN(n18133) );
  INV_X1 U19522 ( .A(n18133), .ZN(n18159) );
  OAI22_X1 U19523 ( .A1(n18162), .A2(n18279), .B1(n17835), .B2(n18159), .ZN(
        n18170) );
  AOI21_X1 U19524 ( .B1(n16538), .B2(n18170), .A(n16537), .ZN(n18056) );
  NOR2_X1 U19525 ( .A1(n18056), .A2(n18289), .ZN(n18075) );
  NOR2_X1 U19526 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16539), .ZN(
        n17645) );
  AOI22_X1 U19527 ( .A1(n18301), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18075), 
        .B2(n17645), .ZN(n16552) );
  INV_X1 U19528 ( .A(n17650), .ZN(n16540) );
  AOI21_X1 U19529 ( .B1(n17871), .B2(n16540), .A(n17651), .ZN(n17642) );
  AOI22_X1 U19530 ( .A1(n17871), .A2(n17638), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17897), .ZN(n17641) );
  NOR2_X1 U19531 ( .A1(n17642), .A2(n17641), .ZN(n17640) );
  AOI211_X1 U19532 ( .C1(n17650), .C2(n16548), .A(n17640), .B(n18137), .ZN(
        n16546) );
  AOI22_X1 U19533 ( .A1(n18767), .A2(n16542), .B1(n18133), .B2(n16541), .ZN(
        n16543) );
  NAND2_X1 U19534 ( .A1(n16544), .A2(n16543), .ZN(n16545) );
  OAI211_X1 U19535 ( .C1(n16546), .C2(n16545), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18199), .ZN(n16551) );
  INV_X1 U19536 ( .A(n17640), .ZN(n16547) );
  NAND4_X1 U19537 ( .A1(n16548), .A2(n18203), .A3(n17638), .A4(n16547), .ZN(
        n16550) );
  NAND3_X1 U19538 ( .A1(n18203), .A2(n17651), .A3(n17641), .ZN(n16549) );
  NAND4_X1 U19539 ( .A1(n16552), .A2(n16551), .A3(n16550), .A4(n16549), .ZN(
        P3_U2834) );
  NOR3_X1 U19540 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16554) );
  NOR4_X1 U19541 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16553) );
  NAND4_X1 U19542 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16554), .A3(n16553), .A4(
        U215), .ZN(U213) );
  INV_X2 U19543 ( .A(U214), .ZN(n16603) );
  NOR2_X1 U19544 ( .A1(n16603), .A2(n16555), .ZN(n16601) );
  AOI222_X1 U19545 ( .A1(n16600), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(n16601), 
        .B2(BUF1_REG_31__SCAN_IN), .C1(n16603), .C2(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n16556) );
  INV_X1 U19546 ( .A(n16556), .ZN(U216) );
  INV_X1 U19547 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19316) );
  INV_X1 U19548 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16640) );
  OAI222_X1 U19549 ( .A1(U212), .A2(n19316), .B1(n16605), .B2(n14628), .C1(
        U214), .C2(n16640), .ZN(U217) );
  AOI22_X1 U19550 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16600), .ZN(n16557) );
  OAI21_X1 U19551 ( .B1(n14636), .B2(n16605), .A(n16557), .ZN(U218) );
  AOI22_X1 U19552 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16600), .ZN(n16558) );
  OAI21_X1 U19553 ( .B1(n16559), .B2(n16605), .A(n16558), .ZN(U219) );
  AOI22_X1 U19554 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16600), .ZN(n16560) );
  OAI21_X1 U19555 ( .B1(n14650), .B2(n16605), .A(n16560), .ZN(U220) );
  AOI22_X1 U19556 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16600), .ZN(n16561) );
  OAI21_X1 U19557 ( .B1(n14656), .B2(n16605), .A(n16561), .ZN(U221) );
  INV_X1 U19558 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16563) );
  AOI22_X1 U19559 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16600), .ZN(n16562) );
  OAI21_X1 U19560 ( .B1(n16563), .B2(n16605), .A(n16562), .ZN(U222) );
  AOI22_X1 U19561 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16600), .ZN(n16564) );
  OAI21_X1 U19562 ( .B1(n16565), .B2(n16605), .A(n16564), .ZN(U223) );
  AOI22_X1 U19563 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16600), .ZN(n16566) );
  OAI21_X1 U19564 ( .B1(n14673), .B2(n16605), .A(n16566), .ZN(U224) );
  INV_X1 U19565 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16568) );
  AOI22_X1 U19566 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16600), .ZN(n16567) );
  OAI21_X1 U19567 ( .B1(n16568), .B2(n16605), .A(n16567), .ZN(U225) );
  AOI222_X1 U19568 ( .A1(n16600), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(n16601), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16603), .C2(P1_DATAO_REG_21__SCAN_IN), 
        .ZN(n16569) );
  INV_X1 U19569 ( .A(n16569), .ZN(U226) );
  INV_X1 U19570 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16571) );
  AOI22_X1 U19571 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16600), .ZN(n16570) );
  OAI21_X1 U19572 ( .B1(n16571), .B2(n16605), .A(n16570), .ZN(U227) );
  AOI222_X1 U19573 ( .A1(n16600), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n16601), 
        .B2(BUF1_REG_19__SCAN_IN), .C1(n16603), .C2(P1_DATAO_REG_19__SCAN_IN), 
        .ZN(n16572) );
  INV_X1 U19574 ( .A(n16572), .ZN(U228) );
  AOI22_X1 U19575 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16600), .ZN(n16573) );
  OAI21_X1 U19576 ( .B1(n14703), .B2(n16605), .A(n16573), .ZN(U229) );
  AOI22_X1 U19577 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16600), .ZN(n16574) );
  OAI21_X1 U19578 ( .B1(n14710), .B2(n16605), .A(n16574), .ZN(U230) );
  AOI22_X1 U19579 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16600), .ZN(n16575) );
  OAI21_X1 U19580 ( .B1(n14718), .B2(n16605), .A(n16575), .ZN(U231) );
  AOI22_X1 U19581 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16600), .ZN(n16576) );
  OAI21_X1 U19582 ( .B1(n12973), .B2(n16605), .A(n16576), .ZN(U232) );
  AOI22_X1 U19583 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16600), .ZN(n16577) );
  OAI21_X1 U19584 ( .B1(n15186), .B2(n16605), .A(n16577), .ZN(U233) );
  AOI22_X1 U19585 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16600), .ZN(n16578) );
  OAI21_X1 U19586 ( .B1(n12659), .B2(n16605), .A(n16578), .ZN(U234) );
  INV_X1 U19587 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16580) );
  AOI22_X1 U19588 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16600), .ZN(n16579) );
  OAI21_X1 U19589 ( .B1(n16580), .B2(n16605), .A(n16579), .ZN(U235) );
  AOI22_X1 U19590 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16600), .ZN(n16581) );
  OAI21_X1 U19591 ( .B1(n12666), .B2(n16605), .A(n16581), .ZN(U236) );
  AOI22_X1 U19592 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16600), .ZN(n16582) );
  OAI21_X1 U19593 ( .B1(n16583), .B2(n16605), .A(n16582), .ZN(U237) );
  AOI22_X1 U19594 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16600), .ZN(n16584) );
  OAI21_X1 U19595 ( .B1(n16585), .B2(n16605), .A(n16584), .ZN(U238) );
  INV_X1 U19596 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16587) );
  AOI22_X1 U19597 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16600), .ZN(n16586) );
  OAI21_X1 U19598 ( .B1(n16587), .B2(n16605), .A(n16586), .ZN(U239) );
  INV_X1 U19599 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16589) );
  AOI22_X1 U19600 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16600), .ZN(n16588) );
  OAI21_X1 U19601 ( .B1(n16589), .B2(n16605), .A(n16588), .ZN(U240) );
  INV_X1 U19602 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16591) );
  AOI22_X1 U19603 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16600), .ZN(n16590) );
  OAI21_X1 U19604 ( .B1(n16591), .B2(n16605), .A(n16590), .ZN(U241) );
  INV_X1 U19605 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U19606 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16600), .ZN(n16592) );
  OAI21_X1 U19607 ( .B1(n16593), .B2(n16605), .A(n16592), .ZN(U242) );
  INV_X1 U19608 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16595) );
  AOI22_X1 U19609 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16600), .ZN(n16594) );
  OAI21_X1 U19610 ( .B1(n16595), .B2(n16605), .A(n16594), .ZN(U243) );
  INV_X1 U19611 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16597) );
  AOI22_X1 U19612 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16600), .ZN(n16596) );
  OAI21_X1 U19613 ( .B1(n16597), .B2(n16605), .A(n16596), .ZN(U244) );
  INV_X1 U19614 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16599) );
  AOI22_X1 U19615 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16600), .ZN(n16598) );
  OAI21_X1 U19616 ( .B1(n16599), .B2(n16605), .A(n16598), .ZN(U245) );
  INV_X1 U19617 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n20972) );
  AOI22_X1 U19618 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16601), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16600), .ZN(n16602) );
  OAI21_X1 U19619 ( .B1(n20972), .B2(U214), .A(n16602), .ZN(U246) );
  INV_X1 U19620 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16606) );
  AOI22_X1 U19621 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16603), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16600), .ZN(n16604) );
  OAI21_X1 U19622 ( .B1(n16606), .B2(n16605), .A(n16604), .ZN(U247) );
  OAI22_X1 U19623 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16638), .ZN(n16607) );
  INV_X1 U19624 ( .A(n16607), .ZN(U251) );
  OAI22_X1 U19625 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16638), .ZN(n16608) );
  INV_X1 U19626 ( .A(n16608), .ZN(U252) );
  OAI22_X1 U19627 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16638), .ZN(n16609) );
  INV_X1 U19628 ( .A(n16609), .ZN(U253) );
  OAI22_X1 U19629 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16638), .ZN(n16610) );
  INV_X1 U19630 ( .A(n16610), .ZN(U254) );
  OAI22_X1 U19631 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16638), .ZN(n16611) );
  INV_X1 U19632 ( .A(n16611), .ZN(U255) );
  OAI22_X1 U19633 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16638), .ZN(n16612) );
  INV_X1 U19634 ( .A(n16612), .ZN(U256) );
  OAI22_X1 U19635 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16638), .ZN(n16613) );
  INV_X1 U19636 ( .A(n16613), .ZN(U257) );
  OAI22_X1 U19637 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16638), .ZN(n16614) );
  INV_X1 U19638 ( .A(n16614), .ZN(U258) );
  OAI22_X1 U19639 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16630), .ZN(n16615) );
  INV_X1 U19640 ( .A(n16615), .ZN(U259) );
  OAI22_X1 U19641 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16630), .ZN(n16616) );
  INV_X1 U19642 ( .A(n16616), .ZN(U260) );
  OAI22_X1 U19643 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16630), .ZN(n16617) );
  INV_X1 U19644 ( .A(n16617), .ZN(U261) );
  OAI22_X1 U19645 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16630), .ZN(n16618) );
  INV_X1 U19646 ( .A(n16618), .ZN(U262) );
  OAI22_X1 U19647 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16630), .ZN(n16619) );
  INV_X1 U19648 ( .A(n16619), .ZN(U263) );
  OAI22_X1 U19649 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16630), .ZN(n16620) );
  INV_X1 U19650 ( .A(n16620), .ZN(U264) );
  OAI22_X1 U19651 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16630), .ZN(n16621) );
  INV_X1 U19652 ( .A(n16621), .ZN(U265) );
  OAI22_X1 U19653 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16638), .ZN(n16622) );
  INV_X1 U19654 ( .A(n16622), .ZN(U266) );
  OAI22_X1 U19655 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16638), .ZN(n16623) );
  INV_X1 U19656 ( .A(n16623), .ZN(U267) );
  OAI22_X1 U19657 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16630), .ZN(n16624) );
  INV_X1 U19658 ( .A(n16624), .ZN(U268) );
  OAI22_X1 U19659 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16638), .ZN(n16625) );
  INV_X1 U19660 ( .A(n16625), .ZN(U269) );
  OAI22_X1 U19661 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16630), .ZN(n16626) );
  INV_X1 U19662 ( .A(n16626), .ZN(U270) );
  OAI22_X1 U19663 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16638), .ZN(n16627) );
  INV_X1 U19664 ( .A(n16627), .ZN(U271) );
  INV_X1 U19665 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16628) );
  INV_X1 U19666 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U19667 ( .A1(n16638), .A2(n16628), .B1(n18345), .B2(U215), .ZN(U272) );
  OAI22_X1 U19668 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16638), .ZN(n16629) );
  INV_X1 U19669 ( .A(n16629), .ZN(U273) );
  OAI22_X1 U19670 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16630), .ZN(n16631) );
  INV_X1 U19671 ( .A(n16631), .ZN(U274) );
  OAI22_X1 U19672 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16638), .ZN(n16632) );
  INV_X1 U19673 ( .A(n16632), .ZN(U275) );
  OAI22_X1 U19674 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16638), .ZN(n16633) );
  INV_X1 U19675 ( .A(n16633), .ZN(U276) );
  OAI22_X1 U19676 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16638), .ZN(n16634) );
  INV_X1 U19677 ( .A(n16634), .ZN(U277) );
  OAI22_X1 U19678 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16638), .ZN(n16635) );
  INV_X1 U19679 ( .A(n16635), .ZN(U278) );
  OAI22_X1 U19680 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16638), .ZN(n16636) );
  INV_X1 U19681 ( .A(n16636), .ZN(U279) );
  OAI22_X1 U19682 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16638), .ZN(n16637) );
  INV_X1 U19683 ( .A(n16637), .ZN(U280) );
  INV_X1 U19684 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U19685 ( .A1(n16638), .A2(n19316), .B1(n18350), .B2(U215), .ZN(U281) );
  INV_X1 U19686 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19310) );
  INV_X1 U19687 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18359) );
  AOI22_X1 U19688 ( .A1(n16638), .A2(n19310), .B1(n18359), .B2(U215), .ZN(U282) );
  INV_X1 U19689 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16639) );
  OAI222_X1 U19690 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n16640), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n19316), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16639), .ZN(n16641) );
  INV_X1 U19691 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18875) );
  INV_X1 U19692 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U19693 ( .A1(n9737), .A2(n18875), .B1(n19987), .B2(n16642), .ZN(
        U347) );
  INV_X1 U19694 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18873) );
  INV_X1 U19695 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19986) );
  AOI22_X1 U19696 ( .A1(n9737), .A2(n18873), .B1(n19986), .B2(n16642), .ZN(
        U348) );
  INV_X1 U19697 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18870) );
  INV_X1 U19698 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n21021) );
  AOI22_X1 U19699 ( .A1(n9737), .A2(n18870), .B1(n21021), .B2(n16642), .ZN(
        U349) );
  INV_X1 U19700 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18869) );
  INV_X1 U19701 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U19702 ( .A1(n9737), .A2(n18869), .B1(n19983), .B2(n16642), .ZN(
        U350) );
  INV_X1 U19703 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18867) );
  INV_X1 U19704 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U19705 ( .A1(n9737), .A2(n18867), .B1(n19981), .B2(n16642), .ZN(
        U351) );
  INV_X1 U19706 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18864) );
  INV_X1 U19707 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19979) );
  AOI22_X1 U19708 ( .A1(n9737), .A2(n18864), .B1(n19979), .B2(n16642), .ZN(
        U352) );
  INV_X1 U19709 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18863) );
  INV_X1 U19710 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19977) );
  AOI22_X1 U19711 ( .A1(n9737), .A2(n18863), .B1(n19977), .B2(n16642), .ZN(
        U353) );
  INV_X1 U19712 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18860) );
  AOI22_X1 U19713 ( .A1(n9737), .A2(n18860), .B1(n19974), .B2(n16642), .ZN(
        U354) );
  INV_X1 U19714 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18915) );
  INV_X1 U19715 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20019) );
  AOI22_X1 U19716 ( .A1(n9737), .A2(n18915), .B1(n20019), .B2(n16641), .ZN(
        U355) );
  INV_X1 U19717 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18913) );
  INV_X1 U19718 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U19719 ( .A1(n9737), .A2(n18913), .B1(n20016), .B2(n16642), .ZN(
        U356) );
  INV_X1 U19720 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18909) );
  INV_X1 U19721 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20014) );
  AOI22_X1 U19722 ( .A1(n9737), .A2(n18909), .B1(n20014), .B2(n16642), .ZN(
        U357) );
  INV_X1 U19723 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18907) );
  INV_X1 U19724 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U19725 ( .A1(n9737), .A2(n18907), .B1(n20012), .B2(n16641), .ZN(
        U358) );
  INV_X1 U19726 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18904) );
  INV_X1 U19727 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20011) );
  AOI22_X1 U19728 ( .A1(n9737), .A2(n18904), .B1(n20011), .B2(n16641), .ZN(
        U359) );
  INV_X1 U19729 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18903) );
  INV_X1 U19730 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20010) );
  AOI22_X1 U19731 ( .A1(n9737), .A2(n18903), .B1(n20010), .B2(n16641), .ZN(
        U360) );
  INV_X1 U19732 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18901) );
  INV_X1 U19733 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20008) );
  AOI22_X1 U19734 ( .A1(n9737), .A2(n18901), .B1(n20008), .B2(n16641), .ZN(
        U361) );
  INV_X1 U19735 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18899) );
  INV_X1 U19736 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U19737 ( .A1(n9737), .A2(n18899), .B1(n20007), .B2(n16642), .ZN(
        U362) );
  INV_X1 U19738 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18897) );
  INV_X1 U19739 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U19740 ( .A1(n9737), .A2(n18897), .B1(n20006), .B2(n16642), .ZN(
        U363) );
  INV_X1 U19741 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18895) );
  INV_X1 U19742 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20004) );
  AOI22_X1 U19743 ( .A1(n9737), .A2(n18895), .B1(n20004), .B2(n16642), .ZN(
        U364) );
  INV_X1 U19744 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18859) );
  INV_X1 U19745 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19972) );
  AOI22_X1 U19746 ( .A1(n9737), .A2(n18859), .B1(n19972), .B2(n16642), .ZN(
        U365) );
  INV_X1 U19747 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18892) );
  INV_X1 U19748 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20003) );
  AOI22_X1 U19749 ( .A1(n9737), .A2(n18892), .B1(n20003), .B2(n16642), .ZN(
        U366) );
  INV_X1 U19750 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18891) );
  INV_X1 U19751 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20001) );
  AOI22_X1 U19752 ( .A1(n9737), .A2(n18891), .B1(n20001), .B2(n16642), .ZN(
        U367) );
  INV_X1 U19753 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18890) );
  INV_X1 U19754 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20907) );
  AOI22_X1 U19755 ( .A1(n9737), .A2(n18890), .B1(n20907), .B2(n16642), .ZN(
        U368) );
  INV_X1 U19756 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18888) );
  INV_X1 U19757 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20825) );
  AOI22_X1 U19758 ( .A1(n9737), .A2(n18888), .B1(n20825), .B2(n16642), .ZN(
        U369) );
  INV_X1 U19759 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18887) );
  INV_X1 U19760 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19998) );
  AOI22_X1 U19761 ( .A1(n9737), .A2(n18887), .B1(n19998), .B2(n16642), .ZN(
        U370) );
  INV_X1 U19762 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18885) );
  INV_X1 U19763 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19996) );
  AOI22_X1 U19764 ( .A1(n9737), .A2(n18885), .B1(n19996), .B2(n16642), .ZN(
        U371) );
  INV_X1 U19765 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18882) );
  INV_X1 U19766 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20915) );
  AOI22_X1 U19767 ( .A1(n9737), .A2(n18882), .B1(n20915), .B2(n16641), .ZN(
        U372) );
  INV_X1 U19768 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18881) );
  INV_X1 U19769 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U19770 ( .A1(n9737), .A2(n18881), .B1(n19993), .B2(n16642), .ZN(
        U373) );
  INV_X1 U19771 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18879) );
  INV_X1 U19772 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19991) );
  AOI22_X1 U19773 ( .A1(n9737), .A2(n18879), .B1(n19991), .B2(n16641), .ZN(
        U374) );
  INV_X1 U19774 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18877) );
  INV_X1 U19775 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19989) );
  AOI22_X1 U19776 ( .A1(n9737), .A2(n18877), .B1(n19989), .B2(n16641), .ZN(
        U375) );
  INV_X1 U19777 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18858) );
  INV_X1 U19778 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U19779 ( .A1(n9737), .A2(n18858), .B1(n19971), .B2(n16642), .ZN(
        U376) );
  INV_X1 U19780 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18857) );
  NAND2_X1 U19781 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18857), .ZN(n16643) );
  INV_X1 U19782 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18845) );
  AOI22_X1 U19783 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n16643), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18845), .ZN(n18925) );
  AOI21_X1 U19784 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18925), .ZN(n16644) );
  INV_X1 U19785 ( .A(n16644), .ZN(P3_U2633) );
  NAND2_X1 U19786 ( .A1(n18987), .A2(n18986), .ZN(n16647) );
  NOR2_X1 U19787 ( .A1(n17580), .A2(n16650), .ZN(n16645) );
  NAND2_X1 U19788 ( .A1(n18977), .A2(n18771), .ZN(n17521) );
  OAI21_X1 U19789 ( .B1(n16645), .B2(n17521), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16646) );
  OAI21_X1 U19790 ( .B1(n16647), .B2(n18974), .A(n16646), .ZN(P3_U2634) );
  AOI21_X1 U19791 ( .B1(n18852), .B2(n18857), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16648) );
  AOI22_X1 U19792 ( .A1(n18983), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16648), 
        .B2(n18984), .ZN(P3_U2635) );
  NOR2_X1 U19793 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18843) );
  OAI21_X1 U19794 ( .B1(n18843), .B2(BS16), .A(n18925), .ZN(n18923) );
  OAI21_X1 U19795 ( .B1(n18925), .B2(n16668), .A(n18923), .ZN(P3_U2636) );
  OAI211_X1 U19796 ( .C1(n17580), .C2(n16650), .A(n16649), .B(n18771), .ZN(
        n16651) );
  INV_X1 U19797 ( .A(n16651), .ZN(n18774) );
  NOR2_X1 U19798 ( .A1(n18774), .A2(n18832), .ZN(n18967) );
  OAI21_X1 U19799 ( .B1(n18967), .B2(n18309), .A(n16652), .ZN(P3_U2637) );
  NOR4_X1 U19800 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16656) );
  NOR4_X1 U19801 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16655) );
  NOR4_X1 U19802 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16654) );
  NOR4_X1 U19803 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16653) );
  NAND4_X1 U19804 ( .A1(n16656), .A2(n16655), .A3(n16654), .A4(n16653), .ZN(
        n16662) );
  NOR4_X1 U19805 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16660) );
  AOI211_X1 U19806 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_7__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16659) );
  NOR4_X1 U19807 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16658) );
  NOR4_X1 U19808 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16657) );
  NAND4_X1 U19809 ( .A1(n16660), .A2(n16659), .A3(n16658), .A4(n16657), .ZN(
        n16661) );
  NOR2_X1 U19810 ( .A1(n16662), .A2(n16661), .ZN(n18965) );
  INV_X1 U19811 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16664) );
  NOR3_X1 U19812 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16665) );
  OAI21_X1 U19813 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16665), .A(n18965), .ZN(
        n16663) );
  OAI21_X1 U19814 ( .B1(n18965), .B2(n16664), .A(n16663), .ZN(P3_U2638) );
  INV_X1 U19815 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18958) );
  INV_X1 U19816 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18924) );
  AOI21_X1 U19817 ( .B1(n18958), .B2(n18924), .A(n16665), .ZN(n16667) );
  INV_X1 U19818 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16666) );
  INV_X1 U19819 ( .A(n18965), .ZN(n18960) );
  AOI22_X1 U19820 ( .A1(n18965), .A2(n16667), .B1(n16666), .B2(n18960), .ZN(
        P3_U2639) );
  NAND3_X1 U19821 ( .A1(n18974), .A2(n18986), .A3(n16668), .ZN(n18841) );
  OR2_X1 U19822 ( .A1(n18937), .A2(n18841), .ZN(n18839) );
  INV_X2 U19823 ( .A(n18839), .ZN(n17014) );
  NOR2_X1 U19824 ( .A1(n21062), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18834) );
  INV_X1 U19825 ( .A(n18834), .ZN(n18706) );
  NOR2_X1 U19826 ( .A1(n18836), .A2(n18706), .ZN(n18827) );
  NOR4_X2 U19827 ( .A1(n18235), .A2(n18989), .A3(n17014), .A4(n18827), .ZN(
        n17030) );
  INV_X1 U19828 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n17052) );
  INV_X1 U19829 ( .A(n18850), .ZN(n18969) );
  OAI211_X1 U19830 ( .C1(n18969), .C2(n18970), .A(n18979), .B(n16668), .ZN(
        n18825) );
  OAI211_X2 U19831 ( .C1(n17052), .C2(n18324), .A(n18825), .B(n16670), .ZN(
        n17033) );
  AOI22_X1 U19832 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16997), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17044), .ZN(n16693) );
  NAND2_X1 U19833 ( .A1(n16668), .A2(n18979), .ZN(n16669) );
  INV_X1 U19834 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16728) );
  NOR2_X1 U19835 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17029) );
  NAND2_X1 U19836 ( .A1(n17029), .A2(n20977), .ZN(n17017) );
  NOR2_X1 U19837 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17017), .ZN(n17002) );
  INV_X1 U19838 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17351) );
  NAND2_X1 U19839 ( .A1(n17002), .A2(n17351), .ZN(n16984) );
  NOR2_X1 U19840 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16984), .ZN(n16972) );
  INV_X1 U19841 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17343) );
  NAND2_X1 U19842 ( .A1(n16972), .A2(n17343), .ZN(n16962) );
  NOR2_X1 U19843 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16962), .ZN(n16951) );
  INV_X1 U19844 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17248) );
  NAND2_X1 U19845 ( .A1(n16951), .A2(n17248), .ZN(n16939) );
  INV_X1 U19846 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20934) );
  NAND2_X1 U19847 ( .A1(n16928), .A2(n20934), .ZN(n16920) );
  NAND2_X1 U19848 ( .A1(n16904), .A2(n17267), .ZN(n16893) );
  INV_X1 U19849 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17250) );
  NAND2_X1 U19850 ( .A1(n16874), .A2(n17250), .ZN(n16868) );
  NAND2_X1 U19851 ( .A1(n16855), .A2(n17218), .ZN(n16840) );
  INV_X1 U19852 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20985) );
  NAND2_X1 U19853 ( .A1(n16829), .A2(n20985), .ZN(n16823) );
  NAND2_X1 U19854 ( .A1(n16811), .A2(n17152), .ZN(n16806) );
  NOR2_X1 U19855 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16806), .ZN(n16794) );
  NAND2_X1 U19856 ( .A1(n16794), .A2(n16788), .ZN(n16787) );
  NOR2_X1 U19857 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16787), .ZN(n16769) );
  NAND2_X1 U19858 ( .A1(n16769), .A2(n16757), .ZN(n16756) );
  NOR2_X1 U19859 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16756), .ZN(n16747) );
  INV_X1 U19860 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n20956) );
  NAND2_X1 U19861 ( .A1(n16747), .A2(n20956), .ZN(n16736) );
  INV_X1 U19862 ( .A(n16736), .ZN(n16727) );
  NAND2_X1 U19863 ( .A1(n16728), .A2(n16727), .ZN(n16726) );
  OR2_X1 U19864 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16717), .ZN(n16695) );
  NOR2_X1 U19865 ( .A1(n16999), .A2(n16695), .ZN(n16696) );
  INV_X1 U19866 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16676) );
  INV_X1 U19867 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18905) );
  INV_X1 U19868 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18900) );
  INV_X1 U19869 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18898) );
  INV_X1 U19870 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18880) );
  INV_X1 U19871 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18876) );
  NAND3_X1 U19872 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n16910) );
  NAND2_X1 U19873 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16912) );
  INV_X1 U19874 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18871) );
  NAND2_X1 U19875 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16955) );
  NOR2_X1 U19876 ( .A1(n18871), .A2(n16955), .ZN(n16917) );
  NAND3_X1 U19877 ( .A1(n16917), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_9__SCAN_IN), .ZN(n16903) );
  NOR4_X1 U19878 ( .A1(n18876), .A2(n16910), .A3(n16912), .A4(n16903), .ZN(
        n16880) );
  NAND2_X1 U19879 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16880), .ZN(n16883) );
  NOR2_X1 U19880 ( .A1(n18880), .A2(n16883), .ZN(n16862) );
  NAND2_X1 U19881 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16862), .ZN(n16779) );
  INV_X1 U19882 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18889) );
  NAND2_X1 U19883 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16839) );
  NOR2_X1 U19884 ( .A1(n18889), .A2(n16839), .ZN(n16780) );
  NAND4_X1 U19885 ( .A1(n16780), .A2(P3_REIP_REG_20__SCAN_IN), .A3(
        P3_REIP_REG_18__SCAN_IN), .A4(P3_REIP_REG_19__SCAN_IN), .ZN(n16793) );
  NAND2_X1 U19886 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16783) );
  OR3_X1 U19887 ( .A1(n16779), .A2(n16793), .A3(n16783), .ZN(n16771) );
  NOR2_X1 U19888 ( .A1(n18898), .A2(n16771), .ZN(n16759) );
  INV_X1 U19889 ( .A(n16759), .ZN(n16746) );
  NOR2_X1 U19890 ( .A1(n18900), .A2(n16746), .ZN(n16751) );
  NAND2_X1 U19891 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16751), .ZN(n16737) );
  OR2_X1 U19892 ( .A1(n18905), .A2(n16737), .ZN(n16672) );
  NOR2_X1 U19893 ( .A1(n17034), .A2(n16672), .ZN(n16730) );
  NAND3_X1 U19894 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16730), .A3(
        P3_REIP_REG_27__SCAN_IN), .ZN(n16715) );
  NOR2_X1 U19895 ( .A1(n18912), .A2(n16715), .ZN(n16689) );
  NAND2_X1 U19896 ( .A1(n16689), .A2(n18916), .ZN(n16701) );
  NAND2_X1 U19897 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16721) );
  NOR2_X1 U19898 ( .A1(n16672), .A2(n17030), .ZN(n16716) );
  INV_X1 U19899 ( .A(n16716), .ZN(n16673) );
  NOR2_X1 U19900 ( .A1(n16721), .A2(n16673), .ZN(n16674) );
  NAND2_X1 U19901 ( .A1(n17034), .A2(n17041), .ZN(n17042) );
  AOI21_X1 U19902 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(n16674), .A(n16913), 
        .ZN(n16694) );
  INV_X1 U19903 ( .A(n16694), .ZN(n16706) );
  AOI21_X1 U19904 ( .B1(n16701), .B2(n16706), .A(n18914), .ZN(n16675) );
  AOI21_X1 U19905 ( .B1(n16696), .B2(n16676), .A(n16675), .ZN(n16692) );
  AOI21_X1 U19906 ( .B1(n16679), .B2(n17634), .A(n16677), .ZN(n16678) );
  INV_X1 U19907 ( .A(n16678), .ZN(n17648) );
  OAI21_X1 U19908 ( .B1(n9871), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16679), .ZN(n17658) );
  AOI21_X1 U19909 ( .B1(n17632), .B2(n17661), .A(n9871), .ZN(n16680) );
  INV_X1 U19910 ( .A(n16680), .ZN(n17662) );
  INV_X1 U19911 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16764) );
  NOR2_X1 U19912 ( .A1(n16683), .A2(n16764), .ZN(n16681) );
  OAI21_X1 U19913 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16681), .A(
        n17632), .ZN(n17676) );
  INV_X1 U19914 ( .A(n16683), .ZN(n16682) );
  AOI22_X1 U19915 ( .A1(n16682), .A2(n16764), .B1(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16683), .ZN(n17685) );
  NOR2_X1 U19916 ( .A1(n9966), .A2(n17701), .ZN(n17671) );
  OAI21_X1 U19917 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17671), .A(
        n16683), .ZN(n17704) );
  INV_X1 U19918 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17716) );
  NAND2_X1 U19919 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17714), .ZN(
        n16685) );
  NOR2_X1 U19920 ( .A1(n17716), .A2(n16685), .ZN(n16684) );
  OAI22_X1 U19921 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16684), .B1(
        n9966), .B2(n17701), .ZN(n17717) );
  XNOR2_X1 U19922 ( .A(n17716), .B(n16685), .ZN(n17723) );
  NAND2_X1 U19923 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17749) );
  NOR2_X1 U19924 ( .A1(n9966), .A2(n9837), .ZN(n17748) );
  INV_X1 U19925 ( .A(n17748), .ZN(n16688) );
  NOR2_X1 U19926 ( .A1(n17749), .A2(n16688), .ZN(n17712) );
  OAI21_X1 U19927 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17712), .A(
        n16685), .ZN(n17739) );
  NAND2_X1 U19928 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17748), .ZN(
        n16687) );
  AOI21_X1 U19929 ( .B1(n9961), .B2(n16687), .A(n17712), .ZN(n16686) );
  INV_X1 U19930 ( .A(n16686), .ZN(n17751) );
  OAI21_X1 U19931 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17748), .A(
        n16687), .ZN(n17760) );
  NOR2_X1 U19932 ( .A1(n9966), .A2(n17773), .ZN(n16843) );
  OAI21_X1 U19933 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16843), .A(
        n16688), .ZN(n17782) );
  INV_X1 U19934 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17790) );
  INV_X1 U19935 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20936) );
  INV_X1 U19936 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17866) );
  INV_X1 U19937 ( .A(n17901), .ZN(n17892) );
  NAND3_X1 U19938 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17892), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16947) );
  NOR2_X1 U19939 ( .A1(n16937), .A2(n16947), .ZN(n16936) );
  NAND2_X1 U19940 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16936), .ZN(
        n16924) );
  NOR2_X1 U19941 ( .A1(n17866), .A2(n16924), .ZN(n16914) );
  NAND2_X1 U19942 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16914), .ZN(
        n17825) );
  NOR2_X1 U19943 ( .A1(n17830), .A2(n17825), .ZN(n16876) );
  NAND2_X1 U19944 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16876), .ZN(
        n17787) );
  NOR2_X1 U19945 ( .A1(n20936), .A2(n17787), .ZN(n16852) );
  INV_X1 U19946 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20933) );
  NAND2_X1 U19947 ( .A1(n16852), .A2(n20933), .ZN(n16845) );
  NAND2_X1 U19948 ( .A1(n17760), .A2(n16822), .ZN(n16821) );
  NAND2_X1 U19949 ( .A1(n16879), .A2(n16821), .ZN(n16814) );
  NAND2_X1 U19950 ( .A1(n17751), .A2(n16814), .ZN(n16813) );
  NAND2_X1 U19951 ( .A1(n16879), .A2(n16813), .ZN(n16805) );
  NAND2_X1 U19952 ( .A1(n17739), .A2(n16805), .ZN(n16804) );
  NAND2_X1 U19953 ( .A1(n16879), .A2(n16804), .ZN(n16798) );
  NAND2_X1 U19954 ( .A1(n17723), .A2(n16798), .ZN(n16797) );
  NAND2_X1 U19955 ( .A1(n16879), .A2(n16797), .ZN(n16786) );
  NAND2_X1 U19956 ( .A1(n17717), .A2(n16786), .ZN(n16785) );
  NAND2_X1 U19957 ( .A1(n16879), .A2(n16785), .ZN(n16775) );
  NAND2_X1 U19958 ( .A1(n17704), .A2(n16775), .ZN(n16774) );
  NAND2_X1 U19959 ( .A1(n16879), .A2(n16774), .ZN(n16761) );
  NAND2_X1 U19960 ( .A1(n17685), .A2(n16761), .ZN(n16760) );
  NAND2_X1 U19961 ( .A1(n16879), .A2(n16760), .ZN(n16750) );
  NAND2_X1 U19962 ( .A1(n17676), .A2(n16750), .ZN(n16749) );
  NAND2_X1 U19963 ( .A1(n16879), .A2(n16749), .ZN(n16742) );
  NAND2_X1 U19964 ( .A1(n17662), .A2(n16742), .ZN(n16741) );
  NAND2_X1 U19965 ( .A1(n16879), .A2(n16741), .ZN(n16732) );
  NAND2_X1 U19966 ( .A1(n17658), .A2(n16732), .ZN(n16731) );
  NAND2_X1 U19967 ( .A1(n16879), .A2(n16731), .ZN(n16720) );
  NAND2_X1 U19968 ( .A1(n17648), .A2(n16720), .ZN(n16719) );
  NAND2_X1 U19969 ( .A1(n16865), .A2(n16719), .ZN(n16712) );
  NAND2_X1 U19970 ( .A1(n16712), .A2(n16711), .ZN(n16710) );
  NAND2_X1 U19971 ( .A1(n16865), .A2(n16710), .ZN(n16700) );
  NAND4_X1 U19972 ( .A1(n17014), .A2(n16879), .A3(n16700), .A4(n16699), .ZN(
        n16691) );
  NAND3_X1 U19973 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16689), .A3(n18914), 
        .ZN(n16690) );
  NAND4_X1 U19974 ( .A1(n16693), .A2(n16692), .A3(n16691), .A4(n16690), .ZN(
        P3_U2640) );
  AOI22_X1 U19975 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16997), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n16694), .ZN(n16704) );
  NAND2_X1 U19976 ( .A1(n16695), .A2(n17043), .ZN(n16705) );
  NOR2_X1 U19977 ( .A1(n17044), .A2(n16696), .ZN(n16697) );
  MUX2_X1 U19978 ( .A(n16705), .B(n16697), .S(P3_EBX_REG_30__SCAN_IN), .Z(
        n16703) );
  AOI21_X1 U19979 ( .B1(n16700), .B2(n16699), .A(n18839), .ZN(n16698) );
  OAI21_X1 U19980 ( .B1(n16700), .B2(n16699), .A(n16698), .ZN(n16702) );
  NAND4_X1 U19981 ( .A1(n16704), .A2(n16703), .A3(n16702), .A4(n16701), .ZN(
        P3_U2641) );
  AOI21_X1 U19982 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16717), .A(n16705), .ZN(
        n16709) );
  OAI22_X1 U19983 ( .A1(n16707), .A2(n17031), .B1(n18912), .B2(n16706), .ZN(
        n16708) );
  AOI211_X1 U19984 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17044), .A(n16709), .B(
        n16708), .ZN(n16714) );
  OAI211_X1 U19985 ( .C1(n16712), .C2(n16711), .A(n17014), .B(n16710), .ZN(
        n16713) );
  OAI211_X1 U19986 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16715), .A(n16714), 
        .B(n16713), .ZN(P3_U2642) );
  AOI22_X1 U19987 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16725) );
  NOR2_X1 U19988 ( .A1(n16913), .A2(n16716), .ZN(n16740) );
  AOI21_X1 U19989 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16726), .A(n16999), .ZN(
        n16718) );
  AOI22_X1 U19990 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16740), .B1(n16718), 
        .B2(n16717), .ZN(n16724) );
  OAI211_X1 U19991 ( .C1(n17648), .C2(n16720), .A(n17014), .B(n16719), .ZN(
        n16723) );
  OAI211_X1 U19992 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16730), .B(n16721), .ZN(n16722) );
  NAND4_X1 U19993 ( .A1(n16725), .A2(n16724), .A3(n16723), .A4(n16722), .ZN(
        P3_U2643) );
  OAI21_X1 U19994 ( .B1(n16727), .B2(n16728), .A(n16726), .ZN(n16735) );
  INV_X1 U19995 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18906) );
  OAI22_X1 U19996 ( .A1(n9967), .A2(n17031), .B1(n17033), .B2(n16728), .ZN(
        n16729) );
  AOI221_X1 U19997 ( .B1(n16730), .B2(n18906), .C1(n16740), .C2(
        P3_REIP_REG_27__SCAN_IN), .A(n16729), .ZN(n16734) );
  OAI211_X1 U19998 ( .C1(n17658), .C2(n16732), .A(n17014), .B(n16731), .ZN(
        n16733) );
  OAI211_X1 U19999 ( .C1(n16735), .C2(n16999), .A(n16734), .B(n16733), .ZN(
        P3_U2644) );
  OAI21_X1 U20000 ( .B1(n16747), .B2(n20956), .A(n16736), .ZN(n16745) );
  NOR2_X1 U20001 ( .A1(n17034), .A2(n16737), .ZN(n16739) );
  OAI22_X1 U20002 ( .A1(n17661), .A2(n17031), .B1(n17033), .B2(n20956), .ZN(
        n16738) );
  AOI221_X1 U20003 ( .B1(n16740), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n16739), 
        .C2(n18905), .A(n16738), .ZN(n16744) );
  OAI211_X1 U20004 ( .C1(n17662), .C2(n16742), .A(n17014), .B(n16741), .ZN(
        n16743) );
  OAI211_X1 U20005 ( .C1(n16745), .C2(n16999), .A(n16744), .B(n16743), .ZN(
        P3_U2645) );
  AOI22_X1 U20006 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16755) );
  NOR2_X1 U20007 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17034), .ZN(n16758) );
  NAND2_X1 U20008 ( .A1(n17024), .A2(n16746), .ZN(n16770) );
  NAND2_X1 U20009 ( .A1(n17041), .A2(n16770), .ZN(n16768) );
  AOI211_X1 U20010 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16756), .A(n16747), .B(
        n16999), .ZN(n16748) );
  AOI221_X1 U20011 ( .B1(n16758), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16768), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16748), .ZN(n16754) );
  OAI211_X1 U20012 ( .C1(n17676), .C2(n16750), .A(n17014), .B(n16749), .ZN(
        n16753) );
  INV_X1 U20013 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18902) );
  NAND3_X1 U20014 ( .A1(n17024), .A2(n16751), .A3(n18902), .ZN(n16752) );
  NAND4_X1 U20015 ( .A1(n16755), .A2(n16754), .A3(n16753), .A4(n16752), .ZN(
        P3_U2646) );
  OAI21_X1 U20016 ( .B1(n16769), .B2(n16757), .A(n16756), .ZN(n16767) );
  AOI22_X1 U20017 ( .A1(n17044), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16759), 
        .B2(n16758), .ZN(n16763) );
  OAI211_X1 U20018 ( .C1(n17685), .C2(n16761), .A(n17014), .B(n16760), .ZN(
        n16762) );
  OAI211_X1 U20019 ( .C1(n17031), .C2(n16764), .A(n16763), .B(n16762), .ZN(
        n16765) );
  AOI21_X1 U20020 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16768), .A(n16765), 
        .ZN(n16766) );
  OAI21_X1 U20021 ( .B1(n16999), .B2(n16767), .A(n16766), .ZN(P3_U2647) );
  INV_X1 U20022 ( .A(n16768), .ZN(n16778) );
  AOI211_X1 U20023 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16787), .A(n16769), .B(
        n16999), .ZN(n16773) );
  OAI22_X1 U20024 ( .A1(n17702), .A2(n17031), .B1(n16771), .B2(n16770), .ZN(
        n16772) );
  AOI211_X1 U20025 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n17044), .A(n16773), .B(
        n16772), .ZN(n16777) );
  OAI211_X1 U20026 ( .C1(n17704), .C2(n16775), .A(n17014), .B(n16774), .ZN(
        n16776) );
  OAI211_X1 U20027 ( .C1(n16778), .C2(n18898), .A(n16777), .B(n16776), .ZN(
        P3_U2648) );
  AOI22_X1 U20028 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16792) );
  INV_X1 U20029 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18893) );
  NAND2_X1 U20030 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16812) );
  NOR2_X1 U20031 ( .A1(n18893), .A2(n16812), .ZN(n16782) );
  AOI21_X1 U20032 ( .B1(n16779), .B2(n17024), .A(n17030), .ZN(n16863) );
  OAI21_X1 U20033 ( .B1(n17034), .B2(n16780), .A(n16863), .ZN(n16781) );
  INV_X1 U20034 ( .A(n16781), .ZN(n16834) );
  OAI21_X1 U20035 ( .B1(n16782), .B2(n16913), .A(n16834), .ZN(n16803) );
  INV_X1 U20036 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18896) );
  INV_X1 U20037 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18894) );
  NAND3_X1 U20038 ( .A1(n17024), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16862), 
        .ZN(n16861) );
  AOI211_X1 U20039 ( .C1(n18896), .C2(n18894), .A(n16793), .B(n16861), .ZN(
        n16784) );
  AOI22_X1 U20040 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16803), .B1(n16784), 
        .B2(n16783), .ZN(n16791) );
  OAI211_X1 U20041 ( .C1(n17717), .C2(n16786), .A(n17014), .B(n16785), .ZN(
        n16790) );
  OAI211_X1 U20042 ( .C1(n16794), .C2(n16788), .A(n17043), .B(n16787), .ZN(
        n16789) );
  NAND4_X1 U20043 ( .A1(n16792), .A2(n16791), .A3(n16790), .A4(n16789), .ZN(
        P3_U2649) );
  OR2_X1 U20044 ( .A1(n16793), .A2(n16861), .ZN(n16801) );
  AOI211_X1 U20045 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16806), .A(n16794), .B(
        n16999), .ZN(n16796) );
  INV_X1 U20046 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17135) );
  OAI22_X1 U20047 ( .A1(n17716), .A2(n17031), .B1(n17033), .B2(n17135), .ZN(
        n16795) );
  AOI211_X1 U20048 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16803), .A(n16796), 
        .B(n16795), .ZN(n16800) );
  OAI211_X1 U20049 ( .C1(n17723), .C2(n16798), .A(n17014), .B(n16797), .ZN(
        n16799) );
  OAI211_X1 U20050 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16801), .A(n16800), 
        .B(n16799), .ZN(P3_U2650) );
  AOI22_X1 U20051 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16810) );
  NOR3_X1 U20052 ( .A1(n18889), .A2(n16839), .A3(n16861), .ZN(n16820) );
  NOR2_X1 U20053 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16812), .ZN(n16802) );
  AOI22_X1 U20054 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16803), .B1(n16820), 
        .B2(n16802), .ZN(n16809) );
  OAI211_X1 U20055 ( .C1(n17739), .C2(n16805), .A(n17014), .B(n16804), .ZN(
        n16808) );
  OAI211_X1 U20056 ( .C1(n16811), .C2(n17152), .A(n17043), .B(n16806), .ZN(
        n16807) );
  NAND4_X1 U20057 ( .A1(n16810), .A2(n16809), .A3(n16808), .A4(n16807), .ZN(
        P3_U2651) );
  AOI211_X1 U20058 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16823), .A(n16811), .B(
        n16999), .ZN(n16819) );
  OAI22_X1 U20059 ( .A1(n9961), .A2(n17031), .B1(n17033), .B2(n17154), .ZN(
        n16818) );
  INV_X1 U20060 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20867) );
  OAI211_X1 U20061 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16820), .B(n16812), .ZN(n16816) );
  OAI211_X1 U20062 ( .C1(n17751), .C2(n16814), .A(n17014), .B(n16813), .ZN(
        n16815) );
  OAI211_X1 U20063 ( .C1(n16834), .C2(n20867), .A(n16816), .B(n16815), .ZN(
        n16817) );
  OR4_X1 U20064 ( .A1(n18301), .A2(n16819), .A3(n16818), .A4(n16817), .ZN(
        P3_U2652) );
  INV_X1 U20065 ( .A(n16820), .ZN(n16828) );
  INV_X1 U20066 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20989) );
  AOI22_X1 U20067 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16826) );
  OAI211_X1 U20068 ( .C1(n17760), .C2(n16822), .A(n17014), .B(n16821), .ZN(
        n16825) );
  OAI211_X1 U20069 ( .C1(n16829), .C2(n20985), .A(n17043), .B(n16823), .ZN(
        n16824) );
  AND4_X1 U20070 ( .A1(n16826), .A2(n18199), .A3(n16825), .A4(n16824), .ZN(
        n16827) );
  OAI221_X1 U20071 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16828), .C1(n20989), 
        .C2(n16834), .A(n16827), .ZN(P3_U2653) );
  AOI211_X1 U20072 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16840), .A(n16829), .B(
        n16999), .ZN(n16838) );
  AOI22_X1 U20073 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16830) );
  INV_X1 U20074 ( .A(n16830), .ZN(n16837) );
  OR2_X1 U20075 ( .A1(n16839), .A2(n16861), .ZN(n16835) );
  OAI211_X1 U20076 ( .C1(n17782), .C2(n16832), .A(n17014), .B(n16831), .ZN(
        n16833) );
  OAI221_X1 U20077 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16835), .C1(n18889), 
        .C2(n16834), .A(n16833), .ZN(n16836) );
  OR4_X1 U20078 ( .A1(n18301), .A2(n16838), .A3(n16837), .A4(n16836), .ZN(
        P3_U2654) );
  OAI21_X1 U20079 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), 
        .A(n16839), .ZN(n16851) );
  OAI211_X1 U20080 ( .C1(n16855), .C2(n17218), .A(n17043), .B(n16840), .ZN(
        n16841) );
  OAI211_X1 U20081 ( .C1(n17033), .C2(n17218), .A(n18199), .B(n16841), .ZN(
        n16842) );
  AOI21_X1 U20082 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16997), .A(
        n16842), .ZN(n16850) );
  INV_X1 U20083 ( .A(n16852), .ZN(n16844) );
  AOI21_X1 U20084 ( .B1(n17790), .B2(n16844), .A(n16843), .ZN(n17788) );
  NAND2_X1 U20085 ( .A1(n16865), .A2(n16845), .ZN(n16846) );
  XNOR2_X1 U20086 ( .A(n17788), .B(n16846), .ZN(n16848) );
  INV_X1 U20087 ( .A(n16863), .ZN(n16847) );
  AOI22_X1 U20088 ( .A1(n17014), .A2(n16848), .B1(P3_REIP_REG_16__SCAN_IN), 
        .B2(n16847), .ZN(n16849) );
  OAI211_X1 U20089 ( .C1(n16861), .C2(n16851), .A(n16850), .B(n16849), .ZN(
        P3_U2655) );
  INV_X1 U20090 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18884) );
  AOI21_X1 U20091 ( .B1(n20936), .B2(n17787), .A(n16852), .ZN(n17802) );
  OAI21_X1 U20092 ( .B1(n17787), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16879), .ZN(n16867) );
  INV_X1 U20093 ( .A(n16867), .ZN(n16854) );
  OAI21_X1 U20094 ( .B1(n17802), .B2(n16854), .A(n17014), .ZN(n16853) );
  AOI21_X1 U20095 ( .B1(n17802), .B2(n16854), .A(n16853), .ZN(n16859) );
  AOI211_X1 U20096 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16868), .A(n16855), .B(
        n16999), .ZN(n16858) );
  OAI22_X1 U20097 ( .A1(n20936), .A2(n17031), .B1(n17033), .B2(n16856), .ZN(
        n16857) );
  NOR4_X1 U20098 ( .A1(n18301), .A2(n16859), .A3(n16858), .A4(n16857), .ZN(
        n16860) );
  OAI221_X1 U20099 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16861), .C1(n18884), 
        .C2(n16863), .A(n16860), .ZN(P3_U2656) );
  INV_X1 U20100 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18883) );
  NAND2_X1 U20101 ( .A1(n17024), .A2(n16862), .ZN(n16864) );
  AOI21_X1 U20102 ( .B1(n18883), .B2(n16864), .A(n16863), .ZN(n16872) );
  OAI21_X1 U20103 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16876), .A(
        n17787), .ZN(n17824) );
  NAND2_X1 U20104 ( .A1(n17014), .A2(n9729), .ZN(n17012) );
  NOR3_X1 U20105 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17830), .A3(
        n17825), .ZN(n16881) );
  OAI21_X1 U20106 ( .B1(n16881), .B2(n17824), .A(n17014), .ZN(n16866) );
  AOI22_X1 U20107 ( .A1(n17824), .A2(n16867), .B1(n17012), .B2(n16866), .ZN(
        n16871) );
  OAI211_X1 U20108 ( .C1(n16874), .C2(n17250), .A(n17043), .B(n16868), .ZN(
        n16869) );
  OAI21_X1 U20109 ( .B1(n17031), .B2(n17810), .A(n16869), .ZN(n16870) );
  NOR3_X1 U20110 ( .A1(n16872), .A2(n16871), .A3(n16870), .ZN(n16873) );
  OAI211_X1 U20111 ( .C1(n17033), .C2(n17250), .A(n16873), .B(n18199), .ZN(
        P3_U2657) );
  INV_X1 U20112 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16890) );
  AOI211_X1 U20113 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16893), .A(n16874), .B(
        n16999), .ZN(n16875) );
  AOI211_X1 U20114 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16997), .A(
        n18301), .B(n16875), .ZN(n16889) );
  INV_X1 U20115 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17846) );
  NOR2_X1 U20116 ( .A1(n17846), .A2(n17825), .ZN(n16878) );
  INV_X1 U20117 ( .A(n16876), .ZN(n16877) );
  OAI21_X1 U20118 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16878), .A(
        n16877), .ZN(n17833) );
  OAI21_X1 U20119 ( .B1(n9729), .B2(n20933), .A(n17014), .ZN(n16965) );
  AOI211_X1 U20120 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16879), .A(
        n17833), .B(n16965), .ZN(n16887) );
  INV_X1 U20121 ( .A(n16880), .ZN(n16896) );
  AOI21_X1 U20122 ( .B1(n17024), .B2(n16896), .A(n17030), .ZN(n16902) );
  INV_X1 U20123 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18878) );
  NAND2_X1 U20124 ( .A1(n17024), .A2(n18878), .ZN(n16895) );
  AOI21_X1 U20125 ( .B1(n16902), .B2(n16895), .A(n18880), .ZN(n16886) );
  INV_X1 U20126 ( .A(n17833), .ZN(n16882) );
  NAND2_X1 U20127 ( .A1(n16879), .A2(n17014), .ZN(n17032) );
  NOR3_X1 U20128 ( .A1(n16882), .A2(n16881), .A3(n17032), .ZN(n16885) );
  NOR3_X1 U20129 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17034), .A3(n16883), 
        .ZN(n16884) );
  NOR4_X1 U20130 ( .A1(n16887), .A2(n16886), .A3(n16885), .A4(n16884), .ZN(
        n16888) );
  OAI211_X1 U20131 ( .C1(n17033), .C2(n16890), .A(n16889), .B(n16888), .ZN(
        P3_U2658) );
  AOI22_X1 U20132 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16900) );
  INV_X1 U20133 ( .A(n17825), .ZN(n16891) );
  AOI22_X1 U20134 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17825), .B1(
        n16891), .B2(n17846), .ZN(n17842) );
  AOI21_X1 U20135 ( .B1(n16891), .B2(n20933), .A(n9729), .ZN(n16892) );
  XNOR2_X1 U20136 ( .A(n17842), .B(n16892), .ZN(n16898) );
  OAI211_X1 U20137 ( .C1(n16904), .C2(n17267), .A(n17043), .B(n16893), .ZN(
        n16894) );
  OAI211_X1 U20138 ( .C1(n16896), .C2(n16895), .A(n18199), .B(n16894), .ZN(
        n16897) );
  AOI21_X1 U20139 ( .B1(n16898), .B2(n17014), .A(n16897), .ZN(n16899) );
  OAI211_X1 U20140 ( .C1(n18878), .C2(n16902), .A(n16900), .B(n16899), .ZN(
        P3_U2659) );
  AOI21_X1 U20141 ( .B1(n16914), .B2(n20933), .A(n9729), .ZN(n16901) );
  OAI21_X1 U20142 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16914), .A(
        n17825), .ZN(n17855) );
  XOR2_X1 U20143 ( .A(n16901), .B(n17855), .Z(n16909) );
  AOI21_X1 U20144 ( .B1(n17044), .B2(P3_EBX_REG_11__SCAN_IN), .A(n18301), .ZN(
        n16908) );
  INV_X1 U20145 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18862) );
  NAND2_X1 U20146 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n17023) );
  NOR2_X1 U20147 ( .A1(n17034), .A2(n17023), .ZN(n17006) );
  NAND2_X1 U20148 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17006), .ZN(n16996) );
  NOR2_X1 U20149 ( .A1(n18862), .A2(n16996), .ZN(n16973) );
  NAND2_X1 U20150 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16973), .ZN(n16971) );
  AOI221_X1 U20151 ( .B1(n16903), .B2(n18876), .C1(n16971), .C2(n18876), .A(
        n16902), .ZN(n16906) );
  AOI211_X1 U20152 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16920), .A(n16904), .B(
        n16999), .ZN(n16905) );
  AOI211_X1 U20153 ( .C1(n16997), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16906), .B(n16905), .ZN(n16907) );
  OAI211_X1 U20154 ( .C1(n18839), .C2(n16909), .A(n16908), .B(n16907), .ZN(
        P3_U2660) );
  AOI22_X1 U20155 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16923) );
  INV_X1 U20156 ( .A(n16910), .ZN(n16911) );
  OAI21_X1 U20157 ( .B1(n16911), .B2(n17034), .A(n17041), .ZN(n17005) );
  AOI21_X1 U20158 ( .B1(n17024), .B2(n16912), .A(n17005), .ZN(n16978) );
  OAI21_X1 U20159 ( .B1(n16917), .B2(n16913), .A(n16978), .ZN(n16941) );
  AOI21_X1 U20160 ( .B1(n17866), .B2(n16924), .A(n16914), .ZN(n17869) );
  OAI21_X1 U20161 ( .B1(n16924), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16879), .ZN(n16927) );
  INV_X1 U20162 ( .A(n16927), .ZN(n16916) );
  OAI21_X1 U20163 ( .B1(n17869), .B2(n16916), .A(n17014), .ZN(n16915) );
  AOI21_X1 U20164 ( .B1(n17869), .B2(n16916), .A(n16915), .ZN(n16919) );
  INV_X1 U20165 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18874) );
  INV_X1 U20166 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18872) );
  INV_X1 U20167 ( .A(n16971), .ZN(n16956) );
  NAND2_X1 U20168 ( .A1(n16917), .A2(n16956), .ZN(n16935) );
  AOI221_X1 U20169 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n18874), .C2(n18872), .A(n16935), .ZN(n16918) );
  AOI211_X1 U20170 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16941), .A(n16919), 
        .B(n16918), .ZN(n16922) );
  OAI211_X1 U20171 ( .C1(n16928), .C2(n20934), .A(n17043), .B(n16920), .ZN(
        n16921) );
  NAND4_X1 U20172 ( .A1(n16923), .A2(n16922), .A3(n18199), .A4(n16921), .ZN(
        P3_U2661) );
  INV_X1 U20173 ( .A(n16941), .ZN(n16934) );
  OAI21_X1 U20174 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16936), .A(
        n16924), .ZN(n17883) );
  NOR2_X1 U20175 ( .A1(n9966), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17016) );
  INV_X1 U20176 ( .A(n17016), .ZN(n16988) );
  NOR2_X1 U20177 ( .A1(n17901), .A2(n16988), .ZN(n16948) );
  OAI221_X1 U20178 ( .B1(n17883), .B2(n16925), .C1(n17883), .C2(n16948), .A(
        n17014), .ZN(n16926) );
  AOI22_X1 U20179 ( .A1(n16927), .A2(n17883), .B1(n17012), .B2(n16926), .ZN(
        n16932) );
  AOI211_X1 U20180 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16939), .A(n16928), .B(
        n16999), .ZN(n16931) );
  AOI22_X1 U20181 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n16929) );
  INV_X1 U20182 ( .A(n16929), .ZN(n16930) );
  NOR4_X1 U20183 ( .A1(n18301), .A2(n16932), .A3(n16931), .A4(n16930), .ZN(
        n16933) );
  OAI221_X1 U20184 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16935), .C1(n18872), 
        .C2(n16934), .A(n16933), .ZN(P3_U2662) );
  OAI21_X1 U20185 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16947), .A(
        n16865), .ZN(n16938) );
  AOI21_X1 U20186 ( .B1(n16937), .B2(n16947), .A(n16936), .ZN(n17893) );
  XOR2_X1 U20187 ( .A(n16938), .B(n17893), .Z(n16946) );
  OAI211_X1 U20188 ( .C1(n16951), .C2(n17248), .A(n17043), .B(n16939), .ZN(
        n16940) );
  OAI211_X1 U20189 ( .C1(n17033), .C2(n17248), .A(n18199), .B(n16940), .ZN(
        n16944) );
  NOR2_X1 U20190 ( .A1(n16955), .A2(n16971), .ZN(n16942) );
  MUX2_X1 U20191 ( .A(n16942), .B(n16941), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n16943) );
  AOI211_X1 U20192 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n16997), .A(
        n16944), .B(n16943), .ZN(n16945) );
  OAI21_X1 U20193 ( .B1(n16946), .B2(n18839), .A(n16945), .ZN(P3_U2663) );
  INV_X1 U20194 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18868) );
  NOR2_X1 U20195 ( .A1(n9966), .A2(n17901), .ZN(n16959) );
  OAI21_X1 U20196 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16959), .A(
        n16947), .ZN(n17920) );
  INV_X1 U20197 ( .A(n17920), .ZN(n16950) );
  NOR2_X1 U20198 ( .A1(n16948), .A2(n9729), .ZN(n16961) );
  INV_X1 U20199 ( .A(n16961), .ZN(n16949) );
  AOI221_X1 U20200 ( .B1(n16950), .B2(n16961), .C1(n17920), .C2(n16949), .A(
        n18839), .ZN(n16954) );
  AOI211_X1 U20201 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16962), .A(n16951), .B(
        n16999), .ZN(n16953) );
  INV_X1 U20202 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17342) );
  OAI22_X1 U20203 ( .A1(n17909), .A2(n17031), .B1(n17033), .B2(n17342), .ZN(
        n16952) );
  NOR4_X1 U20204 ( .A1(n18301), .A2(n16954), .A3(n16953), .A4(n16952), .ZN(
        n16958) );
  OAI211_X1 U20205 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16956), .B(n16955), .ZN(n16957) );
  OAI211_X1 U20206 ( .C1(n16978), .C2(n18868), .A(n16958), .B(n16957), .ZN(
        P3_U2664) );
  INV_X1 U20207 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18866) );
  INV_X1 U20208 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16960) );
  NAND2_X1 U20209 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17928), .ZN(
        n16974) );
  AOI21_X1 U20210 ( .B1(n16960), .B2(n16974), .A(n16959), .ZN(n17929) );
  NAND2_X1 U20211 ( .A1(n17014), .A2(n16961), .ZN(n16964) );
  OAI211_X1 U20212 ( .C1(n16972), .C2(n17343), .A(n17043), .B(n16962), .ZN(
        n16963) );
  OAI211_X1 U20213 ( .C1(n17929), .C2(n16964), .A(n18199), .B(n16963), .ZN(
        n16969) );
  INV_X1 U20214 ( .A(n16974), .ZN(n16966) );
  INV_X1 U20215 ( .A(n16965), .ZN(n17037) );
  OAI211_X1 U20216 ( .C1(n16966), .C2(n9729), .A(n17929), .B(n17037), .ZN(
        n16967) );
  OAI21_X1 U20217 ( .B1(n17343), .B2(n17033), .A(n16967), .ZN(n16968) );
  AOI211_X1 U20218 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16997), .A(
        n16969), .B(n16968), .ZN(n16970) );
  OAI221_X1 U20219 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16971), .C1(n18866), 
        .C2(n16978), .A(n16970), .ZN(P3_U2665) );
  INV_X1 U20220 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16982) );
  AOI211_X1 U20221 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16984), .A(n16972), .B(
        n16999), .ZN(n16980) );
  NOR2_X1 U20222 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16973), .ZN(n16977) );
  NOR2_X1 U20223 ( .A1(n9966), .A2(n17940), .ZN(n16983) );
  OAI21_X1 U20224 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16983), .A(
        n16974), .ZN(n16975) );
  INV_X1 U20225 ( .A(n16975), .ZN(n17942) );
  OAI21_X1 U20226 ( .B1(n17940), .B2(n16988), .A(n16879), .ZN(n16989) );
  XOR2_X1 U20227 ( .A(n17942), .B(n16989), .Z(n16976) );
  OAI22_X1 U20228 ( .A1(n16978), .A2(n16977), .B1(n18839), .B2(n16976), .ZN(
        n16979) );
  AOI211_X1 U20229 ( .C1(n16997), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16980), .B(n16979), .ZN(n16981) );
  OAI211_X1 U20230 ( .C1(n17033), .C2(n16982), .A(n16981), .B(n18199), .ZN(
        P3_U2666) );
  INV_X1 U20231 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16987) );
  NAND2_X1 U20232 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9964), .ZN(
        n16998) );
  AOI21_X1 U20233 ( .B1(n16987), .B2(n16998), .A(n16983), .ZN(n16990) );
  INV_X1 U20234 ( .A(n16990), .ZN(n17959) );
  OAI211_X1 U20235 ( .C1(n17002), .C2(n17351), .A(n17043), .B(n16984), .ZN(
        n16985) );
  OAI21_X1 U20236 ( .B1(n17012), .B2(n17959), .A(n16985), .ZN(n16986) );
  AOI21_X1 U20237 ( .B1(n17044), .B2(P3_EBX_REG_4__SCAN_IN), .A(n16986), .ZN(
        n16995) );
  NAND2_X1 U20238 ( .A1(n9964), .A2(n16987), .ZN(n17951) );
  OAI22_X1 U20239 ( .A1(n16990), .A2(n16989), .B1(n16988), .B2(n17951), .ZN(
        n16993) );
  NAND2_X1 U20240 ( .A1(n18319), .A2(n18989), .ZN(n17040) );
  AOI22_X1 U20241 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16997), .B1(
        P3_REIP_REG_4__SCAN_IN), .B2(n17005), .ZN(n16991) );
  OAI221_X1 U20242 ( .B1(n17040), .B2(n10256), .C1(n17040), .C2(n18777), .A(
        n16991), .ZN(n16992) );
  AOI211_X1 U20243 ( .C1(n17014), .C2(n16993), .A(n18301), .B(n16992), .ZN(
        n16994) );
  OAI211_X1 U20244 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16996), .A(n16995), .B(
        n16994), .ZN(P3_U2667) );
  AOI22_X1 U20245 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16997), .B1(
        n17044), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n17009) );
  INV_X1 U20246 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17020) );
  NOR2_X1 U20247 ( .A1(n9966), .A2(n17020), .ZN(n17011) );
  OAI21_X1 U20248 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17011), .A(
        n16998), .ZN(n17974) );
  AOI21_X1 U20249 ( .B1(n17011), .B2(n20933), .A(n9729), .ZN(n17013) );
  XNOR2_X1 U20250 ( .A(n17974), .B(n17013), .ZN(n17004) );
  AOI21_X1 U20251 ( .B1(n17017), .B2(P3_EBX_REG_3__SCAN_IN), .A(n16999), .ZN(
        n17000) );
  INV_X1 U20252 ( .A(n17000), .ZN(n17001) );
  NOR2_X1 U20253 ( .A1(n18951), .A2(n18944), .ZN(n18790) );
  NAND2_X1 U20254 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18790), .ZN(
        n18787) );
  AOI21_X1 U20255 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18787), .A(
        n17205), .ZN(n18928) );
  OAI22_X1 U20256 ( .A1(n17002), .A2(n17001), .B1(n18928), .B2(n17040), .ZN(
        n17003) );
  AOI21_X1 U20257 ( .B1(n17004), .B2(n17014), .A(n17003), .ZN(n17008) );
  OAI21_X1 U20258 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n17006), .A(n17005), .ZN(
        n17007) );
  NAND3_X1 U20259 ( .A1(n17009), .A2(n17008), .A3(n17007), .ZN(P3_U2668) );
  INV_X1 U20260 ( .A(n18787), .ZN(n17010) );
  AOI21_X1 U20261 ( .B1(n18944), .B2(n18795), .A(n17010), .ZN(n18940) );
  INV_X1 U20262 ( .A(n17040), .ZN(n18991) );
  INV_X1 U20263 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20859) );
  AOI21_X1 U20264 ( .B1(n9966), .B2(n17020), .A(n17011), .ZN(n17979) );
  INV_X1 U20265 ( .A(n17979), .ZN(n17015) );
  OAI22_X1 U20266 ( .A1(n20859), .A2(n17041), .B1(n17015), .B2(n17012), .ZN(
        n17022) );
  OAI211_X1 U20267 ( .C1(n17016), .C2(n17015), .A(n17014), .B(n17013), .ZN(
        n17019) );
  OAI211_X1 U20268 ( .C1(n17029), .C2(n20977), .A(n17043), .B(n17017), .ZN(
        n17018) );
  OAI211_X1 U20269 ( .C1(n17031), .C2(n17020), .A(n17019), .B(n17018), .ZN(
        n17021) );
  AOI211_X1 U20270 ( .C1(n18940), .C2(n18991), .A(n17022), .B(n17021), .ZN(
        n17026) );
  OAI211_X1 U20271 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n17024), .B(n17023), .ZN(n17025) );
  OAI211_X1 U20272 ( .C1(n20977), .C2(n17033), .A(n17026), .B(n17025), .ZN(
        P3_U2669) );
  NAND2_X1 U20273 ( .A1(n17027), .A2(n18795), .ZN(n18945) );
  INV_X1 U20274 ( .A(n17028), .ZN(n17358) );
  NOR2_X1 U20275 ( .A1(n17029), .A2(n17358), .ZN(n17361) );
  AOI22_X1 U20276 ( .A1(n17043), .A2(n17361), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n17030), .ZN(n17039) );
  OAI21_X1 U20277 ( .B1(n20933), .B2(n17032), .A(n17031), .ZN(n17036) );
  INV_X1 U20278 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17363) );
  OAI22_X1 U20279 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17034), .B1(n17033), 
        .B2(n17363), .ZN(n17035) );
  AOI221_X1 U20280 ( .B1(n17037), .B2(n9966), .C1(n17036), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17035), .ZN(n17038) );
  OAI211_X1 U20281 ( .C1(n18945), .C2(n17040), .A(n17039), .B(n17038), .ZN(
        P3_U2670) );
  NAND2_X1 U20282 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17041), .ZN(
        n17047) );
  AOI22_X1 U20283 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17042), .B1(n18991), 
        .B2(n20969), .ZN(n17046) );
  OAI21_X1 U20284 ( .B1(n17044), .B2(n17043), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17045) );
  OAI211_X1 U20285 ( .C1(n18987), .C2(n17047), .A(n17046), .B(n17045), .ZN(
        P3_U2671) );
  INV_X1 U20286 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17050) );
  AND4_X1 U20287 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17048)
         );
  NAND4_X1 U20288 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n17049), .A4(n17048), .ZN(n17080) );
  NAND2_X1 U20289 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17169), .ZN(n17134) );
  NOR3_X1 U20290 ( .A1(n17050), .A2(n17080), .A3(n17134), .ZN(n17075) );
  NAND2_X1 U20291 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17075), .ZN(n17074) );
  INV_X1 U20292 ( .A(n17074), .ZN(n17051) );
  OAI33_X1 U20293 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17074), .A3(n17456), 
        .B1(n17052), .B2(n17366), .B3(n17051), .ZN(P3_U2672) );
  AOI22_X1 U20294 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20295 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20296 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17060) );
  INV_X1 U20297 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21018) );
  OAI22_X1 U20298 ( .A1(n17334), .A2(n17111), .B1(n10256), .B2(n21018), .ZN(
        n17058) );
  AOI22_X1 U20299 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20300 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20301 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17054) );
  NAND2_X1 U20302 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n17053) );
  NAND4_X1 U20303 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        n17057) );
  AOI211_X1 U20304 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17058), .B(n17057), .ZN(n17059) );
  NAND4_X1 U20305 ( .A1(n17062), .A2(n17061), .A3(n17060), .A4(n17059), .ZN(
        n17078) );
  NAND2_X1 U20306 ( .A1(n17079), .A2(n17078), .ZN(n17077) );
  AOI22_X1 U20307 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17202), .ZN(n17072) );
  AOI22_X1 U20308 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17270), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20309 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17326), .ZN(n17063) );
  OAI211_X1 U20310 ( .C1(n18670), .C2(n17275), .A(n17064), .B(n17063), .ZN(
        n17070) );
  AOI22_X1 U20311 ( .A1(n10330), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17290), .ZN(n17068) );
  AOI22_X1 U20312 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17306), .ZN(n17067) );
  AOI22_X1 U20313 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17066) );
  NAND2_X1 U20314 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17313), .ZN(
        n17065) );
  NAND4_X1 U20315 ( .A1(n17068), .A2(n17067), .A3(n17066), .A4(n17065), .ZN(
        n17069) );
  AOI211_X1 U20316 ( .C1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n10289), .A(
        n17070), .B(n17069), .ZN(n17071) );
  OAI211_X1 U20317 ( .C1(n15789), .C2(n18365), .A(n17072), .B(n17071), .ZN(
        n17073) );
  XOR2_X1 U20318 ( .A(n17077), .B(n17073), .Z(n17382) );
  OAI211_X1 U20319 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17075), .A(n17074), .B(
        n17355), .ZN(n17076) );
  OAI21_X1 U20320 ( .B1(n17382), .B2(n17355), .A(n17076), .ZN(P3_U2673) );
  OAI21_X1 U20321 ( .B1(n17079), .B2(n17078), .A(n17077), .ZN(n17386) );
  NOR2_X1 U20322 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17080), .ZN(n17081) );
  AOI22_X1 U20323 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17082), .B1(n17136), 
        .B2(n17081), .ZN(n17083) );
  OAI21_X1 U20324 ( .B1(n17386), .B2(n17355), .A(n17083), .ZN(P3_U2674) );
  OAI21_X1 U20325 ( .B1(n17088), .B2(n17085), .A(n17084), .ZN(n17395) );
  NAND3_X1 U20326 ( .A1(n17087), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17355), 
        .ZN(n17086) );
  OAI221_X1 U20327 ( .B1(n17087), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17355), 
        .C2(n17395), .A(n17086), .ZN(P3_U2676) );
  AOI21_X1 U20328 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17355), .A(n17096), .ZN(
        n17091) );
  AOI21_X1 U20329 ( .B1(n17089), .B2(n17093), .A(n17088), .ZN(n17396) );
  INV_X1 U20330 ( .A(n17396), .ZN(n17090) );
  OAI22_X1 U20331 ( .A1(n17092), .A2(n17091), .B1(n17090), .B2(n17355), .ZN(
        P3_U2677) );
  AOI21_X1 U20332 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17355), .A(n17102), .ZN(
        n17095) );
  OAI21_X1 U20333 ( .B1(n17098), .B2(n17094), .A(n17093), .ZN(n17405) );
  OAI22_X1 U20334 ( .A1(n17096), .A2(n17095), .B1(n17405), .B2(n17355), .ZN(
        P3_U2678) );
  INV_X1 U20335 ( .A(n17097), .ZN(n17108) );
  AOI21_X1 U20336 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17355), .A(n17108), .ZN(
        n17101) );
  AOI21_X1 U20337 ( .B1(n17099), .B2(n17104), .A(n17098), .ZN(n17406) );
  INV_X1 U20338 ( .A(n17406), .ZN(n17100) );
  OAI22_X1 U20339 ( .A1(n17102), .A2(n17101), .B1(n17355), .B2(n17100), .ZN(
        P3_U2679) );
  AOI21_X1 U20340 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17355), .A(n17103), .ZN(
        n17107) );
  OAI21_X1 U20341 ( .B1(n17106), .B2(n17105), .A(n17104), .ZN(n17415) );
  OAI22_X1 U20342 ( .A1(n17108), .A2(n17107), .B1(n17355), .B2(n17415), .ZN(
        P3_U2680) );
  AOI22_X1 U20343 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20344 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20345 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17109) );
  OAI211_X1 U20346 ( .C1(n10404), .C2(n17111), .A(n17110), .B(n17109), .ZN(
        n17117) );
  AOI22_X1 U20347 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20348 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10329), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20349 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17113) );
  NAND2_X1 U20350 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n17112) );
  NAND4_X1 U20351 ( .A1(n17115), .A2(n17114), .A3(n17113), .A4(n17112), .ZN(
        n17116) );
  AOI211_X1 U20352 ( .C1(n10286), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17117), .B(n17116), .ZN(n17118) );
  OAI211_X1 U20353 ( .C1(n17334), .C2(n18355), .A(n17119), .B(n17118), .ZN(
        n17417) );
  INV_X1 U20354 ( .A(n17417), .ZN(n17121) );
  NAND3_X1 U20355 ( .A1(n17122), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17355), 
        .ZN(n17120) );
  OAI221_X1 U20356 ( .B1(n17122), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17355), 
        .C2(n17121), .A(n17120), .ZN(P3_U2681) );
  OAI22_X1 U20357 ( .A1(n9814), .A2(n18584), .B1(n17334), .B2(n20925), .ZN(
        n17133) );
  AOI22_X1 U20358 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20359 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17130) );
  OAI22_X1 U20360 ( .A1(n17263), .A2(n17123), .B1(n17275), .B2(n20824), .ZN(
        n17128) );
  AOI22_X1 U20361 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20362 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20363 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17124) );
  NAND3_X1 U20364 ( .A1(n17126), .A2(n17125), .A3(n17124), .ZN(n17127) );
  AOI211_X1 U20365 ( .C1(n9734), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n17128), .B(n17127), .ZN(n17129) );
  NAND3_X1 U20366 ( .A1(n17131), .A2(n17130), .A3(n17129), .ZN(n17132) );
  AOI211_X1 U20367 ( .C1(n9726), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n17133), .B(n17132), .ZN(n17424) );
  NAND2_X1 U20368 ( .A1(n17355), .A2(n17134), .ZN(n17153) );
  INV_X1 U20369 ( .A(n17153), .ZN(n17137) );
  AOI22_X1 U20370 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17137), .B1(n17136), 
        .B2(n17135), .ZN(n17138) );
  OAI21_X1 U20371 ( .B1(n17424), .B2(n17355), .A(n17138), .ZN(P3_U2682) );
  AOI22_X1 U20372 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20373 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20374 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17205), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17139) );
  OAI211_X1 U20375 ( .C1(n10404), .C2(n17141), .A(n17140), .B(n17139), .ZN(
        n17147) );
  AOI22_X1 U20376 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20377 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20378 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17143) );
  NAND2_X1 U20379 ( .A1(n10289), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n17142) );
  NAND4_X1 U20380 ( .A1(n17145), .A2(n17144), .A3(n17143), .A4(n17142), .ZN(
        n17146) );
  AOI211_X1 U20381 ( .C1(n10286), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17147), .B(n17146), .ZN(n17148) );
  OAI211_X1 U20382 ( .C1(n17334), .C2(n18344), .A(n17149), .B(n17148), .ZN(
        n17427) );
  NAND2_X1 U20383 ( .A1(n17366), .A2(n17427), .ZN(n17150) );
  OAI221_X1 U20384 ( .B1(n17153), .B2(n17152), .C1(n17153), .C2(n17151), .A(
        n17150), .ZN(P3_U2683) );
  AOI21_X1 U20385 ( .B1(n17154), .B2(n17181), .A(n17366), .ZN(n17155) );
  INV_X1 U20386 ( .A(n17155), .ZN(n17168) );
  AOI22_X1 U20387 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17156) );
  OAI21_X1 U20388 ( .B1(n17325), .B2(n17157), .A(n17156), .ZN(n17167) );
  AOI22_X1 U20389 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17164) );
  OAI22_X1 U20390 ( .A1(n17334), .A2(n18338), .B1(n10404), .B2(n17283), .ZN(
        n17162) );
  AOI22_X1 U20391 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20392 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20393 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17158) );
  NAND3_X1 U20394 ( .A1(n17160), .A2(n17159), .A3(n17158), .ZN(n17161) );
  AOI211_X1 U20395 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17162), .B(n17161), .ZN(n17163) );
  OAI211_X1 U20396 ( .C1(n17263), .C2(n17165), .A(n17164), .B(n17163), .ZN(
        n17166) );
  AOI211_X1 U20397 ( .C1(n17205), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17167), .B(n17166), .ZN(n17437) );
  OAI22_X1 U20398 ( .A1(n17169), .A2(n17168), .B1(n17437), .B2(n17355), .ZN(
        P3_U2684) );
  AOI22_X1 U20399 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17170) );
  OAI21_X1 U20400 ( .B1(n10256), .B2(n17171), .A(n17170), .ZN(n17180) );
  AOI22_X1 U20401 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17178) );
  OAI22_X1 U20402 ( .A1(n9813), .A2(n17299), .B1(n17334), .B2(n18333), .ZN(
        n17176) );
  AOI22_X1 U20403 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20404 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20405 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17172) );
  NAND3_X1 U20406 ( .A1(n17174), .A2(n17173), .A3(n17172), .ZN(n17175) );
  AOI211_X1 U20407 ( .C1(n17202), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17176), .B(n17175), .ZN(n17177) );
  OAI211_X1 U20408 ( .C1(n15789), .C2(n18726), .A(n17178), .B(n17177), .ZN(
        n17179) );
  AOI211_X1 U20409 ( .C1(n17205), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n17180), .B(n17179), .ZN(n17441) );
  OAI21_X1 U20410 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17182), .A(n17181), .ZN(
        n17183) );
  AOI22_X1 U20411 ( .A1(n17366), .A2(n17441), .B1(n17183), .B2(n17355), .ZN(
        P3_U2685) );
  AOI22_X1 U20412 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U20413 ( .B1(n10288), .B2(n18650), .A(n17184), .ZN(n17196) );
  AOI22_X1 U20414 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17194) );
  OAI22_X1 U20415 ( .A1(n17334), .A2(n18327), .B1(n17187), .B2(n17186), .ZN(
        n17192) );
  AOI22_X1 U20416 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20417 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20418 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17188) );
  NAND3_X1 U20419 ( .A1(n17190), .A2(n17189), .A3(n17188), .ZN(n17191) );
  AOI211_X1 U20420 ( .C1(n17205), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n17192), .B(n17191), .ZN(n17193) );
  OAI211_X1 U20421 ( .C1(n9813), .C2(n21085), .A(n17194), .B(n17193), .ZN(
        n17195) );
  AOI211_X1 U20422 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n17196), .B(n17195), .ZN(n17447) );
  OAI211_X1 U20423 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17198), .A(n17349), .B(
        n17197), .ZN(n17200) );
  NAND2_X1 U20424 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17365), .ZN(n17199) );
  OAI211_X1 U20425 ( .C1(n17447), .C2(n17355), .A(n17200), .B(n17199), .ZN(
        P3_U2686) );
  AOI22_X1 U20426 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17201) );
  OAI21_X1 U20427 ( .B1(n15789), .B2(n18713), .A(n17201), .ZN(n17214) );
  AOI22_X1 U20428 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17202), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17212) );
  OAI22_X1 U20429 ( .A1(n17334), .A2(n18322), .B1(n17204), .B2(n17203), .ZN(
        n17210) );
  AOI22_X1 U20430 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20431 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U20432 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17206) );
  NAND3_X1 U20433 ( .A1(n17208), .A2(n17207), .A3(n17206), .ZN(n17209) );
  AOI211_X1 U20434 ( .C1(n17326), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17210), .B(n17209), .ZN(n17211) );
  OAI211_X1 U20435 ( .C1(n10288), .C2(n18646), .A(n17212), .B(n17211), .ZN(
        n17213) );
  AOI211_X1 U20436 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17214), .B(n17213), .ZN(n17454) );
  NOR2_X1 U20437 ( .A1(n17216), .A2(n17215), .ZN(n17232) );
  NAND2_X1 U20438 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17232), .ZN(n17231) );
  OAI21_X1 U20439 ( .B1(n17366), .B2(n17218), .A(n17231), .ZN(n17217) );
  OAI221_X1 U20440 ( .B1(n18361), .B2(n17231), .C1(n17231), .C2(n17218), .A(
        n17217), .ZN(n17219) );
  OAI21_X1 U20441 ( .B1(n17454), .B2(n17355), .A(n17219), .ZN(P3_U2687) );
  AOI22_X1 U20442 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17290), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n15818), .ZN(n17230) );
  AOI22_X1 U20443 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17326), .ZN(n17229) );
  OAI22_X1 U20444 ( .A1(n18593), .A2(n9771), .B1(n17334), .B2(n18765), .ZN(
        n17227) );
  AOI22_X1 U20445 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10327), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20446 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20447 ( .A1(n9726), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17306), .ZN(n17220) );
  OAI211_X1 U20448 ( .C1(n10404), .C2(n18365), .A(n17221), .B(n17220), .ZN(
        n17222) );
  AOI21_X1 U20449 ( .B1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n10286), .A(
        n17222), .ZN(n17223) );
  OAI211_X1 U20450 ( .C1(n15789), .C2(n17225), .A(n17224), .B(n17223), .ZN(
        n17226) );
  AOI211_X1 U20451 ( .C1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n10331), .A(
        n17227), .B(n17226), .ZN(n17228) );
  NAND3_X1 U20452 ( .A1(n17230), .A2(n17229), .A3(n17228), .ZN(n17459) );
  INV_X1 U20453 ( .A(n17459), .ZN(n17234) );
  OAI211_X1 U20454 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17232), .A(n17231), .B(
        n17355), .ZN(n17233) );
  OAI21_X1 U20455 ( .B1(n17234), .B2(n17355), .A(n17233), .ZN(P3_U2688) );
  AOI22_X1 U20456 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10286), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20457 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20458 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17235) );
  OAI211_X1 U20459 ( .C1(n10404), .C2(n18355), .A(n17236), .B(n17235), .ZN(
        n17243) );
  AOI22_X1 U20460 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20461 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U20462 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17239) );
  NAND2_X1 U20463 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n17238) );
  NAND4_X1 U20464 ( .A1(n17241), .A2(n17240), .A3(n17239), .A4(n17238), .ZN(
        n17242) );
  AOI211_X1 U20465 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17243), .B(n17242), .ZN(n17244) );
  OAI211_X1 U20466 ( .C1(n17334), .C2(n20886), .A(n17245), .B(n17244), .ZN(
        n17463) );
  INV_X1 U20467 ( .A(n17463), .ZN(n17253) );
  OAI21_X1 U20468 ( .B1(n17247), .B2(n17246), .A(P3_EBX_REG_14__SCAN_IN), .ZN(
        n17252) );
  NOR2_X1 U20469 ( .A1(n17365), .A2(n17352), .ZN(n17347) );
  NAND2_X1 U20470 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17347), .ZN(n17346) );
  NOR3_X1 U20471 ( .A1(n17248), .A2(n17342), .A3(n17339), .ZN(n17304) );
  INV_X1 U20472 ( .A(n17304), .ZN(n17337) );
  NOR2_X1 U20473 ( .A1(n17249), .A2(n17337), .ZN(n17320) );
  NAND2_X1 U20474 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17320), .ZN(n17301) );
  INV_X1 U20475 ( .A(n17301), .ZN(n17285) );
  NAND2_X1 U20476 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17285), .ZN(n17266) );
  NOR2_X1 U20477 ( .A1(n17456), .A2(n17266), .ZN(n17268) );
  NAND4_X1 U20478 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17268), .A4(n17250), .ZN(n17251) );
  OAI211_X1 U20479 ( .C1(n17253), .C2(n17355), .A(n17252), .B(n17251), .ZN(
        P3_U2689) );
  AOI22_X1 U20480 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17254) );
  OAI21_X1 U20481 ( .B1(n17325), .B2(n18659), .A(n17254), .ZN(n17265) );
  AOI22_X1 U20482 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17261) );
  AOI22_X1 U20483 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U20484 ( .B1(n17334), .B2(n18739), .A(n17255), .ZN(n17259) );
  AOI22_X1 U20485 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U20486 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10331), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17256) );
  OAI211_X1 U20487 ( .C1(n10404), .C2(n18344), .A(n17257), .B(n17256), .ZN(
        n17258) );
  AOI211_X1 U20488 ( .C1(n10286), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17259), .B(n17258), .ZN(n17260) );
  OAI211_X1 U20489 ( .C1(n17263), .C2(n17262), .A(n17261), .B(n17260), .ZN(
        n17264) );
  AOI211_X1 U20490 ( .C1(n17205), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n17265), .B(n17264), .ZN(n17470) );
  AND2_X1 U20491 ( .A1(n17355), .A2(n17266), .ZN(n17284) );
  AOI22_X1 U20492 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17284), .B1(n17268), 
        .B2(n17267), .ZN(n17269) );
  OAI21_X1 U20493 ( .B1(n17470), .B2(n17355), .A(n17269), .ZN(P3_U2691) );
  AOI22_X1 U20494 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20495 ( .A1(n17270), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17271) );
  OAI21_X1 U20496 ( .B1(n9771), .B2(n18578), .A(n17271), .ZN(n17280) );
  AOI22_X1 U20497 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10327), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U20498 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U20499 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17272) );
  OAI211_X1 U20500 ( .C1(n17275), .C2(n17274), .A(n17273), .B(n17272), .ZN(
        n17276) );
  AOI21_X1 U20501 ( .B1(n10289), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17276), .ZN(n17277) );
  OAI211_X1 U20502 ( .C1(n10404), .C2(n18338), .A(n17278), .B(n17277), .ZN(
        n17279) );
  AOI211_X1 U20503 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17280), .B(n17279), .ZN(n17281) );
  OAI211_X1 U20504 ( .C1(n10256), .C2(n17283), .A(n17282), .B(n17281), .ZN(
        n17474) );
  INV_X1 U20505 ( .A(n17474), .ZN(n17287) );
  OAI21_X1 U20506 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17285), .A(n17284), .ZN(
        n17286) );
  OAI21_X1 U20507 ( .B1(n17287), .B2(n17355), .A(n17286), .ZN(P3_U2692) );
  AOI22_X1 U20508 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17313), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20509 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17237), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U20510 ( .A1(n17205), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17288) );
  OAI211_X1 U20511 ( .C1(n10404), .C2(n18333), .A(n17289), .B(n17288), .ZN(
        n17296) );
  AOI22_X1 U20512 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U20513 ( .A1(n10330), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U20514 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17290), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17292) );
  NAND2_X1 U20515 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n17291) );
  NAND4_X1 U20516 ( .A1(n17294), .A2(n17293), .A3(n17292), .A4(n17291), .ZN(
        n17295) );
  AOI211_X1 U20517 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17296), .B(n17295), .ZN(n17297) );
  OAI211_X1 U20518 ( .C1(n17300), .C2(n17299), .A(n17298), .B(n17297), .ZN(
        n17477) );
  INV_X1 U20519 ( .A(n17477), .ZN(n17303) );
  OAI21_X1 U20520 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17320), .A(n17301), .ZN(
        n17302) );
  AOI22_X1 U20521 ( .A1(n17366), .A2(n17303), .B1(n17302), .B2(n17355), .ZN(
        P3_U2693) );
  OAI21_X1 U20522 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17304), .A(n17355), .ZN(
        n17319) );
  AOI22_X1 U20523 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10330), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17305) );
  OAI21_X1 U20524 ( .B1(n17325), .B2(n18650), .A(n17305), .ZN(n17318) );
  AOI22_X1 U20525 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17315) );
  OAI22_X1 U20526 ( .A1(n10404), .A2(n18327), .B1(n9771), .B2(n18573), .ZN(
        n17312) );
  AOI22_X1 U20527 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20528 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20529 ( .A1(n10286), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10289), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17308) );
  NAND3_X1 U20530 ( .A1(n17310), .A2(n17309), .A3(n17308), .ZN(n17311) );
  AOI211_X1 U20531 ( .C1(n17313), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n17312), .B(n17311), .ZN(n17314) );
  OAI211_X1 U20532 ( .C1(n9814), .C2(n17316), .A(n17315), .B(n17314), .ZN(
        n17317) );
  AOI211_X1 U20533 ( .C1(n17323), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n17318), .B(n17317), .ZN(n17481) );
  OAI22_X1 U20534 ( .A1(n17320), .A2(n17319), .B1(n17481), .B2(n17355), .ZN(
        P3_U2694) );
  AOI22_X1 U20535 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15818), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17321) );
  OAI21_X1 U20536 ( .B1(n9771), .B2(n18570), .A(n17321), .ZN(n17336) );
  AOI22_X1 U20537 ( .A1(n17323), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10330), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U20538 ( .A1(n10327), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10286), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17324) );
  OAI21_X1 U20539 ( .B1(n17325), .B2(n18646), .A(n17324), .ZN(n17331) );
  AOI22_X1 U20540 ( .A1(n17327), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20541 ( .A1(n10331), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17328) );
  OAI211_X1 U20542 ( .C1(n10404), .C2(n18322), .A(n17329), .B(n17328), .ZN(
        n17330) );
  AOI211_X1 U20543 ( .C1(n10289), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17331), .B(n17330), .ZN(n17332) );
  OAI211_X1 U20544 ( .C1(n17334), .C2(n18713), .A(n17333), .B(n17332), .ZN(
        n17335) );
  AOI211_X1 U20545 ( .C1(n17205), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n17336), .B(n17335), .ZN(n17487) );
  NOR2_X1 U20546 ( .A1(n17456), .A2(n17339), .ZN(n17340) );
  OAI221_X1 U20547 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17340), .A(n17337), .ZN(n17338) );
  AOI22_X1 U20548 ( .A1(n17366), .A2(n17487), .B1(n17338), .B2(n17355), .ZN(
        P3_U2695) );
  NAND2_X1 U20549 ( .A1(n17355), .A2(n17339), .ZN(n17344) );
  AOI22_X1 U20550 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17366), .B1(
        n17340), .B2(n17342), .ZN(n17341) );
  OAI21_X1 U20551 ( .B1(n17342), .B2(n17344), .A(n17341), .ZN(P3_U2696) );
  AND2_X1 U20552 ( .A1(n17343), .A2(n17346), .ZN(n17345) );
  OAI22_X1 U20553 ( .A1(n17345), .A2(n17344), .B1(n18355), .B2(n17355), .ZN(
        P3_U2697) );
  OAI21_X1 U20554 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17347), .A(n17346), .ZN(
        n17348) );
  AOI22_X1 U20555 ( .A1(n17366), .A2(n20925), .B1(n17348), .B2(n17355), .ZN(
        P3_U2698) );
  AND2_X1 U20556 ( .A1(n17350), .A2(n17349), .ZN(n17359) );
  AND2_X1 U20557 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17359), .ZN(n17357) );
  NOR2_X1 U20558 ( .A1(n17366), .A2(n17351), .ZN(n17353) );
  OAI22_X1 U20559 ( .A1(n17357), .A2(n17353), .B1(n17352), .B2(n17368), .ZN(
        n17354) );
  OAI21_X1 U20560 ( .B1(n17355), .B2(n18344), .A(n17354), .ZN(P3_U2699) );
  AOI21_X1 U20561 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17355), .A(n17359), .ZN(
        n17356) );
  OAI22_X1 U20562 ( .A1(n17357), .A2(n17356), .B1(n18338), .B2(n17355), .ZN(
        P3_U2700) );
  AOI221_X1 U20563 ( .B1(n17358), .B2(n17362), .C1(n17456), .C2(n17362), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17360) );
  AOI211_X1 U20564 ( .C1(n17366), .C2(n18333), .A(n17360), .B(n17359), .ZN(
        P3_U2701) );
  INV_X1 U20565 ( .A(n17361), .ZN(n17364) );
  OAI222_X1 U20566 ( .A1(n17364), .A2(n17368), .B1(n17363), .B2(n17362), .C1(
        n18327), .C2(n17355), .ZN(P3_U2702) );
  AOI22_X1 U20567 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17366), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17365), .ZN(n17367) );
  OAI21_X1 U20568 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17368), .A(n17367), .ZN(
        P3_U2703) );
  INV_X1 U20569 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17529) );
  INV_X1 U20570 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17532) );
  INV_X1 U20571 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17630) );
  NAND2_X1 U20572 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17369), .ZN(n17516) );
  NAND3_X1 U20573 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17371) );
  NAND4_X1 U20574 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17370) );
  NOR3_X2 U20575 ( .A1(n17516), .A2(n17371), .A3(n17370), .ZN(n17455) );
  NAND3_X1 U20576 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .ZN(n17462) );
  NAND4_X1 U20577 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n17372)
         );
  NOR2_X1 U20578 ( .A1(n17462), .A2(n17372), .ZN(n17457) );
  NAND2_X1 U20579 ( .A1(n17455), .A2(n17457), .ZN(n17458) );
  NAND2_X1 U20580 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n17416) );
  NAND4_X1 U20581 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17373)
         );
  NAND2_X1 U20582 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17412), .ZN(n17411) );
  NAND2_X1 U20583 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17408), .ZN(n17407) );
  NAND2_X1 U20584 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17397), .ZN(n17392) );
  NOR2_X2 U20585 ( .A1(n17529), .A2(n17392), .ZN(n17388) );
  NAND2_X1 U20586 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17388), .ZN(n17383) );
  NAND2_X1 U20587 ( .A1(n17379), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17378) );
  NAND2_X1 U20588 ( .A1(n17374), .A2(n17432), .ZN(n17423) );
  OAI22_X1 U20589 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17515), .B1(n17432), 
        .B2(n17379), .ZN(n17375) );
  AOI22_X1 U20590 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17448), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17375), .ZN(n17376) );
  OAI21_X1 U20591 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17378), .A(n17376), .ZN(
        P3_U2704) );
  NOR2_X2 U20592 ( .A1(n17377), .A2(n17506), .ZN(n17449) );
  AOI22_X1 U20593 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17448), .ZN(n17381) );
  OAI211_X1 U20594 ( .C1(n17379), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17506), .B(
        n17378), .ZN(n17380) );
  OAI211_X1 U20595 ( .C1(n17382), .C2(n17508), .A(n17381), .B(n17380), .ZN(
        P3_U2705) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17448), .ZN(n17385) );
  OAI211_X1 U20597 ( .C1(n17388), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17506), .B(
        n17383), .ZN(n17384) );
  OAI211_X1 U20598 ( .C1(n17386), .C2(n17508), .A(n17385), .B(n17384), .ZN(
        P3_U2706) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17449), .B1(n17513), .B2(
        n17387), .ZN(n17391) );
  AOI211_X1 U20600 ( .C1(n17529), .C2(n17392), .A(n17388), .B(n17432), .ZN(
        n17389) );
  INV_X1 U20601 ( .A(n17389), .ZN(n17390) );
  OAI211_X1 U20602 ( .C1(n17423), .C2(n20975), .A(n17391), .B(n17390), .ZN(
        P3_U2707) );
  AOI22_X1 U20603 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17448), .ZN(n17394) );
  OAI211_X1 U20604 ( .C1(n17397), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17506), .B(
        n17392), .ZN(n17393) );
  OAI211_X1 U20605 ( .C1(n17395), .C2(n17508), .A(n17394), .B(n17393), .ZN(
        P3_U2708) );
  INV_X1 U20606 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17449), .B1(n17513), .B2(
        n17396), .ZN(n17400) );
  AOI211_X1 U20608 ( .C1(n17532), .C2(n17401), .A(n17397), .B(n17432), .ZN(
        n17398) );
  INV_X1 U20609 ( .A(n17398), .ZN(n17399) );
  OAI211_X1 U20610 ( .C1(n17423), .C2(n18328), .A(n17400), .B(n17399), .ZN(
        P3_U2709) );
  AOI22_X1 U20611 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17448), .ZN(n17404) );
  OAI211_X1 U20612 ( .C1(n17402), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17506), .B(
        n17401), .ZN(n17403) );
  OAI211_X1 U20613 ( .C1(n17405), .C2(n17508), .A(n17404), .B(n17403), .ZN(
        P3_U2710) );
  AOI22_X1 U20614 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17449), .B1(n17513), .B2(
        n17406), .ZN(n17410) );
  OAI211_X1 U20615 ( .C1(n17408), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17506), .B(
        n17407), .ZN(n17409) );
  OAI211_X1 U20616 ( .C1(n17423), .C2(n18316), .A(n17410), .B(n17409), .ZN(
        P3_U2711) );
  AOI22_X1 U20617 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17448), .ZN(n17414) );
  OAI211_X1 U20618 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17412), .A(n17506), .B(
        n17411), .ZN(n17413) );
  OAI211_X1 U20619 ( .C1(n17415), .C2(n17508), .A(n17414), .B(n17413), .ZN(
        P3_U2712) );
  INV_X1 U20620 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17583) );
  NAND2_X1 U20621 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17442), .ZN(n17438) );
  NOR2_X1 U20622 ( .A1(n17416), .A2(n17438), .ZN(n17418) );
  NAND2_X1 U20623 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17418), .ZN(n17422) );
  AOI22_X1 U20624 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17448), .B1(n17513), .B2(
        n17417), .ZN(n17421) );
  INV_X1 U20625 ( .A(n17418), .ZN(n17428) );
  NAND2_X1 U20626 ( .A1(n17506), .A2(n17428), .ZN(n17431) );
  OAI21_X1 U20627 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17515), .A(n17431), .ZN(
        n17419) );
  AOI22_X1 U20628 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17449), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17419), .ZN(n17420) );
  OAI211_X1 U20629 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17422), .A(n17421), .B(
        n17420), .ZN(P3_U2713) );
  INV_X1 U20630 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17540) );
  OAI22_X1 U20631 ( .A1(n17424), .A2(n17508), .B1(n18345), .B2(n17423), .ZN(
        n17425) );
  AOI21_X1 U20632 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17449), .A(n17425), .ZN(
        n17426) );
  OAI221_X1 U20633 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17428), .C1(n17540), 
        .C2(n17431), .A(n17426), .ZN(P3_U2714) );
  INV_X1 U20634 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17448), .B1(n17513), .B2(
        n17427), .ZN(n17430) );
  INV_X1 U20636 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17544) );
  NOR2_X1 U20637 ( .A1(n17544), .A2(n17438), .ZN(n17433) );
  AOI22_X1 U20638 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17449), .B1(n17433), .B2(
        n17428), .ZN(n17429) );
  OAI211_X1 U20639 ( .C1(n17542), .C2(n17431), .A(n17430), .B(n17429), .ZN(
        P3_U2715) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17448), .ZN(n17436) );
  AOI211_X1 U20641 ( .C1(n17544), .C2(n17438), .A(n17433), .B(n17432), .ZN(
        n17434) );
  INV_X1 U20642 ( .A(n17434), .ZN(n17435) );
  OAI211_X1 U20643 ( .C1(n17437), .C2(n17508), .A(n17436), .B(n17435), .ZN(
        P3_U2716) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17448), .ZN(n17440) );
  OAI211_X1 U20645 ( .C1(n17442), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17506), .B(
        n17438), .ZN(n17439) );
  OAI211_X1 U20646 ( .C1(n17441), .C2(n17508), .A(n17440), .B(n17439), .ZN(
        P3_U2717) );
  AOI22_X1 U20647 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17448), .ZN(n17446) );
  INV_X1 U20648 ( .A(n17450), .ZN(n17444) );
  INV_X1 U20649 ( .A(n17442), .ZN(n17443) );
  OAI211_X1 U20650 ( .C1(n17444), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17506), .B(
        n17443), .ZN(n17445) );
  OAI211_X1 U20651 ( .C1(n17447), .C2(n17508), .A(n17446), .B(n17445), .ZN(
        P3_U2718) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17449), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17448), .ZN(n17453) );
  OAI211_X1 U20653 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17451), .A(n17506), .B(
        n17450), .ZN(n17452) );
  OAI211_X1 U20654 ( .C1(n17454), .C2(n17508), .A(n17453), .B(n17452), .ZN(
        P3_U2719) );
  INV_X1 U20655 ( .A(n17455), .ZN(n17484) );
  NAND2_X1 U20656 ( .A1(n17457), .A2(n17490), .ZN(n17461) );
  NAND2_X1 U20657 ( .A1(n17506), .A2(n17458), .ZN(n17465) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17514), .B1(n17513), .B2(
        n17459), .ZN(n17460) );
  OAI221_X1 U20659 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17461), .C1(n17630), 
        .C2(n17465), .A(n17460), .ZN(P3_U2720) );
  NAND3_X1 U20660 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17490), .ZN(n17480) );
  NOR2_X1 U20661 ( .A1(n17462), .A2(n17480), .ZN(n17472) );
  NAND2_X1 U20662 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17472), .ZN(n17466) );
  INV_X1 U20663 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17625) );
  AOI22_X1 U20664 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17514), .B1(n17513), .B2(
        n17463), .ZN(n17464) );
  OAI221_X1 U20665 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17466), .C1(n17625), 
        .C2(n17465), .A(n17464), .ZN(P3_U2721) );
  INV_X1 U20666 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17623) );
  INV_X1 U20667 ( .A(n17466), .ZN(n17469) );
  AOI21_X1 U20668 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17506), .A(n17472), .ZN(
        n17468) );
  OAI222_X1 U20669 ( .A1(n17511), .A2(n17623), .B1(n17469), .B2(n17468), .C1(
        n17508), .C2(n17467), .ZN(P3_U2722) );
  INV_X1 U20670 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17618) );
  INV_X1 U20671 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17557) );
  NOR2_X1 U20672 ( .A1(n17557), .A2(n17480), .ZN(n17473) );
  AOI22_X1 U20673 ( .A1(n17473), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17506), .ZN(n17471) );
  OAI222_X1 U20674 ( .A1(n17511), .A2(n17618), .B1(n17472), .B2(n17471), .C1(
        n17508), .C2(n17470), .ZN(P3_U2723) );
  INV_X1 U20675 ( .A(n17473), .ZN(n17476) );
  INV_X1 U20676 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17616) );
  NAND2_X1 U20677 ( .A1(n17506), .A2(n17476), .ZN(n17479) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17514), .B1(n17513), .B2(
        n17474), .ZN(n17475) );
  OAI221_X1 U20679 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17476), .C1(n17616), 
        .C2(n17479), .A(n17475), .ZN(P3_U2724) );
  AOI22_X1 U20680 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17514), .B1(n17513), .B2(
        n17477), .ZN(n17478) );
  OAI221_X1 U20681 ( .B1(n17479), .B2(n17557), .C1(n17479), .C2(n17480), .A(
        n17478), .ZN(P3_U2725) );
  INV_X1 U20682 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17612) );
  INV_X1 U20683 ( .A(n17480), .ZN(n17483) );
  AOI22_X1 U20684 ( .A1(n17490), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17506), .ZN(n17482) );
  OAI222_X1 U20685 ( .A1(n17511), .A2(n17612), .B1(n17483), .B2(n17482), .C1(
        n17508), .C2(n17481), .ZN(P3_U2726) );
  INV_X1 U20686 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17610) );
  AOI22_X1 U20687 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17514), .B1(n17490), .B2(
        n17610), .ZN(n17486) );
  NAND3_X1 U20688 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17506), .A3(n17484), .ZN(
        n17485) );
  OAI211_X1 U20689 ( .C1(n17487), .C2(n17508), .A(n17486), .B(n17485), .ZN(
        P3_U2727) );
  INV_X1 U20690 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18356) );
  INV_X1 U20691 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17565) );
  INV_X1 U20692 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17570) );
  INV_X1 U20693 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17602) );
  NOR3_X1 U20694 ( .A1(n17602), .A2(n17578), .A3(n17515), .ZN(n17505) );
  NAND2_X1 U20695 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17510), .ZN(n17498) );
  NOR2_X1 U20696 ( .A1(n17570), .A2(n17498), .ZN(n17501) );
  NAND2_X1 U20697 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17501), .ZN(n17491) );
  NOR2_X1 U20698 ( .A1(n17565), .A2(n17491), .ZN(n17494) );
  AOI21_X1 U20699 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17506), .A(n17494), .ZN(
        n17489) );
  OAI222_X1 U20700 ( .A1(n17511), .A2(n18356), .B1(n17490), .B2(n17489), .C1(
        n17508), .C2(n17488), .ZN(P3_U2728) );
  INV_X1 U20701 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18351) );
  INV_X1 U20702 ( .A(n17491), .ZN(n17497) );
  AOI21_X1 U20703 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17506), .A(n17497), .ZN(
        n17493) );
  OAI222_X1 U20704 ( .A1(n17511), .A2(n18351), .B1(n17494), .B2(n17493), .C1(
        n17508), .C2(n17492), .ZN(P3_U2729) );
  INV_X1 U20705 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18346) );
  AOI21_X1 U20706 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17506), .A(n17501), .ZN(
        n17496) );
  OAI222_X1 U20707 ( .A1(n17511), .A2(n18346), .B1(n17497), .B2(n17496), .C1(
        n17508), .C2(n17495), .ZN(P3_U2730) );
  INV_X1 U20708 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18339) );
  INV_X1 U20709 ( .A(n17498), .ZN(n17504) );
  AOI21_X1 U20710 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17506), .A(n17504), .ZN(
        n17500) );
  OAI222_X1 U20711 ( .A1(n17511), .A2(n18339), .B1(n17501), .B2(n17500), .C1(
        n17508), .C2(n17499), .ZN(P3_U2731) );
  INV_X1 U20712 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18334) );
  AOI21_X1 U20713 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17506), .A(n17510), .ZN(
        n17503) );
  OAI222_X1 U20714 ( .A1(n17511), .A2(n18334), .B1(n17504), .B2(n17503), .C1(
        n17508), .C2(n17502), .ZN(P3_U2732) );
  INV_X1 U20715 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18329) );
  AOI21_X1 U20716 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17506), .A(n17505), .ZN(
        n17509) );
  OAI222_X1 U20717 ( .A1(n17511), .A2(n18329), .B1(n17510), .B2(n17509), .C1(
        n17508), .C2(n17507), .ZN(P3_U2733) );
  AOI22_X1 U20718 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17514), .B1(n17513), .B2(
        n17512), .ZN(n17520) );
  NOR2_X1 U20719 ( .A1(n17578), .A2(n17515), .ZN(n17518) );
  NOR2_X1 U20720 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17515), .ZN(n17517) );
  OAI22_X1 U20721 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17518), .B1(n17517), .B2(
        n17516), .ZN(n17519) );
  NAND2_X1 U20722 ( .A1(n17520), .A2(n17519), .ZN(P3_U2734) );
  NOR2_X1 U20723 ( .A1(n18937), .A2(n17995), .ZN(n17563) );
  NOR2_X4 U20724 ( .A1(n18980), .A2(n17524), .ZN(n17566) );
  AND2_X1 U20725 ( .A1(n17566), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20726 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U20727 ( .A1(n18980), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U20728 ( .B1(n17599), .B2(n17548), .A(n17525), .ZN(P3_U2737) );
  INV_X1 U20729 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17527) );
  AOI22_X1 U20730 ( .A1(n18980), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17526) );
  OAI21_X1 U20731 ( .B1(n17527), .B2(n17548), .A(n17526), .ZN(P3_U2738) );
  AOI22_X1 U20732 ( .A1(n18980), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17528) );
  OAI21_X1 U20733 ( .B1(n17529), .B2(n17548), .A(n17528), .ZN(P3_U2739) );
  INV_X1 U20734 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U20735 ( .A1(n18980), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17530) );
  OAI21_X1 U20736 ( .B1(n17595), .B2(n17548), .A(n17530), .ZN(P3_U2740) );
  AOI22_X1 U20737 ( .A1(n18980), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U20738 ( .B1(n17532), .B2(n17548), .A(n17531), .ZN(P3_U2741) );
  INV_X1 U20739 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20953) );
  AOI22_X1 U20740 ( .A1(n18980), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U20741 ( .B1(n20953), .B2(n17548), .A(n17533), .ZN(P3_U2742) );
  INV_X1 U20742 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17591) );
  AOI22_X1 U20743 ( .A1(n18980), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17534) );
  OAI21_X1 U20744 ( .B1(n17591), .B2(n17548), .A(n17534), .ZN(P3_U2743) );
  INV_X1 U20745 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17536) );
  AOI22_X1 U20746 ( .A1(n18980), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U20747 ( .B1(n17536), .B2(n17548), .A(n17535), .ZN(P3_U2744) );
  INV_X1 U20748 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U20749 ( .A1(n18980), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17537) );
  OAI21_X1 U20750 ( .B1(n17538), .B2(n17548), .A(n17537), .ZN(P3_U2745) );
  AOI22_X1 U20751 ( .A1(n17563), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17539) );
  OAI21_X1 U20752 ( .B1(n17540), .B2(n17548), .A(n17539), .ZN(P3_U2746) );
  AOI22_X1 U20753 ( .A1(n17563), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17541) );
  OAI21_X1 U20754 ( .B1(n17542), .B2(n17548), .A(n17541), .ZN(P3_U2747) );
  AOI22_X1 U20755 ( .A1(n17563), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17543) );
  OAI21_X1 U20756 ( .B1(n17544), .B2(n17548), .A(n17543), .ZN(P3_U2748) );
  INV_X1 U20757 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20851) );
  AOI22_X1 U20758 ( .A1(n17563), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17545) );
  OAI21_X1 U20759 ( .B1(n20851), .B2(n17548), .A(n17545), .ZN(P3_U2749) );
  AOI22_X1 U20760 ( .A1(n17563), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17546) );
  OAI21_X1 U20761 ( .B1(n17583), .B2(n17548), .A(n17546), .ZN(P3_U2750) );
  INV_X1 U20762 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U20763 ( .A1(n17563), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17547) );
  OAI21_X1 U20764 ( .B1(n20990), .B2(n17548), .A(n17547), .ZN(P3_U2751) );
  AOI22_X1 U20765 ( .A1(n17563), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17549) );
  OAI21_X1 U20766 ( .B1(n17630), .B2(n17577), .A(n17549), .ZN(P3_U2752) );
  AOI22_X1 U20767 ( .A1(n17563), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17550) );
  OAI21_X1 U20768 ( .B1(n17625), .B2(n17577), .A(n17550), .ZN(P3_U2753) );
  INV_X1 U20769 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17552) );
  AOI22_X1 U20770 ( .A1(n17563), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17551) );
  OAI21_X1 U20771 ( .B1(n17552), .B2(n17577), .A(n17551), .ZN(P3_U2754) );
  INV_X1 U20772 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20773 ( .A1(n17563), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17553) );
  OAI21_X1 U20774 ( .B1(n17554), .B2(n17577), .A(n17553), .ZN(P3_U2755) );
  AOI22_X1 U20775 ( .A1(n18980), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17555) );
  OAI21_X1 U20776 ( .B1(n17616), .B2(n17577), .A(n17555), .ZN(P3_U2756) );
  AOI22_X1 U20777 ( .A1(n18980), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17556) );
  OAI21_X1 U20778 ( .B1(n17557), .B2(n17577), .A(n17556), .ZN(P3_U2757) );
  INV_X1 U20779 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17559) );
  AOI22_X1 U20780 ( .A1(n18980), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17558) );
  OAI21_X1 U20781 ( .B1(n17559), .B2(n17577), .A(n17558), .ZN(P3_U2758) );
  AOI22_X1 U20782 ( .A1(n18980), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17560) );
  OAI21_X1 U20783 ( .B1(n17610), .B2(n17577), .A(n17560), .ZN(P3_U2759) );
  INV_X1 U20784 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17562) );
  AOI22_X1 U20785 ( .A1(n18980), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17561) );
  OAI21_X1 U20786 ( .B1(n17562), .B2(n17577), .A(n17561), .ZN(P3_U2760) );
  AOI22_X1 U20787 ( .A1(n17563), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17564) );
  OAI21_X1 U20788 ( .B1(n17565), .B2(n17577), .A(n17564), .ZN(P3_U2761) );
  INV_X1 U20789 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17568) );
  AOI22_X1 U20790 ( .A1(n18980), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17567) );
  OAI21_X1 U20791 ( .B1(n17568), .B2(n17577), .A(n17567), .ZN(P3_U2762) );
  AOI22_X1 U20792 ( .A1(n18980), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17569) );
  OAI21_X1 U20793 ( .B1(n17570), .B2(n17577), .A(n17569), .ZN(P3_U2763) );
  INV_X1 U20794 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17572) );
  AOI22_X1 U20795 ( .A1(n18980), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17571) );
  OAI21_X1 U20796 ( .B1(n17572), .B2(n17577), .A(n17571), .ZN(P3_U2764) );
  INV_X1 U20797 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U20798 ( .A1(n18980), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17573) );
  OAI21_X1 U20799 ( .B1(n17574), .B2(n17577), .A(n17573), .ZN(P3_U2765) );
  AOI22_X1 U20800 ( .A1(n18980), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17575) );
  OAI21_X1 U20801 ( .B1(n17602), .B2(n17577), .A(n17575), .ZN(P3_U2766) );
  AOI22_X1 U20802 ( .A1(n18980), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17566), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17576) );
  OAI21_X1 U20803 ( .B1(n17578), .B2(n17577), .A(n17576), .ZN(P3_U2767) );
  INV_X1 U20804 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n20888) );
  NAND3_X1 U20805 ( .A1(n18324), .A2(n17580), .A3(n17579), .ZN(n17629) );
  AOI22_X1 U20806 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17626), .ZN(n17581) );
  OAI21_X1 U20807 ( .B1(n20888), .B2(n17622), .A(n17581), .ZN(P3_U2768) );
  AOI22_X1 U20808 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17627), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17626), .ZN(n17582) );
  OAI21_X1 U20809 ( .B1(n17583), .B2(n17629), .A(n17582), .ZN(P3_U2769) );
  AOI22_X1 U20810 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17626), .ZN(n17584) );
  OAI21_X1 U20811 ( .B1(n18329), .B2(n17622), .A(n17584), .ZN(P3_U2770) );
  AOI22_X1 U20812 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17626), .ZN(n17585) );
  OAI21_X1 U20813 ( .B1(n18334), .B2(n17622), .A(n17585), .ZN(P3_U2771) );
  AOI22_X1 U20814 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17626), .ZN(n17586) );
  OAI21_X1 U20815 ( .B1(n18339), .B2(n17622), .A(n17586), .ZN(P3_U2772) );
  AOI22_X1 U20816 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17626), .ZN(n17587) );
  OAI21_X1 U20817 ( .B1(n18346), .B2(n17622), .A(n17587), .ZN(P3_U2773) );
  AOI22_X1 U20818 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17626), .ZN(n17588) );
  OAI21_X1 U20819 ( .B1(n18351), .B2(n17622), .A(n17588), .ZN(P3_U2774) );
  AOI22_X1 U20820 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17626), .ZN(n17589) );
  OAI21_X1 U20821 ( .B1(n18356), .B2(n17622), .A(n17589), .ZN(P3_U2775) );
  AOI22_X1 U20822 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17627), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17626), .ZN(n17590) );
  OAI21_X1 U20823 ( .B1(n17591), .B2(n17629), .A(n17590), .ZN(P3_U2776) );
  AOI22_X1 U20824 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17626), .ZN(n17592) );
  OAI21_X1 U20825 ( .B1(n17612), .B2(n17622), .A(n17592), .ZN(P3_U2777) );
  INV_X1 U20826 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U20827 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17626), .ZN(n17593) );
  OAI21_X1 U20828 ( .B1(n17614), .B2(n17622), .A(n17593), .ZN(P3_U2778) );
  AOI22_X1 U20829 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17627), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17626), .ZN(n17594) );
  OAI21_X1 U20830 ( .B1(n17595), .B2(n17629), .A(n17594), .ZN(P3_U2779) );
  AOI22_X1 U20831 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17626), .ZN(n17596) );
  OAI21_X1 U20832 ( .B1(n17618), .B2(n17622), .A(n17596), .ZN(P3_U2780) );
  AOI22_X1 U20833 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17620), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17626), .ZN(n17597) );
  OAI21_X1 U20834 ( .B1(n17623), .B2(n17622), .A(n17597), .ZN(P3_U2781) );
  AOI22_X1 U20835 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17627), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17626), .ZN(n17598) );
  OAI21_X1 U20836 ( .B1(n17599), .B2(n17629), .A(n17598), .ZN(P3_U2782) );
  AOI22_X1 U20837 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17626), .ZN(n17600) );
  OAI21_X1 U20838 ( .B1(n20888), .B2(n17622), .A(n17600), .ZN(P3_U2783) );
  AOI22_X1 U20839 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17627), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17626), .ZN(n17601) );
  OAI21_X1 U20840 ( .B1(n17602), .B2(n17629), .A(n17601), .ZN(P3_U2784) );
  AOI22_X1 U20841 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17619), .ZN(n17603) );
  OAI21_X1 U20842 ( .B1(n18329), .B2(n17622), .A(n17603), .ZN(P3_U2785) );
  AOI22_X1 U20843 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17619), .ZN(n17604) );
  OAI21_X1 U20844 ( .B1(n18334), .B2(n17622), .A(n17604), .ZN(P3_U2786) );
  AOI22_X1 U20845 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17619), .ZN(n17605) );
  OAI21_X1 U20846 ( .B1(n18339), .B2(n17622), .A(n17605), .ZN(P3_U2787) );
  AOI22_X1 U20847 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17619), .ZN(n17606) );
  OAI21_X1 U20848 ( .B1(n18346), .B2(n17622), .A(n17606), .ZN(P3_U2788) );
  AOI22_X1 U20849 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17619), .ZN(n17607) );
  OAI21_X1 U20850 ( .B1(n18351), .B2(n17622), .A(n17607), .ZN(P3_U2789) );
  AOI22_X1 U20851 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17619), .ZN(n17608) );
  OAI21_X1 U20852 ( .B1(n18356), .B2(n17622), .A(n17608), .ZN(P3_U2790) );
  AOI22_X1 U20853 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17627), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17626), .ZN(n17609) );
  OAI21_X1 U20854 ( .B1(n17610), .B2(n17629), .A(n17609), .ZN(P3_U2791) );
  AOI22_X1 U20855 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17619), .ZN(n17611) );
  OAI21_X1 U20856 ( .B1(n17612), .B2(n17622), .A(n17611), .ZN(P3_U2792) );
  AOI22_X1 U20857 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17619), .ZN(n17613) );
  OAI21_X1 U20858 ( .B1(n17614), .B2(n17622), .A(n17613), .ZN(P3_U2793) );
  AOI22_X1 U20859 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17627), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17626), .ZN(n17615) );
  OAI21_X1 U20860 ( .B1(n17616), .B2(n17629), .A(n17615), .ZN(P3_U2794) );
  AOI22_X1 U20861 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17619), .ZN(n17617) );
  OAI21_X1 U20862 ( .B1(n17618), .B2(n17622), .A(n17617), .ZN(P3_U2795) );
  AOI22_X1 U20863 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17620), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17619), .ZN(n17621) );
  OAI21_X1 U20864 ( .B1(n17623), .B2(n17622), .A(n17621), .ZN(P3_U2796) );
  AOI22_X1 U20865 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17627), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17626), .ZN(n17624) );
  OAI21_X1 U20866 ( .B1(n17625), .B2(n17629), .A(n17624), .ZN(P3_U2797) );
  AOI22_X1 U20867 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17627), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17626), .ZN(n17628) );
  OAI21_X1 U20868 ( .B1(n17630), .B2(n17629), .A(n17628), .ZN(P3_U2798) );
  INV_X1 U20869 ( .A(n17995), .ZN(n17826) );
  INV_X1 U20870 ( .A(n17968), .ZN(n17956) );
  OAI21_X1 U20871 ( .B1(n17633), .B2(n17956), .A(n17996), .ZN(n17631) );
  AOI21_X1 U20872 ( .B1(n17826), .B2(n17632), .A(n17631), .ZN(n17659) );
  OAI21_X1 U20873 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17770), .A(
        n17659), .ZN(n17649) );
  NAND2_X1 U20874 ( .A1(n17633), .A2(n17785), .ZN(n17653) );
  AOI221_X1 U20875 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(n9967), .C2(n17634), .A(n17653), .ZN(n17636) );
  INV_X1 U20876 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18911) );
  NOR2_X1 U20877 ( .A1(n18199), .A2(n18911), .ZN(n17635) );
  AOI211_X1 U20878 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17649), .A(
        n17636), .B(n17635), .ZN(n17647) );
  NOR2_X1 U20879 ( .A1(n17900), .A2(n9775), .ZN(n17742) );
  OAI22_X1 U20880 ( .A1(n18006), .A2(n17691), .B1(n17637), .B2(n18000), .ZN(
        n17667) );
  NOR2_X1 U20881 ( .A1(n18009), .A2(n17667), .ZN(n17639) );
  NOR3_X1 U20882 ( .A1(n17742), .A2(n17639), .A3(n17638), .ZN(n17644) );
  AOI211_X1 U20883 ( .C1(n17642), .C2(n17641), .A(n17640), .B(n17898), .ZN(
        n17643) );
  AOI211_X1 U20884 ( .C1(n17779), .C2(n17645), .A(n17644), .B(n17643), .ZN(
        n17646) );
  OAI211_X1 U20885 ( .C1(n17843), .C2(n17648), .A(n17647), .B(n17646), .ZN(
        P3_U2802) );
  AOI22_X1 U20886 ( .A1(n18301), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17649), .ZN(n17657) );
  NOR2_X1 U20887 ( .A1(n18007), .A2(n17795), .ZN(n17655) );
  NOR2_X1 U20888 ( .A1(n17651), .A2(n17650), .ZN(n17652) );
  XOR2_X1 U20889 ( .A(n17652), .B(n17871), .Z(n18012) );
  OAI22_X1 U20890 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17653), .B1(
        n18012), .B2(n17898), .ZN(n17654) );
  AOI221_X1 U20891 ( .B1(n17655), .B2(n18009), .C1(n17667), .C2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n17654), .ZN(n17656) );
  OAI211_X1 U20892 ( .C1(n17843), .C2(n17658), .A(n17657), .B(n17656), .ZN(
        P3_U2803) );
  INV_X1 U20893 ( .A(n18023), .ZN(n18025) );
  NAND4_X1 U20894 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18021), .A3(
        n18025), .A4(n18013), .ZN(n18019) );
  AOI221_X1 U20895 ( .B1(n18358), .B2(n17661), .C1(n17660), .C2(n17661), .A(
        n17659), .ZN(n17664) );
  AOI21_X1 U20896 ( .B1(n17843), .B2(n17770), .A(n17662), .ZN(n17663) );
  AOI211_X1 U20897 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n18301), .A(n17664), 
        .B(n17663), .ZN(n17669) );
  OAI21_X1 U20898 ( .B1(n17666), .B2(n18013), .A(n17665), .ZN(n18015) );
  AOI22_X1 U20899 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17667), .B1(
        n17888), .B2(n18015), .ZN(n17668) );
  OAI211_X1 U20900 ( .C1(n17795), .C2(n18019), .A(n17669), .B(n17668), .ZN(
        P3_U2804) );
  XOR2_X1 U20901 ( .A(n17670), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18035) );
  OR2_X1 U20902 ( .A1(n17673), .A2(n18358), .ZN(n17700) );
  OAI211_X1 U20903 ( .C1(n17995), .C2(n17671), .A(n17996), .B(n17700), .ZN(
        n17672) );
  INV_X1 U20904 ( .A(n17672), .ZN(n17703) );
  OAI21_X1 U20905 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17770), .A(
        n17703), .ZN(n17689) );
  NOR2_X1 U20906 ( .A1(n18199), .A2(n18902), .ZN(n18030) );
  NAND2_X1 U20907 ( .A1(n17673), .A2(n17785), .ZN(n17686) );
  OAI21_X1 U20908 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17674), .ZN(n17675) );
  OAI22_X1 U20909 ( .A1(n17843), .A2(n17676), .B1(n17686), .B2(n17675), .ZN(
        n17677) );
  AOI211_X1 U20910 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17689), .A(
        n18030), .B(n17677), .ZN(n17683) );
  XOR2_X1 U20911 ( .A(n17678), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18032) );
  OAI21_X1 U20912 ( .B1(n17871), .B2(n17680), .A(n17679), .ZN(n17681) );
  XOR2_X1 U20913 ( .A(n17681), .B(n18022), .Z(n18031) );
  AOI22_X1 U20914 ( .A1(n9775), .A2(n18032), .B1(n17888), .B2(n18031), .ZN(
        n17682) );
  OAI211_X1 U20915 ( .C1(n17691), .C2(n18035), .A(n17683), .B(n17682), .ZN(
        P3_U2805) );
  OR2_X1 U20916 ( .A1(n17684), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18048) );
  NOR2_X1 U20917 ( .A1(n18199), .A2(n18900), .ZN(n17688) );
  OAI22_X1 U20918 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17686), .B1(
        n17843), .B2(n17685), .ZN(n17687) );
  AOI211_X1 U20919 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17689), .A(
        n17688), .B(n17687), .ZN(n17696) );
  OAI22_X1 U20920 ( .A1(n18041), .A2(n17691), .B1(n17690), .B2(n18000), .ZN(
        n17707) );
  OAI21_X1 U20921 ( .B1(n17694), .B2(n17693), .A(n17692), .ZN(n18037) );
  AOI22_X1 U20922 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17707), .B1(
        n17888), .B2(n18037), .ZN(n17695) );
  OAI211_X1 U20923 ( .C1(n17795), .C2(n18048), .A(n17696), .B(n17695), .ZN(
        P3_U2806) );
  OAI22_X1 U20924 ( .A1(n17697), .A2(n17710), .B1(n17871), .B2(n18058), .ZN(
        n17698) );
  NOR2_X1 U20925 ( .A1(n17698), .A2(n17743), .ZN(n17699) );
  XOR2_X1 U20926 ( .A(n17699), .B(n20822), .Z(n18054) );
  OAI22_X1 U20927 ( .A1(n17703), .A2(n17702), .B1(n17701), .B2(n17700), .ZN(
        n17706) );
  NAND2_X1 U20928 ( .A1(n18235), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18052) );
  OAI221_X1 U20929 ( .B1(n17704), .B2(n17843), .C1(n17704), .C2(n17770), .A(
        n18052), .ZN(n17705) );
  AOI211_X1 U20930 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17707), .A(
        n17706), .B(n17705), .ZN(n17709) );
  NAND3_X1 U20931 ( .A1(n18021), .A2(n17779), .A3(n20822), .ZN(n17708) );
  OAI211_X1 U20932 ( .C1(n18054), .C2(n17898), .A(n17709), .B(n17708), .ZN(
        P3_U2807) );
  OAI221_X1 U20933 ( .B1(n17710), .B2(n9820), .C1(n17710), .C2(n18066), .A(
        n9977), .ZN(n17711) );
  XOR2_X1 U20934 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17711), .Z(
        n18074) );
  OAI22_X1 U20935 ( .A1(n17714), .A2(n17956), .B1(n17712), .B2(n17995), .ZN(
        n17713) );
  NOR2_X1 U20936 ( .A1(n17941), .A2(n17713), .ZN(n17736) );
  OAI21_X1 U20937 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17770), .A(
        n17736), .ZN(n17727) );
  INV_X1 U20938 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17715) );
  NAND2_X1 U20939 ( .A1(n17714), .A2(n17785), .ZN(n17724) );
  AOI221_X1 U20940 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17716), .C2(n17715), .A(
        n17724), .ZN(n17719) );
  NAND2_X1 U20941 ( .A1(n18301), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18072) );
  OAI21_X1 U20942 ( .B1(n17717), .B2(n17843), .A(n18072), .ZN(n17718) );
  AOI211_X1 U20943 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17727), .A(
        n17719), .B(n17718), .ZN(n17722) );
  AOI22_X1 U20944 ( .A1(n17900), .A2(n18132), .B1(n9775), .B2(n18057), .ZN(
        n17794) );
  OAI21_X1 U20945 ( .B1(n18066), .B2(n17742), .A(n17794), .ZN(n17732) );
  OAI21_X1 U20946 ( .B1(n18055), .B2(n17795), .A(n18058), .ZN(n17720) );
  OAI21_X1 U20947 ( .B1(n18058), .B2(n17732), .A(n17720), .ZN(n17721) );
  OAI211_X1 U20948 ( .C1(n17898), .C2(n18074), .A(n17722), .B(n17721), .ZN(
        P3_U2808) );
  INV_X1 U20949 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18067) );
  NAND2_X1 U20950 ( .A1(n18082), .A2(n18067), .ZN(n18087) );
  NOR2_X1 U20951 ( .A1(n18062), .A2(n17769), .ZN(n18077) );
  NAND2_X1 U20952 ( .A1(n17779), .A2(n18077), .ZN(n17758) );
  NOR2_X1 U20953 ( .A1(n18199), .A2(n18894), .ZN(n17726) );
  OAI22_X1 U20954 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17724), .B1(
        n17843), .B2(n17723), .ZN(n17725) );
  AOI211_X1 U20955 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17727), .A(
        n17726), .B(n17725), .ZN(n17734) );
  NAND3_X1 U20956 ( .A1(n17871), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17728), .ZN(n17753) );
  INV_X1 U20957 ( .A(n17729), .ZN(n17765) );
  OAI22_X1 U20958 ( .A1(n18060), .A2(n17753), .B1(n17765), .B2(n17730), .ZN(
        n17731) );
  XNOR2_X1 U20959 ( .A(n18067), .B(n17731), .ZN(n18076) );
  AOI22_X1 U20960 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17732), .B1(
        n17888), .B2(n18076), .ZN(n17733) );
  OAI211_X1 U20961 ( .C1(n18087), .C2(n17758), .A(n17734), .B(n17733), .ZN(
        P3_U2809) );
  NAND2_X1 U20962 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17735), .ZN(
        n18094) );
  AOI221_X1 U20963 ( .B1(n17737), .B2(n21028), .C1(n18358), .C2(n21028), .A(
        n17736), .ZN(n17741) );
  AOI21_X1 U20964 ( .B1(n17843), .B2(n17770), .A(n17739), .ZN(n17740) );
  AOI211_X1 U20965 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n18301), .A(n17741), 
        .B(n17740), .ZN(n17747) );
  NAND2_X1 U20966 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18077), .ZN(
        n18063) );
  INV_X1 U20967 ( .A(n18063), .ZN(n18089) );
  OAI21_X1 U20968 ( .B1(n17742), .B2(n18089), .A(n17794), .ZN(n17755) );
  INV_X1 U20969 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17744) );
  AOI221_X1 U20970 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17753), 
        .C1(n17744), .C2(n17764), .A(n17743), .ZN(n17745) );
  XOR2_X1 U20971 ( .A(n17745), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n18088) );
  AOI22_X1 U20972 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17755), .B1(
        n17888), .B2(n18088), .ZN(n17746) );
  OAI211_X1 U20973 ( .C1(n18094), .C2(n17758), .A(n17747), .B(n17746), .ZN(
        P3_U2810) );
  INV_X1 U20974 ( .A(n17991), .ZN(n17882) );
  OAI21_X1 U20975 ( .B1(n17941), .B2(n9837), .A(n17882), .ZN(n17771) );
  OAI21_X1 U20976 ( .B1(n17748), .B2(n17995), .A(n17771), .ZN(n17762) );
  NAND2_X1 U20977 ( .A1(n18235), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18097) );
  NOR2_X1 U20978 ( .A1(n17829), .A2(n9837), .ZN(n17763) );
  OAI211_X1 U20979 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17763), .B(n17749), .ZN(n17750) );
  OAI211_X1 U20980 ( .C1(n17751), .C2(n17843), .A(n18097), .B(n17750), .ZN(
        n17752) );
  AOI21_X1 U20981 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17762), .A(
        n17752), .ZN(n17757) );
  OAI21_X1 U20982 ( .B1(n17765), .B2(n17764), .A(n17753), .ZN(n17754) );
  XOR2_X1 U20983 ( .A(n17754), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18095) );
  AOI22_X1 U20984 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17755), .B1(
        n17888), .B2(n18095), .ZN(n17756) );
  OAI211_X1 U20985 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17758), .A(
        n17757), .B(n17756), .ZN(P3_U2811) );
  INV_X1 U20986 ( .A(n17794), .ZN(n17759) );
  AOI21_X1 U20987 ( .B1(n17779), .B2(n18062), .A(n17759), .ZN(n17777) );
  OAI22_X1 U20988 ( .A1(n18199), .A2(n20989), .B1(n17843), .B2(n17760), .ZN(
        n17761) );
  AOI221_X1 U20989 ( .B1(n17763), .B2(n9960), .C1(n17762), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17761), .ZN(n17768) );
  OAI21_X1 U20990 ( .B1(n17897), .B2(n17769), .A(n17764), .ZN(n17766) );
  XOR2_X1 U20991 ( .A(n17766), .B(n17765), .Z(n18112) );
  NOR2_X1 U20992 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18062), .ZN(
        n18111) );
  AOI22_X1 U20993 ( .A1(n17888), .A2(n18112), .B1(n17779), .B2(n18111), .ZN(
        n17767) );
  OAI211_X1 U20994 ( .C1(n17777), .C2(n17769), .A(n17768), .B(n17767), .ZN(
        P3_U2812) );
  NAND2_X2 U20995 ( .A1(n17843), .A2(n17770), .ZN(n17988) );
  AOI221_X1 U20996 ( .B1(n17773), .B2(n17772), .C1(n18358), .C2(n17772), .A(
        n17771), .ZN(n17774) );
  AOI21_X1 U20997 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n18301), .A(n17774), 
        .ZN(n17781) );
  NOR2_X1 U20998 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18125), .ZN(
        n18115) );
  AOI21_X1 U20999 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17776), .A(
        n17775), .ZN(n18119) );
  OAI22_X1 U21000 ( .A1(n18119), .A2(n17898), .B1(n17777), .B2(n18106), .ZN(
        n17778) );
  AOI21_X1 U21001 ( .B1(n17779), .B2(n18115), .A(n17778), .ZN(n17780) );
  OAI211_X1 U21002 ( .C1(n17975), .C2(n17782), .A(n17781), .B(n17780), .ZN(
        P3_U2813) );
  OAI21_X1 U21003 ( .B1(n17897), .B2(n9820), .A(n17783), .ZN(n17784) );
  XOR2_X1 U21004 ( .A(n17784), .B(n18125), .Z(n18127) );
  NAND2_X1 U21005 ( .A1(n17786), .A2(n17785), .ZN(n17800) );
  AOI221_X1 U21006 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n20936), .C2(n17790), .A(
        n17800), .ZN(n17792) );
  OAI21_X1 U21007 ( .B1(n17786), .B2(n17956), .A(n17996), .ZN(n17813) );
  AOI21_X1 U21008 ( .B1(n17826), .B2(n17787), .A(n17813), .ZN(n17799) );
  AOI22_X1 U21009 ( .A1(n18301), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17803), 
        .B2(n17788), .ZN(n17789) );
  OAI21_X1 U21010 ( .B1(n17799), .B2(n17790), .A(n17789), .ZN(n17791) );
  AOI211_X1 U21011 ( .C1(n18127), .C2(n17888), .A(n17792), .B(n17791), .ZN(
        n17793) );
  OAI221_X1 U21012 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17795), 
        .C1(n18125), .C2(n17794), .A(n17793), .ZN(P3_U2814) );
  INV_X1 U21013 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17854) );
  NAND3_X1 U21014 ( .A1(n17814), .A2(n17897), .A3(n17854), .ZN(n17848) );
  OAI22_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17848), .B1(
        n17815), .B2(n17796), .ZN(n17797) );
  OAI221_X1 U21016 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n10354), 
        .C1(n18178), .C2(n17871), .A(n17797), .ZN(n17798) );
  XOR2_X1 U21017 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17798), .Z(
        n18138) );
  NAND2_X1 U21018 ( .A1(n18235), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18141) );
  OAI221_X1 U21019 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17800), .C1(
        n20936), .C2(n17799), .A(n18141), .ZN(n17801) );
  AOI21_X1 U21020 ( .B1(n17803), .B2(n17802), .A(n17801), .ZN(n17809) );
  AOI21_X1 U21021 ( .B1(n18143), .B2(n17819), .A(n17804), .ZN(n18139) );
  AND2_X1 U21022 ( .A1(n18132), .A2(n17900), .ZN(n17807) );
  NAND2_X1 U21023 ( .A1(n17805), .A2(n18143), .ZN(n17806) );
  AOI22_X1 U21024 ( .A1(n9775), .A2(n18139), .B1(n17807), .B2(n17806), .ZN(
        n17808) );
  OAI211_X1 U21025 ( .C1(n17898), .C2(n18138), .A(n17809), .B(n17808), .ZN(
        P3_U2815) );
  NAND3_X1 U21026 ( .A1(n17928), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18704), .ZN(n17907) );
  NOR2_X1 U21027 ( .A1(n17902), .A2(n17907), .ZN(n17881) );
  NAND2_X1 U21028 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17881), .ZN(
        n17880) );
  NOR2_X1 U21029 ( .A1(n17866), .A2(n17880), .ZN(n17865) );
  NAND2_X1 U21030 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17865), .ZN(
        n17811) );
  OAI21_X1 U21031 ( .B1(n17830), .B2(n17811), .A(n17810), .ZN(n17812) );
  AOI22_X1 U21032 ( .A1(n18301), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17813), 
        .B2(n17812), .ZN(n17823) );
  NAND2_X1 U21033 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18187), .ZN(
        n18163) );
  INV_X1 U21034 ( .A(n18163), .ZN(n17836) );
  NAND2_X1 U21035 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17836), .ZN(
        n18144) );
  AOI221_X1 U21036 ( .B1(n17835), .B2(n10354), .C1(n18144), .C2(n10354), .A(
        n18134), .ZN(n18153) );
  NAND2_X1 U21037 ( .A1(n17814), .A2(n17897), .ZN(n17860) );
  INV_X1 U21038 ( .A(n17860), .ZN(n17816) );
  NOR2_X1 U21039 ( .A1(n17897), .A2(n17815), .ZN(n17877) );
  INV_X1 U21040 ( .A(n18144), .ZN(n18146) );
  AOI22_X1 U21041 ( .A1(n17817), .A2(n17816), .B1(n17877), .B2(n18146), .ZN(
        n17818) );
  XOR2_X1 U21042 ( .A(n17818), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18151) );
  OAI221_X1 U21043 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18146), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17820), .A(n17819), .ZN(
        n18156) );
  OAI22_X1 U21044 ( .A1(n18151), .A2(n17898), .B1(n18000), .B2(n18156), .ZN(
        n17821) );
  AOI21_X1 U21045 ( .B1(n17900), .B2(n18153), .A(n17821), .ZN(n17822) );
  OAI211_X1 U21046 ( .C1(n17975), .C2(n17824), .A(n17823), .B(n17822), .ZN(
        P3_U2816) );
  INV_X1 U21047 ( .A(n17841), .ZN(n17891) );
  OR2_X1 U21048 ( .A1(n18163), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18168) );
  AOI22_X1 U21049 ( .A1(n17968), .A2(n17828), .B1(n17826), .B2(n17825), .ZN(
        n17827) );
  NAND2_X1 U21050 ( .A1(n17827), .A2(n17996), .ZN(n17845) );
  NOR2_X1 U21051 ( .A1(n17829), .A2(n17828), .ZN(n17847) );
  OAI211_X1 U21052 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17847), .B(n17830), .ZN(n17832) );
  NAND2_X1 U21053 ( .A1(n18235), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17831) );
  OAI211_X1 U21054 ( .C1(n17843), .C2(n17833), .A(n17832), .B(n17831), .ZN(
        n17834) );
  AOI21_X1 U21055 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17845), .A(
        n17834), .ZN(n17840) );
  AOI22_X1 U21056 ( .A1(n17900), .A2(n17835), .B1(n9775), .B2(n18162), .ZN(
        n17890) );
  OAI21_X1 U21057 ( .B1(n17891), .B2(n17836), .A(n17890), .ZN(n17850) );
  INV_X1 U21058 ( .A(n17877), .ZN(n17837) );
  OAI22_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17848), .B1(
        n17837), .B2(n18163), .ZN(n17838) );
  XOR2_X1 U21060 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17838), .Z(
        n18157) );
  AOI22_X1 U21061 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17850), .B1(
        n17888), .B2(n18157), .ZN(n17839) );
  OAI211_X1 U21062 ( .C1(n17891), .C2(n18168), .A(n17840), .B(n17839), .ZN(
        P3_U2817) );
  NAND2_X1 U21063 ( .A1(n17841), .A2(n18163), .ZN(n17853) );
  OAI22_X1 U21064 ( .A1(n18199), .A2(n18878), .B1(n17843), .B2(n17842), .ZN(
        n17844) );
  AOI221_X1 U21065 ( .B1(n17847), .B2(n17846), .C1(n17845), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17844), .ZN(n17852) );
  NAND2_X1 U21066 ( .A1(n18180), .A2(n17877), .ZN(n17859) );
  OAI21_X1 U21067 ( .B1(n17854), .B2(n17859), .A(n17848), .ZN(n17849) );
  XOR2_X1 U21068 ( .A(n17849), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18169) );
  AOI22_X1 U21069 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17850), .B1(
        n17888), .B2(n18169), .ZN(n17851) );
  OAI211_X1 U21070 ( .C1(n18172), .C2(n17853), .A(n17852), .B(n17851), .ZN(
        P3_U2818) );
  NAND2_X1 U21071 ( .A1(n18180), .A2(n17854), .ZN(n18192) );
  INV_X1 U21072 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17857) );
  NOR2_X1 U21073 ( .A1(n17857), .A2(n17865), .ZN(n17858) );
  OAI22_X1 U21074 ( .A1(n17975), .A2(n17855), .B1(n18199), .B2(n18876), .ZN(
        n17856) );
  AOI221_X1 U21075 ( .B1(n17882), .B2(n17858), .C1(n17857), .C2(n17865), .A(
        n17856), .ZN(n17864) );
  OAI21_X1 U21076 ( .B1(n18180), .B2(n17891), .A(n17890), .ZN(n17862) );
  NAND2_X1 U21077 ( .A1(n17860), .A2(n17859), .ZN(n17861) );
  XOR2_X1 U21078 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17861), .Z(
        n18179) );
  AOI22_X1 U21079 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17862), .B1(
        n17888), .B2(n18179), .ZN(n17863) );
  OAI211_X1 U21080 ( .C1(n17891), .C2(n18192), .A(n17864), .B(n17863), .ZN(
        P3_U2819) );
  AOI211_X1 U21081 ( .C1(n17880), .C2(n17866), .A(n17991), .B(n17865), .ZN(
        n17868) );
  NOR2_X1 U21082 ( .A1(n18199), .A2(n18874), .ZN(n17867) );
  AOI211_X1 U21083 ( .C1(n17869), .C2(n17988), .A(n17868), .B(n17867), .ZN(
        n17876) );
  NOR2_X1 U21084 ( .A1(n17871), .A2(n17870), .ZN(n17878) );
  AOI22_X1 U21085 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17877), .B1(
        n17878), .B2(n18206), .ZN(n17872) );
  XOR2_X1 U21086 ( .A(n21002), .B(n17872), .Z(n18195) );
  NOR2_X1 U21087 ( .A1(n18180), .A2(n17891), .ZN(n17874) );
  NAND2_X1 U21088 ( .A1(n21002), .A2(n18206), .ZN(n17873) );
  AOI22_X1 U21089 ( .A1(n17888), .A2(n18195), .B1(n17874), .B2(n17873), .ZN(
        n17875) );
  OAI211_X1 U21090 ( .C1(n17890), .C2(n21002), .A(n17876), .B(n17875), .ZN(
        P3_U2820) );
  NOR2_X1 U21091 ( .A1(n17878), .A2(n17877), .ZN(n17879) );
  XOR2_X1 U21092 ( .A(n17879), .B(n18206), .Z(n18202) );
  NOR2_X1 U21093 ( .A1(n18199), .A2(n18872), .ZN(n17887) );
  INV_X1 U21094 ( .A(n17880), .ZN(n17885) );
  AOI21_X1 U21095 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17882), .A(
        n17881), .ZN(n17884) );
  OAI22_X1 U21096 ( .A1(n17885), .A2(n17884), .B1(n17975), .B2(n17883), .ZN(
        n17886) );
  AOI211_X1 U21097 ( .C1(n17888), .C2(n18202), .A(n17887), .B(n17886), .ZN(
        n17889) );
  OAI221_X1 U21098 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17891), .C1(
        n18206), .C2(n17890), .A(n17889), .ZN(P3_U2821) );
  OAI21_X1 U21099 ( .B1(n17892), .B2(n17956), .A(n17996), .ZN(n17908) );
  AOI22_X1 U21100 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17908), .B1(
        n17893), .B2(n17988), .ZN(n17906) );
  OAI21_X1 U21101 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17895), .A(
        n17894), .ZN(n18210) );
  OAI21_X1 U21102 ( .B1(n18213), .B2(n17897), .A(n17896), .ZN(n18208) );
  OAI22_X1 U21103 ( .A1(n18000), .A2(n18210), .B1(n17898), .B2(n18208), .ZN(
        n17899) );
  AOI21_X1 U21104 ( .B1(n17900), .B2(n18213), .A(n17899), .ZN(n17905) );
  NAND2_X1 U21105 ( .A1(n18301), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18224) );
  NOR2_X1 U21106 ( .A1(n17901), .A2(n17909), .ZN(n17903) );
  OAI211_X1 U21107 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17903), .A(
        n18704), .B(n17902), .ZN(n17904) );
  NAND4_X1 U21108 ( .A1(n17906), .A2(n17905), .A3(n18224), .A4(n17904), .ZN(
        P3_U2822) );
  INV_X1 U21109 ( .A(n17907), .ZN(n17910) );
  NOR2_X1 U21110 ( .A1(n18199), .A2(n18868), .ZN(n18226) );
  AOI221_X1 U21111 ( .B1(n17910), .B2(n17909), .C1(n17908), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18226), .ZN(n17919) );
  AOI21_X1 U21112 ( .B1(n17913), .B2(n17912), .A(n17911), .ZN(n18228) );
  AOI21_X1 U21113 ( .B1(n17916), .B2(n17915), .A(n17914), .ZN(n17917) );
  XOR2_X1 U21114 ( .A(n17917), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18227) );
  AOI22_X1 U21115 ( .A1(n17994), .A2(n18228), .B1(n9775), .B2(n18227), .ZN(
        n17918) );
  OAI211_X1 U21116 ( .C1(n17975), .C2(n17920), .A(n17919), .B(n17918), .ZN(
        P3_U2823) );
  OAI21_X1 U21117 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17922), .A(
        n17921), .ZN(n18240) );
  AOI21_X1 U21118 ( .B1(n17925), .B2(n17924), .A(n17923), .ZN(n18237) );
  NAND2_X1 U21119 ( .A1(n17928), .A2(n18704), .ZN(n17926) );
  OAI22_X1 U21120 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17926), .B1(
        n18199), .B2(n18866), .ZN(n17927) );
  AOI21_X1 U21121 ( .B1(n17994), .B2(n18237), .A(n17927), .ZN(n17931) );
  AOI21_X1 U21122 ( .B1(n17928), .B2(n18704), .A(n17991), .ZN(n17944) );
  AOI22_X1 U21123 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17944), .B1(
        n17929), .B2(n17988), .ZN(n17930) );
  OAI211_X1 U21124 ( .C1(n18000), .C2(n18240), .A(n17931), .B(n17930), .ZN(
        P3_U2824) );
  OAI21_X1 U21125 ( .B1(n17934), .B2(n17933), .A(n17932), .ZN(n18247) );
  OAI21_X1 U21126 ( .B1(n17937), .B2(n17936), .A(n17935), .ZN(n17938) );
  XOR2_X1 U21127 ( .A(n17938), .B(n10348), .Z(n18244) );
  AOI22_X1 U21128 ( .A1(n17994), .A2(n18244), .B1(n18235), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17946) );
  OAI21_X1 U21129 ( .B1(n17941), .B2(n17940), .A(n17939), .ZN(n17943) );
  AOI22_X1 U21130 ( .A1(n17944), .A2(n17943), .B1(n17942), .B2(n17988), .ZN(
        n17945) );
  OAI211_X1 U21131 ( .C1(n18000), .C2(n18247), .A(n17946), .B(n17945), .ZN(
        P3_U2825) );
  OAI21_X1 U21132 ( .B1(n17949), .B2(n17948), .A(n17947), .ZN(n17950) );
  XOR2_X1 U21133 ( .A(n17950), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18257) );
  OAI22_X1 U21134 ( .A1(n18000), .A2(n18257), .B1(n18358), .B2(n17951), .ZN(
        n17952) );
  AOI21_X1 U21135 ( .B1(n18301), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17952), .ZN(
        n17958) );
  AOI21_X1 U21136 ( .B1(n17955), .B2(n17954), .A(n17953), .ZN(n18255) );
  OAI21_X1 U21137 ( .B1(n9964), .B2(n17956), .A(n17996), .ZN(n17971) );
  AOI22_X1 U21138 ( .A1(n17994), .A2(n18255), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17971), .ZN(n17957) );
  OAI211_X1 U21139 ( .C1(n17975), .C2(n17959), .A(n17958), .B(n17957), .ZN(
        P3_U2826) );
  OAI21_X1 U21140 ( .B1(n17962), .B2(n17961), .A(n17960), .ZN(n17963) );
  XOR2_X1 U21141 ( .A(n17963), .B(n10344), .Z(n18261) );
  AOI22_X1 U21142 ( .A1(n17994), .A2(n18261), .B1(n18235), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17973) );
  OAI21_X1 U21143 ( .B1(n17966), .B2(n17965), .A(n17964), .ZN(n18258) );
  NAND2_X1 U21144 ( .A1(n17968), .A2(n17967), .ZN(n17969) );
  NAND2_X1 U21145 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17996), .ZN(
        n17980) );
  OAI22_X1 U21146 ( .A1(n18000), .A2(n18258), .B1(n17969), .B2(n17980), .ZN(
        n17970) );
  AOI21_X1 U21147 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17971), .A(
        n17970), .ZN(n17972) );
  OAI211_X1 U21148 ( .C1(n17975), .C2(n17974), .A(n17973), .B(n17972), .ZN(
        P3_U2827) );
  AOI21_X1 U21149 ( .B1(n17978), .B2(n17977), .A(n17976), .ZN(n18273) );
  AOI22_X1 U21150 ( .A1(n17994), .A2(n18273), .B1(n17979), .B2(n17988), .ZN(
        n17983) );
  OAI21_X1 U21151 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18704), .A(
        n17980), .ZN(n17982) );
  NAND2_X1 U21152 ( .A1(n18235), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18284) );
  OAI211_X1 U21153 ( .C1(n18272), .C2(n18271), .A(n9775), .B(n18270), .ZN(
        n17981) );
  NAND4_X1 U21154 ( .A1(n17983), .A2(n17982), .A3(n18284), .A4(n17981), .ZN(
        P3_U2828) );
  NOR2_X1 U21155 ( .A1(n17993), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17984) );
  XNOR2_X1 U21156 ( .A(n17984), .B(n17987), .ZN(n18286) );
  AOI22_X1 U21157 ( .A1(n9775), .A2(n18286), .B1(n18235), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17990) );
  AOI21_X1 U21158 ( .B1(n17992), .B2(n17987), .A(n17986), .ZN(n18288) );
  AOI22_X1 U21159 ( .A1(n17994), .A2(n18288), .B1(n9966), .B2(n17988), .ZN(
        n17989) );
  OAI211_X1 U21160 ( .C1(n17991), .C2(n9966), .A(n17990), .B(n17989), .ZN(
        P3_U2829) );
  OAI21_X1 U21161 ( .B1(n17993), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17992), .ZN(n18304) );
  INV_X1 U21162 ( .A(n18304), .ZN(n18306) );
  INV_X1 U21163 ( .A(n17994), .ZN(n17999) );
  NAND3_X1 U21164 ( .A1(n18937), .A2(n17996), .A3(n17995), .ZN(n17997) );
  AOI22_X1 U21165 ( .A1(n18301), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17997), .ZN(n17998) );
  OAI221_X1 U21166 ( .B1(n18306), .B2(n18000), .C1(n18304), .C2(n17999), .A(
        n17998), .ZN(P3_U2830) );
  INV_X1 U21167 ( .A(n18203), .ZN(n18209) );
  AOI22_X1 U21168 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18291), .B1(
        n18235), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n18011) );
  INV_X1 U21169 ( .A(n9773), .ZN(n18188) );
  NAND2_X1 U21170 ( .A1(n18188), .A2(n18805), .ZN(n18266) );
  INV_X1 U21171 ( .A(n18266), .ZN(n18214) );
  NAND2_X1 U21172 ( .A1(n9773), .A2(n18954), .ZN(n18268) );
  NAND3_X1 U21173 ( .A1(n18100), .A2(n18021), .A3(n18268), .ZN(n18038) );
  OAI21_X1 U21174 ( .B1(n18023), .B2(n18038), .A(n18266), .ZN(n18027) );
  OAI211_X1 U21175 ( .C1(n18002), .C2(n18214), .A(n18027), .B(n18001), .ZN(
        n18003) );
  AOI21_X1 U21176 ( .B1(n18767), .B2(n18004), .A(n18003), .ZN(n18005) );
  OAI21_X1 U21177 ( .B1(n18006), .B2(n18159), .A(n18005), .ZN(n18016) );
  INV_X1 U21178 ( .A(n18075), .ZN(n18047) );
  OAI22_X1 U21179 ( .A1(n18009), .A2(n18289), .B1(n18007), .B2(n18047), .ZN(
        n18008) );
  OAI21_X1 U21180 ( .B1(n18009), .B2(n18016), .A(n18008), .ZN(n18010) );
  OAI211_X1 U21181 ( .C1(n18012), .C2(n18209), .A(n18011), .B(n18010), .ZN(
        P3_U2835) );
  OAI22_X1 U21182 ( .A1(n18013), .A2(n18285), .B1(n18199), .B2(n18905), .ZN(
        n18014) );
  AOI21_X1 U21183 ( .B1(n18203), .B2(n18015), .A(n18014), .ZN(n18018) );
  NAND3_X1 U21184 ( .A1(n18298), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n18016), .ZN(n18017) );
  OAI211_X1 U21185 ( .C1(n18019), .C2(n18047), .A(n18018), .B(n18017), .ZN(
        P3_U2836) );
  AOI21_X1 U21186 ( .B1(n18021), .B2(n18020), .A(n18798), .ZN(n18042) );
  AOI211_X1 U21187 ( .C1(n18780), .C2(n18023), .A(n18042), .B(n18022), .ZN(
        n18028) );
  AOI21_X1 U21188 ( .B1(n18025), .B2(n18024), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18026) );
  AOI211_X1 U21189 ( .C1(n18028), .C2(n18027), .A(n18026), .B(n18289), .ZN(
        n18029) );
  AOI211_X1 U21190 ( .C1(n18291), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18030), .B(n18029), .ZN(n18034) );
  AOI22_X1 U21191 ( .A1(n18287), .A2(n18032), .B1(n18203), .B2(n18031), .ZN(
        n18033) );
  OAI211_X1 U21192 ( .C1(n18036), .C2(n18035), .A(n18034), .B(n18033), .ZN(
        P3_U2837) );
  AOI22_X1 U21193 ( .A1(n18301), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18203), 
        .B2(n18037), .ZN(n18046) );
  AOI22_X1 U21194 ( .A1(n18767), .A2(n18039), .B1(n18266), .B2(n18038), .ZN(
        n18040) );
  OAI211_X1 U21195 ( .C1(n18041), .C2(n18159), .A(n18040), .B(n18285), .ZN(
        n18044) );
  NOR3_X1 U21196 ( .A1(n18042), .A2(n20822), .A3(n18044), .ZN(n18043) );
  NOR2_X1 U21197 ( .A1(n18043), .A2(n18301), .ZN(n18050) );
  OAI211_X1 U21198 ( .C1(n18145), .C2(n18044), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18050), .ZN(n18045) );
  OAI211_X1 U21199 ( .C1(n18048), .C2(n18047), .A(n18046), .B(n18045), .ZN(
        P3_U2838) );
  NOR3_X1 U21200 ( .A1(n18291), .A2(n18056), .A3(n18049), .ZN(n18051) );
  OAI21_X1 U21201 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18051), .A(
        n18050), .ZN(n18053) );
  OAI211_X1 U21202 ( .C1(n18209), .C2(n18054), .A(n18053), .B(n18052), .ZN(
        P3_U2839) );
  AOI221_X1 U21203 ( .B1(n18056), .B2(n18058), .C1(n18055), .C2(n18058), .A(
        n18289), .ZN(n18071) );
  AOI22_X1 U21204 ( .A1(n18767), .A2(n18057), .B1(n18133), .B2(n18132), .ZN(
        n18079) );
  INV_X1 U21205 ( .A(n18122), .ZN(n18078) );
  AOI21_X1 U21206 ( .B1(n18066), .B2(n18078), .A(n18188), .ZN(n18059) );
  AOI211_X1 U21207 ( .C1(n18780), .C2(n18060), .A(n18059), .B(n18058), .ZN(
        n18069) );
  OAI21_X1 U21208 ( .B1(n18062), .B2(n18061), .A(n18780), .ZN(n18102) );
  OAI21_X1 U21209 ( .B1(n18064), .B2(n18063), .A(n18778), .ZN(n18065) );
  OAI211_X1 U21210 ( .C1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n18798), .A(
        n18102), .B(n18065), .ZN(n18080) );
  NAND2_X1 U21211 ( .A1(n18279), .A2(n18159), .ZN(n18182) );
  INV_X1 U21212 ( .A(n18182), .ZN(n18104) );
  OAI22_X1 U21213 ( .A1(n18805), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18066), .B2(n18104), .ZN(n18084) );
  AOI211_X1 U21214 ( .C1(n18067), .C2(n18193), .A(n18080), .B(n18084), .ZN(
        n18068) );
  NAND3_X1 U21215 ( .A1(n18079), .A2(n18069), .A3(n18068), .ZN(n18070) );
  AOI22_X1 U21216 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18291), .B1(
        n18071), .B2(n18070), .ZN(n18073) );
  OAI211_X1 U21217 ( .C1(n18074), .C2(n18209), .A(n18073), .B(n18072), .ZN(
        P3_U2840) );
  NAND2_X1 U21218 ( .A1(n18075), .A2(n18077), .ZN(n18099) );
  AOI22_X1 U21219 ( .A1(n18301), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18203), 
        .B2(n18076), .ZN(n18086) );
  AOI21_X1 U21220 ( .B1(n18078), .B2(n18077), .A(n18188), .ZN(n18081) );
  NAND2_X1 U21221 ( .A1(n18298), .A2(n18079), .ZN(n18124) );
  NOR3_X1 U21222 ( .A1(n18081), .A2(n18124), .A3(n18080), .ZN(n18090) );
  OAI21_X1 U21223 ( .B1(n18290), .B2(n18082), .A(n18090), .ZN(n18083) );
  OAI211_X1 U21224 ( .C1(n18084), .C2(n18083), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18199), .ZN(n18085) );
  OAI211_X1 U21225 ( .C1(n18087), .C2(n18099), .A(n18086), .B(n18085), .ZN(
        P3_U2841) );
  AOI22_X1 U21226 ( .A1(n18301), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18203), 
        .B2(n18088), .ZN(n18093) );
  AOI221_X1 U21227 ( .B1(n18104), .B2(n18090), .C1(n18089), .C2(n18090), .A(
        n18301), .ZN(n18096) );
  NOR3_X1 U21228 ( .A1(n18290), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n18986), .ZN(n18091) );
  OAI21_X1 U21229 ( .B1(n18096), .B2(n18091), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18092) );
  OAI211_X1 U21230 ( .C1(n18094), .C2(n18099), .A(n18093), .B(n18092), .ZN(
        P3_U2842) );
  AOI22_X1 U21231 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18096), .B1(
        n18203), .B2(n18095), .ZN(n18098) );
  OAI211_X1 U21232 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18099), .A(
        n18098), .B(n18097), .ZN(P3_U2843) );
  NAND2_X1 U21233 ( .A1(n18100), .A2(n18268), .ZN(n18101) );
  AOI221_X1 U21234 ( .B1(n18125), .B2(n18266), .C1(n18101), .C2(n18266), .A(
        n18124), .ZN(n18103) );
  OAI211_X1 U21235 ( .C1(n18105), .C2(n18104), .A(n18103), .B(n18102), .ZN(
        n18116) );
  OAI221_X1 U21236 ( .B1(n18116), .B2(n18106), .C1(n18116), .C2(n18266), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18114) );
  INV_X1 U21237 ( .A(n18107), .ZN(n18108) );
  OAI22_X1 U21238 ( .A1(n18275), .A2(n18798), .B1(n18248), .B2(n18276), .ZN(
        n18263) );
  NAND2_X1 U21239 ( .A1(n18108), .A2(n18263), .ZN(n18219) );
  NOR2_X1 U21240 ( .A1(n18109), .A2(n18219), .ZN(n18171) );
  OAI21_X1 U21241 ( .B1(n18171), .B2(n18170), .A(n18298), .ZN(n18207) );
  NOR2_X1 U21242 ( .A1(n18110), .A2(n18207), .ZN(n18126) );
  AOI22_X1 U21243 ( .A1(n18203), .A2(n18112), .B1(n18126), .B2(n18111), .ZN(
        n18113) );
  OAI221_X1 U21244 ( .B1(n18301), .B2(n18114), .C1(n18199), .C2(n20989), .A(
        n18113), .ZN(P3_U2844) );
  AOI22_X1 U21245 ( .A1(n18301), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18126), 
        .B2(n18115), .ZN(n18118) );
  NAND3_X1 U21246 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18199), .A3(
        n18116), .ZN(n18117) );
  OAI211_X1 U21247 ( .C1(n18119), .C2(n18209), .A(n18118), .B(n18117), .ZN(
        P3_U2845) );
  AOI22_X1 U21248 ( .A1(n18780), .A2(n18121), .B1(n18778), .B2(n18120), .ZN(
        n18158) );
  OAI21_X1 U21249 ( .B1(n18143), .B2(n9773), .A(n18122), .ZN(n18123) );
  OAI211_X1 U21250 ( .C1(n18131), .C2(n18186), .A(n18158), .B(n18123), .ZN(
        n18130) );
  OAI221_X1 U21251 ( .B1(n18124), .B2(n18145), .C1(n18124), .C2(n18130), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18129) );
  INV_X1 U21252 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18886) );
  AOI22_X1 U21253 ( .A1(n18127), .A2(n18203), .B1(n18126), .B2(n18125), .ZN(
        n18128) );
  OAI221_X1 U21254 ( .B1(n18301), .B2(n18129), .C1(n18199), .C2(n18886), .A(
        n18128), .ZN(P3_U2846) );
  OAI221_X1 U21255 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18131), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18171), .A(n18130), .ZN(
        n18136) );
  OAI211_X1 U21256 ( .C1(n18134), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18133), .B(n18132), .ZN(n18135) );
  OAI211_X1 U21257 ( .C1(n18138), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        n18140) );
  AOI22_X1 U21258 ( .A1(n18298), .A2(n18140), .B1(n18287), .B2(n18139), .ZN(
        n18142) );
  OAI211_X1 U21259 ( .C1(n18285), .C2(n18143), .A(n18142), .B(n18141), .ZN(
        P3_U2847) );
  NOR2_X1 U21260 ( .A1(n18199), .A2(n18883), .ZN(n18150) );
  NOR2_X1 U21261 ( .A1(n18188), .A2(n18185), .ZN(n18201) );
  AOI211_X1 U21262 ( .C1(n18145), .C2(n18144), .A(n18201), .B(n10354), .ZN(
        n18148) );
  AOI21_X1 U21263 ( .B1(n18171), .B2(n18146), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18147) );
  AOI211_X1 U21264 ( .C1(n18158), .C2(n18148), .A(n18147), .B(n18289), .ZN(
        n18149) );
  AOI211_X1 U21265 ( .C1(n18291), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18150), .B(n18149), .ZN(n18155) );
  INV_X1 U21266 ( .A(n18151), .ZN(n18152) );
  AOI22_X1 U21267 ( .A1(n18212), .A2(n18153), .B1(n18203), .B2(n18152), .ZN(
        n18154) );
  OAI211_X1 U21268 ( .C1(n18305), .C2(n18156), .A(n18155), .B(n18154), .ZN(
        P3_U2848) );
  AOI22_X1 U21269 ( .A1(n18301), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18203), 
        .B2(n18157), .ZN(n18167) );
  OAI21_X1 U21270 ( .B1(n18160), .B2(n18159), .A(n18158), .ZN(n18161) );
  AOI21_X1 U21271 ( .B1(n18767), .B2(n18162), .A(n18161), .ZN(n18181) );
  OAI22_X1 U21272 ( .A1(n18163), .A2(n18201), .B1(n18182), .B2(n9773), .ZN(
        n18164) );
  OAI211_X1 U21273 ( .C1(n18187), .C2(n18186), .A(n18181), .B(n18164), .ZN(
        n18174) );
  OAI21_X1 U21274 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18186), .A(
        n18285), .ZN(n18165) );
  OAI211_X1 U21275 ( .C1(n18174), .C2(n18165), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18199), .ZN(n18166) );
  OAI211_X1 U21276 ( .C1(n18207), .C2(n18168), .A(n18167), .B(n18166), .ZN(
        P3_U2849) );
  AOI22_X1 U21277 ( .A1(n18301), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18203), 
        .B2(n18169), .ZN(n18177) );
  NOR2_X1 U21278 ( .A1(n18171), .A2(n18170), .ZN(n18173) );
  NOR2_X1 U21279 ( .A1(n18173), .A2(n18172), .ZN(n18175) );
  OAI221_X1 U21280 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18175), 
        .C1(n18178), .C2(n18174), .A(n18298), .ZN(n18176) );
  OAI211_X1 U21281 ( .C1(n18285), .C2(n18178), .A(n18177), .B(n18176), .ZN(
        P3_U2850) );
  AOI22_X1 U21282 ( .A1(n18301), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18203), 
        .B2(n18179), .ZN(n18191) );
  INV_X1 U21283 ( .A(n18180), .ZN(n18183) );
  NAND2_X1 U21284 ( .A1(n18298), .A2(n18181), .ZN(n18200) );
  AOI21_X1 U21285 ( .B1(n18183), .B2(n18182), .A(n18200), .ZN(n18184) );
  OAI221_X1 U21286 ( .B1(n18188), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18188), .C2(n18185), .A(n18184), .ZN(n18194) );
  OAI22_X1 U21287 ( .A1(n18188), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18187), .B2(n18186), .ZN(n18189) );
  OAI211_X1 U21288 ( .C1(n18194), .C2(n18189), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18199), .ZN(n18190) );
  OAI211_X1 U21289 ( .C1(n18192), .C2(n18207), .A(n18191), .B(n18190), .ZN(
        P3_U2851) );
  OAI221_X1 U21290 ( .B1(n18194), .B2(n18206), .C1(n18194), .C2(n18193), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18198) );
  NOR2_X1 U21291 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18207), .ZN(
        n18196) );
  AOI22_X1 U21292 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18196), .B1(
        n18203), .B2(n18195), .ZN(n18197) );
  OAI221_X1 U21293 ( .B1(n18301), .B2(n18198), .C1(n18199), .C2(n18874), .A(
        n18197), .ZN(P3_U2852) );
  OAI21_X1 U21294 ( .B1(n18201), .B2(n18200), .A(n18199), .ZN(n18205) );
  AOI22_X1 U21295 ( .A1(n18301), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18203), 
        .B2(n18202), .ZN(n18204) );
  OAI221_X1 U21296 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18207), .C1(
        n18206), .C2(n18205), .A(n18204), .ZN(P3_U2853) );
  OAI22_X1 U21297 ( .A1(n18305), .A2(n18210), .B1(n18209), .B2(n18208), .ZN(
        n18211) );
  AOI21_X1 U21298 ( .B1(n18213), .B2(n18212), .A(n18211), .ZN(n18225) );
  OAI21_X1 U21299 ( .B1(n18215), .B2(n18214), .A(n18268), .ZN(n18216) );
  AOI21_X1 U21300 ( .B1(n18780), .B2(n18217), .A(n18216), .ZN(n18234) );
  OAI211_X1 U21301 ( .C1(n18218), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18234), .ZN(n18229) );
  OAI221_X1 U21302 ( .B1(n18291), .B2(n18292), .C1(n18291), .C2(n18229), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18223) );
  NOR2_X1 U21303 ( .A1(n18220), .A2(n18219), .ZN(n18230) );
  NAND4_X1 U21304 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18298), .A3(
        n18230), .A4(n18221), .ZN(n18222) );
  NAND4_X1 U21305 ( .A1(n18225), .A2(n18224), .A3(n18223), .A4(n18222), .ZN(
        P3_U2854) );
  AOI21_X1 U21306 ( .B1(n18291), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18226), .ZN(n18233) );
  AOI22_X1 U21307 ( .A1(n18297), .A2(n18228), .B1(n18287), .B2(n18227), .ZN(
        n18232) );
  OAI211_X1 U21308 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18230), .A(
        n18298), .B(n18229), .ZN(n18231) );
  NAND3_X1 U21309 ( .A1(n18233), .A2(n18232), .A3(n18231), .ZN(P3_U2855) );
  OAI21_X1 U21310 ( .B1(n18234), .B2(n18289), .A(n18285), .ZN(n18241) );
  AOI22_X1 U21311 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18241), .B1(
        n18235), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18239) );
  NAND3_X1 U21312 ( .A1(n18298), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18263), .ZN(n18251) );
  NOR4_X1 U21313 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18250), .A3(
        n10348), .A4(n18251), .ZN(n18236) );
  AOI21_X1 U21314 ( .B1(n18237), .B2(n18297), .A(n18236), .ZN(n18238) );
  OAI211_X1 U21315 ( .C1(n18305), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        P3_U2856) );
  NOR2_X1 U21316 ( .A1(n18250), .A2(n18251), .ZN(n18242) );
  MUX2_X1 U21317 ( .A(n18242), .B(n18241), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18243) );
  AOI21_X1 U21318 ( .B1(n18297), .B2(n18244), .A(n18243), .ZN(n18246) );
  NAND2_X1 U21319 ( .A1(n18301), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18245) );
  OAI211_X1 U21320 ( .C1(n18247), .C2(n18305), .A(n18246), .B(n18245), .ZN(
        P3_U2857) );
  NOR2_X1 U21321 ( .A1(n18199), .A2(n18862), .ZN(n18254) );
  AOI22_X1 U21322 ( .A1(n18780), .A2(n18275), .B1(n18248), .B2(n18266), .ZN(
        n18249) );
  NAND3_X1 U21323 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18249), .A3(
        n18268), .ZN(n18262) );
  AOI21_X1 U21324 ( .B1(n18292), .B2(n18262), .A(n18291), .ZN(n18252) );
  AOI22_X1 U21325 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18252), .B1(
        n18251), .B2(n18250), .ZN(n18253) );
  AOI211_X1 U21326 ( .C1(n18255), .C2(n18297), .A(n18254), .B(n18253), .ZN(
        n18256) );
  OAI21_X1 U21327 ( .B1(n18305), .B2(n18257), .A(n18256), .ZN(P3_U2858) );
  INV_X1 U21328 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18861) );
  NOR2_X1 U21329 ( .A1(n18199), .A2(n18861), .ZN(n18260) );
  OAI22_X1 U21330 ( .A1(n10344), .A2(n18285), .B1(n18305), .B2(n18258), .ZN(
        n18259) );
  AOI211_X1 U21331 ( .C1(n18297), .C2(n18261), .A(n18260), .B(n18259), .ZN(
        n18265) );
  OAI211_X1 U21332 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18263), .A(
        n18298), .B(n18262), .ZN(n18264) );
  NAND2_X1 U21333 ( .A1(n18265), .A2(n18264), .ZN(P3_U2859) );
  NOR2_X1 U21334 ( .A1(n18938), .A2(n18954), .ZN(n18267) );
  AOI22_X1 U21335 ( .A1(n18780), .A2(n18267), .B1(n18938), .B2(n18266), .ZN(
        n18269) );
  AOI21_X1 U21336 ( .B1(n18269), .B2(n18268), .A(n20943), .ZN(n18282) );
  OAI21_X1 U21337 ( .B1(n18272), .B2(n18271), .A(n18270), .ZN(n18280) );
  AOI22_X1 U21338 ( .A1(n18780), .A2(n18275), .B1(n18274), .B2(n18273), .ZN(
        n18278) );
  OR3_X1 U21339 ( .A1(n18938), .A2(n18276), .A3(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18277) );
  OAI211_X1 U21340 ( .C1(n18280), .C2(n18279), .A(n18278), .B(n18277), .ZN(
        n18281) );
  OAI21_X1 U21341 ( .B1(n18282), .B2(n18281), .A(n18298), .ZN(n18283) );
  OAI211_X1 U21342 ( .C1(n18285), .C2(n20943), .A(n18284), .B(n18283), .ZN(
        P3_U2860) );
  AOI22_X1 U21343 ( .A1(n18297), .A2(n18288), .B1(n18287), .B2(n18286), .ZN(
        n18296) );
  NAND2_X1 U21344 ( .A1(n18301), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18295) );
  NOR3_X1 U21345 ( .A1(n18290), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18289), .ZN(n18299) );
  OAI21_X1 U21346 ( .B1(n18291), .B2(n18299), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18294) );
  OAI211_X1 U21347 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18778), .A(
        n18292), .B(n18938), .ZN(n18293) );
  NAND4_X1 U21348 ( .A1(n18296), .A2(n18295), .A3(n18294), .A4(n18293), .ZN(
        P3_U2861) );
  INV_X1 U21349 ( .A(n18297), .ZN(n18303) );
  AOI21_X1 U21350 ( .B1(n18805), .B2(n18298), .A(n18954), .ZN(n18300) );
  AOI221_X1 U21351 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18301), .C1(n18300), 
        .C2(n18199), .A(n18299), .ZN(n18302) );
  OAI221_X1 U21352 ( .B1(n18306), .B2(n18305), .C1(n18304), .C2(n18303), .A(
        n18302), .ZN(P3_U2862) );
  AOI21_X1 U21353 ( .B1(n18309), .B2(n18308), .A(n18307), .ZN(n18828) );
  OAI21_X1 U21354 ( .B1(n18828), .B2(n18366), .A(n18314), .ZN(n18310) );
  OAI221_X1 U21355 ( .B1(n18565), .B2(n18976), .C1(n18565), .C2(n18314), .A(
        n18310), .ZN(P3_U2863) );
  INV_X1 U21356 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18817) );
  NAND2_X1 U21357 ( .A1(n18814), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18595) );
  INV_X1 U21358 ( .A(n18595), .ZN(n18544) );
  NAND2_X1 U21359 ( .A1(n18817), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18498) );
  INV_X1 U21360 ( .A(n18498), .ZN(n18500) );
  NOR2_X1 U21361 ( .A1(n18544), .A2(n18500), .ZN(n18312) );
  OAI22_X1 U21362 ( .A1(n18313), .A2(n18817), .B1(n18312), .B2(n18311), .ZN(
        P3_U2866) );
  NOR2_X1 U21363 ( .A1(n18818), .A2(n18314), .ZN(P3_U2867) );
  NOR2_X1 U21364 ( .A1(n18814), .A2(n18817), .ZN(n18640) );
  NOR2_X1 U21365 ( .A1(n18565), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18543) );
  NAND2_X1 U21366 ( .A1(n18640), .A2(n18543), .ZN(n18665) );
  INV_X1 U21367 ( .A(n18665), .ZN(n18757) );
  NOR2_X1 U21368 ( .A1(n18817), .A2(n18474), .ZN(n18705) );
  NAND2_X1 U21369 ( .A1(n18565), .A2(n18705), .ZN(n18701) );
  INV_X1 U21370 ( .A(n18701), .ZN(n18676) );
  NOR2_X1 U21371 ( .A1(n18757), .A2(n18676), .ZN(n18671) );
  NAND2_X1 U21372 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18808) );
  INV_X1 U21373 ( .A(n18640), .ZN(n18643) );
  NAND2_X1 U21374 ( .A1(n18809), .A2(n18565), .ZN(n18810) );
  NOR2_X1 U21375 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18410) );
  INV_X1 U21376 ( .A(n18410), .ZN(n18408) );
  NOR2_X1 U21377 ( .A1(n18810), .A2(n18408), .ZN(n18427) );
  NOR2_X1 U21378 ( .A1(n18761), .A2(n18423), .ZN(n18387) );
  INV_X1 U21379 ( .A(n18367), .ZN(n18675) );
  OAI21_X1 U21380 ( .B1(n18565), .B2(n21062), .A(n18675), .ZN(n18566) );
  OAI22_X1 U21381 ( .A1(n18671), .A2(n18358), .B1(n18387), .B2(n18566), .ZN(
        n18364) );
  INV_X1 U21382 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18315) );
  NOR2_X2 U21383 ( .A1(n18358), .A2(n18315), .ZN(n18710) );
  NOR2_X2 U21384 ( .A1(n18367), .A2(n20888), .ZN(n18707) );
  NOR2_X1 U21385 ( .A1(n18834), .A2(n18387), .ZN(n18357) );
  AOI22_X1 U21386 ( .A1(n18676), .A2(n18710), .B1(n18707), .B2(n18357), .ZN(
        n18321) );
  NOR2_X2 U21387 ( .A1(n18316), .A2(n18358), .ZN(n18708) );
  NAND2_X1 U21388 ( .A1(n18318), .A2(n18317), .ZN(n18360) );
  NOR2_X1 U21389 ( .A1(n18319), .A2(n18360), .ZN(n18709) );
  AOI22_X1 U21390 ( .A1(n18757), .A2(n18708), .B1(n18423), .B2(n18709), .ZN(
        n18320) );
  OAI211_X1 U21391 ( .C1(n18322), .C2(n18364), .A(n18321), .B(n18320), .ZN(
        P3_U2868) );
  AND2_X1 U21392 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18704), .ZN(n18714) );
  AND2_X1 U21393 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18675), .ZN(n18715) );
  AOI22_X1 U21394 ( .A1(n18757), .A2(n18714), .B1(n18357), .B2(n18715), .ZN(
        n18326) );
  INV_X1 U21395 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18323) );
  NOR2_X2 U21396 ( .A1(n18323), .A2(n18358), .ZN(n18716) );
  NOR2_X1 U21397 ( .A1(n18324), .A2(n18360), .ZN(n18647) );
  AOI22_X1 U21398 ( .A1(n18676), .A2(n18716), .B1(n18423), .B2(n18647), .ZN(
        n18325) );
  OAI211_X1 U21399 ( .C1(n18327), .C2(n18364), .A(n18326), .B(n18325), .ZN(
        P3_U2869) );
  NOR2_X2 U21400 ( .A1(n18328), .A2(n18358), .ZN(n18721) );
  NOR2_X2 U21401 ( .A1(n18329), .A2(n18367), .ZN(n18720) );
  AOI22_X1 U21402 ( .A1(n18757), .A2(n18721), .B1(n18357), .B2(n18720), .ZN(
        n18332) );
  AND2_X1 U21403 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18704), .ZN(n18723) );
  NOR2_X1 U21404 ( .A1(n18330), .A2(n18360), .ZN(n18722) );
  AOI22_X1 U21405 ( .A1(n18676), .A2(n18723), .B1(n18427), .B2(n18722), .ZN(
        n18331) );
  OAI211_X1 U21406 ( .C1(n18333), .C2(n18364), .A(n18332), .B(n18331), .ZN(
        P3_U2870) );
  AND2_X1 U21407 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n18704), .ZN(n18729) );
  NOR2_X2 U21408 ( .A1(n18334), .A2(n18367), .ZN(n18727) );
  AOI22_X1 U21409 ( .A1(n18676), .A2(n18729), .B1(n18357), .B2(n18727), .ZN(
        n18337) );
  INV_X1 U21410 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19419) );
  NOR2_X2 U21411 ( .A1(n19419), .A2(n18358), .ZN(n18728) );
  NOR2_X1 U21412 ( .A1(n18335), .A2(n18360), .ZN(n18653) );
  AOI22_X1 U21413 ( .A1(n18757), .A2(n18728), .B1(n18427), .B2(n18653), .ZN(
        n18336) );
  OAI211_X1 U21414 ( .C1(n18338), .C2(n18364), .A(n18337), .B(n18336), .ZN(
        P3_U2871) );
  NOR2_X2 U21415 ( .A1(n20975), .A2(n18358), .ZN(n18735) );
  NOR2_X2 U21416 ( .A1(n18339), .A2(n18367), .ZN(n18733) );
  AOI22_X1 U21417 ( .A1(n18757), .A2(n18735), .B1(n18357), .B2(n18733), .ZN(
        n18343) );
  INV_X1 U21418 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18340) );
  NOR2_X2 U21419 ( .A1(n18340), .A2(n18358), .ZN(n18734) );
  NOR2_X1 U21420 ( .A1(n18341), .A2(n18360), .ZN(n18736) );
  AOI22_X1 U21421 ( .A1(n18676), .A2(n18734), .B1(n18427), .B2(n18736), .ZN(
        n18342) );
  OAI211_X1 U21422 ( .C1(n18344), .C2(n18364), .A(n18343), .B(n18342), .ZN(
        P3_U2872) );
  NOR2_X2 U21423 ( .A1(n18345), .A2(n18358), .ZN(n18742) );
  NOR2_X2 U21424 ( .A1(n18346), .A2(n18367), .ZN(n18740) );
  AOI22_X1 U21425 ( .A1(n18676), .A2(n18742), .B1(n18357), .B2(n18740), .ZN(
        n18349) );
  AND2_X1 U21426 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18704), .ZN(n18741) );
  NOR2_X1 U21427 ( .A1(n9752), .A2(n18360), .ZN(n18581) );
  AOI22_X1 U21428 ( .A1(n18757), .A2(n18741), .B1(n18427), .B2(n18581), .ZN(
        n18348) );
  OAI211_X1 U21429 ( .C1(n20925), .C2(n18364), .A(n18349), .B(n18348), .ZN(
        P3_U2873) );
  NOR2_X2 U21430 ( .A1(n18350), .A2(n18358), .ZN(n18748) );
  NOR2_X2 U21431 ( .A1(n18351), .A2(n18367), .ZN(n18749) );
  AOI22_X1 U21432 ( .A1(n18757), .A2(n18748), .B1(n18357), .B2(n18749), .ZN(
        n18354) );
  AND2_X1 U21433 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18704), .ZN(n18751) );
  NOR2_X1 U21434 ( .A1(n18352), .A2(n18360), .ZN(n18750) );
  AOI22_X1 U21435 ( .A1(n18676), .A2(n18751), .B1(n18427), .B2(n18750), .ZN(
        n18353) );
  OAI211_X1 U21436 ( .C1(n18355), .C2(n18364), .A(n18354), .B(n18353), .ZN(
        P3_U2874) );
  AND2_X1 U21437 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18704), .ZN(n18756) );
  NOR2_X2 U21438 ( .A1(n18356), .A2(n18367), .ZN(n18755) );
  AOI22_X1 U21439 ( .A1(n18676), .A2(n18756), .B1(n18357), .B2(n18755), .ZN(
        n18363) );
  NOR2_X2 U21440 ( .A1(n18359), .A2(n18358), .ZN(n18759) );
  NOR2_X1 U21441 ( .A1(n18361), .A2(n18360), .ZN(n18760) );
  AOI22_X1 U21442 ( .A1(n18757), .A2(n18759), .B1(n18427), .B2(n18760), .ZN(
        n18362) );
  OAI211_X1 U21443 ( .C1(n18365), .C2(n18364), .A(n18363), .B(n18362), .ZN(
        P3_U2875) );
  NAND2_X1 U21444 ( .A1(n18543), .A2(n18410), .ZN(n18386) );
  NAND2_X1 U21445 ( .A1(n18809), .A2(n18706), .ZN(n18642) );
  NOR2_X1 U21446 ( .A1(n18408), .A2(n18642), .ZN(n18382) );
  AOI22_X1 U21447 ( .A1(n18676), .A2(n18708), .B1(n18707), .B2(n18382), .ZN(
        n18369) );
  NOR2_X1 U21448 ( .A1(n18367), .A2(n18366), .ZN(n18702) );
  INV_X1 U21449 ( .A(n18702), .ZN(n18409) );
  NOR2_X1 U21450 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18409), .ZN(
        n18639) );
  AOI22_X1 U21451 ( .A1(n18704), .A2(n18705), .B1(n18410), .B2(n18639), .ZN(
        n18383) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18383), .B1(
        n18761), .B2(n18710), .ZN(n18368) );
  OAI211_X1 U21453 ( .C1(n18679), .C2(n18386), .A(n18369), .B(n18368), .ZN(
        P3_U2876) );
  INV_X1 U21454 ( .A(n18647), .ZN(n18719) );
  AOI22_X1 U21455 ( .A1(n18761), .A2(n18716), .B1(n18715), .B2(n18382), .ZN(
        n18371) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18383), .B1(
        n18676), .B2(n18714), .ZN(n18370) );
  OAI211_X1 U21457 ( .C1(n18719), .C2(n18386), .A(n18371), .B(n18370), .ZN(
        P3_U2877) );
  AOI22_X1 U21458 ( .A1(n18761), .A2(n18723), .B1(n18720), .B2(n18382), .ZN(
        n18373) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18383), .B1(
        n18676), .B2(n18721), .ZN(n18372) );
  OAI211_X1 U21460 ( .C1(n18684), .C2(n18386), .A(n18373), .B(n18372), .ZN(
        P3_U2878) );
  INV_X1 U21461 ( .A(n18653), .ZN(n18732) );
  AOI22_X1 U21462 ( .A1(n18761), .A2(n18729), .B1(n18727), .B2(n18382), .ZN(
        n18375) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18383), .B1(
        n18676), .B2(n18728), .ZN(n18374) );
  OAI211_X1 U21464 ( .C1(n18732), .C2(n18386), .A(n18375), .B(n18374), .ZN(
        P3_U2879) );
  INV_X1 U21465 ( .A(n18736), .ZN(n18689) );
  AOI22_X1 U21466 ( .A1(n18676), .A2(n18735), .B1(n18733), .B2(n18382), .ZN(
        n18377) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18383), .B1(
        n18761), .B2(n18734), .ZN(n18376) );
  OAI211_X1 U21468 ( .C1(n18689), .C2(n18386), .A(n18377), .B(n18376), .ZN(
        P3_U2880) );
  AOI22_X1 U21469 ( .A1(n18761), .A2(n18742), .B1(n18740), .B2(n18382), .ZN(
        n18379) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18383), .B1(
        n18676), .B2(n18741), .ZN(n18378) );
  OAI211_X1 U21471 ( .C1(n18746), .C2(n18386), .A(n18379), .B(n18378), .ZN(
        P3_U2881) );
  INV_X1 U21472 ( .A(n18750), .ZN(n18694) );
  AOI22_X1 U21473 ( .A1(n18761), .A2(n18751), .B1(n18749), .B2(n18382), .ZN(
        n18381) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18383), .B1(
        n18676), .B2(n18748), .ZN(n18380) );
  OAI211_X1 U21475 ( .C1(n18694), .C2(n18386), .A(n18381), .B(n18380), .ZN(
        P3_U2882) );
  INV_X1 U21476 ( .A(n18760), .ZN(n18700) );
  AOI22_X1 U21477 ( .A1(n18761), .A2(n18756), .B1(n18755), .B2(n18382), .ZN(
        n18385) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18383), .B1(
        n18676), .B2(n18759), .ZN(n18384) );
  OAI211_X1 U21479 ( .C1(n18700), .C2(n18386), .A(n18385), .B(n18384), .ZN(
        P3_U2883) );
  NOR2_X1 U21480 ( .A1(n18809), .A2(n18408), .ZN(n18454) );
  NAND2_X1 U21481 ( .A1(n18454), .A2(n18565), .ZN(n18407) );
  INV_X1 U21482 ( .A(n18386), .ZN(n18449) );
  NOR2_X1 U21483 ( .A1(n18449), .A2(n18470), .ZN(n18432) );
  OAI21_X1 U21484 ( .B1(n18387), .B2(n18672), .A(n18432), .ZN(n18388) );
  OAI211_X1 U21485 ( .C1(n18470), .C2(n21062), .A(n18675), .B(n18388), .ZN(
        n18404) );
  NOR2_X1 U21486 ( .A1(n18834), .A2(n18432), .ZN(n18403) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18404), .B1(
        n18707), .B2(n18403), .ZN(n18390) );
  AOI22_X1 U21488 ( .A1(n18761), .A2(n18708), .B1(n18423), .B2(n18710), .ZN(
        n18389) );
  OAI211_X1 U21489 ( .C1(n18679), .C2(n18407), .A(n18390), .B(n18389), .ZN(
        P3_U2884) );
  AOI22_X1 U21490 ( .A1(n18761), .A2(n18714), .B1(n18715), .B2(n18403), .ZN(
        n18392) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18404), .B1(
        n18427), .B2(n18716), .ZN(n18391) );
  OAI211_X1 U21492 ( .C1(n18719), .C2(n18407), .A(n18392), .B(n18391), .ZN(
        P3_U2885) );
  AOI22_X1 U21493 ( .A1(n18761), .A2(n18721), .B1(n18720), .B2(n18403), .ZN(
        n18394) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18404), .B1(
        n18427), .B2(n18723), .ZN(n18393) );
  OAI211_X1 U21495 ( .C1(n18684), .C2(n18407), .A(n18394), .B(n18393), .ZN(
        P3_U2886) );
  AOI22_X1 U21496 ( .A1(n18761), .A2(n18728), .B1(n18727), .B2(n18403), .ZN(
        n18396) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18404), .B1(
        n18427), .B2(n18729), .ZN(n18395) );
  OAI211_X1 U21498 ( .C1(n18732), .C2(n18407), .A(n18396), .B(n18395), .ZN(
        P3_U2887) );
  AOI22_X1 U21499 ( .A1(n18761), .A2(n18735), .B1(n18733), .B2(n18403), .ZN(
        n18398) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18404), .B1(
        n18427), .B2(n18734), .ZN(n18397) );
  OAI211_X1 U21501 ( .C1(n18689), .C2(n18407), .A(n18398), .B(n18397), .ZN(
        P3_U2888) );
  AOI22_X1 U21502 ( .A1(n18423), .A2(n18742), .B1(n18740), .B2(n18403), .ZN(
        n18400) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18404), .B1(
        n18761), .B2(n18741), .ZN(n18399) );
  OAI211_X1 U21504 ( .C1(n18746), .C2(n18407), .A(n18400), .B(n18399), .ZN(
        P3_U2889) );
  AOI22_X1 U21505 ( .A1(n18761), .A2(n18748), .B1(n18749), .B2(n18403), .ZN(
        n18402) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18404), .B1(
        n18423), .B2(n18751), .ZN(n18401) );
  OAI211_X1 U21507 ( .C1(n18694), .C2(n18407), .A(n18402), .B(n18401), .ZN(
        P3_U2890) );
  AOI22_X1 U21508 ( .A1(n18423), .A2(n18756), .B1(n18755), .B2(n18403), .ZN(
        n18406) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18404), .B1(
        n18761), .B2(n18759), .ZN(n18405) );
  OAI211_X1 U21510 ( .C1(n18700), .C2(n18407), .A(n18406), .B(n18405), .ZN(
        P3_U2891) );
  NOR2_X2 U21511 ( .A1(n18808), .A2(n18408), .ZN(n18493) );
  INV_X1 U21512 ( .A(n18493), .ZN(n18431) );
  AND2_X1 U21513 ( .A1(n18706), .A2(n18454), .ZN(n18426) );
  AOI22_X1 U21514 ( .A1(n18710), .A2(n18449), .B1(n18707), .B2(n18426), .ZN(
        n18412) );
  AOI21_X1 U21515 ( .B1(n18809), .B2(n18672), .A(n18409), .ZN(n18499) );
  NAND2_X1 U21516 ( .A1(n18410), .A2(n18499), .ZN(n18428) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18428), .B1(
        n18423), .B2(n18708), .ZN(n18411) );
  OAI211_X1 U21518 ( .C1(n18679), .C2(n18431), .A(n18412), .B(n18411), .ZN(
        P3_U2892) );
  AOI22_X1 U21519 ( .A1(n18423), .A2(n18714), .B1(n18715), .B2(n18426), .ZN(
        n18414) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18428), .B1(
        n18716), .B2(n18449), .ZN(n18413) );
  OAI211_X1 U21521 ( .C1(n18719), .C2(n18431), .A(n18414), .B(n18413), .ZN(
        P3_U2893) );
  AOI22_X1 U21522 ( .A1(n18723), .A2(n18449), .B1(n18720), .B2(n18426), .ZN(
        n18416) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18428), .B1(
        n18423), .B2(n18721), .ZN(n18415) );
  OAI211_X1 U21524 ( .C1(n18684), .C2(n18431), .A(n18416), .B(n18415), .ZN(
        P3_U2894) );
  AOI22_X1 U21525 ( .A1(n18729), .A2(n18449), .B1(n18727), .B2(n18426), .ZN(
        n18418) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18428), .B1(
        n18423), .B2(n18728), .ZN(n18417) );
  OAI211_X1 U21527 ( .C1(n18732), .C2(n18431), .A(n18418), .B(n18417), .ZN(
        P3_U2895) );
  AOI22_X1 U21528 ( .A1(n18734), .A2(n18449), .B1(n18733), .B2(n18426), .ZN(
        n18420) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18428), .B1(
        n18423), .B2(n18735), .ZN(n18419) );
  OAI211_X1 U21530 ( .C1(n18689), .C2(n18431), .A(n18420), .B(n18419), .ZN(
        P3_U2896) );
  AOI22_X1 U21531 ( .A1(n18740), .A2(n18426), .B1(n18742), .B2(n18449), .ZN(
        n18422) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18428), .B1(
        n18423), .B2(n18741), .ZN(n18421) );
  OAI211_X1 U21533 ( .C1(n18746), .C2(n18431), .A(n18422), .B(n18421), .ZN(
        P3_U2897) );
  AOI22_X1 U21534 ( .A1(n18423), .A2(n18748), .B1(n18749), .B2(n18426), .ZN(
        n18425) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18428), .B1(
        n18751), .B2(n18449), .ZN(n18424) );
  OAI211_X1 U21536 ( .C1(n18694), .C2(n18431), .A(n18425), .B(n18424), .ZN(
        P3_U2898) );
  AOI22_X1 U21537 ( .A1(n18756), .A2(n18449), .B1(n18755), .B2(n18426), .ZN(
        n18430) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18428), .B1(
        n18427), .B2(n18759), .ZN(n18429) );
  OAI211_X1 U21539 ( .C1(n18700), .C2(n18431), .A(n18430), .B(n18429), .ZN(
        P3_U2899) );
  NOR2_X2 U21540 ( .A1(n18810), .A2(n18498), .ZN(n18516) );
  INV_X1 U21541 ( .A(n18516), .ZN(n18453) );
  NOR2_X1 U21542 ( .A1(n18493), .A2(n18516), .ZN(n18476) );
  NOR2_X1 U21543 ( .A1(n18834), .A2(n18476), .ZN(n18448) );
  AOI22_X1 U21544 ( .A1(n18708), .A2(n18449), .B1(n18707), .B2(n18448), .ZN(
        n18435) );
  OAI21_X1 U21545 ( .B1(n18432), .B2(n18672), .A(n18476), .ZN(n18433) );
  OAI211_X1 U21546 ( .C1(n18516), .C2(n21062), .A(n18675), .B(n18433), .ZN(
        n18450) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18450), .B1(
        n18710), .B2(n18470), .ZN(n18434) );
  OAI211_X1 U21548 ( .C1(n18679), .C2(n18453), .A(n18435), .B(n18434), .ZN(
        P3_U2900) );
  AOI22_X1 U21549 ( .A1(n18716), .A2(n18470), .B1(n18715), .B2(n18448), .ZN(
        n18437) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18450), .B1(
        n18714), .B2(n18449), .ZN(n18436) );
  OAI211_X1 U21551 ( .C1(n18719), .C2(n18453), .A(n18437), .B(n18436), .ZN(
        P3_U2901) );
  AOI22_X1 U21552 ( .A1(n18723), .A2(n18470), .B1(n18720), .B2(n18448), .ZN(
        n18439) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18450), .B1(
        n18721), .B2(n18449), .ZN(n18438) );
  OAI211_X1 U21554 ( .C1(n18684), .C2(n18453), .A(n18439), .B(n18438), .ZN(
        P3_U2902) );
  AOI22_X1 U21555 ( .A1(n18729), .A2(n18470), .B1(n18727), .B2(n18448), .ZN(
        n18441) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18450), .B1(
        n18728), .B2(n18449), .ZN(n18440) );
  OAI211_X1 U21557 ( .C1(n18732), .C2(n18453), .A(n18441), .B(n18440), .ZN(
        P3_U2903) );
  AOI22_X1 U21558 ( .A1(n18735), .A2(n18449), .B1(n18733), .B2(n18448), .ZN(
        n18443) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18450), .B1(
        n18734), .B2(n18470), .ZN(n18442) );
  OAI211_X1 U21560 ( .C1(n18689), .C2(n18453), .A(n18443), .B(n18442), .ZN(
        P3_U2904) );
  AOI22_X1 U21561 ( .A1(n18741), .A2(n18449), .B1(n18740), .B2(n18448), .ZN(
        n18445) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18450), .B1(
        n18742), .B2(n18470), .ZN(n18444) );
  OAI211_X1 U21563 ( .C1(n18746), .C2(n18453), .A(n18445), .B(n18444), .ZN(
        P3_U2905) );
  AOI22_X1 U21564 ( .A1(n18749), .A2(n18448), .B1(n18748), .B2(n18449), .ZN(
        n18447) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18450), .B1(
        n18751), .B2(n18470), .ZN(n18446) );
  OAI211_X1 U21566 ( .C1(n18694), .C2(n18453), .A(n18447), .B(n18446), .ZN(
        P3_U2906) );
  AOI22_X1 U21567 ( .A1(n18759), .A2(n18449), .B1(n18755), .B2(n18448), .ZN(
        n18452) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18450), .B1(
        n18756), .B2(n18470), .ZN(n18451) );
  OAI211_X1 U21569 ( .C1(n18700), .C2(n18453), .A(n18452), .B(n18451), .ZN(
        P3_U2907) );
  NAND2_X1 U21570 ( .A1(n18500), .A2(n18543), .ZN(n18475) );
  NOR2_X1 U21571 ( .A1(n18498), .A2(n18642), .ZN(n18469) );
  AOI22_X1 U21572 ( .A1(n18708), .A2(n18470), .B1(n18707), .B2(n18469), .ZN(
        n18456) );
  AOI22_X1 U21573 ( .A1(n18704), .A2(n18454), .B1(n18500), .B2(n18639), .ZN(
        n18471) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18471), .B1(
        n18710), .B2(n18493), .ZN(n18455) );
  OAI211_X1 U21575 ( .C1(n18679), .C2(n18475), .A(n18456), .B(n18455), .ZN(
        P3_U2908) );
  AOI22_X1 U21576 ( .A1(n18715), .A2(n18469), .B1(n18714), .B2(n18470), .ZN(
        n18458) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18471), .B1(
        n18716), .B2(n18493), .ZN(n18457) );
  OAI211_X1 U21578 ( .C1(n18719), .C2(n18475), .A(n18458), .B(n18457), .ZN(
        P3_U2909) );
  AOI22_X1 U21579 ( .A1(n18723), .A2(n18493), .B1(n18720), .B2(n18469), .ZN(
        n18460) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18471), .B1(
        n18721), .B2(n18470), .ZN(n18459) );
  OAI211_X1 U21581 ( .C1(n18684), .C2(n18475), .A(n18460), .B(n18459), .ZN(
        P3_U2910) );
  AOI22_X1 U21582 ( .A1(n18729), .A2(n18493), .B1(n18727), .B2(n18469), .ZN(
        n18462) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18471), .B1(
        n18728), .B2(n18470), .ZN(n18461) );
  OAI211_X1 U21584 ( .C1(n18732), .C2(n18475), .A(n18462), .B(n18461), .ZN(
        P3_U2911) );
  AOI22_X1 U21585 ( .A1(n18734), .A2(n18493), .B1(n18733), .B2(n18469), .ZN(
        n18464) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18471), .B1(
        n18735), .B2(n18470), .ZN(n18463) );
  OAI211_X1 U21587 ( .C1(n18689), .C2(n18475), .A(n18464), .B(n18463), .ZN(
        P3_U2912) );
  AOI22_X1 U21588 ( .A1(n18741), .A2(n18470), .B1(n18740), .B2(n18469), .ZN(
        n18466) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18471), .B1(
        n18742), .B2(n18493), .ZN(n18465) );
  OAI211_X1 U21590 ( .C1(n18746), .C2(n18475), .A(n18466), .B(n18465), .ZN(
        P3_U2913) );
  AOI22_X1 U21591 ( .A1(n18749), .A2(n18469), .B1(n18748), .B2(n18470), .ZN(
        n18468) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18471), .B1(
        n18751), .B2(n18493), .ZN(n18467) );
  OAI211_X1 U21593 ( .C1(n18694), .C2(n18475), .A(n18468), .B(n18467), .ZN(
        P3_U2914) );
  AOI22_X1 U21594 ( .A1(n18759), .A2(n18470), .B1(n18755), .B2(n18469), .ZN(
        n18473) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18471), .B1(
        n18756), .B2(n18493), .ZN(n18472) );
  OAI211_X1 U21596 ( .C1(n18700), .C2(n18475), .A(n18473), .B(n18472), .ZN(
        P3_U2915) );
  NOR2_X1 U21597 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18474), .ZN(
        n18545) );
  NAND2_X1 U21598 ( .A1(n18545), .A2(n18565), .ZN(n18497) );
  INV_X1 U21599 ( .A(n18475), .ZN(n18538) );
  INV_X1 U21600 ( .A(n18497), .ZN(n18560) );
  NOR2_X1 U21601 ( .A1(n18538), .A2(n18560), .ZN(n18521) );
  NOR2_X1 U21602 ( .A1(n18834), .A2(n18521), .ZN(n18492) );
  AOI22_X1 U21603 ( .A1(n18708), .A2(n18493), .B1(n18707), .B2(n18492), .ZN(
        n18479) );
  AOI221_X1 U21604 ( .B1(n18521), .B2(n18672), .C1(n18521), .C2(n18476), .A(
        n18566), .ZN(n18477) );
  INV_X1 U21605 ( .A(n18477), .ZN(n18494) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18494), .B1(
        n18710), .B2(n18516), .ZN(n18478) );
  OAI211_X1 U21607 ( .C1(n18679), .C2(n18497), .A(n18479), .B(n18478), .ZN(
        P3_U2916) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18494), .B1(
        n18715), .B2(n18492), .ZN(n18481) );
  AOI22_X1 U21609 ( .A1(n18716), .A2(n18516), .B1(n18714), .B2(n18493), .ZN(
        n18480) );
  OAI211_X1 U21610 ( .C1(n18719), .C2(n18497), .A(n18481), .B(n18480), .ZN(
        P3_U2917) );
  AOI22_X1 U21611 ( .A1(n18723), .A2(n18516), .B1(n18720), .B2(n18492), .ZN(
        n18483) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18494), .B1(
        n18721), .B2(n18493), .ZN(n18482) );
  OAI211_X1 U21613 ( .C1(n18684), .C2(n18497), .A(n18483), .B(n18482), .ZN(
        P3_U2918) );
  AOI22_X1 U21614 ( .A1(n18729), .A2(n18516), .B1(n18727), .B2(n18492), .ZN(
        n18485) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18494), .B1(
        n18728), .B2(n18493), .ZN(n18484) );
  OAI211_X1 U21616 ( .C1(n18732), .C2(n18497), .A(n18485), .B(n18484), .ZN(
        P3_U2919) );
  AOI22_X1 U21617 ( .A1(n18735), .A2(n18493), .B1(n18733), .B2(n18492), .ZN(
        n18487) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18494), .B1(
        n18734), .B2(n18516), .ZN(n18486) );
  OAI211_X1 U21619 ( .C1(n18689), .C2(n18497), .A(n18487), .B(n18486), .ZN(
        P3_U2920) );
  AOI22_X1 U21620 ( .A1(n18740), .A2(n18492), .B1(n18742), .B2(n18516), .ZN(
        n18489) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18494), .B1(
        n18741), .B2(n18493), .ZN(n18488) );
  OAI211_X1 U21622 ( .C1(n18746), .C2(n18497), .A(n18489), .B(n18488), .ZN(
        P3_U2921) );
  AOI22_X1 U21623 ( .A1(n18751), .A2(n18516), .B1(n18749), .B2(n18492), .ZN(
        n18491) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18494), .B1(
        n18748), .B2(n18493), .ZN(n18490) );
  OAI211_X1 U21625 ( .C1(n18694), .C2(n18497), .A(n18491), .B(n18490), .ZN(
        P3_U2922) );
  AOI22_X1 U21626 ( .A1(n18759), .A2(n18493), .B1(n18755), .B2(n18492), .ZN(
        n18496) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18494), .B1(
        n18756), .B2(n18516), .ZN(n18495) );
  OAI211_X1 U21628 ( .C1(n18700), .C2(n18497), .A(n18496), .B(n18495), .ZN(
        P3_U2923) );
  NOR2_X2 U21629 ( .A1(n18808), .A2(n18498), .ZN(n18590) );
  INV_X1 U21630 ( .A(n18590), .ZN(n18520) );
  AND2_X1 U21631 ( .A1(n18706), .A2(n18545), .ZN(n18515) );
  AOI22_X1 U21632 ( .A1(n18708), .A2(n18516), .B1(n18707), .B2(n18515), .ZN(
        n18502) );
  NAND2_X1 U21633 ( .A1(n18500), .A2(n18499), .ZN(n18517) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18517), .B1(
        n18710), .B2(n18538), .ZN(n18501) );
  OAI211_X1 U21635 ( .C1(n18679), .C2(n18520), .A(n18502), .B(n18501), .ZN(
        P3_U2924) );
  AOI22_X1 U21636 ( .A1(n18716), .A2(n18538), .B1(n18715), .B2(n18515), .ZN(
        n18504) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18517), .B1(
        n18714), .B2(n18516), .ZN(n18503) );
  OAI211_X1 U21638 ( .C1(n18719), .C2(n18520), .A(n18504), .B(n18503), .ZN(
        P3_U2925) );
  AOI22_X1 U21639 ( .A1(n18723), .A2(n18538), .B1(n18720), .B2(n18515), .ZN(
        n18506) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18517), .B1(
        n18721), .B2(n18516), .ZN(n18505) );
  OAI211_X1 U21641 ( .C1(n18684), .C2(n18520), .A(n18506), .B(n18505), .ZN(
        P3_U2926) );
  AOI22_X1 U21642 ( .A1(n18728), .A2(n18516), .B1(n18727), .B2(n18515), .ZN(
        n18508) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18517), .B1(
        n18729), .B2(n18538), .ZN(n18507) );
  OAI211_X1 U21644 ( .C1(n18732), .C2(n18520), .A(n18508), .B(n18507), .ZN(
        P3_U2927) );
  AOI22_X1 U21645 ( .A1(n18735), .A2(n18516), .B1(n18733), .B2(n18515), .ZN(
        n18510) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18517), .B1(
        n18734), .B2(n18538), .ZN(n18509) );
  OAI211_X1 U21647 ( .C1(n18689), .C2(n18520), .A(n18510), .B(n18509), .ZN(
        P3_U2928) );
  AOI22_X1 U21648 ( .A1(n18741), .A2(n18516), .B1(n18740), .B2(n18515), .ZN(
        n18512) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18517), .B1(
        n18742), .B2(n18538), .ZN(n18511) );
  OAI211_X1 U21650 ( .C1(n18746), .C2(n18520), .A(n18512), .B(n18511), .ZN(
        P3_U2929) );
  AOI22_X1 U21651 ( .A1(n18751), .A2(n18538), .B1(n18749), .B2(n18515), .ZN(
        n18514) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18517), .B1(
        n18748), .B2(n18516), .ZN(n18513) );
  OAI211_X1 U21653 ( .C1(n18694), .C2(n18520), .A(n18514), .B(n18513), .ZN(
        P3_U2930) );
  AOI22_X1 U21654 ( .A1(n18759), .A2(n18516), .B1(n18755), .B2(n18515), .ZN(
        n18519) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18517), .B1(
        n18756), .B2(n18538), .ZN(n18518) );
  OAI211_X1 U21656 ( .C1(n18700), .C2(n18520), .A(n18519), .B(n18518), .ZN(
        P3_U2931) );
  NOR2_X2 U21657 ( .A1(n18810), .A2(n18595), .ZN(n18612) );
  INV_X1 U21658 ( .A(n18612), .ZN(n18542) );
  NOR2_X1 U21659 ( .A1(n18590), .A2(n18612), .ZN(n18567) );
  NOR2_X1 U21660 ( .A1(n18834), .A2(n18567), .ZN(n18537) );
  AOI22_X1 U21661 ( .A1(n18710), .A2(n18560), .B1(n18707), .B2(n18537), .ZN(
        n18524) );
  OAI21_X1 U21662 ( .B1(n18521), .B2(n18672), .A(n18567), .ZN(n18522) );
  OAI211_X1 U21663 ( .C1(n18612), .C2(n21062), .A(n18675), .B(n18522), .ZN(
        n18539) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18539), .B1(
        n18708), .B2(n18538), .ZN(n18523) );
  OAI211_X1 U21665 ( .C1(n18679), .C2(n18542), .A(n18524), .B(n18523), .ZN(
        P3_U2932) );
  AOI22_X1 U21666 ( .A1(n18715), .A2(n18537), .B1(n18714), .B2(n18538), .ZN(
        n18526) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18539), .B1(
        n18716), .B2(n18560), .ZN(n18525) );
  OAI211_X1 U21668 ( .C1(n18719), .C2(n18542), .A(n18526), .B(n18525), .ZN(
        P3_U2933) );
  AOI22_X1 U21669 ( .A1(n18721), .A2(n18538), .B1(n18720), .B2(n18537), .ZN(
        n18528) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18539), .B1(
        n18723), .B2(n18560), .ZN(n18527) );
  OAI211_X1 U21671 ( .C1(n18684), .C2(n18542), .A(n18528), .B(n18527), .ZN(
        P3_U2934) );
  AOI22_X1 U21672 ( .A1(n18728), .A2(n18538), .B1(n18727), .B2(n18537), .ZN(
        n18530) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18539), .B1(
        n18729), .B2(n18560), .ZN(n18529) );
  OAI211_X1 U21674 ( .C1(n18732), .C2(n18542), .A(n18530), .B(n18529), .ZN(
        P3_U2935) );
  AOI22_X1 U21675 ( .A1(n18734), .A2(n18560), .B1(n18733), .B2(n18537), .ZN(
        n18532) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18539), .B1(
        n18735), .B2(n18538), .ZN(n18531) );
  OAI211_X1 U21677 ( .C1(n18689), .C2(n18542), .A(n18532), .B(n18531), .ZN(
        P3_U2936) );
  AOI22_X1 U21678 ( .A1(n18741), .A2(n18538), .B1(n18740), .B2(n18537), .ZN(
        n18534) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18539), .B1(
        n18742), .B2(n18560), .ZN(n18533) );
  OAI211_X1 U21680 ( .C1(n18746), .C2(n18542), .A(n18534), .B(n18533), .ZN(
        P3_U2937) );
  AOI22_X1 U21681 ( .A1(n18749), .A2(n18537), .B1(n18748), .B2(n18538), .ZN(
        n18536) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18539), .B1(
        n18751), .B2(n18560), .ZN(n18535) );
  OAI211_X1 U21683 ( .C1(n18694), .C2(n18542), .A(n18536), .B(n18535), .ZN(
        P3_U2938) );
  AOI22_X1 U21684 ( .A1(n18756), .A2(n18560), .B1(n18755), .B2(n18537), .ZN(
        n18541) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18539), .B1(
        n18759), .B2(n18538), .ZN(n18540) );
  OAI211_X1 U21686 ( .C1(n18700), .C2(n18542), .A(n18541), .B(n18540), .ZN(
        P3_U2939) );
  NAND2_X1 U21687 ( .A1(n18544), .A2(n18543), .ZN(n18564) );
  NOR2_X1 U21688 ( .A1(n18595), .A2(n18642), .ZN(n18596) );
  AOI22_X1 U21689 ( .A1(n18710), .A2(n18590), .B1(n18707), .B2(n18596), .ZN(
        n18547) );
  AOI22_X1 U21690 ( .A1(n18704), .A2(n18545), .B1(n18544), .B2(n18639), .ZN(
        n18561) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18561), .B1(
        n18708), .B2(n18560), .ZN(n18546) );
  OAI211_X1 U21692 ( .C1(n18679), .C2(n18564), .A(n18547), .B(n18546), .ZN(
        P3_U2940) );
  AOI22_X1 U21693 ( .A1(n18715), .A2(n18596), .B1(n18714), .B2(n18560), .ZN(
        n18549) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18561), .B1(
        n18716), .B2(n18590), .ZN(n18548) );
  OAI211_X1 U21695 ( .C1(n18719), .C2(n18564), .A(n18549), .B(n18548), .ZN(
        P3_U2941) );
  AOI22_X1 U21696 ( .A1(n18721), .A2(n18560), .B1(n18720), .B2(n18596), .ZN(
        n18551) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18561), .B1(
        n18723), .B2(n18590), .ZN(n18550) );
  OAI211_X1 U21698 ( .C1(n18684), .C2(n18564), .A(n18551), .B(n18550), .ZN(
        P3_U2942) );
  AOI22_X1 U21699 ( .A1(n18728), .A2(n18560), .B1(n18727), .B2(n18596), .ZN(
        n18553) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18561), .B1(
        n18729), .B2(n18590), .ZN(n18552) );
  OAI211_X1 U21701 ( .C1(n18732), .C2(n18564), .A(n18553), .B(n18552), .ZN(
        P3_U2943) );
  AOI22_X1 U21702 ( .A1(n18735), .A2(n18560), .B1(n18733), .B2(n18596), .ZN(
        n18555) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18561), .B1(
        n18734), .B2(n18590), .ZN(n18554) );
  OAI211_X1 U21704 ( .C1(n18689), .C2(n18564), .A(n18555), .B(n18554), .ZN(
        P3_U2944) );
  AOI22_X1 U21705 ( .A1(n18741), .A2(n18560), .B1(n18740), .B2(n18596), .ZN(
        n18557) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18561), .B1(
        n18742), .B2(n18590), .ZN(n18556) );
  OAI211_X1 U21707 ( .C1(n18746), .C2(n18564), .A(n18557), .B(n18556), .ZN(
        P3_U2945) );
  AOI22_X1 U21708 ( .A1(n18749), .A2(n18596), .B1(n18748), .B2(n18560), .ZN(
        n18559) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18561), .B1(
        n18751), .B2(n18590), .ZN(n18558) );
  OAI211_X1 U21710 ( .C1(n18694), .C2(n18564), .A(n18559), .B(n18558), .ZN(
        P3_U2946) );
  AOI22_X1 U21711 ( .A1(n18759), .A2(n18560), .B1(n18755), .B2(n18596), .ZN(
        n18563) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18561), .B1(
        n18756), .B2(n18590), .ZN(n18562) );
  OAI211_X1 U21713 ( .C1(n18700), .C2(n18564), .A(n18563), .B(n18562), .ZN(
        P3_U2947) );
  INV_X1 U21714 ( .A(n18564), .ZN(n18634) );
  NOR2_X1 U21715 ( .A1(n18809), .A2(n18595), .ZN(n18641) );
  NAND2_X1 U21716 ( .A1(n18565), .A2(n18641), .ZN(n18588) );
  NOR2_X1 U21717 ( .A1(n18634), .A2(n18666), .ZN(n18617) );
  AOI221_X1 U21718 ( .B1(n18567), .B2(n18617), .C1(n18672), .C2(n18617), .A(
        n18566), .ZN(n18594) );
  NOR2_X1 U21719 ( .A1(n18834), .A2(n18617), .ZN(n18589) );
  AOI22_X1 U21720 ( .A1(n18710), .A2(n18612), .B1(n18707), .B2(n18589), .ZN(
        n18569) );
  AOI22_X1 U21721 ( .A1(n18708), .A2(n18590), .B1(n18709), .B2(n18666), .ZN(
        n18568) );
  OAI211_X1 U21722 ( .C1(n18594), .C2(n18570), .A(n18569), .B(n18568), .ZN(
        P3_U2948) );
  AOI22_X1 U21723 ( .A1(n18716), .A2(n18612), .B1(n18715), .B2(n18589), .ZN(
        n18572) );
  AOI22_X1 U21724 ( .A1(n18647), .A2(n18666), .B1(n18714), .B2(n18590), .ZN(
        n18571) );
  OAI211_X1 U21725 ( .C1(n18594), .C2(n18573), .A(n18572), .B(n18571), .ZN(
        P3_U2949) );
  AOI22_X1 U21726 ( .A1(n18723), .A2(n18612), .B1(n18720), .B2(n18589), .ZN(
        n18575) );
  INV_X1 U21727 ( .A(n18594), .ZN(n18585) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18585), .B1(
        n18721), .B2(n18590), .ZN(n18574) );
  OAI211_X1 U21729 ( .C1(n18684), .C2(n18588), .A(n18575), .B(n18574), .ZN(
        P3_U2950) );
  AOI22_X1 U21730 ( .A1(n18728), .A2(n18590), .B1(n18727), .B2(n18589), .ZN(
        n18577) );
  AOI22_X1 U21731 ( .A1(n18653), .A2(n18666), .B1(n18729), .B2(n18612), .ZN(
        n18576) );
  OAI211_X1 U21732 ( .C1(n18594), .C2(n18578), .A(n18577), .B(n18576), .ZN(
        P3_U2951) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18585), .B1(
        n18733), .B2(n18589), .ZN(n18580) );
  AOI22_X1 U21734 ( .A1(n18734), .A2(n18612), .B1(n18735), .B2(n18590), .ZN(
        n18579) );
  OAI211_X1 U21735 ( .C1(n18689), .C2(n18588), .A(n18580), .B(n18579), .ZN(
        P3_U2952) );
  AOI22_X1 U21736 ( .A1(n18741), .A2(n18590), .B1(n18740), .B2(n18589), .ZN(
        n18583) );
  AOI22_X1 U21737 ( .A1(n18581), .A2(n18666), .B1(n18742), .B2(n18612), .ZN(
        n18582) );
  OAI211_X1 U21738 ( .C1(n18594), .C2(n18584), .A(n18583), .B(n18582), .ZN(
        P3_U2953) );
  AOI22_X1 U21739 ( .A1(n18749), .A2(n18589), .B1(n18748), .B2(n18590), .ZN(
        n18587) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18585), .B1(
        n18751), .B2(n18612), .ZN(n18586) );
  OAI211_X1 U21741 ( .C1(n18694), .C2(n18588), .A(n18587), .B(n18586), .ZN(
        P3_U2954) );
  AOI22_X1 U21742 ( .A1(n18756), .A2(n18612), .B1(n18755), .B2(n18589), .ZN(
        n18592) );
  AOI22_X1 U21743 ( .A1(n18759), .A2(n18590), .B1(n18760), .B2(n18666), .ZN(
        n18591) );
  OAI211_X1 U21744 ( .C1(n18594), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P3_U2955) );
  NOR2_X2 U21745 ( .A1(n18808), .A2(n18595), .ZN(n18697) );
  INV_X1 U21746 ( .A(n18697), .ZN(n18616) );
  AND2_X1 U21747 ( .A1(n18706), .A2(n18641), .ZN(n18611) );
  AOI22_X1 U21748 ( .A1(n18708), .A2(n18612), .B1(n18707), .B2(n18611), .ZN(
        n18598) );
  AOI22_X1 U21749 ( .A1(n18704), .A2(n18596), .B1(n18702), .B2(n18641), .ZN(
        n18613) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18613), .B1(
        n18710), .B2(n18634), .ZN(n18597) );
  OAI211_X1 U21751 ( .C1(n18679), .C2(n18616), .A(n18598), .B(n18597), .ZN(
        P3_U2956) );
  AOI22_X1 U21752 ( .A1(n18716), .A2(n18634), .B1(n18715), .B2(n18611), .ZN(
        n18600) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18613), .B1(
        n18714), .B2(n18612), .ZN(n18599) );
  OAI211_X1 U21754 ( .C1(n18719), .C2(n18616), .A(n18600), .B(n18599), .ZN(
        P3_U2957) );
  AOI22_X1 U21755 ( .A1(n18723), .A2(n18634), .B1(n18720), .B2(n18611), .ZN(
        n18602) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18613), .B1(
        n18721), .B2(n18612), .ZN(n18601) );
  OAI211_X1 U21757 ( .C1(n18684), .C2(n18616), .A(n18602), .B(n18601), .ZN(
        P3_U2958) );
  AOI22_X1 U21758 ( .A1(n18729), .A2(n18634), .B1(n18727), .B2(n18611), .ZN(
        n18604) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18613), .B1(
        n18728), .B2(n18612), .ZN(n18603) );
  OAI211_X1 U21760 ( .C1(n18732), .C2(n18616), .A(n18604), .B(n18603), .ZN(
        P3_U2959) );
  AOI22_X1 U21761 ( .A1(n18735), .A2(n18612), .B1(n18733), .B2(n18611), .ZN(
        n18606) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18613), .B1(
        n18734), .B2(n18634), .ZN(n18605) );
  OAI211_X1 U21763 ( .C1(n18689), .C2(n18616), .A(n18606), .B(n18605), .ZN(
        P3_U2960) );
  AOI22_X1 U21764 ( .A1(n18740), .A2(n18611), .B1(n18742), .B2(n18634), .ZN(
        n18608) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18613), .B1(
        n18741), .B2(n18612), .ZN(n18607) );
  OAI211_X1 U21766 ( .C1(n18746), .C2(n18616), .A(n18608), .B(n18607), .ZN(
        P3_U2961) );
  AOI22_X1 U21767 ( .A1(n18751), .A2(n18634), .B1(n18749), .B2(n18611), .ZN(
        n18610) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18613), .B1(
        n18748), .B2(n18612), .ZN(n18609) );
  OAI211_X1 U21769 ( .C1(n18694), .C2(n18616), .A(n18610), .B(n18609), .ZN(
        P3_U2962) );
  AOI22_X1 U21770 ( .A1(n18756), .A2(n18634), .B1(n18755), .B2(n18611), .ZN(
        n18615) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18613), .B1(
        n18759), .B2(n18612), .ZN(n18614) );
  OAI211_X1 U21772 ( .C1(n18700), .C2(n18616), .A(n18615), .B(n18614), .ZN(
        P3_U2963) );
  NOR2_X2 U21773 ( .A1(n18810), .A2(n18643), .ZN(n18758) );
  INV_X1 U21774 ( .A(n18758), .ZN(n18638) );
  NOR2_X1 U21775 ( .A1(n18697), .A2(n18758), .ZN(n18673) );
  NOR2_X1 U21776 ( .A1(n18834), .A2(n18673), .ZN(n18633) );
  AOI22_X1 U21777 ( .A1(n18710), .A2(n18666), .B1(n18707), .B2(n18633), .ZN(
        n18620) );
  OAI21_X1 U21778 ( .B1(n18617), .B2(n18672), .A(n18673), .ZN(n18618) );
  OAI211_X1 U21779 ( .C1(n18758), .C2(n21062), .A(n18675), .B(n18618), .ZN(
        n18635) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18635), .B1(
        n18708), .B2(n18634), .ZN(n18619) );
  OAI211_X1 U21781 ( .C1(n18679), .C2(n18638), .A(n18620), .B(n18619), .ZN(
        P3_U2964) );
  AOI22_X1 U21782 ( .A1(n18715), .A2(n18633), .B1(n18714), .B2(n18634), .ZN(
        n18622) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18635), .B1(
        n18716), .B2(n18666), .ZN(n18621) );
  OAI211_X1 U21784 ( .C1(n18719), .C2(n18638), .A(n18622), .B(n18621), .ZN(
        P3_U2965) );
  AOI22_X1 U21785 ( .A1(n18721), .A2(n18634), .B1(n18720), .B2(n18633), .ZN(
        n18624) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18635), .B1(
        n18723), .B2(n18666), .ZN(n18623) );
  OAI211_X1 U21787 ( .C1(n18684), .C2(n18638), .A(n18624), .B(n18623), .ZN(
        P3_U2966) );
  AOI22_X1 U21788 ( .A1(n18728), .A2(n18634), .B1(n18727), .B2(n18633), .ZN(
        n18626) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18635), .B1(
        n18729), .B2(n18666), .ZN(n18625) );
  OAI211_X1 U21790 ( .C1(n18732), .C2(n18638), .A(n18626), .B(n18625), .ZN(
        P3_U2967) );
  AOI22_X1 U21791 ( .A1(n18734), .A2(n18666), .B1(n18733), .B2(n18633), .ZN(
        n18628) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18635), .B1(
        n18735), .B2(n18634), .ZN(n18627) );
  OAI211_X1 U21793 ( .C1(n18689), .C2(n18638), .A(n18628), .B(n18627), .ZN(
        P3_U2968) );
  AOI22_X1 U21794 ( .A1(n18741), .A2(n18634), .B1(n18740), .B2(n18633), .ZN(
        n18630) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18635), .B1(
        n18742), .B2(n18666), .ZN(n18629) );
  OAI211_X1 U21796 ( .C1(n18746), .C2(n18638), .A(n18630), .B(n18629), .ZN(
        P3_U2969) );
  AOI22_X1 U21797 ( .A1(n18751), .A2(n18666), .B1(n18749), .B2(n18633), .ZN(
        n18632) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18635), .B1(
        n18748), .B2(n18634), .ZN(n18631) );
  OAI211_X1 U21799 ( .C1(n18694), .C2(n18638), .A(n18632), .B(n18631), .ZN(
        P3_U2970) );
  AOI22_X1 U21800 ( .A1(n18756), .A2(n18666), .B1(n18755), .B2(n18633), .ZN(
        n18637) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18635), .B1(
        n18759), .B2(n18634), .ZN(n18636) );
  OAI211_X1 U21802 ( .C1(n18700), .C2(n18638), .A(n18637), .B(n18636), .ZN(
        P3_U2971) );
  AOI22_X1 U21803 ( .A1(n18704), .A2(n18641), .B1(n18640), .B2(n18639), .ZN(
        n18662) );
  INV_X1 U21804 ( .A(n18662), .ZN(n18669) );
  NOR2_X1 U21805 ( .A1(n18643), .A2(n18642), .ZN(n18703) );
  AOI22_X1 U21806 ( .A1(n18708), .A2(n18666), .B1(n18707), .B2(n18703), .ZN(
        n18645) );
  AOI22_X1 U21807 ( .A1(n18757), .A2(n18709), .B1(n18710), .B2(n18697), .ZN(
        n18644) );
  OAI211_X1 U21808 ( .C1(n18646), .C2(n18669), .A(n18645), .B(n18644), .ZN(
        P3_U2972) );
  AOI22_X1 U21809 ( .A1(n18715), .A2(n18703), .B1(n18714), .B2(n18666), .ZN(
        n18649) );
  AOI22_X1 U21810 ( .A1(n18757), .A2(n18647), .B1(n18716), .B2(n18697), .ZN(
        n18648) );
  OAI211_X1 U21811 ( .C1(n18650), .C2(n18669), .A(n18649), .B(n18648), .ZN(
        P3_U2973) );
  AOI22_X1 U21812 ( .A1(n18721), .A2(n18666), .B1(n18720), .B2(n18703), .ZN(
        n18652) );
  AOI22_X1 U21813 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18662), .B1(
        n18723), .B2(n18697), .ZN(n18651) );
  OAI211_X1 U21814 ( .C1(n18665), .C2(n18684), .A(n18652), .B(n18651), .ZN(
        P3_U2974) );
  AOI22_X1 U21815 ( .A1(n18728), .A2(n18666), .B1(n18727), .B2(n18703), .ZN(
        n18655) );
  AOI22_X1 U21816 ( .A1(n18757), .A2(n18653), .B1(n18729), .B2(n18697), .ZN(
        n18654) );
  OAI211_X1 U21817 ( .C1(n18656), .C2(n18669), .A(n18655), .B(n18654), .ZN(
        P3_U2975) );
  AOI22_X1 U21818 ( .A1(n18734), .A2(n18697), .B1(n18733), .B2(n18703), .ZN(
        n18658) );
  AOI22_X1 U21819 ( .A1(n18757), .A2(n18736), .B1(n18735), .B2(n18666), .ZN(
        n18657) );
  OAI211_X1 U21820 ( .C1(n18659), .C2(n18669), .A(n18658), .B(n18657), .ZN(
        P3_U2976) );
  AOI22_X1 U21821 ( .A1(n18740), .A2(n18703), .B1(n18742), .B2(n18697), .ZN(
        n18661) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18662), .B1(
        n18741), .B2(n18666), .ZN(n18660) );
  OAI211_X1 U21823 ( .C1(n18665), .C2(n18746), .A(n18661), .B(n18660), .ZN(
        P3_U2977) );
  AOI22_X1 U21824 ( .A1(n18749), .A2(n18703), .B1(n18748), .B2(n18666), .ZN(
        n18664) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18662), .B1(
        n18751), .B2(n18697), .ZN(n18663) );
  OAI211_X1 U21826 ( .C1(n18665), .C2(n18694), .A(n18664), .B(n18663), .ZN(
        P3_U2978) );
  AOI22_X1 U21827 ( .A1(n18759), .A2(n18666), .B1(n18755), .B2(n18703), .ZN(
        n18668) );
  AOI22_X1 U21828 ( .A1(n18757), .A2(n18760), .B1(n18756), .B2(n18697), .ZN(
        n18667) );
  OAI211_X1 U21829 ( .C1(n18670), .C2(n18669), .A(n18668), .B(n18667), .ZN(
        P3_U2979) );
  NOR2_X1 U21830 ( .A1(n18834), .A2(n18671), .ZN(n18695) );
  AOI22_X1 U21831 ( .A1(n18710), .A2(n18758), .B1(n18707), .B2(n18695), .ZN(
        n18678) );
  OAI21_X1 U21832 ( .B1(n18673), .B2(n18672), .A(n18671), .ZN(n18674) );
  OAI211_X1 U21833 ( .C1(n18676), .C2(n21062), .A(n18675), .B(n18674), .ZN(
        n18696) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18696), .B1(
        n18708), .B2(n18697), .ZN(n18677) );
  OAI211_X1 U21835 ( .C1(n18701), .C2(n18679), .A(n18678), .B(n18677), .ZN(
        P3_U2980) );
  AOI22_X1 U21836 ( .A1(n18716), .A2(n18758), .B1(n18715), .B2(n18695), .ZN(
        n18681) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18696), .B1(
        n18714), .B2(n18697), .ZN(n18680) );
  OAI211_X1 U21838 ( .C1(n18701), .C2(n18719), .A(n18681), .B(n18680), .ZN(
        P3_U2981) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18696), .B1(
        n18720), .B2(n18695), .ZN(n18683) );
  AOI22_X1 U21840 ( .A1(n18723), .A2(n18758), .B1(n18721), .B2(n18697), .ZN(
        n18682) );
  OAI211_X1 U21841 ( .C1(n18701), .C2(n18684), .A(n18683), .B(n18682), .ZN(
        P3_U2982) );
  AOI22_X1 U21842 ( .A1(n18729), .A2(n18758), .B1(n18727), .B2(n18695), .ZN(
        n18686) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18696), .B1(
        n18728), .B2(n18697), .ZN(n18685) );
  OAI211_X1 U21844 ( .C1(n18701), .C2(n18732), .A(n18686), .B(n18685), .ZN(
        P3_U2983) );
  AOI22_X1 U21845 ( .A1(n18734), .A2(n18758), .B1(n18733), .B2(n18695), .ZN(
        n18688) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18696), .B1(
        n18735), .B2(n18697), .ZN(n18687) );
  OAI211_X1 U21847 ( .C1(n18701), .C2(n18689), .A(n18688), .B(n18687), .ZN(
        P3_U2984) );
  AOI22_X1 U21848 ( .A1(n18741), .A2(n18697), .B1(n18740), .B2(n18695), .ZN(
        n18691) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18696), .B1(
        n18742), .B2(n18758), .ZN(n18690) );
  OAI211_X1 U21850 ( .C1(n18701), .C2(n18746), .A(n18691), .B(n18690), .ZN(
        P3_U2985) );
  AOI22_X1 U21851 ( .A1(n18751), .A2(n18758), .B1(n18749), .B2(n18695), .ZN(
        n18693) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18696), .B1(
        n18748), .B2(n18697), .ZN(n18692) );
  OAI211_X1 U21853 ( .C1(n18701), .C2(n18694), .A(n18693), .B(n18692), .ZN(
        P3_U2986) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18696), .B1(
        n18755), .B2(n18695), .ZN(n18699) );
  AOI22_X1 U21855 ( .A1(n18759), .A2(n18697), .B1(n18756), .B2(n18758), .ZN(
        n18698) );
  OAI211_X1 U21856 ( .C1(n18701), .C2(n18700), .A(n18699), .B(n18698), .ZN(
        P3_U2987) );
  AOI22_X1 U21857 ( .A1(n18704), .A2(n18703), .B1(n18705), .B2(n18702), .ZN(
        n18743) );
  INV_X1 U21858 ( .A(n18743), .ZN(n18764) );
  AND2_X1 U21859 ( .A1(n18706), .A2(n18705), .ZN(n18754) );
  AOI22_X1 U21860 ( .A1(n18708), .A2(n18758), .B1(n18707), .B2(n18754), .ZN(
        n18712) );
  AOI22_X1 U21861 ( .A1(n18757), .A2(n18710), .B1(n18761), .B2(n18709), .ZN(
        n18711) );
  OAI211_X1 U21862 ( .C1(n18713), .C2(n18764), .A(n18712), .B(n18711), .ZN(
        P3_U2988) );
  INV_X1 U21863 ( .A(n18761), .ZN(n18747) );
  AOI22_X1 U21864 ( .A1(n18715), .A2(n18754), .B1(n18714), .B2(n18758), .ZN(
        n18718) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18743), .B1(
        n18757), .B2(n18716), .ZN(n18717) );
  OAI211_X1 U21866 ( .C1(n18747), .C2(n18719), .A(n18718), .B(n18717), .ZN(
        P3_U2989) );
  AOI22_X1 U21867 ( .A1(n18721), .A2(n18758), .B1(n18720), .B2(n18754), .ZN(
        n18725) );
  AOI22_X1 U21868 ( .A1(n18757), .A2(n18723), .B1(n18761), .B2(n18722), .ZN(
        n18724) );
  OAI211_X1 U21869 ( .C1(n18726), .C2(n18764), .A(n18725), .B(n18724), .ZN(
        P3_U2990) );
  AOI22_X1 U21870 ( .A1(n18728), .A2(n18758), .B1(n18727), .B2(n18754), .ZN(
        n18731) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18743), .B1(
        n18757), .B2(n18729), .ZN(n18730) );
  OAI211_X1 U21872 ( .C1(n18747), .C2(n18732), .A(n18731), .B(n18730), .ZN(
        P3_U2991) );
  AOI22_X1 U21873 ( .A1(n18757), .A2(n18734), .B1(n18733), .B2(n18754), .ZN(
        n18738) );
  AOI22_X1 U21874 ( .A1(n18761), .A2(n18736), .B1(n18735), .B2(n18758), .ZN(
        n18737) );
  OAI211_X1 U21875 ( .C1(n18739), .C2(n18764), .A(n18738), .B(n18737), .ZN(
        P3_U2992) );
  AOI22_X1 U21876 ( .A1(n18741), .A2(n18758), .B1(n18740), .B2(n18754), .ZN(
        n18745) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18743), .B1(
        n18757), .B2(n18742), .ZN(n18744) );
  OAI211_X1 U21878 ( .C1(n18747), .C2(n18746), .A(n18745), .B(n18744), .ZN(
        P3_U2993) );
  AOI22_X1 U21879 ( .A1(n18749), .A2(n18754), .B1(n18748), .B2(n18758), .ZN(
        n18753) );
  AOI22_X1 U21880 ( .A1(n18757), .A2(n18751), .B1(n18761), .B2(n18750), .ZN(
        n18752) );
  OAI211_X1 U21881 ( .C1(n20886), .C2(n18764), .A(n18753), .B(n18752), .ZN(
        P3_U2994) );
  AOI22_X1 U21882 ( .A1(n18757), .A2(n18756), .B1(n18755), .B2(n18754), .ZN(
        n18763) );
  AOI22_X1 U21883 ( .A1(n18761), .A2(n18760), .B1(n18759), .B2(n18758), .ZN(
        n18762) );
  OAI211_X1 U21884 ( .C1(n18765), .C2(n18764), .A(n18763), .B(n18762), .ZN(
        P3_U2995) );
  AND2_X1 U21885 ( .A1(n18766), .A2(n18789), .ZN(n18770) );
  NOR2_X1 U21886 ( .A1(n18780), .A2(n18767), .ZN(n18769) );
  OAI222_X1 U21887 ( .A1(n18773), .A2(n18772), .B1(n18771), .B2(n18770), .C1(
        n18769), .C2(n18768), .ZN(n18968) );
  OAI21_X1 U21888 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18774), .ZN(n18775) );
  OAI211_X1 U21889 ( .C1(n18777), .C2(n18802), .A(n18776), .B(n18775), .ZN(
        n18823) );
  NAND2_X1 U21890 ( .A1(n18944), .A2(n18795), .ZN(n18785) );
  NOR2_X1 U21891 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18778), .ZN(
        n18806) );
  INV_X1 U21892 ( .A(n18806), .ZN(n18779) );
  AOI22_X1 U21893 ( .A1(n18780), .A2(n18785), .B1(n18790), .B2(n18779), .ZN(
        n18781) );
  NOR2_X1 U21894 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18781), .ZN(
        n18930) );
  OAI21_X1 U21895 ( .B1(n18784), .B2(n18783), .A(n18782), .ZN(n18793) );
  OAI21_X1 U21896 ( .B1(n18805), .B2(n18790), .A(n18785), .ZN(n18786) );
  AOI21_X1 U21897 ( .B1(n18787), .B2(n18793), .A(n18786), .ZN(n18931) );
  NAND2_X1 U21898 ( .A1(n18802), .A2(n18931), .ZN(n18788) );
  AOI22_X1 U21899 ( .A1(n18802), .A2(n18930), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18788), .ZN(n18821) );
  INV_X1 U21900 ( .A(n18802), .ZN(n18812) );
  AOI211_X1 U21901 ( .C1(n18951), .C2(n18944), .A(n18790), .B(n18789), .ZN(
        n18801) );
  NAND2_X1 U21902 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n9773), .ZN(
        n18791) );
  AOI211_X1 U21903 ( .C1(n18792), .C2(n18791), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18951), .ZN(n18800) );
  AOI21_X1 U21904 ( .B1(n18951), .B2(n18794), .A(n18793), .ZN(n18797) );
  NAND2_X1 U21905 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18795), .ZN(
        n18796) );
  OAI22_X1 U21906 ( .A1(n18940), .A2(n18798), .B1(n18797), .B2(n18796), .ZN(
        n18799) );
  NOR3_X1 U21907 ( .A1(n18801), .A2(n18800), .A3(n18799), .ZN(n18936) );
  AOI22_X1 U21908 ( .A1(n18812), .A2(n18944), .B1(n18936), .B2(n18802), .ZN(
        n18816) );
  NOR2_X1 U21909 ( .A1(n18804), .A2(n9773), .ZN(n18807) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18805), .B1(
        n18807), .B2(n20969), .ZN(n18953) );
  OAI22_X1 U21911 ( .A1(n18807), .A2(n18945), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18806), .ZN(n18949) );
  AOI222_X1 U21912 ( .A1(n18953), .A2(n18949), .B1(n18953), .B2(n18809), .C1(
        n18949), .C2(n18808), .ZN(n18811) );
  OAI21_X1 U21913 ( .B1(n18812), .B2(n18811), .A(n18810), .ZN(n18815) );
  AND2_X1 U21914 ( .A1(n18816), .A2(n18815), .ZN(n18813) );
  OAI221_X1 U21915 ( .B1(n18816), .B2(n18815), .C1(n18814), .C2(n18813), .A(
        n18818), .ZN(n18820) );
  AOI21_X1 U21916 ( .B1(n18818), .B2(n18817), .A(n18816), .ZN(n18819) );
  AOI222_X1 U21917 ( .A1(n18821), .A2(n18820), .B1(n18821), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18820), .C2(n18819), .ZN(
        n18822) );
  NOR4_X1 U21918 ( .A1(n18824), .A2(n18968), .A3(n18823), .A4(n18822), .ZN(
        n18833) );
  OAI211_X1 U21919 ( .C1(n18826), .C2(n18825), .A(n18977), .B(n18833), .ZN(
        n18927) );
  OAI21_X1 U21920 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18979), .A(n18927), 
        .ZN(n18835) );
  AOI221_X1 U21921 ( .B1(n18828), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18835), 
        .C2(P3_STATE2_REG_0__SCAN_IN), .A(n18827), .ZN(n18831) );
  NAND2_X1 U21922 ( .A1(n18971), .A2(n18980), .ZN(n18838) );
  OAI211_X1 U21923 ( .C1(n18829), .C2(n18973), .A(n18974), .B(n18838), .ZN(
        n18830) );
  OAI211_X1 U21924 ( .C1(n18833), .C2(n18832), .A(n18831), .B(n18830), .ZN(
        P3_U2996) );
  NAND4_X1 U21925 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18971), .A4(n18986), .ZN(n18840) );
  OR3_X1 U21926 ( .A1(n18836), .A2(n18835), .A3(n18834), .ZN(n18837) );
  NAND4_X1 U21927 ( .A1(n18839), .A2(n18838), .A3(n18840), .A4(n18837), .ZN(
        P3_U2997) );
  AND4_X1 U21928 ( .A1(n18973), .A2(n18841), .A3(n18840), .A4(n18926), .ZN(
        P3_U2998) );
  INV_X1 U21929 ( .A(n18925), .ZN(n18842) );
  AND2_X1 U21930 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18842), .ZN(
        P3_U2999) );
  AND2_X1 U21931 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18842), .ZN(
        P3_U3000) );
  AND2_X1 U21932 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18842), .ZN(
        P3_U3001) );
  AND2_X1 U21933 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18842), .ZN(
        P3_U3002) );
  AND2_X1 U21934 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18842), .ZN(
        P3_U3003) );
  AND2_X1 U21935 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18842), .ZN(
        P3_U3004) );
  AND2_X1 U21936 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18842), .ZN(
        P3_U3005) );
  AND2_X1 U21937 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18842), .ZN(
        P3_U3006) );
  AND2_X1 U21938 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18842), .ZN(
        P3_U3007) );
  AND2_X1 U21939 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18842), .ZN(
        P3_U3008) );
  AND2_X1 U21940 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18842), .ZN(
        P3_U3009) );
  AND2_X1 U21941 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18842), .ZN(
        P3_U3010) );
  AND2_X1 U21942 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18842), .ZN(
        P3_U3011) );
  AND2_X1 U21943 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18842), .ZN(
        P3_U3012) );
  AND2_X1 U21944 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18842), .ZN(
        P3_U3013) );
  AND2_X1 U21945 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18842), .ZN(
        P3_U3014) );
  AND2_X1 U21946 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18842), .ZN(
        P3_U3015) );
  AND2_X1 U21947 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18842), .ZN(
        P3_U3016) );
  AND2_X1 U21948 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18842), .ZN(
        P3_U3017) );
  AND2_X1 U21949 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18842), .ZN(
        P3_U3018) );
  AND2_X1 U21950 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18842), .ZN(
        P3_U3019) );
  AND2_X1 U21951 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18842), .ZN(
        P3_U3020) );
  AND2_X1 U21952 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18842), .ZN(P3_U3021) );
  AND2_X1 U21953 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18842), .ZN(P3_U3022) );
  AND2_X1 U21954 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18842), .ZN(P3_U3023) );
  AND2_X1 U21955 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18842), .ZN(P3_U3024) );
  AND2_X1 U21956 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18842), .ZN(P3_U3025) );
  AND2_X1 U21957 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18842), .ZN(P3_U3026) );
  AND2_X1 U21958 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18842), .ZN(P3_U3027) );
  AND2_X1 U21959 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18842), .ZN(P3_U3028) );
  NOR2_X1 U21960 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18845), .ZN(n18848) );
  OAI21_X1 U21961 ( .B1(n18843), .B2(n20852), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18844) );
  AOI22_X1 U21962 ( .A1(n18971), .A2(n18848), .B1(n18984), .B2(n18844), .ZN(
        n18847) );
  NAND3_X1 U21963 ( .A1(NA), .A2(n18852), .A3(n18845), .ZN(n18846) );
  OAI211_X1 U21964 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18847), .B(n18846), .ZN(P3_U3029) );
  NAND2_X1 U21965 ( .A1(HOLD), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18849) );
  AOI22_X1 U21966 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18849), .B1(HOLD), 
        .B2(n18848), .ZN(n18851) );
  NAND2_X1 U21967 ( .A1(n18971), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18856) );
  OAI211_X1 U21968 ( .C1(n18851), .C2(n18852), .A(n18856), .B(n18850), .ZN(
        P3_U3030) );
  INV_X1 U21969 ( .A(NA), .ZN(n20906) );
  OAI21_X1 U21970 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n20906), .A(n18852), 
        .ZN(n18855) );
  OAI222_X1 U21971 ( .A1(n18857), .A2(n20852), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n18856), .C2(NA), .ZN(n18853)
         );
  OAI211_X1 U21972 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n18853), .ZN(n18854) );
  OAI221_X1 U21973 ( .B1(n18857), .B2(n18856), .C1(n18857), .C2(n18855), .A(
        n18854), .ZN(P3_U3031) );
  OAI222_X1 U21974 ( .A1(n18908), .A2(n20859), .B1(n18858), .B2(n18983), .C1(
        n18958), .C2(n18910), .ZN(P3_U3032) );
  OAI222_X1 U21975 ( .A1(n18908), .A2(n18861), .B1(n18859), .B2(n18983), .C1(
        n20859), .C2(n18910), .ZN(P3_U3033) );
  OAI222_X1 U21976 ( .A1(n18861), .A2(n18910), .B1(n18860), .B2(n18983), .C1(
        n18862), .C2(n18908), .ZN(P3_U3034) );
  INV_X1 U21977 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18865) );
  OAI222_X1 U21978 ( .A1(n18908), .A2(n18865), .B1(n18863), .B2(n18983), .C1(
        n18862), .C2(n18910), .ZN(P3_U3035) );
  OAI222_X1 U21979 ( .A1(n18865), .A2(n18910), .B1(n18864), .B2(n18983), .C1(
        n18866), .C2(n18908), .ZN(P3_U3036) );
  OAI222_X1 U21980 ( .A1(n18908), .A2(n18868), .B1(n18867), .B2(n18983), .C1(
        n18866), .C2(n18910), .ZN(P3_U3037) );
  OAI222_X1 U21981 ( .A1(n18908), .A2(n18871), .B1(n18869), .B2(n18983), .C1(
        n18868), .C2(n18910), .ZN(P3_U3038) );
  OAI222_X1 U21982 ( .A1(n18871), .A2(n18910), .B1(n18870), .B2(n18983), .C1(
        n18872), .C2(n18908), .ZN(P3_U3039) );
  OAI222_X1 U21983 ( .A1(n18908), .A2(n18874), .B1(n18873), .B2(n18983), .C1(
        n18872), .C2(n18910), .ZN(P3_U3040) );
  OAI222_X1 U21984 ( .A1(n18908), .A2(n18876), .B1(n18875), .B2(n18983), .C1(
        n18874), .C2(n18910), .ZN(P3_U3041) );
  OAI222_X1 U21985 ( .A1(n18908), .A2(n18878), .B1(n18877), .B2(n18983), .C1(
        n18876), .C2(n18910), .ZN(P3_U3042) );
  OAI222_X1 U21986 ( .A1(n18908), .A2(n18880), .B1(n18879), .B2(n18983), .C1(
        n18878), .C2(n18910), .ZN(P3_U3043) );
  OAI222_X1 U21987 ( .A1(n18908), .A2(n18883), .B1(n18881), .B2(n18983), .C1(
        n18880), .C2(n18910), .ZN(P3_U3044) );
  OAI222_X1 U21988 ( .A1(n18883), .A2(n18910), .B1(n18882), .B2(n18983), .C1(
        n18884), .C2(n18908), .ZN(P3_U3045) );
  OAI222_X1 U21989 ( .A1(n18908), .A2(n18886), .B1(n18885), .B2(n18983), .C1(
        n18884), .C2(n18917), .ZN(P3_U3046) );
  OAI222_X1 U21990 ( .A1(n18908), .A2(n18889), .B1(n18887), .B2(n18983), .C1(
        n18886), .C2(n18917), .ZN(P3_U3047) );
  OAI222_X1 U21991 ( .A1(n18889), .A2(n18910), .B1(n18888), .B2(n18983), .C1(
        n20989), .C2(n18908), .ZN(P3_U3048) );
  OAI222_X1 U21992 ( .A1(n20989), .A2(n18910), .B1(n18890), .B2(n18983), .C1(
        n20867), .C2(n18908), .ZN(P3_U3049) );
  OAI222_X1 U21993 ( .A1(n18908), .A2(n18893), .B1(n18891), .B2(n18983), .C1(
        n20867), .C2(n18917), .ZN(P3_U3050) );
  OAI222_X1 U21994 ( .A1(n18893), .A2(n18910), .B1(n18892), .B2(n18983), .C1(
        n18894), .C2(n18908), .ZN(P3_U3051) );
  OAI222_X1 U21995 ( .A1(n18908), .A2(n18896), .B1(n18895), .B2(n18983), .C1(
        n18894), .C2(n18917), .ZN(P3_U3052) );
  OAI222_X1 U21996 ( .A1(n18908), .A2(n18898), .B1(n18897), .B2(n18983), .C1(
        n18896), .C2(n18917), .ZN(P3_U3053) );
  OAI222_X1 U21997 ( .A1(n18908), .A2(n18900), .B1(n18899), .B2(n18983), .C1(
        n18898), .C2(n18917), .ZN(P3_U3054) );
  OAI222_X1 U21998 ( .A1(n18908), .A2(n18902), .B1(n18901), .B2(n18983), .C1(
        n18900), .C2(n18917), .ZN(P3_U3055) );
  OAI222_X1 U21999 ( .A1(n18908), .A2(n18905), .B1(n18903), .B2(n18983), .C1(
        n18902), .C2(n18917), .ZN(P3_U3056) );
  OAI222_X1 U22000 ( .A1(n18905), .A2(n18910), .B1(n18904), .B2(n18983), .C1(
        n18906), .C2(n18908), .ZN(P3_U3057) );
  OAI222_X1 U22001 ( .A1(n18908), .A2(n18911), .B1(n18907), .B2(n18983), .C1(
        n18906), .C2(n18910), .ZN(P3_U3058) );
  OAI222_X1 U22002 ( .A1(n18911), .A2(n18910), .B1(n18909), .B2(n18983), .C1(
        n18912), .C2(n18908), .ZN(P3_U3059) );
  OAI222_X1 U22003 ( .A1(n18908), .A2(n18916), .B1(n18913), .B2(n18983), .C1(
        n18912), .C2(n18917), .ZN(P3_U3060) );
  OAI222_X1 U22004 ( .A1(n18917), .A2(n18916), .B1(n18915), .B2(n18983), .C1(
        n18914), .C2(n18908), .ZN(P3_U3061) );
  OAI22_X1 U22005 ( .A1(n18984), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18983), .ZN(n18918) );
  INV_X1 U22006 ( .A(n18918), .ZN(P3_U3274) );
  OAI22_X1 U22007 ( .A1(n18984), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18983), .ZN(n18919) );
  INV_X1 U22008 ( .A(n18919), .ZN(P3_U3275) );
  OAI22_X1 U22009 ( .A1(n18984), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18983), .ZN(n18920) );
  INV_X1 U22010 ( .A(n18920), .ZN(P3_U3276) );
  OAI22_X1 U22011 ( .A1(n18984), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18983), .ZN(n18921) );
  INV_X1 U22012 ( .A(n18921), .ZN(P3_U3277) );
  OAI21_X1 U22013 ( .B1(n18925), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18923), 
        .ZN(n18922) );
  INV_X1 U22014 ( .A(n18922), .ZN(P3_U3280) );
  OAI21_X1 U22015 ( .B1(n18925), .B2(n18924), .A(n18923), .ZN(P3_U3281) );
  OAI221_X1 U22016 ( .B1(n21062), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21062), 
        .C2(n18927), .A(n18926), .ZN(P3_U3282) );
  INV_X1 U22017 ( .A(n18928), .ZN(n18929) );
  AOI22_X1 U22018 ( .A1(n18987), .A2(n18930), .B1(n18952), .B2(n18929), .ZN(
        n18935) );
  INV_X1 U22019 ( .A(n18931), .ZN(n18932) );
  AOI21_X1 U22020 ( .B1(n18987), .B2(n18932), .A(n18957), .ZN(n18934) );
  OAI22_X1 U22021 ( .A1(n18957), .A2(n18935), .B1(n18934), .B2(n18933), .ZN(
        P3_U3285) );
  INV_X1 U22022 ( .A(n18936), .ZN(n18942) );
  NOR2_X1 U22023 ( .A1(n18937), .A2(n18954), .ZN(n18946) );
  OAI22_X1 U22024 ( .A1(n18939), .A2(n18938), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18947) );
  INV_X1 U22025 ( .A(n18947), .ZN(n18941) );
  AOI222_X1 U22026 ( .A1(n18942), .A2(n18987), .B1(n18946), .B2(n18941), .C1(
        n18952), .C2(n18940), .ZN(n18943) );
  AOI22_X1 U22027 ( .A1(n18957), .A2(n18944), .B1(n18943), .B2(n18955), .ZN(
        P3_U3288) );
  INV_X1 U22028 ( .A(n18945), .ZN(n18948) );
  AOI222_X1 U22029 ( .A1(n18949), .A2(n18987), .B1(n18952), .B2(n18948), .C1(
        n18947), .C2(n18946), .ZN(n18950) );
  AOI22_X1 U22030 ( .A1(n18957), .A2(n18951), .B1(n18950), .B2(n18955), .ZN(
        P3_U3289) );
  AOI222_X1 U22031 ( .A1(n18954), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18987), 
        .B2(n18953), .C1(n20969), .C2(n18952), .ZN(n18956) );
  AOI22_X1 U22032 ( .A1(n18957), .A2(n20969), .B1(n18956), .B2(n18955), .ZN(
        P3_U3290) );
  AOI21_X1 U22033 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18959) );
  AOI22_X1 U22034 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18959), .B2(n18958), .ZN(n18962) );
  INV_X1 U22035 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18961) );
  AOI22_X1 U22036 ( .A1(n18965), .A2(n18962), .B1(n18961), .B2(n18960), .ZN(
        P3_U3292) );
  INV_X1 U22037 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18964) );
  OAI21_X1 U22038 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18965), .ZN(n18963) );
  OAI21_X1 U22039 ( .B1(n18965), .B2(n18964), .A(n18963), .ZN(P3_U3293) );
  INV_X1 U22040 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18990) );
  OAI22_X1 U22041 ( .A1(n18984), .A2(n18990), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18983), .ZN(n18966) );
  INV_X1 U22042 ( .A(n18966), .ZN(P3_U3294) );
  MUX2_X1 U22043 ( .A(P3_MORE_REG_SCAN_IN), .B(n18968), .S(n18967), .Z(
        P3_U3295) );
  OAI21_X1 U22044 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18970), .A(n18969), 
        .ZN(n18972) );
  AOI211_X1 U22045 ( .C1(n18988), .C2(n18972), .A(n18971), .B(n18986), .ZN(
        n18975) );
  OAI21_X1 U22046 ( .B1(n18975), .B2(n18974), .A(n18973), .ZN(n18982) );
  NOR2_X1 U22047 ( .A1(n18977), .A2(n18976), .ZN(n18978) );
  AOI211_X1 U22048 ( .C1(n18980), .C2(n18979), .A(n18978), .B(n18989), .ZN(
        n18981) );
  MUX2_X1 U22049 ( .A(n18982), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18981), 
        .Z(P3_U3296) );
  OAI22_X1 U22050 ( .A1(n18984), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18983), .ZN(n18985) );
  INV_X1 U22051 ( .A(n18985), .ZN(P3_U3297) );
  AOI21_X1 U22052 ( .B1(n18987), .B2(n18986), .A(n18989), .ZN(n18993) );
  AOI22_X1 U22053 ( .A1(n18993), .A2(n18990), .B1(n18989), .B2(n18988), .ZN(
        P3_U3298) );
  INV_X1 U22054 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18992) );
  AOI21_X1 U22055 ( .B1(n18993), .B2(n18992), .A(n18991), .ZN(P3_U3299) );
  INV_X1 U22056 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19960) );
  NOR2_X1 U22057 ( .A1(n19960), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19964) );
  NOR2_X1 U22058 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19965) );
  AOI21_X1 U22059 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19964), .A(n19965), 
        .ZN(n19958) );
  INV_X1 U22060 ( .A(n19958), .ZN(n20027) );
  AOI21_X1 U22061 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20027), .ZN(n18994) );
  INV_X1 U22062 ( .A(n18994), .ZN(P2_U2815) );
  INV_X1 U22063 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18996) );
  OAI22_X1 U22064 ( .A1(n20074), .A2(n18996), .B1(n19309), .B2(n18995), .ZN(
        P2_U2816) );
  INV_X1 U22065 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19966) );
  NAND2_X1 U22066 ( .A1(n19966), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20089) );
  OAI21_X1 U22067 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n20753), .A(n19966), 
        .ZN(n18997) );
  AOI22_X1 U22068 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(n20088), .B1(n18998), 
        .B2(n18997), .ZN(P2_U2817) );
  OAI21_X1 U22069 ( .B1(n20753), .B2(BS16), .A(n20027), .ZN(n20025) );
  OAI21_X1 U22070 ( .B1(n20027), .B2(n19770), .A(n20025), .ZN(P2_U2818) );
  AND2_X1 U22071 ( .A1(n19304), .A2(n18999), .ZN(n20070) );
  OAI21_X1 U22072 ( .B1(n20070), .B2(n19001), .A(n19000), .ZN(P2_U2819) );
  NOR4_X1 U22073 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19005) );
  NOR4_X1 U22074 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_14__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n19004) );
  NOR4_X1 U22075 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19003) );
  NOR4_X1 U22076 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19002) );
  NAND4_X1 U22077 ( .A1(n19005), .A2(n19004), .A3(n19003), .A4(n19002), .ZN(
        n19011) );
  NOR4_X1 U22078 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19009) );
  AOI211_X1 U22079 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_15__SCAN_IN), .B(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19008) );
  NOR4_X1 U22080 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_10__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19007) );
  NOR4_X1 U22081 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19006) );
  NAND4_X1 U22082 ( .A1(n19009), .A2(n19008), .A3(n19007), .A4(n19006), .ZN(
        n19010) );
  NOR2_X1 U22083 ( .A1(n19011), .A2(n19010), .ZN(n19021) );
  INV_X1 U22084 ( .A(n19021), .ZN(n19019) );
  NOR2_X1 U22085 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19019), .ZN(n19014) );
  INV_X1 U22086 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19012) );
  AOI22_X1 U22087 ( .A1(n19014), .A2(n20901), .B1(n19019), .B2(n19012), .ZN(
        P2_U2820) );
  OR3_X1 U22088 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19018) );
  INV_X1 U22089 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19013) );
  AOI22_X1 U22090 ( .A1(n19014), .A2(n19018), .B1(n19019), .B2(n19013), .ZN(
        P2_U2821) );
  INV_X1 U22091 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20026) );
  NAND2_X1 U22092 ( .A1(n19014), .A2(n20026), .ZN(n19017) );
  OAI21_X1 U22093 ( .B1(n20901), .B2(n19970), .A(n19021), .ZN(n19015) );
  OAI21_X1 U22094 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19021), .A(n19015), 
        .ZN(n19016) );
  OAI221_X1 U22095 ( .B1(n19017), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19017), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19016), .ZN(P2_U2822) );
  INV_X1 U22096 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19020) );
  OAI221_X1 U22097 ( .B1(n19021), .B2(n19020), .C1(n19019), .C2(n19018), .A(
        n19017), .ZN(P2_U2823) );
  INV_X1 U22098 ( .A(n19027), .ZN(n19022) );
  AOI22_X1 U22099 ( .A1(n19023), .A2(n19194), .B1(n19022), .B2(n19235), .ZN(
        n19032) );
  OAI22_X1 U22100 ( .A1(n20002), .A2(n19178), .B1(n11049), .B2(n19197), .ZN(
        n19024) );
  AOI21_X1 U22101 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19236), .A(
        n19024), .ZN(n19031) );
  AOI22_X1 U22102 ( .A1(n10220), .A2(n19224), .B1(n19025), .B2(n16282), .ZN(
        n19030) );
  OAI211_X1 U22103 ( .C1(n19028), .C2(n19027), .A(n19185), .B(n19026), .ZN(
        n19029) );
  NAND4_X1 U22104 ( .A1(n19032), .A2(n19031), .A3(n19030), .A4(n19029), .ZN(
        P2_U2835) );
  NAND2_X1 U22105 ( .A1(n19190), .A2(n19033), .ZN(n19034) );
  XOR2_X1 U22106 ( .A(n19035), .B(n19034), .Z(n19043) );
  AOI22_X1 U22107 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19223), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19236), .ZN(n19036) );
  OAI21_X1 U22108 ( .B1(n19037), .B2(n19228), .A(n19036), .ZN(n19038) );
  AOI211_X1 U22109 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19222), .A(n11600), .B(
        n19038), .ZN(n19042) );
  AOI22_X1 U22110 ( .A1(n19040), .A2(n19224), .B1(n19039), .B2(n16282), .ZN(
        n19041) );
  OAI211_X1 U22111 ( .C1(n19955), .C2(n19043), .A(n19042), .B(n19041), .ZN(
        P2_U2836) );
  NOR2_X1 U22112 ( .A1(n19206), .A2(n19044), .ZN(n19046) );
  XOR2_X1 U22113 ( .A(n19046), .B(n19045), .Z(n19056) );
  INV_X1 U22114 ( .A(n19047), .ZN(n19049) );
  AOI22_X1 U22115 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19236), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19223), .ZN(n19048) );
  OAI21_X1 U22116 ( .B1(n19049), .B2(n19228), .A(n19048), .ZN(n19050) );
  AOI211_X1 U22117 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19222), .A(n11600), .B(
        n19050), .ZN(n19055) );
  OAI22_X1 U22118 ( .A1(n19052), .A2(n19213), .B1(n19051), .B2(n19200), .ZN(
        n19053) );
  INV_X1 U22119 ( .A(n19053), .ZN(n19054) );
  OAI211_X1 U22120 ( .C1(n19955), .C2(n19056), .A(n19055), .B(n19054), .ZN(
        P2_U2837) );
  NAND2_X1 U22121 ( .A1(n19190), .A2(n19057), .ZN(n19058) );
  XNOR2_X1 U22122 ( .A(n19059), .B(n19058), .ZN(n19068) );
  AOI22_X1 U22123 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19236), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19223), .ZN(n19060) );
  OAI21_X1 U22124 ( .B1(n19061), .B2(n19228), .A(n19060), .ZN(n19062) );
  AOI211_X1 U22125 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19222), .A(n11600), .B(
        n19062), .ZN(n19067) );
  INV_X1 U22126 ( .A(n19063), .ZN(n19064) );
  AOI22_X1 U22127 ( .A1(n19065), .A2(n19224), .B1(n19064), .B2(n16282), .ZN(
        n19066) );
  OAI211_X1 U22128 ( .C1(n19955), .C2(n19068), .A(n19067), .B(n19066), .ZN(
        P2_U2838) );
  NOR2_X1 U22129 ( .A1(n19206), .A2(n19069), .ZN(n19071) );
  XOR2_X1 U22130 ( .A(n19071), .B(n19070), .Z(n19079) );
  OAI21_X1 U22131 ( .B1(n11062), .B2(n19197), .A(n19210), .ZN(n19075) );
  INV_X1 U22132 ( .A(n19072), .ZN(n19073) );
  OAI22_X1 U22133 ( .A1(n19073), .A2(n19228), .B1(n19997), .B2(n19178), .ZN(
        n19074) );
  AOI211_X1 U22134 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19236), .A(
        n19075), .B(n19074), .ZN(n19078) );
  AOI22_X1 U22135 ( .A1(n19251), .A2(n19224), .B1(n19076), .B2(n16282), .ZN(
        n19077) );
  OAI211_X1 U22136 ( .C1(n19955), .C2(n19079), .A(n19078), .B(n19077), .ZN(
        P2_U2839) );
  OAI22_X1 U22137 ( .A1(n19080), .A2(n19228), .B1(n19995), .B2(n19178), .ZN(
        n19081) );
  AOI211_X1 U22138 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19222), .A(n11600), .B(
        n19081), .ZN(n19089) );
  NAND2_X1 U22139 ( .A1(n19190), .A2(n19082), .ZN(n19083) );
  XNOR2_X1 U22140 ( .A(n19084), .B(n19083), .ZN(n19087) );
  OAI22_X1 U22141 ( .A1(n19256), .A2(n19213), .B1(n19085), .B2(n19200), .ZN(
        n19086) );
  AOI21_X1 U22142 ( .B1(n19185), .B2(n19087), .A(n19086), .ZN(n19088) );
  OAI211_X1 U22143 ( .C1(n19090), .C2(n19174), .A(n19089), .B(n19088), .ZN(
        P2_U2840) );
  NOR2_X1 U22144 ( .A1(n19206), .A2(n19091), .ZN(n19093) );
  XOR2_X1 U22145 ( .A(n19093), .B(n19092), .Z(n19100) );
  AOI22_X1 U22146 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19223), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19236), .ZN(n19094) );
  OAI21_X1 U22147 ( .B1(n19095), .B2(n19228), .A(n19094), .ZN(n19096) );
  AOI211_X1 U22148 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19222), .A(n11600), .B(
        n19096), .ZN(n19099) );
  AOI22_X1 U22149 ( .A1(n19257), .A2(n19224), .B1(n19097), .B2(n16282), .ZN(
        n19098) );
  OAI211_X1 U22150 ( .C1(n19955), .C2(n19100), .A(n19099), .B(n19098), .ZN(
        P2_U2841) );
  OAI21_X1 U22151 ( .B1(n11293), .B2(n19197), .A(n19210), .ZN(n19105) );
  INV_X1 U22152 ( .A(n19101), .ZN(n19103) );
  OAI22_X1 U22153 ( .A1(n19103), .A2(n19228), .B1(n19174), .B2(n19102), .ZN(
        n19104) );
  AOI211_X1 U22154 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19223), .A(n19105), 
        .B(n19104), .ZN(n19112) );
  NAND2_X1 U22155 ( .A1(n19190), .A2(n19106), .ZN(n19107) );
  XNOR2_X1 U22156 ( .A(n19108), .B(n19107), .ZN(n19110) );
  AOI22_X1 U22157 ( .A1(n19110), .A2(n19185), .B1(n19109), .B2(n16282), .ZN(
        n19111) );
  OAI211_X1 U22158 ( .C1(n19261), .C2(n19213), .A(n19112), .B(n19111), .ZN(
        P2_U2842) );
  OAI21_X1 U22159 ( .B1(n19113), .B2(n19197), .A(n19210), .ZN(n19117) );
  OAI22_X1 U22160 ( .A1(n19115), .A2(n19228), .B1(n19174), .B2(n19114), .ZN(
        n19116) );
  AOI211_X1 U22161 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19223), .A(n19117), 
        .B(n19116), .ZN(n19124) );
  NAND2_X1 U22162 ( .A1(n19190), .A2(n19118), .ZN(n19119) );
  XNOR2_X1 U22163 ( .A(n19120), .B(n19119), .ZN(n19122) );
  AOI22_X1 U22164 ( .A1(n19122), .A2(n19185), .B1(n19121), .B2(n16282), .ZN(
        n19123) );
  OAI211_X1 U22165 ( .C1(n19265), .C2(n19213), .A(n19124), .B(n19123), .ZN(
        P2_U2844) );
  NOR2_X1 U22166 ( .A1(n19206), .A2(n19125), .ZN(n19127) );
  XOR2_X1 U22167 ( .A(n19127), .B(n19126), .Z(n19137) );
  INV_X1 U22168 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19130) );
  AOI22_X1 U22169 ( .A1(n19128), .A2(n19194), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19236), .ZN(n19129) );
  OAI211_X1 U22170 ( .C1(n19130), .C2(n19197), .A(n19129), .B(n19210), .ZN(
        n19131) );
  AOI21_X1 U22171 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n19223), .A(n19131), 
        .ZN(n19136) );
  INV_X1 U22172 ( .A(n19132), .ZN(n19133) );
  AOI22_X1 U22173 ( .A1(n19134), .A2(n19224), .B1(n19133), .B2(n16282), .ZN(
        n19135) );
  OAI211_X1 U22174 ( .C1(n19955), .C2(n19137), .A(n19136), .B(n19135), .ZN(
        P2_U2845) );
  INV_X1 U22175 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19985) );
  INV_X1 U22176 ( .A(n19138), .ZN(n19140) );
  OAI22_X1 U22177 ( .A1(n19140), .A2(n19228), .B1(n19174), .B2(n19139), .ZN(
        n19141) );
  AOI211_X1 U22178 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19222), .A(n11600), .B(
        n19141), .ZN(n19150) );
  NAND2_X1 U22179 ( .A1(n19190), .A2(n19142), .ZN(n19143) );
  XNOR2_X1 U22180 ( .A(n19144), .B(n19143), .ZN(n19148) );
  INV_X1 U22181 ( .A(n19145), .ZN(n19146) );
  OAI22_X1 U22182 ( .A1(n19271), .A2(n19213), .B1(n19146), .B2(n19200), .ZN(
        n19147) );
  AOI21_X1 U22183 ( .B1(n19185), .B2(n19148), .A(n19147), .ZN(n19149) );
  OAI211_X1 U22184 ( .C1(n19985), .C2(n19178), .A(n19150), .B(n19149), .ZN(
        P2_U2846) );
  NOR2_X1 U22185 ( .A1(n19206), .A2(n19151), .ZN(n19153) );
  XOR2_X1 U22186 ( .A(n19153), .B(n19152), .Z(n19162) );
  INV_X1 U22187 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19984) );
  AOI22_X1 U22188 ( .A1(n19154), .A2(n19194), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19236), .ZN(n19155) );
  OAI21_X1 U22189 ( .B1(n19984), .B2(n19178), .A(n19155), .ZN(n19156) );
  AOI211_X1 U22190 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19222), .A(n11600), .B(
        n19156), .ZN(n19161) );
  INV_X1 U22191 ( .A(n19157), .ZN(n19273) );
  OAI22_X1 U22192 ( .A1(n19158), .A2(n19200), .B1(n19213), .B2(n19273), .ZN(
        n19159) );
  INV_X1 U22193 ( .A(n19159), .ZN(n19160) );
  OAI211_X1 U22194 ( .C1(n19955), .C2(n19162), .A(n19161), .B(n19160), .ZN(
        P2_U2847) );
  NAND2_X1 U22195 ( .A1(n19190), .A2(n19163), .ZN(n19165) );
  XOR2_X1 U22196 ( .A(n19165), .B(n19164), .Z(n19173) );
  AOI22_X1 U22197 ( .A1(n19166), .A2(n19194), .B1(P2_REIP_REG_7__SCAN_IN), 
        .B2(n19223), .ZN(n19167) );
  OAI211_X1 U22198 ( .C1(n19168), .C2(n19197), .A(n19167), .B(n19210), .ZN(
        n19171) );
  OAI22_X1 U22199 ( .A1(n19274), .A2(n19213), .B1(n19169), .B2(n19200), .ZN(
        n19170) );
  AOI211_X1 U22200 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19236), .A(
        n19171), .B(n19170), .ZN(n19172) );
  OAI21_X1 U22201 ( .B1(n19173), .B2(n19955), .A(n19172), .ZN(P2_U2848) );
  OAI22_X1 U22202 ( .A1(n19175), .A2(n19228), .B1(n19174), .B2(n10101), .ZN(
        n19176) );
  INV_X1 U22203 ( .A(n19176), .ZN(n19177) );
  OAI21_X1 U22204 ( .B1(n19980), .B2(n19178), .A(n19177), .ZN(n19179) );
  AOI211_X1 U22205 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19222), .A(n19180), .B(
        n19179), .ZN(n19188) );
  NOR2_X1 U22206 ( .A1(n19206), .A2(n19181), .ZN(n19183) );
  XNOR2_X1 U22207 ( .A(n19183), .B(n19182), .ZN(n19186) );
  AOI22_X1 U22208 ( .A1(n19186), .A2(n19185), .B1(n19184), .B2(n16282), .ZN(
        n19187) );
  OAI211_X1 U22209 ( .C1(n19213), .C2(n19276), .A(n19188), .B(n19187), .ZN(
        P2_U2849) );
  NAND2_X1 U22210 ( .A1(n19190), .A2(n19189), .ZN(n19192) );
  XOR2_X1 U22211 ( .A(n19192), .B(n19191), .Z(n19204) );
  INV_X1 U22212 ( .A(n19193), .ZN(n19195) );
  AOI22_X1 U22213 ( .A1(n19195), .A2(n19194), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19236), .ZN(n19196) );
  OAI211_X1 U22214 ( .C1(n19198), .C2(n19197), .A(n19196), .B(n19210), .ZN(
        n19202) );
  OAI22_X1 U22215 ( .A1(n19285), .A2(n19213), .B1(n19200), .B2(n19199), .ZN(
        n19201) );
  AOI211_X1 U22216 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19223), .A(n19202), .B(
        n19201), .ZN(n19203) );
  OAI21_X1 U22217 ( .B1(n19204), .B2(n19955), .A(n19203), .ZN(P2_U2850) );
  NOR2_X1 U22218 ( .A1(n19206), .A2(n19205), .ZN(n19208) );
  XOR2_X1 U22219 ( .A(n19208), .B(n19207), .Z(n19221) );
  NOR2_X1 U22220 ( .A1(n19209), .A2(n19228), .ZN(n19215) );
  AOI22_X1 U22221 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19223), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19222), .ZN(n19211) );
  OAI211_X1 U22222 ( .C1(n19213), .C2(n19212), .A(n19211), .B(n19210), .ZN(
        n19214) );
  AOI211_X1 U22223 ( .C1(n19236), .C2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19215), .B(n19214), .ZN(n19220) );
  INV_X1 U22224 ( .A(n19216), .ZN(n19281) );
  AOI22_X1 U22225 ( .A1(n19281), .A2(n19218), .B1(n16282), .B2(n19217), .ZN(
        n19219) );
  OAI211_X1 U22226 ( .C1(n19955), .C2(n19221), .A(n19220), .B(n19219), .ZN(
        P2_U2851) );
  AOI22_X1 U22227 ( .A1(n19223), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19222), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n19227) );
  NAND2_X1 U22228 ( .A1(n19225), .A2(n19224), .ZN(n19226) );
  OAI211_X1 U22229 ( .C1(n19229), .C2(n19228), .A(n19227), .B(n19226), .ZN(
        n19230) );
  AOI21_X1 U22230 ( .B1(n19231), .B2(n16282), .A(n19230), .ZN(n19232) );
  OAI21_X1 U22231 ( .B1(n20059), .B2(n19233), .A(n19232), .ZN(n19234) );
  INV_X1 U22232 ( .A(n19234), .ZN(n19238) );
  OAI21_X1 U22233 ( .B1(n19236), .B2(n19235), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19237) );
  OAI211_X1 U22234 ( .C1(n19240), .C2(n19239), .A(n19238), .B(n19237), .ZN(
        P2_U2855) );
  AOI22_X1 U22235 ( .A1(n19241), .A2(n19295), .B1(BUF2_REG_31__SCAN_IN), .B2(
        n19248), .ZN(n19243) );
  AOI22_X1 U22236 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19294), .B1(n19247), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19242) );
  NAND2_X1 U22237 ( .A1(n19243), .A2(n19242), .ZN(P2_U2888) );
  INV_X1 U22238 ( .A(n19244), .ZN(n19245) );
  AOI22_X1 U22239 ( .A1(n19246), .A2(n19245), .B1(n19294), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19254) );
  AOI22_X1 U22240 ( .A1(n19248), .A2(BUF2_REG_16__SCAN_IN), .B1(n19247), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19253) );
  NOR2_X1 U22241 ( .A1(n19249), .A2(n19299), .ZN(n19250) );
  AOI21_X1 U22242 ( .B1(n19251), .B2(n19295), .A(n19250), .ZN(n19252) );
  NAND3_X1 U22243 ( .A1(n19254), .A2(n19253), .A3(n19252), .ZN(P2_U2903) );
  OAI222_X1 U22244 ( .A1(n19256), .A2(n19286), .B1(n19347), .B2(n19275), .C1(
        n19255), .C2(n19303), .ZN(P2_U2904) );
  INV_X1 U22245 ( .A(n19257), .ZN(n19259) );
  AOI22_X1 U22246 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19294), .B1(n19377), 
        .B2(n19278), .ZN(n19258) );
  OAI21_X1 U22247 ( .B1(n19286), .B2(n19259), .A(n19258), .ZN(P2_U2905) );
  OAI222_X1 U22248 ( .A1(n19261), .A2(n19286), .B1(n12678), .B2(n19275), .C1(
        n19303), .C2(n19260), .ZN(P2_U2906) );
  OAI222_X1 U22249 ( .A1(n19263), .A2(n19286), .B1(n12673), .B2(n19275), .C1(
        n19303), .C2(n19262), .ZN(P2_U2907) );
  INV_X1 U22250 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19353) );
  OAI222_X1 U22251 ( .A1(n19265), .A2(n19286), .B1(n19353), .B2(n19275), .C1(
        n19303), .C2(n19264), .ZN(P2_U2908) );
  AOI22_X1 U22252 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19294), .B1(n19266), 
        .B2(n19278), .ZN(n19267) );
  OAI21_X1 U22253 ( .B1(n19286), .B2(n19268), .A(n19267), .ZN(P2_U2909) );
  AOI22_X1 U22254 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19294), .B1(n19269), .B2(
        n19278), .ZN(n19270) );
  OAI21_X1 U22255 ( .B1(n19286), .B2(n19271), .A(n19270), .ZN(P2_U2910) );
  INV_X1 U22256 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19359) );
  OAI222_X1 U22257 ( .A1(n19273), .A2(n19286), .B1(n19359), .B2(n19275), .C1(
        n19303), .C2(n19272), .ZN(P2_U2911) );
  INV_X1 U22258 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19361) );
  OAI222_X1 U22259 ( .A1(n19274), .A2(n19286), .B1(n19361), .B2(n19275), .C1(
        n19303), .C2(n19433), .ZN(P2_U2912) );
  INV_X1 U22260 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19364) );
  OAI222_X1 U22261 ( .A1(n19276), .A2(n19286), .B1(n19364), .B2(n19275), .C1(
        n19303), .C2(n19426), .ZN(P2_U2913) );
  INV_X1 U22262 ( .A(n19277), .ZN(n19279) );
  AOI22_X1 U22263 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19294), .B1(n19279), .B2(
        n19278), .ZN(n19284) );
  NAND3_X1 U22264 ( .A1(n19282), .A2(n19281), .A3(n19280), .ZN(n19283) );
  OAI211_X1 U22265 ( .C1(n19286), .C2(n19285), .A(n19284), .B(n19283), .ZN(
        P2_U2914) );
  AOI22_X1 U22266 ( .A1(n19295), .A2(n19287), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19294), .ZN(n19293) );
  AOI21_X1 U22267 ( .B1(n19290), .B2(n19289), .A(n19288), .ZN(n19291) );
  OR2_X1 U22268 ( .A1(n19291), .A2(n19299), .ZN(n19292) );
  OAI211_X1 U22269 ( .C1(n19422), .C2(n19303), .A(n19293), .B(n19292), .ZN(
        P2_U2916) );
  AOI22_X1 U22270 ( .A1(n19295), .A2(n20055), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19294), .ZN(n19302) );
  AOI21_X1 U22271 ( .B1(n19298), .B2(n19297), .A(n19296), .ZN(n19300) );
  OR2_X1 U22272 ( .A1(n19300), .A2(n19299), .ZN(n19301) );
  OAI211_X1 U22273 ( .C1(n19410), .C2(n19303), .A(n19302), .B(n19301), .ZN(
        P2_U2918) );
  NAND2_X1 U22274 ( .A1(n19305), .A2(n19304), .ZN(n19307) );
  NAND2_X1 U22275 ( .A1(n19307), .A2(n19306), .ZN(n19308) );
  NAND2_X1 U22276 ( .A1(n20072), .A2(n19309), .ZN(n19313) );
  NAND2_X1 U22277 ( .A1(n19376), .A2(n19313), .ZN(n19317) );
  NOR2_X1 U22278 ( .A1(n19317), .A2(n19310), .ZN(P2_U2920) );
  INV_X1 U22279 ( .A(n19311), .ZN(n19312) );
  INV_X1 U22280 ( .A(n19344), .ZN(n19314) );
  INV_X1 U22281 ( .A(n19313), .ZN(n19338) );
  CLKBUF_X1 U22282 ( .A(n19338), .Z(n20076) );
  AOI22_X1 U22283 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19314), .B1(n20076), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19315) );
  OAI21_X1 U22284 ( .B1(n19317), .B2(n19316), .A(n19315), .ZN(P2_U2921) );
  AOI22_X1 U22285 ( .A1(n19338), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19318) );
  OAI21_X1 U22286 ( .B1(n20903), .B2(n19344), .A(n19318), .ZN(P2_U2922) );
  AOI22_X1 U22287 ( .A1(n19338), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19319) );
  OAI21_X1 U22288 ( .B1(n19320), .B2(n19344), .A(n19319), .ZN(P2_U2923) );
  AOI22_X1 U22289 ( .A1(n19338), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19321) );
  OAI21_X1 U22290 ( .B1(n19322), .B2(n19344), .A(n19321), .ZN(P2_U2924) );
  AOI22_X1 U22291 ( .A1(n19338), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19323) );
  OAI21_X1 U22292 ( .B1(n19324), .B2(n19344), .A(n19323), .ZN(P2_U2925) );
  AOI22_X1 U22293 ( .A1(n19338), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19325) );
  OAI21_X1 U22294 ( .B1(n19326), .B2(n19344), .A(n19325), .ZN(P2_U2926) );
  AOI22_X1 U22295 ( .A1(n19338), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19327) );
  OAI21_X1 U22296 ( .B1(n19328), .B2(n19344), .A(n19327), .ZN(P2_U2927) );
  INV_X1 U22297 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19330) );
  AOI22_X1 U22298 ( .A1(n19338), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19329) );
  OAI21_X1 U22299 ( .B1(n19330), .B2(n19344), .A(n19329), .ZN(P2_U2928) );
  INV_X1 U22300 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19332) );
  AOI22_X1 U22301 ( .A1(n19338), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19331) );
  OAI21_X1 U22302 ( .B1(n19332), .B2(n19344), .A(n19331), .ZN(P2_U2929) );
  AOI22_X1 U22303 ( .A1(n19338), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19333) );
  OAI21_X1 U22304 ( .B1(n20873), .B2(n19344), .A(n19333), .ZN(P2_U2930) );
  INV_X1 U22305 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19335) );
  AOI22_X1 U22306 ( .A1(n19338), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19334) );
  OAI21_X1 U22307 ( .B1(n19335), .B2(n19344), .A(n19334), .ZN(P2_U2931) );
  AOI22_X1 U22308 ( .A1(n19338), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19336) );
  OAI21_X1 U22309 ( .B1(n19337), .B2(n19344), .A(n19336), .ZN(P2_U2932) );
  INV_X1 U22310 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19340) );
  AOI22_X1 U22311 ( .A1(n19338), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19339) );
  OAI21_X1 U22312 ( .B1(n19340), .B2(n19344), .A(n19339), .ZN(P2_U2933) );
  AOI22_X1 U22313 ( .A1(n20076), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19341) );
  OAI21_X1 U22314 ( .B1(n19342), .B2(n19344), .A(n19341), .ZN(P2_U2934) );
  AOI22_X1 U22315 ( .A1(n20076), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19343) );
  OAI21_X1 U22316 ( .B1(n19345), .B2(n19344), .A(n19343), .ZN(P2_U2935) );
  AOI22_X1 U22317 ( .A1(n20076), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19346) );
  OAI21_X1 U22318 ( .B1(n19347), .B2(n19376), .A(n19346), .ZN(P2_U2936) );
  INV_X1 U22319 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19349) );
  AOI22_X1 U22320 ( .A1(n20076), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19348) );
  OAI21_X1 U22321 ( .B1(n19349), .B2(n19376), .A(n19348), .ZN(P2_U2937) );
  AOI22_X1 U22322 ( .A1(n20076), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19350) );
  OAI21_X1 U22323 ( .B1(n12678), .B2(n19376), .A(n19350), .ZN(P2_U2938) );
  AOI22_X1 U22324 ( .A1(n20076), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19351) );
  OAI21_X1 U22325 ( .B1(n12673), .B2(n19376), .A(n19351), .ZN(P2_U2939) );
  AOI22_X1 U22326 ( .A1(n20076), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19352) );
  OAI21_X1 U22327 ( .B1(n19353), .B2(n19376), .A(n19352), .ZN(P2_U2940) );
  AOI22_X1 U22328 ( .A1(n20076), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19354) );
  OAI21_X1 U22329 ( .B1(n19355), .B2(n19376), .A(n19354), .ZN(P2_U2941) );
  AOI22_X1 U22330 ( .A1(n20076), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19356) );
  OAI21_X1 U22331 ( .B1(n19357), .B2(n19376), .A(n19356), .ZN(P2_U2942) );
  AOI22_X1 U22332 ( .A1(n20076), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19358) );
  OAI21_X1 U22333 ( .B1(n19359), .B2(n19376), .A(n19358), .ZN(P2_U2943) );
  AOI22_X1 U22334 ( .A1(n20076), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19360) );
  OAI21_X1 U22335 ( .B1(n19361), .B2(n19376), .A(n19360), .ZN(P2_U2944) );
  AOI22_X1 U22336 ( .A1(n20076), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19363) );
  OAI21_X1 U22337 ( .B1(n19364), .B2(n19376), .A(n19363), .ZN(P2_U2945) );
  INV_X1 U22338 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19366) );
  AOI22_X1 U22339 ( .A1(n20076), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19365) );
  OAI21_X1 U22340 ( .B1(n19366), .B2(n19376), .A(n19365), .ZN(P2_U2946) );
  INV_X1 U22341 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19368) );
  AOI22_X1 U22342 ( .A1(n20076), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19367) );
  OAI21_X1 U22343 ( .B1(n19368), .B2(n19376), .A(n19367), .ZN(P2_U2947) );
  INV_X1 U22344 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19370) );
  AOI22_X1 U22345 ( .A1(n20076), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19369) );
  OAI21_X1 U22346 ( .B1(n19370), .B2(n19376), .A(n19369), .ZN(P2_U2948) );
  INV_X1 U22347 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19372) );
  AOI22_X1 U22348 ( .A1(n20076), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19371) );
  OAI21_X1 U22349 ( .B1(n19372), .B2(n19376), .A(n19371), .ZN(P2_U2949) );
  INV_X1 U22350 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19374) );
  AOI22_X1 U22351 ( .A1(n20076), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19373) );
  OAI21_X1 U22352 ( .B1(n19374), .B2(n19376), .A(n19373), .ZN(P2_U2950) );
  AOI22_X1 U22353 ( .A1(n20076), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19362), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19375) );
  OAI21_X1 U22354 ( .B1(n12723), .B2(n19376), .A(n19375), .ZN(P2_U2951) );
  AOI22_X1 U22355 ( .A1(n19381), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19380), .ZN(n19379) );
  NAND2_X1 U22356 ( .A1(n19378), .A2(n19377), .ZN(n19382) );
  NAND2_X1 U22357 ( .A1(n19379), .A2(n19382), .ZN(P2_U2966) );
  AOI22_X1 U22358 ( .A1(n19381), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19380), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19383) );
  NAND2_X1 U22359 ( .A1(n19383), .A2(n19382), .ZN(P2_U2981) );
  NAND2_X1 U22360 ( .A1(n19384), .A2(n19388), .ZN(n19386) );
  OAI211_X1 U22361 ( .C1(n19388), .C2(n19387), .A(n19386), .B(n19385), .ZN(
        n19389) );
  INV_X1 U22362 ( .A(n19389), .ZN(n19409) );
  INV_X1 U22363 ( .A(n19390), .ZN(n19394) );
  AOI22_X1 U22364 ( .A1(n19394), .A2(n19393), .B1(n19392), .B2(n19391), .ZN(
        n19407) );
  NAND2_X1 U22365 ( .A1(n19396), .A2(n19395), .ZN(n19403) );
  NAND2_X1 U22366 ( .A1(n19180), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19397) );
  OAI211_X1 U22367 ( .C1(n19400), .C2(n19399), .A(n19398), .B(n19397), .ZN(
        n19401) );
  INV_X1 U22368 ( .A(n19401), .ZN(n19402) );
  OAI211_X1 U22369 ( .C1(n10769), .C2(n19404), .A(n19403), .B(n19402), .ZN(
        n19405) );
  INV_X1 U22370 ( .A(n19405), .ZN(n19406) );
  OAI211_X1 U22371 ( .C1(n19409), .C2(n19408), .A(n19407), .B(n19406), .ZN(
        P2_U3044) );
  AOI22_X1 U22372 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19435), .ZN(n19905) );
  INV_X1 U22373 ( .A(n19905), .ZN(n19786) );
  NOR2_X2 U22374 ( .A1(n11377), .A2(n19414), .ZN(n19900) );
  AOI22_X1 U22375 ( .A1(n19786), .A2(n19927), .B1(n19432), .B2(n19900), .ZN(
        n19412) );
  NOR2_X2 U22376 ( .A1(n19410), .A2(n9715), .ZN(n19901) );
  AOI22_X1 U22377 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19435), .ZN(n19789) );
  INV_X1 U22378 ( .A(n19789), .ZN(n19902) );
  AOI22_X1 U22379 ( .A1(n19901), .A2(n19436), .B1(n19465), .B2(n19902), .ZN(
        n19411) );
  OAI211_X1 U22380 ( .C1(n19439), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P2_U3049) );
  AOI22_X1 U22381 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19435), .ZN(n19911) );
  INV_X1 U22382 ( .A(n19911), .ZN(n19685) );
  NOR2_X2 U22383 ( .A1(n10668), .A2(n19414), .ZN(n19906) );
  AOI22_X1 U22384 ( .A1(n19685), .A2(n19927), .B1(n19432), .B2(n19906), .ZN(
        n19417) );
  NOR2_X2 U22385 ( .A1(n19415), .A2(n9715), .ZN(n19907) );
  AOI22_X1 U22386 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19435), .ZN(n19688) );
  AOI22_X1 U22387 ( .A1(n19907), .A2(n19436), .B1(n19465), .B2(n19908), .ZN(
        n19416) );
  OAI211_X1 U22388 ( .C1(n19439), .C2(n12337), .A(n19417), .B(n19416), .ZN(
        P2_U3050) );
  OAI22_X2 U22389 ( .A1(n14650), .A2(n19420), .B1(n19419), .B2(n19418), .ZN(
        n19914) );
  AND2_X1 U22390 ( .A1(n19421), .A2(n19430), .ZN(n19912) );
  AOI22_X1 U22391 ( .A1(n19914), .A2(n19927), .B1(n19432), .B2(n19912), .ZN(
        n19425) );
  NOR2_X2 U22392 ( .A1(n19422), .A2(n9715), .ZN(n19913) );
  AOI22_X2 U22393 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19435), .ZN(n19917) );
  INV_X1 U22394 ( .A(n19917), .ZN(n19423) );
  AOI22_X1 U22395 ( .A1(n19913), .A2(n19436), .B1(n19465), .B2(n19423), .ZN(
        n19424) );
  OAI211_X1 U22396 ( .C1(n19439), .C2(n12320), .A(n19425), .B(n19424), .ZN(
        P2_U3051) );
  AOI22_X1 U22397 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19435), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19434), .ZN(n19802) );
  AND2_X1 U22398 ( .A1(n10656), .A2(n19430), .ZN(n19932) );
  AOI22_X1 U22399 ( .A1(n19934), .A2(n19927), .B1(n19432), .B2(n19932), .ZN(
        n19428) );
  NOR2_X2 U22400 ( .A1(n19426), .A2(n9715), .ZN(n19933) );
  AOI22_X1 U22401 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19435), .ZN(n19937) );
  INV_X1 U22402 ( .A(n19937), .ZN(n19798) );
  AOI22_X1 U22403 ( .A1(n19933), .A2(n19436), .B1(n19465), .B2(n19798), .ZN(
        n19427) );
  OAI211_X1 U22404 ( .C1(n19439), .C2(n19429), .A(n19428), .B(n19427), .ZN(
        P2_U3054) );
  AOI22_X1 U22405 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19434), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19435), .ZN(n19845) );
  AOI22_X1 U22406 ( .A1(n19942), .A2(n19927), .B1(n19432), .B2(n19938), .ZN(
        n19438) );
  NOR2_X2 U22407 ( .A1(n19433), .A2(n9715), .ZN(n19940) );
  INV_X1 U22408 ( .A(n19948), .ZN(n19840) );
  AOI22_X1 U22409 ( .A1(n19940), .A2(n19436), .B1(n19465), .B2(n19840), .ZN(
        n19437) );
  OAI211_X1 U22410 ( .C1(n19439), .C2(n10185), .A(n19438), .B(n19437), .ZN(
        P2_U3055) );
  NOR2_X1 U22411 ( .A1(n19671), .A2(n19501), .ZN(n19463) );
  INV_X1 U22412 ( .A(n19463), .ZN(n19444) );
  NAND2_X1 U22413 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19444), .ZN(n19440) );
  OR2_X1 U22414 ( .A1(n19441), .A2(n19440), .ZN(n19446) );
  OAI21_X1 U22415 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19443), .A(n12754), 
        .ZN(n19442) );
  AND2_X1 U22416 ( .A1(n19446), .A2(n19442), .ZN(n19464) );
  AOI22_X1 U22417 ( .A1(n19464), .A2(n19887), .B1(n19886), .B2(n19463), .ZN(
        n19449) );
  AND2_X1 U22418 ( .A1(n19672), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19611) );
  INV_X1 U22419 ( .A(n19611), .ZN(n19550) );
  OAI21_X1 U22420 ( .B1(n19550), .B2(n19673), .A(n19443), .ZN(n19447) );
  NAND2_X1 U22421 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19444), .ZN(n19445) );
  NAND4_X1 U22422 ( .A1(n19447), .A2(n19889), .A3(n19446), .A4(n19445), .ZN(
        n19466) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19820), .ZN(n19448) );
  OAI211_X1 U22424 ( .C1(n19749), .C2(n19492), .A(n19449), .B(n19448), .ZN(
        P2_U3056) );
  AOI22_X1 U22425 ( .A1(n19464), .A2(n19901), .B1(n19900), .B2(n19463), .ZN(
        n19451) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19786), .ZN(n19450) );
  OAI211_X1 U22427 ( .C1(n19789), .C2(n19492), .A(n19451), .B(n19450), .ZN(
        P2_U3057) );
  AOI22_X1 U22428 ( .A1(n19464), .A2(n19907), .B1(n19906), .B2(n19463), .ZN(
        n19453) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19685), .ZN(n19452) );
  OAI211_X1 U22430 ( .C1(n19688), .C2(n19492), .A(n19453), .B(n19452), .ZN(
        P2_U3058) );
  AOI22_X1 U22431 ( .A1(n19464), .A2(n19913), .B1(n19912), .B2(n19463), .ZN(
        n19455) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19914), .ZN(n19454) );
  OAI211_X1 U22433 ( .C1(n19917), .C2(n19492), .A(n19455), .B(n19454), .ZN(
        P2_U3059) );
  AOI22_X1 U22434 ( .A1(n19464), .A2(n19919), .B1(n19918), .B2(n19463), .ZN(
        n19457) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19867), .ZN(n19456) );
  OAI211_X1 U22436 ( .C1(n19870), .C2(n19492), .A(n19457), .B(n19456), .ZN(
        P2_U3060) );
  AOI22_X1 U22437 ( .A1(n19464), .A2(n19925), .B1(n19924), .B2(n19463), .ZN(
        n19460) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19832), .ZN(n19459) );
  OAI211_X1 U22439 ( .C1(n19598), .C2(n19492), .A(n19460), .B(n19459), .ZN(
        P2_U3061) );
  AOI22_X1 U22440 ( .A1(n19464), .A2(n19933), .B1(n19932), .B2(n19463), .ZN(
        n19462) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19934), .ZN(n19461) );
  OAI211_X1 U22442 ( .C1(n19937), .C2(n19492), .A(n19462), .B(n19461), .ZN(
        P2_U3062) );
  AOI22_X1 U22443 ( .A1(n19464), .A2(n19940), .B1(n19938), .B2(n19463), .ZN(
        n19468) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19942), .ZN(n19467) );
  OAI211_X1 U22445 ( .C1(n19948), .C2(n19492), .A(n19468), .B(n19467), .ZN(
        P2_U3063) );
  INV_X1 U22446 ( .A(n19474), .ZN(n19469) );
  NOR2_X1 U22447 ( .A1(n19705), .A2(n19501), .ZN(n19495) );
  OAI21_X1 U22448 ( .B1(n19469), .B2(n19495), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19472) );
  INV_X1 U22449 ( .A(n19501), .ZN(n19470) );
  NAND2_X1 U22450 ( .A1(n19471), .A2(n19470), .ZN(n19475) );
  NAND2_X1 U22451 ( .A1(n19472), .A2(n19475), .ZN(n19496) );
  AOI22_X1 U22452 ( .A1(n19496), .A2(n19887), .B1(n19886), .B2(n19495), .ZN(
        n19481) );
  INV_X1 U22453 ( .A(n19495), .ZN(n19473) );
  OAI21_X1 U22454 ( .B1(n19474), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19473), 
        .ZN(n19478) );
  OAI21_X1 U22455 ( .B1(n19526), .B2(n19497), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19476) );
  NAND2_X1 U22456 ( .A1(n19476), .A2(n19475), .ZN(n19477) );
  MUX2_X1 U22457 ( .A(n19478), .B(n19477), .S(n20029), .Z(n19479) );
  NAND2_X1 U22458 ( .A1(n19479), .A2(n19889), .ZN(n19498) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19498), .B1(
        n19526), .B2(n19896), .ZN(n19480) );
  OAI211_X1 U22460 ( .C1(n19899), .C2(n19492), .A(n19481), .B(n19480), .ZN(
        P2_U3064) );
  AOI22_X1 U22461 ( .A1(n19496), .A2(n19901), .B1(n19900), .B2(n19495), .ZN(
        n19483) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19498), .B1(
        n19526), .B2(n19902), .ZN(n19482) );
  OAI211_X1 U22463 ( .C1(n19905), .C2(n19492), .A(n19483), .B(n19482), .ZN(
        P2_U3065) );
  AOI22_X1 U22464 ( .A1(n19496), .A2(n19907), .B1(n19906), .B2(n19495), .ZN(
        n19485) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19498), .B1(
        n19526), .B2(n19908), .ZN(n19484) );
  OAI211_X1 U22466 ( .C1(n19911), .C2(n19492), .A(n19485), .B(n19484), .ZN(
        P2_U3066) );
  AOI22_X1 U22467 ( .A1(n19496), .A2(n19913), .B1(n19912), .B2(n19495), .ZN(
        n19487) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19914), .ZN(n19486) );
  OAI211_X1 U22469 ( .C1(n19917), .C2(n19524), .A(n19487), .B(n19486), .ZN(
        P2_U3067) );
  AOI22_X1 U22470 ( .A1(n19496), .A2(n19919), .B1(n19918), .B2(n19495), .ZN(
        n19489) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19867), .ZN(n19488) );
  OAI211_X1 U22472 ( .C1(n19870), .C2(n19524), .A(n19489), .B(n19488), .ZN(
        P2_U3068) );
  AOI22_X1 U22473 ( .A1(n19496), .A2(n19925), .B1(n19924), .B2(n19495), .ZN(
        n19491) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19498), .B1(
        n19526), .B2(n19926), .ZN(n19490) );
  OAI211_X1 U22475 ( .C1(n19931), .C2(n19492), .A(n19491), .B(n19490), .ZN(
        P2_U3069) );
  AOI22_X1 U22476 ( .A1(n19496), .A2(n19933), .B1(n19932), .B2(n19495), .ZN(
        n19494) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19934), .ZN(n19493) );
  OAI211_X1 U22478 ( .C1(n19937), .C2(n19524), .A(n19494), .B(n19493), .ZN(
        P2_U3070) );
  AOI22_X1 U22479 ( .A1(n19496), .A2(n19940), .B1(n19938), .B2(n19495), .ZN(
        n19500) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19498), .B1(
        n19497), .B2(n19942), .ZN(n19499) );
  OAI211_X1 U22481 ( .C1(n19948), .C2(n19524), .A(n19500), .B(n19499), .ZN(
        P2_U3071) );
  NOR2_X1 U22482 ( .A1(n19739), .A2(n19501), .ZN(n19525) );
  AOI22_X1 U22483 ( .A1(n19896), .A2(n19546), .B1(n19886), .B2(n19525), .ZN(
        n19511) );
  OAI21_X1 U22484 ( .B1(n19550), .B2(n20030), .A(n20029), .ZN(n19509) );
  NOR2_X1 U22485 ( .A1(n10880), .A2(n19501), .ZN(n19505) );
  OAI21_X1 U22486 ( .B1(n19506), .B2(n12754), .A(n20037), .ZN(n19503) );
  INV_X1 U22487 ( .A(n19525), .ZN(n19502) );
  AOI21_X1 U22488 ( .B1(n19503), .B2(n19502), .A(n9715), .ZN(n19504) );
  OAI21_X1 U22489 ( .B1(n19509), .B2(n19505), .A(n19504), .ZN(n19528) );
  INV_X1 U22490 ( .A(n19505), .ZN(n19508) );
  OAI21_X1 U22491 ( .B1(n19506), .B2(n19525), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19507) );
  OAI21_X1 U22492 ( .B1(n19509), .B2(n19508), .A(n19507), .ZN(n19527) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19528), .B1(
        n19887), .B2(n19527), .ZN(n19510) );
  OAI211_X1 U22494 ( .C1(n19899), .C2(n19524), .A(n19511), .B(n19510), .ZN(
        P2_U3072) );
  AOI22_X1 U22495 ( .A1(n19786), .A2(n19526), .B1(n19525), .B2(n19900), .ZN(
        n19513) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19528), .B1(
        n19901), .B2(n19527), .ZN(n19512) );
  OAI211_X1 U22497 ( .C1(n19789), .C2(n19541), .A(n19513), .B(n19512), .ZN(
        P2_U3073) );
  AOI22_X1 U22498 ( .A1(n19908), .A2(n19546), .B1(n19525), .B2(n19906), .ZN(
        n19515) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19528), .B1(
        n19907), .B2(n19527), .ZN(n19514) );
  OAI211_X1 U22500 ( .C1(n19911), .C2(n19524), .A(n19515), .B(n19514), .ZN(
        P2_U3074) );
  AOI22_X1 U22501 ( .A1(n19914), .A2(n19526), .B1(n19525), .B2(n19912), .ZN(
        n19517) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19528), .B1(
        n19913), .B2(n19527), .ZN(n19516) );
  OAI211_X1 U22503 ( .C1(n19917), .C2(n19541), .A(n19517), .B(n19516), .ZN(
        P2_U3075) );
  AOI22_X1 U22504 ( .A1(n19867), .A2(n19526), .B1(n19918), .B2(n19525), .ZN(
        n19519) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19528), .B1(
        n19919), .B2(n19527), .ZN(n19518) );
  OAI211_X1 U22506 ( .C1(n19870), .C2(n19541), .A(n19519), .B(n19518), .ZN(
        P2_U3076) );
  AOI22_X1 U22507 ( .A1(n19832), .A2(n19526), .B1(n19924), .B2(n19525), .ZN(
        n19521) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19528), .B1(
        n19925), .B2(n19527), .ZN(n19520) );
  OAI211_X1 U22509 ( .C1(n19598), .C2(n19541), .A(n19521), .B(n19520), .ZN(
        P2_U3077) );
  AOI22_X1 U22510 ( .A1(n19798), .A2(n19546), .B1(n19525), .B2(n19932), .ZN(
        n19523) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19528), .B1(
        n19933), .B2(n19527), .ZN(n19522) );
  OAI211_X1 U22512 ( .C1(n19802), .C2(n19524), .A(n19523), .B(n19522), .ZN(
        P2_U3078) );
  AOI22_X1 U22513 ( .A1(n19942), .A2(n19526), .B1(n19525), .B2(n19938), .ZN(
        n19530) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19528), .B1(
        n19940), .B2(n19527), .ZN(n19529) );
  OAI211_X1 U22515 ( .C1(n19948), .C2(n19541), .A(n19530), .B(n19529), .ZN(
        P2_U3079) );
  AOI22_X1 U22516 ( .A1(n19545), .A2(n19901), .B1(n19900), .B2(n19544), .ZN(
        n19532) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19547), .B1(
        n19564), .B2(n19902), .ZN(n19531) );
  OAI211_X1 U22518 ( .C1(n19905), .C2(n19541), .A(n19532), .B(n19531), .ZN(
        P2_U3081) );
  AOI22_X1 U22519 ( .A1(n19545), .A2(n19907), .B1(n19906), .B2(n19544), .ZN(
        n19534) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19547), .B1(
        n19564), .B2(n19908), .ZN(n19533) );
  OAI211_X1 U22521 ( .C1(n19911), .C2(n19541), .A(n19534), .B(n19533), .ZN(
        P2_U3082) );
  AOI22_X1 U22522 ( .A1(n19545), .A2(n19913), .B1(n19912), .B2(n19544), .ZN(
        n19536) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19547), .B1(
        n19546), .B2(n19914), .ZN(n19535) );
  OAI211_X1 U22524 ( .C1(n19917), .C2(n19578), .A(n19536), .B(n19535), .ZN(
        P2_U3083) );
  AOI22_X1 U22525 ( .A1(n19545), .A2(n19919), .B1(n19918), .B2(n19544), .ZN(
        n19538) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19547), .B1(
        n19564), .B2(n19920), .ZN(n19537) );
  OAI211_X1 U22527 ( .C1(n19923), .C2(n19541), .A(n19538), .B(n19537), .ZN(
        P2_U3084) );
  AOI22_X1 U22528 ( .A1(n19545), .A2(n19925), .B1(n19924), .B2(n19544), .ZN(
        n19540) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19547), .B1(
        n19564), .B2(n19926), .ZN(n19539) );
  OAI211_X1 U22530 ( .C1(n19931), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3085) );
  AOI22_X1 U22531 ( .A1(n19545), .A2(n19933), .B1(n19932), .B2(n19544), .ZN(
        n19543) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19547), .B1(
        n19546), .B2(n19934), .ZN(n19542) );
  OAI211_X1 U22533 ( .C1(n19937), .C2(n19578), .A(n19543), .B(n19542), .ZN(
        P2_U3086) );
  AOI22_X1 U22534 ( .A1(n19545), .A2(n19940), .B1(n19938), .B2(n19544), .ZN(
        n19549) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19547), .B1(
        n19546), .B2(n19942), .ZN(n19548) );
  OAI211_X1 U22536 ( .C1(n19948), .C2(n19578), .A(n19549), .B(n19548), .ZN(
        P2_U3087) );
  NOR2_X1 U22537 ( .A1(n21022), .A2(n19556), .ZN(n19580) );
  AOI22_X1 U22538 ( .A1(n19820), .A2(n19564), .B1(n19886), .B2(n19580), .ZN(
        n19559) );
  OAI21_X1 U22539 ( .B1(n19550), .B2(n19817), .A(n20029), .ZN(n19557) );
  INV_X1 U22540 ( .A(n19556), .ZN(n19554) );
  INV_X1 U22541 ( .A(n10941), .ZN(n19552) );
  INV_X1 U22542 ( .A(n20029), .ZN(n19852) );
  INV_X1 U22543 ( .A(n19580), .ZN(n19551) );
  OAI211_X1 U22544 ( .C1(n19552), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19852), 
        .B(n19551), .ZN(n19553) );
  OAI211_X1 U22545 ( .C1(n19557), .C2(n19554), .A(n19889), .B(n19553), .ZN(
        n19575) );
  OAI21_X1 U22546 ( .B1(n10941), .B2(n19580), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19555) );
  OAI21_X1 U22547 ( .B1(n19557), .B2(n19556), .A(n19555), .ZN(n19574) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19575), .B1(
        n19887), .B2(n19574), .ZN(n19558) );
  OAI211_X1 U22549 ( .C1(n19749), .C2(n19567), .A(n19559), .B(n19558), .ZN(
        P2_U3088) );
  AOI22_X1 U22550 ( .A1(n19786), .A2(n19564), .B1(n19580), .B2(n19900), .ZN(
        n19561) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19575), .B1(
        n19901), .B2(n19574), .ZN(n19560) );
  OAI211_X1 U22552 ( .C1(n19789), .C2(n19567), .A(n19561), .B(n19560), .ZN(
        P2_U3089) );
  AOI22_X1 U22553 ( .A1(n19685), .A2(n19564), .B1(n19906), .B2(n19580), .ZN(
        n19563) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19575), .B1(
        n19907), .B2(n19574), .ZN(n19562) );
  OAI211_X1 U22555 ( .C1(n19688), .C2(n19567), .A(n19563), .B(n19562), .ZN(
        P2_U3090) );
  AOI22_X1 U22556 ( .A1(n19914), .A2(n19564), .B1(n19580), .B2(n19912), .ZN(
        n19566) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19575), .B1(
        n19913), .B2(n19574), .ZN(n19565) );
  OAI211_X1 U22558 ( .C1(n19917), .C2(n19567), .A(n19566), .B(n19565), .ZN(
        P2_U3091) );
  AOI22_X1 U22559 ( .A1(n19920), .A2(n19603), .B1(n19918), .B2(n19580), .ZN(
        n19569) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19575), .B1(
        n19919), .B2(n19574), .ZN(n19568) );
  OAI211_X1 U22561 ( .C1(n19923), .C2(n19578), .A(n19569), .B(n19568), .ZN(
        P2_U3092) );
  AOI22_X1 U22562 ( .A1(n19926), .A2(n19603), .B1(n19924), .B2(n19580), .ZN(
        n19571) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19575), .B1(
        n19925), .B2(n19574), .ZN(n19570) );
  OAI211_X1 U22564 ( .C1(n19931), .C2(n19578), .A(n19571), .B(n19570), .ZN(
        P2_U3093) );
  AOI22_X1 U22565 ( .A1(n19798), .A2(n19603), .B1(n19932), .B2(n19580), .ZN(
        n19573) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19575), .B1(
        n19933), .B2(n19574), .ZN(n19572) );
  OAI211_X1 U22567 ( .C1(n19802), .C2(n19578), .A(n19573), .B(n19572), .ZN(
        P2_U3094) );
  AOI22_X1 U22568 ( .A1(n19840), .A2(n19603), .B1(n19580), .B2(n19938), .ZN(
        n19577) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19575), .B1(
        n19940), .B2(n19574), .ZN(n19576) );
  OAI211_X1 U22570 ( .C1(n19845), .C2(n19578), .A(n19577), .B(n19576), .ZN(
        P2_U3095) );
  NAND2_X1 U22571 ( .A1(n12315), .A2(n19883), .ZN(n19609) );
  NOR2_X1 U22572 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19609), .ZN(
        n19601) );
  NOR2_X1 U22573 ( .A1(n19580), .A2(n19601), .ZN(n19583) );
  OAI21_X1 U22574 ( .B1(n10939), .B2(n19601), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19581) );
  OAI21_X1 U22575 ( .B1(n19583), .B2(n19852), .A(n19581), .ZN(n19602) );
  AOI22_X1 U22576 ( .A1(n19602), .A2(n19887), .B1(n19886), .B2(n19601), .ZN(
        n19587) );
  OAI21_X1 U22577 ( .B1(n19603), .B2(n19630), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19584) );
  AOI211_X1 U22578 ( .C1(n10939), .C2(n20037), .A(n20029), .B(n19601), .ZN(
        n19582) );
  AOI211_X1 U22579 ( .C1(n19584), .C2(n19583), .A(n9715), .B(n19582), .ZN(
        n19585) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19820), .ZN(n19586) );
  OAI211_X1 U22581 ( .C1(n19749), .C2(n19637), .A(n19587), .B(n19586), .ZN(
        P2_U3096) );
  AOI22_X1 U22582 ( .A1(n19602), .A2(n19901), .B1(n19900), .B2(n19601), .ZN(
        n19589) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19786), .ZN(n19588) );
  OAI211_X1 U22584 ( .C1(n19789), .C2(n19637), .A(n19589), .B(n19588), .ZN(
        P2_U3097) );
  AOI22_X1 U22585 ( .A1(n19602), .A2(n19907), .B1(n19906), .B2(n19601), .ZN(
        n19591) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19685), .ZN(n19590) );
  OAI211_X1 U22587 ( .C1(n19688), .C2(n19637), .A(n19591), .B(n19590), .ZN(
        P2_U3098) );
  AOI22_X1 U22588 ( .A1(n19602), .A2(n19913), .B1(n19912), .B2(n19601), .ZN(
        n19593) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19914), .ZN(n19592) );
  OAI211_X1 U22590 ( .C1(n19917), .C2(n19637), .A(n19593), .B(n19592), .ZN(
        P2_U3099) );
  AOI22_X1 U22591 ( .A1(n19602), .A2(n19919), .B1(n19918), .B2(n19601), .ZN(
        n19595) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19867), .ZN(n19594) );
  OAI211_X1 U22593 ( .C1(n19870), .C2(n19637), .A(n19595), .B(n19594), .ZN(
        P2_U3100) );
  AOI22_X1 U22594 ( .A1(n19602), .A2(n19925), .B1(n19924), .B2(n19601), .ZN(
        n19597) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19832), .ZN(n19596) );
  OAI211_X1 U22596 ( .C1(n19598), .C2(n19637), .A(n19597), .B(n19596), .ZN(
        P2_U3101) );
  AOI22_X1 U22597 ( .A1(n19602), .A2(n19933), .B1(n19932), .B2(n19601), .ZN(
        n19600) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19934), .ZN(n19599) );
  OAI211_X1 U22599 ( .C1(n19937), .C2(n19637), .A(n19600), .B(n19599), .ZN(
        P2_U3102) );
  AOI22_X1 U22600 ( .A1(n19602), .A2(n19940), .B1(n19938), .B2(n19601), .ZN(
        n19606) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19942), .ZN(n19605) );
  OAI211_X1 U22602 ( .C1(n19948), .C2(n19637), .A(n19606), .B(n19605), .ZN(
        P2_U3103) );
  NOR2_X1 U22603 ( .A1(n21022), .A2(n19609), .ZN(n19645) );
  INV_X1 U22604 ( .A(n19645), .ZN(n19642) );
  NAND2_X1 U22605 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19642), .ZN(n19607) );
  NOR2_X1 U22606 ( .A1(n19608), .A2(n19607), .ZN(n19614) );
  INV_X1 U22607 ( .A(n19609), .ZN(n19616) );
  AOI21_X1 U22608 ( .B1(n20037), .B2(n19616), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19610) );
  NOR2_X1 U22609 ( .A1(n19614), .A2(n19610), .ZN(n19633) );
  AOI22_X1 U22610 ( .A1(n19633), .A2(n19887), .B1(n19886), .B2(n19645), .ZN(
        n19619) );
  INV_X1 U22611 ( .A(n19893), .ZN(n19846) );
  AND2_X1 U22612 ( .A1(n19611), .A2(n19846), .ZN(n20028) );
  AND2_X1 U22613 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19642), .ZN(n19612) );
  NOR3_X1 U22614 ( .A1(n19614), .A2(n9715), .A3(n19612), .ZN(n19615) );
  OAI21_X1 U22615 ( .B1(n19616), .B2(n20028), .A(n19615), .ZN(n19634) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19634), .B1(
        n19665), .B2(n19896), .ZN(n19618) );
  OAI211_X1 U22617 ( .C1(n19899), .C2(n19637), .A(n19619), .B(n19618), .ZN(
        P2_U3104) );
  AOI22_X1 U22618 ( .A1(n19633), .A2(n19901), .B1(n19900), .B2(n19645), .ZN(
        n19621) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19634), .B1(
        n19665), .B2(n19902), .ZN(n19620) );
  OAI211_X1 U22620 ( .C1(n19905), .C2(n19637), .A(n19621), .B(n19620), .ZN(
        P2_U3105) );
  AOI22_X1 U22621 ( .A1(n19633), .A2(n19907), .B1(n19906), .B2(n19645), .ZN(
        n19623) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19634), .B1(
        n19665), .B2(n19908), .ZN(n19622) );
  OAI211_X1 U22623 ( .C1(n19911), .C2(n19637), .A(n19623), .B(n19622), .ZN(
        P2_U3106) );
  AOI22_X1 U22624 ( .A1(n19633), .A2(n19913), .B1(n19912), .B2(n19645), .ZN(
        n19625) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19634), .B1(
        n19630), .B2(n19914), .ZN(n19624) );
  OAI211_X1 U22626 ( .C1(n19917), .C2(n19661), .A(n19625), .B(n19624), .ZN(
        P2_U3107) );
  AOI22_X1 U22627 ( .A1(n19633), .A2(n19919), .B1(n19918), .B2(n19645), .ZN(
        n19627) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19634), .B1(
        n19665), .B2(n19920), .ZN(n19626) );
  OAI211_X1 U22629 ( .C1(n19923), .C2(n19637), .A(n19627), .B(n19626), .ZN(
        P2_U3108) );
  AOI22_X1 U22630 ( .A1(n19633), .A2(n19925), .B1(n19924), .B2(n19645), .ZN(
        n19629) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19634), .B1(
        n19665), .B2(n19926), .ZN(n19628) );
  OAI211_X1 U22632 ( .C1(n19931), .C2(n19637), .A(n19629), .B(n19628), .ZN(
        P2_U3109) );
  AOI22_X1 U22633 ( .A1(n19633), .A2(n19933), .B1(n19932), .B2(n19645), .ZN(
        n19632) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19634), .B1(
        n19630), .B2(n19934), .ZN(n19631) );
  OAI211_X1 U22635 ( .C1(n19937), .C2(n19661), .A(n19632), .B(n19631), .ZN(
        P2_U3110) );
  AOI22_X1 U22636 ( .A1(n19633), .A2(n19940), .B1(n19938), .B2(n19645), .ZN(
        n19636) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19634), .B1(
        n19665), .B2(n19840), .ZN(n19635) );
  OAI211_X1 U22638 ( .C1(n19845), .C2(n19637), .A(n19636), .B(n19635), .ZN(
        P2_U3111) );
  NAND2_X1 U22639 ( .A1(n20047), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19744) );
  INV_X1 U22640 ( .A(n19744), .ZN(n19738) );
  NAND2_X1 U22641 ( .A1(n19738), .A2(n10880), .ZN(n19679) );
  NOR2_X1 U22642 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19679), .ZN(
        n19664) );
  AOI22_X1 U22643 ( .A1(n19699), .A2(n19896), .B1(n19886), .B2(n19664), .ZN(
        n19650) );
  AOI21_X1 U22644 ( .B1(n19697), .B2(n19661), .A(n19770), .ZN(n19639) );
  NOR2_X1 U22645 ( .A1(n19639), .A2(n19852), .ZN(n19644) );
  INV_X1 U22646 ( .A(n19640), .ZN(n19646) );
  AOI21_X1 U22647 ( .B1(n19646), .B2(n20037), .A(n20029), .ZN(n19641) );
  AOI21_X1 U22648 ( .B1(n19644), .B2(n19642), .A(n19641), .ZN(n19643) );
  OAI21_X1 U22649 ( .B1(n19664), .B2(n19643), .A(n19889), .ZN(n19667) );
  OAI21_X1 U22650 ( .B1(n19664), .B2(n19645), .A(n19644), .ZN(n19648) );
  OAI21_X1 U22651 ( .B1(n19646), .B2(n19664), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19647) );
  NAND2_X1 U22652 ( .A1(n19648), .A2(n19647), .ZN(n19666) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19667), .B1(
        n19887), .B2(n19666), .ZN(n19649) );
  OAI211_X1 U22654 ( .C1(n19899), .C2(n19661), .A(n19650), .B(n19649), .ZN(
        P2_U3112) );
  AOI22_X1 U22655 ( .A1(n19902), .A2(n19699), .B1(n19900), .B2(n19664), .ZN(
        n19652) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19901), .ZN(n19651) );
  OAI211_X1 U22657 ( .C1(n19905), .C2(n19661), .A(n19652), .B(n19651), .ZN(
        P2_U3113) );
  AOI22_X1 U22658 ( .A1(n19685), .A2(n19665), .B1(n19906), .B2(n19664), .ZN(
        n19654) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19907), .ZN(n19653) );
  OAI211_X1 U22660 ( .C1(n19688), .C2(n19697), .A(n19654), .B(n19653), .ZN(
        P2_U3114) );
  AOI22_X1 U22661 ( .A1(n19914), .A2(n19665), .B1(n19912), .B2(n19664), .ZN(
        n19656) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19913), .ZN(n19655) );
  OAI211_X1 U22663 ( .C1(n19917), .C2(n19697), .A(n19656), .B(n19655), .ZN(
        P2_U3115) );
  AOI22_X1 U22664 ( .A1(n19920), .A2(n19699), .B1(n19918), .B2(n19664), .ZN(
        n19658) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19919), .ZN(n19657) );
  OAI211_X1 U22666 ( .C1(n19923), .C2(n19661), .A(n19658), .B(n19657), .ZN(
        P2_U3116) );
  AOI22_X1 U22667 ( .A1(n19699), .A2(n19926), .B1(n19924), .B2(n19664), .ZN(
        n19660) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19925), .ZN(n19659) );
  OAI211_X1 U22669 ( .C1(n19931), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P2_U3117) );
  AOI22_X1 U22670 ( .A1(n19934), .A2(n19665), .B1(n19932), .B2(n19664), .ZN(
        n19663) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19933), .ZN(n19662) );
  OAI211_X1 U22672 ( .C1(n19937), .C2(n19697), .A(n19663), .B(n19662), .ZN(
        P2_U3118) );
  AOI22_X1 U22673 ( .A1(n19942), .A2(n19665), .B1(n19938), .B2(n19664), .ZN(
        n19669) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19667), .B1(
        n19666), .B2(n19940), .ZN(n19668) );
  OAI211_X1 U22675 ( .C1(n19948), .C2(n19697), .A(n19669), .B(n19668), .ZN(
        P2_U3119) );
  NOR2_X1 U22676 ( .A1(n19671), .A2(n19744), .ZN(n19698) );
  AOI22_X1 U22677 ( .A1(n19820), .A2(n19699), .B1(n19886), .B2(n19698), .ZN(
        n19682) );
  OR2_X1 U22678 ( .A1(n19672), .A2(n19770), .ZN(n19892) );
  OAI21_X1 U22679 ( .B1(n19892), .B2(n19673), .A(n20029), .ZN(n19680) );
  INV_X1 U22680 ( .A(n19679), .ZN(n19677) );
  INV_X1 U22681 ( .A(n10943), .ZN(n19675) );
  INV_X1 U22682 ( .A(n19698), .ZN(n19674) );
  OAI211_X1 U22683 ( .C1(n19675), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19852), 
        .B(n19674), .ZN(n19676) );
  OAI211_X1 U22684 ( .C1(n19680), .C2(n19677), .A(n19889), .B(n19676), .ZN(
        n19701) );
  OAI21_X1 U22685 ( .B1(n10943), .B2(n19698), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19678) );
  OAI21_X1 U22686 ( .B1(n19680), .B2(n19679), .A(n19678), .ZN(n19700) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19701), .B1(
        n19887), .B2(n19700), .ZN(n19681) );
  OAI211_X1 U22688 ( .C1(n19749), .C2(n19736), .A(n19682), .B(n19681), .ZN(
        P2_U3120) );
  AOI22_X1 U22689 ( .A1(n19786), .A2(n19699), .B1(n19900), .B2(n19698), .ZN(
        n19684) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19701), .B1(
        n19901), .B2(n19700), .ZN(n19683) );
  OAI211_X1 U22691 ( .C1(n19789), .C2(n19736), .A(n19684), .B(n19683), .ZN(
        P2_U3121) );
  AOI22_X1 U22692 ( .A1(n19685), .A2(n19699), .B1(n19906), .B2(n19698), .ZN(
        n19687) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19701), .B1(
        n19907), .B2(n19700), .ZN(n19686) );
  OAI211_X1 U22694 ( .C1(n19688), .C2(n19736), .A(n19687), .B(n19686), .ZN(
        P2_U3122) );
  AOI22_X1 U22695 ( .A1(n19914), .A2(n19699), .B1(n19912), .B2(n19698), .ZN(
        n19690) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19701), .B1(
        n19913), .B2(n19700), .ZN(n19689) );
  OAI211_X1 U22697 ( .C1(n19917), .C2(n19736), .A(n19690), .B(n19689), .ZN(
        P2_U3123) );
  AOI22_X1 U22698 ( .A1(n19867), .A2(n19699), .B1(n19918), .B2(n19698), .ZN(
        n19692) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19701), .B1(
        n19919), .B2(n19700), .ZN(n19691) );
  OAI211_X1 U22700 ( .C1(n19870), .C2(n19736), .A(n19692), .B(n19691), .ZN(
        P2_U3124) );
  INV_X1 U22701 ( .A(n19736), .ZN(n19722) );
  AOI22_X1 U22702 ( .A1(n19722), .A2(n19926), .B1(n19924), .B2(n19698), .ZN(
        n19694) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19701), .B1(
        n19925), .B2(n19700), .ZN(n19693) );
  OAI211_X1 U22704 ( .C1(n19931), .C2(n19697), .A(n19694), .B(n19693), .ZN(
        P2_U3125) );
  AOI22_X1 U22705 ( .A1(n19798), .A2(n19722), .B1(n19932), .B2(n19698), .ZN(
        n19696) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19701), .B1(
        n19933), .B2(n19700), .ZN(n19695) );
  OAI211_X1 U22707 ( .C1(n19802), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U3126) );
  AOI22_X1 U22708 ( .A1(n19699), .A2(n19942), .B1(n19938), .B2(n19698), .ZN(
        n19703) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19701), .B1(
        n19940), .B2(n19700), .ZN(n19702) );
  OAI211_X1 U22710 ( .C1(n19948), .C2(n19736), .A(n19703), .B(n19702), .ZN(
        P2_U3127) );
  INV_X1 U22711 ( .A(n20030), .ZN(n19704) );
  NOR2_X1 U22712 ( .A1(n19705), .A2(n19744), .ZN(n19731) );
  AOI22_X1 U22713 ( .A1(n19820), .A2(n19722), .B1(n19886), .B2(n19731), .ZN(
        n19717) );
  AOI21_X1 U22714 ( .B1(n19711), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19709) );
  AOI21_X1 U22715 ( .B1(n19760), .B2(n19736), .A(n19770), .ZN(n19706) );
  NOR2_X1 U22716 ( .A1(n19706), .A2(n19852), .ZN(n19710) );
  NAND2_X1 U22717 ( .A1(n19707), .A2(n19738), .ZN(n19714) );
  NAND2_X1 U22718 ( .A1(n19710), .A2(n19714), .ZN(n19708) );
  OAI211_X1 U22719 ( .C1(n19731), .C2(n19709), .A(n19708), .B(n19889), .ZN(
        n19733) );
  INV_X1 U22720 ( .A(n19710), .ZN(n19715) );
  INV_X1 U22721 ( .A(n19711), .ZN(n19712) );
  OAI21_X1 U22722 ( .B1(n19712), .B2(n19731), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19713) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19733), .B1(
        n19887), .B2(n19732), .ZN(n19716) );
  OAI211_X1 U22724 ( .C1(n19749), .C2(n19760), .A(n19717), .B(n19716), .ZN(
        P2_U3128) );
  AOI22_X1 U22725 ( .A1(n19786), .A2(n19722), .B1(n19900), .B2(n19731), .ZN(
        n19719) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19733), .B1(
        n19901), .B2(n19732), .ZN(n19718) );
  OAI211_X1 U22727 ( .C1(n19789), .C2(n19760), .A(n19719), .B(n19718), .ZN(
        P2_U3129) );
  AOI22_X1 U22728 ( .A1(n19765), .A2(n19908), .B1(n19906), .B2(n19731), .ZN(
        n19721) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19733), .B1(
        n19907), .B2(n19732), .ZN(n19720) );
  OAI211_X1 U22730 ( .C1(n19911), .C2(n19736), .A(n19721), .B(n19720), .ZN(
        P2_U3130) );
  AOI22_X1 U22731 ( .A1(n19914), .A2(n19722), .B1(n19912), .B2(n19731), .ZN(
        n19724) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19733), .B1(
        n19913), .B2(n19732), .ZN(n19723) );
  OAI211_X1 U22733 ( .C1(n19917), .C2(n19760), .A(n19724), .B(n19723), .ZN(
        P2_U3131) );
  AOI22_X1 U22734 ( .A1(n19920), .A2(n19765), .B1(n19918), .B2(n19731), .ZN(
        n19726) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19733), .B1(
        n19919), .B2(n19732), .ZN(n19725) );
  OAI211_X1 U22736 ( .C1(n19923), .C2(n19736), .A(n19726), .B(n19725), .ZN(
        P2_U3132) );
  AOI22_X1 U22737 ( .A1(n19765), .A2(n19926), .B1(n19924), .B2(n19731), .ZN(
        n19728) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19733), .B1(
        n19925), .B2(n19732), .ZN(n19727) );
  OAI211_X1 U22739 ( .C1(n19931), .C2(n19736), .A(n19728), .B(n19727), .ZN(
        P2_U3133) );
  AOI22_X1 U22740 ( .A1(n19798), .A2(n19765), .B1(n19932), .B2(n19731), .ZN(
        n19730) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19733), .B1(
        n19933), .B2(n19732), .ZN(n19729) );
  OAI211_X1 U22742 ( .C1(n19802), .C2(n19736), .A(n19730), .B(n19729), .ZN(
        P2_U3134) );
  AOI22_X1 U22743 ( .A1(n19840), .A2(n19765), .B1(n19938), .B2(n19731), .ZN(
        n19735) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19733), .B1(
        n19940), .B2(n19732), .ZN(n19734) );
  OAI211_X1 U22745 ( .C1(n19845), .C2(n19736), .A(n19735), .B(n19734), .ZN(
        P2_U3135) );
  NAND2_X1 U22746 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19738), .ZN(
        n19741) );
  NOR2_X1 U22747 ( .A1(n19739), .A2(n19744), .ZN(n19763) );
  OAI21_X1 U22748 ( .B1(n19742), .B2(n19763), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19740) );
  OAI21_X1 U22749 ( .B1(n19741), .B2(n19852), .A(n19740), .ZN(n19764) );
  AOI22_X1 U22750 ( .A1(n19764), .A2(n19887), .B1(n19886), .B2(n19763), .ZN(
        n19748) );
  INV_X1 U22751 ( .A(n19742), .ZN(n19743) );
  AOI21_X1 U22752 ( .B1(n19743), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19746) );
  OAI22_X1 U22753 ( .A1(n19892), .A2(n20030), .B1(n10880), .B2(n19744), .ZN(
        n19745) );
  OAI211_X1 U22754 ( .C1(n19763), .C2(n19746), .A(n19745), .B(n19889), .ZN(
        n19766) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19766), .B1(
        n19765), .B2(n19820), .ZN(n19747) );
  OAI211_X1 U22756 ( .C1(n19749), .C2(n19801), .A(n19748), .B(n19747), .ZN(
        P2_U3136) );
  AOI22_X1 U22757 ( .A1(n19764), .A2(n19901), .B1(n19900), .B2(n19763), .ZN(
        n19751) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19766), .B1(
        n19765), .B2(n19786), .ZN(n19750) );
  OAI211_X1 U22759 ( .C1(n19789), .C2(n19801), .A(n19751), .B(n19750), .ZN(
        P2_U3137) );
  AOI22_X1 U22760 ( .A1(n19764), .A2(n19907), .B1(n19906), .B2(n19763), .ZN(
        n19753) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19766), .B1(
        n19805), .B2(n19908), .ZN(n19752) );
  OAI211_X1 U22762 ( .C1(n19911), .C2(n19760), .A(n19753), .B(n19752), .ZN(
        P2_U3138) );
  AOI22_X1 U22763 ( .A1(n19764), .A2(n19913), .B1(n19912), .B2(n19763), .ZN(
        n19755) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19766), .B1(
        n19765), .B2(n19914), .ZN(n19754) );
  OAI211_X1 U22765 ( .C1(n19917), .C2(n19801), .A(n19755), .B(n19754), .ZN(
        P2_U3139) );
  AOI22_X1 U22766 ( .A1(n19764), .A2(n19919), .B1(n19918), .B2(n19763), .ZN(
        n19757) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19766), .B1(
        n19765), .B2(n19867), .ZN(n19756) );
  OAI211_X1 U22768 ( .C1(n19870), .C2(n19801), .A(n19757), .B(n19756), .ZN(
        P2_U3140) );
  AOI22_X1 U22769 ( .A1(n19764), .A2(n19925), .B1(n19924), .B2(n19763), .ZN(
        n19759) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19766), .B1(
        n19805), .B2(n19926), .ZN(n19758) );
  OAI211_X1 U22771 ( .C1(n19931), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P2_U3141) );
  AOI22_X1 U22772 ( .A1(n19764), .A2(n19933), .B1(n19932), .B2(n19763), .ZN(
        n19762) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19766), .B1(
        n19765), .B2(n19934), .ZN(n19761) );
  OAI211_X1 U22774 ( .C1(n19937), .C2(n19801), .A(n19762), .B(n19761), .ZN(
        P2_U3142) );
  AOI22_X1 U22775 ( .A1(n19764), .A2(n19940), .B1(n19938), .B2(n19763), .ZN(
        n19768) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19766), .B1(
        n19765), .B2(n19942), .ZN(n19767) );
  OAI211_X1 U22777 ( .C1(n19948), .C2(n19801), .A(n19768), .B(n19767), .ZN(
        P2_U3143) );
  AOI21_X1 U22778 ( .B1(n19801), .B2(n19844), .A(n19770), .ZN(n19771) );
  AOI21_X1 U22779 ( .B1(n19778), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19771), .ZN(n19776) );
  NAND2_X1 U22780 ( .A1(n10940), .A2(n20037), .ZN(n19773) );
  NAND3_X1 U22781 ( .A1(n10880), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19814) );
  NOR2_X1 U22782 ( .A1(n19814), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19803) );
  INV_X1 U22783 ( .A(n19803), .ZN(n19772) );
  NAND3_X1 U22784 ( .A1(n19773), .A2(n19772), .A3(n19852), .ZN(n19774) );
  NAND2_X1 U22785 ( .A1(n19774), .A2(n19889), .ZN(n19775) );
  INV_X1 U22786 ( .A(n19806), .ZN(n19785) );
  INV_X1 U22787 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n19784) );
  INV_X1 U22788 ( .A(n19777), .ZN(n19781) );
  INV_X1 U22789 ( .A(n19778), .ZN(n19780) );
  OAI21_X1 U22790 ( .B1(n10940), .B2(n19803), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19779) );
  OAI21_X1 U22791 ( .B1(n19781), .B2(n19780), .A(n19779), .ZN(n19804) );
  AOI22_X1 U22792 ( .A1(n19804), .A2(n19887), .B1(n19886), .B2(n19803), .ZN(
        n19783) );
  AOI22_X1 U22793 ( .A1(n19836), .A2(n19896), .B1(n19805), .B2(n19820), .ZN(
        n19782) );
  OAI211_X1 U22794 ( .C1(n19785), .C2(n19784), .A(n19783), .B(n19782), .ZN(
        P2_U3144) );
  AOI22_X1 U22795 ( .A1(n19804), .A2(n19901), .B1(n19900), .B2(n19803), .ZN(
        n19788) );
  AOI22_X1 U22796 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19806), .B1(
        n19805), .B2(n19786), .ZN(n19787) );
  OAI211_X1 U22797 ( .C1(n19789), .C2(n19844), .A(n19788), .B(n19787), .ZN(
        P2_U3145) );
  AOI22_X1 U22798 ( .A1(n19804), .A2(n19907), .B1(n19906), .B2(n19803), .ZN(
        n19791) );
  AOI22_X1 U22799 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19806), .B1(
        n19836), .B2(n19908), .ZN(n19790) );
  OAI211_X1 U22800 ( .C1(n19911), .C2(n19801), .A(n19791), .B(n19790), .ZN(
        P2_U3146) );
  AOI22_X1 U22801 ( .A1(n19804), .A2(n19913), .B1(n19912), .B2(n19803), .ZN(
        n19793) );
  AOI22_X1 U22802 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19806), .B1(
        n19805), .B2(n19914), .ZN(n19792) );
  OAI211_X1 U22803 ( .C1(n19917), .C2(n19844), .A(n19793), .B(n19792), .ZN(
        P2_U3147) );
  AOI22_X1 U22804 ( .A1(n19804), .A2(n19919), .B1(n19918), .B2(n19803), .ZN(
        n19795) );
  AOI22_X1 U22805 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19806), .B1(
        n19805), .B2(n19867), .ZN(n19794) );
  OAI211_X1 U22806 ( .C1(n19870), .C2(n19844), .A(n19795), .B(n19794), .ZN(
        P2_U3148) );
  AOI22_X1 U22807 ( .A1(n19804), .A2(n19925), .B1(n19924), .B2(n19803), .ZN(
        n19797) );
  AOI22_X1 U22808 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19806), .B1(
        n19836), .B2(n19926), .ZN(n19796) );
  OAI211_X1 U22809 ( .C1(n19931), .C2(n19801), .A(n19797), .B(n19796), .ZN(
        P2_U3149) );
  AOI22_X1 U22810 ( .A1(n19804), .A2(n19933), .B1(n19932), .B2(n19803), .ZN(
        n19800) );
  AOI22_X1 U22811 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19806), .B1(
        n19836), .B2(n19798), .ZN(n19799) );
  OAI211_X1 U22812 ( .C1(n19802), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P2_U3150) );
  AOI22_X1 U22813 ( .A1(n19804), .A2(n19940), .B1(n19938), .B2(n19803), .ZN(
        n19808) );
  AOI22_X1 U22814 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19806), .B1(
        n19805), .B2(n19942), .ZN(n19807) );
  OAI211_X1 U22815 ( .C1(n19948), .C2(n19844), .A(n19808), .B(n19807), .ZN(
        P2_U3151) );
  OAI21_X1 U22816 ( .B1(n19892), .B2(n19817), .A(n19814), .ZN(n19813) );
  NOR2_X1 U22817 ( .A1(n21022), .A2(n19814), .ZN(n19850) );
  INV_X1 U22818 ( .A(n19850), .ZN(n19809) );
  NAND2_X1 U22819 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19809), .ZN(n19810) );
  OR2_X1 U22820 ( .A1(n10942), .A2(n19810), .ZN(n19816) );
  OAI211_X1 U22821 ( .C1(n19850), .C2(n20037), .A(n19816), .B(n19889), .ZN(
        n19811) );
  INV_X1 U22822 ( .A(n19811), .ZN(n19812) );
  INV_X1 U22823 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19823) );
  OAI21_X1 U22824 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19814), .A(n12754), 
        .ZN(n19815) );
  AND2_X1 U22825 ( .A1(n19816), .A2(n19815), .ZN(n19839) );
  AOI22_X1 U22826 ( .A1(n19839), .A2(n19887), .B1(n19886), .B2(n19850), .ZN(
        n19822) );
  INV_X1 U22827 ( .A(n19817), .ZN(n19818) );
  AOI22_X1 U22828 ( .A1(n19877), .A2(n19896), .B1(n19836), .B2(n19820), .ZN(
        n19821) );
  OAI211_X1 U22829 ( .C1(n19835), .C2(n19823), .A(n19822), .B(n19821), .ZN(
        P2_U3152) );
  AOI22_X1 U22830 ( .A1(n19839), .A2(n19901), .B1(n19900), .B2(n19850), .ZN(
        n19825) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19841), .B1(
        n19877), .B2(n19902), .ZN(n19824) );
  OAI211_X1 U22832 ( .C1(n19905), .C2(n19844), .A(n19825), .B(n19824), .ZN(
        P2_U3153) );
  AOI22_X1 U22833 ( .A1(n19839), .A2(n19907), .B1(n19906), .B2(n19850), .ZN(
        n19827) );
  AOI22_X1 U22834 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19841), .B1(
        n19877), .B2(n19908), .ZN(n19826) );
  OAI211_X1 U22835 ( .C1(n19911), .C2(n19844), .A(n19827), .B(n19826), .ZN(
        P2_U3154) );
  AOI22_X1 U22836 ( .A1(n19839), .A2(n19913), .B1(n19912), .B2(n19850), .ZN(
        n19829) );
  AOI22_X1 U22837 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19841), .B1(
        n19836), .B2(n19914), .ZN(n19828) );
  OAI211_X1 U22838 ( .C1(n19917), .C2(n19873), .A(n19829), .B(n19828), .ZN(
        P2_U3155) );
  AOI22_X1 U22839 ( .A1(n19839), .A2(n19919), .B1(n19918), .B2(n19850), .ZN(
        n19831) );
  AOI22_X1 U22840 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19841), .B1(
        n19877), .B2(n19920), .ZN(n19830) );
  OAI211_X1 U22841 ( .C1(n19923), .C2(n19844), .A(n19831), .B(n19830), .ZN(
        P2_U3156) );
  AOI22_X1 U22842 ( .A1(n19839), .A2(n19925), .B1(n19924), .B2(n19850), .ZN(
        n19834) );
  AOI22_X1 U22843 ( .A1(n19877), .A2(n19926), .B1(n19836), .B2(n19832), .ZN(
        n19833) );
  OAI211_X1 U22844 ( .C1(n19835), .C2(n20860), .A(n19834), .B(n19833), .ZN(
        P2_U3157) );
  AOI22_X1 U22845 ( .A1(n19839), .A2(n19933), .B1(n19932), .B2(n19850), .ZN(
        n19838) );
  AOI22_X1 U22846 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19841), .B1(
        n19836), .B2(n19934), .ZN(n19837) );
  OAI211_X1 U22847 ( .C1(n19937), .C2(n19873), .A(n19838), .B(n19837), .ZN(
        P2_U3158) );
  AOI22_X1 U22848 ( .A1(n19839), .A2(n19940), .B1(n19938), .B2(n19850), .ZN(
        n19843) );
  AOI22_X1 U22849 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19841), .B1(
        n19877), .B2(n19840), .ZN(n19842) );
  OAI211_X1 U22850 ( .C1(n19845), .C2(n19844), .A(n19843), .B(n19842), .ZN(
        P2_U3159) );
  INV_X1 U22851 ( .A(n19883), .ZN(n19848) );
  NOR3_X2 U22852 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12315), .A3(
        n19848), .ZN(n19876) );
  AOI22_X1 U22853 ( .A1(n19943), .A2(n19896), .B1(n19886), .B2(n19876), .ZN(
        n19860) );
  OAI21_X1 U22854 ( .B1(n19943), .B2(n19877), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19849) );
  NAND2_X1 U22855 ( .A1(n19849), .A2(n20029), .ZN(n19858) );
  NOR2_X1 U22856 ( .A1(n19876), .A2(n19850), .ZN(n19857) );
  INV_X1 U22857 ( .A(n19857), .ZN(n19855) );
  INV_X1 U22858 ( .A(n10938), .ZN(n19853) );
  INV_X1 U22859 ( .A(n19876), .ZN(n19851) );
  OAI211_X1 U22860 ( .C1(n19853), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19852), 
        .B(n19851), .ZN(n19854) );
  OAI211_X1 U22861 ( .C1(n19858), .C2(n19855), .A(n19889), .B(n19854), .ZN(
        n19879) );
  OAI21_X1 U22862 ( .B1(n10938), .B2(n19876), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19856) );
  AOI22_X1 U22863 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19879), .B1(
        n19887), .B2(n19878), .ZN(n19859) );
  OAI211_X1 U22864 ( .C1(n19899), .C2(n19873), .A(n19860), .B(n19859), .ZN(
        P2_U3160) );
  AOI22_X1 U22865 ( .A1(n19902), .A2(n19943), .B1(n19900), .B2(n19876), .ZN(
        n19862) );
  AOI22_X1 U22866 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19879), .B1(
        n19901), .B2(n19878), .ZN(n19861) );
  OAI211_X1 U22867 ( .C1(n19905), .C2(n19873), .A(n19862), .B(n19861), .ZN(
        P2_U3161) );
  AOI22_X1 U22868 ( .A1(n19943), .A2(n19908), .B1(n19906), .B2(n19876), .ZN(
        n19864) );
  AOI22_X1 U22869 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19879), .B1(
        n19907), .B2(n19878), .ZN(n19863) );
  OAI211_X1 U22870 ( .C1(n19911), .C2(n19873), .A(n19864), .B(n19863), .ZN(
        P2_U3162) );
  AOI22_X1 U22871 ( .A1(n19914), .A2(n19877), .B1(n19912), .B2(n19876), .ZN(
        n19866) );
  AOI22_X1 U22872 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19879), .B1(
        n19913), .B2(n19878), .ZN(n19865) );
  OAI211_X1 U22873 ( .C1(n19917), .C2(n19930), .A(n19866), .B(n19865), .ZN(
        P2_U3163) );
  AOI22_X1 U22874 ( .A1(n19867), .A2(n19877), .B1(n19918), .B2(n19876), .ZN(
        n19869) );
  AOI22_X1 U22875 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19879), .B1(
        n19919), .B2(n19878), .ZN(n19868) );
  OAI211_X1 U22876 ( .C1(n19870), .C2(n19930), .A(n19869), .B(n19868), .ZN(
        P2_U3164) );
  AOI22_X1 U22877 ( .A1(n19943), .A2(n19926), .B1(n19924), .B2(n19876), .ZN(
        n19872) );
  AOI22_X1 U22878 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19879), .B1(
        n19925), .B2(n19878), .ZN(n19871) );
  OAI211_X1 U22879 ( .C1(n19931), .C2(n19873), .A(n19872), .B(n19871), .ZN(
        P2_U3165) );
  AOI22_X1 U22880 ( .A1(n19877), .A2(n19934), .B1(n19932), .B2(n19876), .ZN(
        n19875) );
  AOI22_X1 U22881 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19879), .B1(
        n19933), .B2(n19878), .ZN(n19874) );
  OAI211_X1 U22882 ( .C1(n19937), .C2(n19930), .A(n19875), .B(n19874), .ZN(
        P2_U3166) );
  AOI22_X1 U22883 ( .A1(n19877), .A2(n19942), .B1(n19938), .B2(n19876), .ZN(
        n19881) );
  AOI22_X1 U22884 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19879), .B1(
        n19940), .B2(n19878), .ZN(n19880) );
  OAI211_X1 U22885 ( .C1(n19948), .C2(n19930), .A(n19881), .B(n19880), .ZN(
        P2_U3167) );
  INV_X1 U22886 ( .A(n19882), .ZN(n19939) );
  NOR3_X1 U22887 ( .A1(n10944), .A2(n19939), .A3(n12754), .ZN(n19888) );
  NAND2_X1 U22888 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19883), .ZN(
        n19894) );
  INV_X1 U22889 ( .A(n19894), .ZN(n19884) );
  AOI21_X1 U22890 ( .B1(n20037), .B2(n19884), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19885) );
  NOR2_X1 U22891 ( .A1(n19888), .A2(n19885), .ZN(n19941) );
  AOI22_X1 U22892 ( .A1(n19941), .A2(n19887), .B1(n19939), .B2(n19886), .ZN(
        n19898) );
  INV_X1 U22893 ( .A(n19888), .ZN(n19890) );
  OAI211_X1 U22894 ( .C1(n19939), .C2(n20037), .A(n19890), .B(n19889), .ZN(
        n19891) );
  AOI221_X1 U22895 ( .B1(n19894), .B2(n19893), .C1(n19894), .C2(n19892), .A(
        n19891), .ZN(n19895) );
  AOI22_X1 U22896 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19944), .B1(
        n19927), .B2(n19896), .ZN(n19897) );
  OAI211_X1 U22897 ( .C1(n19899), .C2(n19930), .A(n19898), .B(n19897), .ZN(
        P2_U3168) );
  AOI22_X1 U22898 ( .A1(n19941), .A2(n19901), .B1(n19939), .B2(n19900), .ZN(
        n19904) );
  AOI22_X1 U22899 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19944), .B1(
        n19927), .B2(n19902), .ZN(n19903) );
  OAI211_X1 U22900 ( .C1(n19905), .C2(n19930), .A(n19904), .B(n19903), .ZN(
        P2_U3169) );
  AOI22_X1 U22901 ( .A1(n19941), .A2(n19907), .B1(n19939), .B2(n19906), .ZN(
        n19910) );
  AOI22_X1 U22902 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19944), .B1(
        n19927), .B2(n19908), .ZN(n19909) );
  OAI211_X1 U22903 ( .C1(n19911), .C2(n19930), .A(n19910), .B(n19909), .ZN(
        P2_U3170) );
  AOI22_X1 U22904 ( .A1(n19941), .A2(n19913), .B1(n19939), .B2(n19912), .ZN(
        n19916) );
  AOI22_X1 U22905 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19944), .B1(
        n19943), .B2(n19914), .ZN(n19915) );
  OAI211_X1 U22906 ( .C1(n19917), .C2(n19947), .A(n19916), .B(n19915), .ZN(
        P2_U3171) );
  AOI22_X1 U22907 ( .A1(n19941), .A2(n19919), .B1(n19939), .B2(n19918), .ZN(
        n19922) );
  AOI22_X1 U22908 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19944), .B1(
        n19927), .B2(n19920), .ZN(n19921) );
  OAI211_X1 U22909 ( .C1(n19923), .C2(n19930), .A(n19922), .B(n19921), .ZN(
        P2_U3172) );
  AOI22_X1 U22910 ( .A1(n19941), .A2(n19925), .B1(n19939), .B2(n19924), .ZN(
        n19929) );
  AOI22_X1 U22911 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19944), .B1(
        n19927), .B2(n19926), .ZN(n19928) );
  OAI211_X1 U22912 ( .C1(n19931), .C2(n19930), .A(n19929), .B(n19928), .ZN(
        P2_U3173) );
  AOI22_X1 U22913 ( .A1(n19941), .A2(n19933), .B1(n19939), .B2(n19932), .ZN(
        n19936) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19944), .B1(
        n19943), .B2(n19934), .ZN(n19935) );
  OAI211_X1 U22915 ( .C1(n19937), .C2(n19947), .A(n19936), .B(n19935), .ZN(
        P2_U3174) );
  AOI22_X1 U22916 ( .A1(n19941), .A2(n19940), .B1(n19939), .B2(n19938), .ZN(
        n19946) );
  AOI22_X1 U22917 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19944), .B1(
        n19943), .B2(n19942), .ZN(n19945) );
  OAI211_X1 U22918 ( .C1(n19948), .C2(n19947), .A(n19946), .B(n19945), .ZN(
        P2_U3175) );
  INV_X1 U22919 ( .A(n19949), .ZN(n19951) );
  OAI221_X1 U22920 ( .B1(n20073), .B2(n19951), .C1(n20073), .C2(n20756), .A(
        n19950), .ZN(n19956) );
  OAI211_X1 U22921 ( .C1(n19953), .C2(n19957), .A(n19952), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19954) );
  OAI211_X1 U22922 ( .C1(n19957), .C2(n19956), .A(n19955), .B(n19954), .ZN(
        P2_U3177) );
  AND2_X1 U22923 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19958), .ZN(
        P2_U3179) );
  AND2_X1 U22924 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19958), .ZN(
        P2_U3180) );
  INV_X1 U22925 ( .A(n20027), .ZN(n19959) );
  AND2_X1 U22926 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19959), .ZN(
        P2_U3181) );
  AND2_X1 U22927 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19958), .ZN(
        P2_U3182) );
  AND2_X1 U22928 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19959), .ZN(
        P2_U3183) );
  AND2_X1 U22929 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19958), .ZN(
        P2_U3184) );
  AND2_X1 U22930 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19959), .ZN(
        P2_U3185) );
  AND2_X1 U22931 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19958), .ZN(
        P2_U3186) );
  AND2_X1 U22932 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19959), .ZN(
        P2_U3187) );
  AND2_X1 U22933 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19959), .ZN(
        P2_U3188) );
  AND2_X1 U22934 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19959), .ZN(
        P2_U3189) );
  AND2_X1 U22935 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19959), .ZN(
        P2_U3190) );
  AND2_X1 U22936 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19959), .ZN(
        P2_U3191) );
  AND2_X1 U22937 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19959), .ZN(
        P2_U3192) );
  AND2_X1 U22938 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19958), .ZN(
        P2_U3193) );
  AND2_X1 U22939 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19958), .ZN(
        P2_U3194) );
  AND2_X1 U22940 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19958), .ZN(
        P2_U3195) );
  AND2_X1 U22941 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19958), .ZN(
        P2_U3196) );
  AND2_X1 U22942 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19958), .ZN(
        P2_U3197) );
  AND2_X1 U22943 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19958), .ZN(
        P2_U3198) );
  AND2_X1 U22944 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19958), .ZN(
        P2_U3199) );
  AND2_X1 U22945 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19958), .ZN(
        P2_U3200) );
  AND2_X1 U22946 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19959), .ZN(P2_U3201) );
  AND2_X1 U22947 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19959), .ZN(P2_U3202) );
  AND2_X1 U22948 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19959), .ZN(P2_U3203) );
  AND2_X1 U22949 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19959), .ZN(P2_U3204) );
  AND2_X1 U22950 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19959), .ZN(P2_U3205) );
  AND2_X1 U22951 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19959), .ZN(P2_U3206) );
  AND2_X1 U22952 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19959), .ZN(P2_U3207) );
  AND2_X1 U22953 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19959), .ZN(P2_U3208) );
  NOR2_X1 U22954 ( .A1(n20756), .A2(n19960), .ZN(n20752) );
  INV_X1 U22955 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20904) );
  NOR3_X1 U22956 ( .A1(n20752), .A2(n20904), .A3(n19966), .ZN(n19963) );
  NOR2_X1 U22957 ( .A1(n20753), .A2(n20088), .ZN(n19961) );
  OAI21_X1 U22958 ( .B1(HOLD), .B2(n20904), .A(n19961), .ZN(n19962) );
  NAND2_X1 U22959 ( .A1(n19965), .A2(NA), .ZN(n20759) );
  OAI211_X1 U22960 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19963), .A(n19962), 
        .B(n20759), .ZN(P2_U3209) );
  INV_X1 U22961 ( .A(n19964), .ZN(n19969) );
  NOR2_X1 U22962 ( .A1(n19965), .A2(n20904), .ZN(n19967) );
  OAI21_X1 U22963 ( .B1(HOLD), .B2(n19966), .A(P2_STATE_REG_2__SCAN_IN), .ZN(
        n20755) );
  AOI211_X1 U22964 ( .C1(n19967), .C2(n20755), .A(n20082), .B(n20752), .ZN(
        n19968) );
  OAI21_X1 U22965 ( .B1(n20852), .B2(n19969), .A(n19968), .ZN(P2_U3210) );
  OAI222_X1 U22966 ( .A1(n20020), .A2(n19973), .B1(n19971), .B2(n20088), .C1(
        n19970), .C2(n20017), .ZN(P2_U3212) );
  OAI222_X1 U22967 ( .A1(n20017), .A2(n19973), .B1(n19972), .B2(n20088), .C1(
        n19975), .C2(n20020), .ZN(P2_U3213) );
  OAI222_X1 U22968 ( .A1(n20017), .A2(n19975), .B1(n19974), .B2(n20088), .C1(
        n19976), .C2(n20020), .ZN(P2_U3214) );
  OAI222_X1 U22969 ( .A1(n20020), .A2(n19978), .B1(n19977), .B2(n20088), .C1(
        n19976), .C2(n20017), .ZN(P2_U3215) );
  OAI222_X1 U22970 ( .A1(n20020), .A2(n19980), .B1(n19979), .B2(n20088), .C1(
        n19978), .C2(n20017), .ZN(P2_U3216) );
  OAI222_X1 U22971 ( .A1(n20020), .A2(n19982), .B1(n19981), .B2(n20088), .C1(
        n19980), .C2(n20017), .ZN(P2_U3217) );
  OAI222_X1 U22972 ( .A1(n20020), .A2(n19984), .B1(n19983), .B2(n20088), .C1(
        n19982), .C2(n20017), .ZN(P2_U3218) );
  OAI222_X1 U22973 ( .A1(n20020), .A2(n19985), .B1(n21021), .B2(n20088), .C1(
        n19984), .C2(n20017), .ZN(P2_U3219) );
  OAI222_X1 U22974 ( .A1(n20020), .A2(n20870), .B1(n19986), .B2(n20088), .C1(
        n19985), .C2(n20017), .ZN(P2_U3220) );
  INV_X1 U22975 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19988) );
  OAI222_X1 U22976 ( .A1(n20020), .A2(n19988), .B1(n19987), .B2(n20088), .C1(
        n20870), .C2(n20017), .ZN(P2_U3221) );
  INV_X1 U22977 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19990) );
  OAI222_X1 U22978 ( .A1(n20020), .A2(n19990), .B1(n19989), .B2(n20088), .C1(
        n19988), .C2(n20017), .ZN(P2_U3222) );
  OAI222_X1 U22979 ( .A1(n20020), .A2(n19992), .B1(n19991), .B2(n20088), .C1(
        n19990), .C2(n20017), .ZN(P2_U3223) );
  INV_X1 U22980 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19994) );
  OAI222_X1 U22981 ( .A1(n20020), .A2(n19994), .B1(n19993), .B2(n20088), .C1(
        n19992), .C2(n20017), .ZN(P2_U3224) );
  OAI222_X1 U22982 ( .A1(n20020), .A2(n19995), .B1(n20915), .B2(n20088), .C1(
        n19994), .C2(n20017), .ZN(P2_U3225) );
  OAI222_X1 U22983 ( .A1(n20020), .A2(n19997), .B1(n19996), .B2(n20088), .C1(
        n19995), .C2(n20017), .ZN(P2_U3226) );
  OAI222_X1 U22984 ( .A1(n20020), .A2(n19999), .B1(n19998), .B2(n20088), .C1(
        n19997), .C2(n20017), .ZN(P2_U3227) );
  INV_X1 U22985 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n21056) );
  OAI222_X1 U22986 ( .A1(n20020), .A2(n21056), .B1(n20825), .B2(n20088), .C1(
        n19999), .C2(n20017), .ZN(P2_U3228) );
  INV_X1 U22987 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20000) );
  OAI222_X1 U22988 ( .A1(n20020), .A2(n20000), .B1(n20907), .B2(n20088), .C1(
        n21056), .C2(n20017), .ZN(P2_U3229) );
  OAI222_X1 U22989 ( .A1(n20020), .A2(n20002), .B1(n20001), .B2(n20088), .C1(
        n20000), .C2(n20017), .ZN(P2_U3230) );
  OAI222_X1 U22990 ( .A1(n20020), .A2(n21000), .B1(n20003), .B2(n20088), .C1(
        n20002), .C2(n20017), .ZN(P2_U3231) );
  OAI222_X1 U22991 ( .A1(n20020), .A2(n20005), .B1(n20004), .B2(n20088), .C1(
        n21000), .C2(n20017), .ZN(P2_U3232) );
  OAI222_X1 U22992 ( .A1(n20020), .A2(n21070), .B1(n20006), .B2(n20088), .C1(
        n20005), .C2(n20017), .ZN(P2_U3233) );
  OAI222_X1 U22993 ( .A1(n20020), .A2(n11542), .B1(n20007), .B2(n20088), .C1(
        n21070), .C2(n20017), .ZN(P2_U3234) );
  OAI222_X1 U22994 ( .A1(n20020), .A2(n20009), .B1(n20008), .B2(n20088), .C1(
        n11542), .C2(n20017), .ZN(P2_U3235) );
  OAI222_X1 U22995 ( .A1(n20020), .A2(n20937), .B1(n20010), .B2(n20088), .C1(
        n20009), .C2(n20017), .ZN(P2_U3236) );
  INV_X1 U22996 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20013) );
  OAI222_X1 U22997 ( .A1(n20020), .A2(n20013), .B1(n20011), .B2(n20088), .C1(
        n20937), .C2(n20017), .ZN(P2_U3237) );
  OAI222_X1 U22998 ( .A1(n20017), .A2(n20013), .B1(n20012), .B2(n20088), .C1(
        n11551), .C2(n20020), .ZN(P2_U3238) );
  OAI222_X1 U22999 ( .A1(n20020), .A2(n20015), .B1(n20014), .B2(n20088), .C1(
        n11551), .C2(n20017), .ZN(P2_U3239) );
  INV_X1 U23000 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20018) );
  OAI222_X1 U23001 ( .A1(n20020), .A2(n20018), .B1(n20016), .B2(n20088), .C1(
        n20015), .C2(n20017), .ZN(P2_U3240) );
  OAI222_X1 U23002 ( .A1(n20020), .A2(n16276), .B1(n20019), .B2(n20088), .C1(
        n20018), .C2(n20017), .ZN(P2_U3241) );
  OAI22_X1 U23003 ( .A1(n20089), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20088), .ZN(n20021) );
  INV_X1 U23004 ( .A(n20021), .ZN(P2_U3585) );
  MUX2_X1 U23005 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20089), .Z(P2_U3586) );
  OAI22_X1 U23006 ( .A1(n20089), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20088), .ZN(n20022) );
  INV_X1 U23007 ( .A(n20022), .ZN(P2_U3587) );
  OAI22_X1 U23008 ( .A1(n20089), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20088), .ZN(n20023) );
  INV_X1 U23009 ( .A(n20023), .ZN(P2_U3588) );
  OAI21_X1 U23010 ( .B1(n20027), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20025), 
        .ZN(n20024) );
  INV_X1 U23011 ( .A(n20024), .ZN(P2_U3591) );
  OAI21_X1 U23012 ( .B1(n20027), .B2(n20026), .A(n20025), .ZN(P2_U3592) );
  INV_X1 U23013 ( .A(n20062), .ZN(n20064) );
  NAND2_X1 U23014 ( .A1(n20028), .A2(n20029), .ZN(n20036) );
  NAND2_X1 U23015 ( .A1(n20029), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20052) );
  OR2_X1 U23016 ( .A1(n20030), .A2(n20052), .ZN(n20041) );
  NAND3_X1 U23017 ( .A1(n20053), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20031), 
        .ZN(n20032) );
  NAND2_X1 U23018 ( .A1(n20032), .A2(n20048), .ZN(n20042) );
  NAND2_X1 U23019 ( .A1(n20041), .A2(n20042), .ZN(n20033) );
  NAND2_X1 U23020 ( .A1(n20034), .A2(n20033), .ZN(n20035) );
  OAI211_X1 U23021 ( .C1(n20038), .C2(n20037), .A(n20036), .B(n20035), .ZN(
        n20039) );
  INV_X1 U23022 ( .A(n20039), .ZN(n20040) );
  AOI22_X1 U23023 ( .A1(n20064), .A2(n12315), .B1(n20040), .B2(n20062), .ZN(
        P2_U3602) );
  OAI21_X1 U23024 ( .B1(n20043), .B2(n20042), .A(n20041), .ZN(n20044) );
  AOI21_X1 U23025 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20045), .A(n20044), 
        .ZN(n20046) );
  AOI22_X1 U23026 ( .A1(n20064), .A2(n20047), .B1(n20046), .B2(n20062), .ZN(
        P2_U3603) );
  INV_X1 U23027 ( .A(n20048), .ZN(n20058) );
  OR3_X1 U23028 ( .A1(n20050), .A2(n20058), .A3(n20049), .ZN(n20051) );
  OAI21_X1 U23029 ( .B1(n20053), .B2(n20052), .A(n20051), .ZN(n20054) );
  AOI21_X1 U23030 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20055), .A(n20054), 
        .ZN(n20056) );
  AOI22_X1 U23031 ( .A1(n20064), .A2(n10880), .B1(n20056), .B2(n20062), .ZN(
        P2_U3604) );
  OAI21_X1 U23032 ( .B1(n20059), .B2(n20058), .A(n20057), .ZN(n20060) );
  AOI21_X1 U23033 ( .B1(n20072), .B2(n20061), .A(n20060), .ZN(n20063) );
  AOI22_X1 U23034 ( .A1(n20064), .A2(n21022), .B1(n20063), .B2(n20062), .ZN(
        P2_U3605) );
  AOI22_X1 U23035 ( .A1(n20088), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20065), 
        .B2(n20089), .ZN(P2_U3608) );
  INV_X1 U23036 ( .A(n20066), .ZN(n20067) );
  OAI21_X1 U23037 ( .B1(n20069), .B2(n20068), .A(n20067), .ZN(n20071) );
  MUX2_X1 U23038 ( .A(P2_MORE_REG_SCAN_IN), .B(n20071), .S(n20070), .Z(
        P2_U3609) );
  NOR3_X1 U23039 ( .A1(n20073), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n20072), 
        .ZN(n20075) );
  AOI211_X1 U23040 ( .C1(n20756), .C2(n20076), .A(n20075), .B(n20074), .ZN(
        n20087) );
  NAND2_X1 U23041 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20756), .ZN(n20079) );
  NOR4_X1 U23042 ( .A1(n20082), .A2(n11377), .A3(n20077), .A4(n19309), .ZN(
        n20078) );
  AOI21_X1 U23043 ( .B1(n20080), .B2(n20079), .A(n20078), .ZN(n20086) );
  AND2_X1 U23044 ( .A1(n20081), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20084) );
  NAND2_X1 U23045 ( .A1(n20082), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20083) );
  AOI21_X1 U23046 ( .B1(n20084), .B2(n20083), .A(n20087), .ZN(n20085) );
  AOI22_X1 U23047 ( .A1(n20904), .A2(n20087), .B1(n20086), .B2(n20085), .ZN(
        P2_U3610) );
  OAI22_X1 U23048 ( .A1(n20089), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20088), .ZN(n20090) );
  INV_X1 U23049 ( .A(n20090), .ZN(P2_U3611) );
  OAI21_X1 U23050 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20091), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20672) );
  NAND2_X1 U23051 ( .A1(n12089), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20736) );
  OAI21_X1 U23052 ( .B1(n20672), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20751), .ZN(
        n20092) );
  INV_X1 U23053 ( .A(n20092), .ZN(P1_U2802) );
  INV_X1 U23054 ( .A(n20093), .ZN(n20095) );
  OAI21_X1 U23055 ( .B1(n20095), .B2(n20094), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20096) );
  OAI21_X1 U23056 ( .B1(n20097), .B2(n11886), .A(n20096), .ZN(P1_U2803) );
  NAND2_X1 U23057 ( .A1(n20680), .A2(n12089), .ZN(n20669) );
  INV_X1 U23058 ( .A(n20669), .ZN(n20099) );
  OAI21_X1 U23059 ( .B1(n20099), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20751), .ZN(
        n20098) );
  OAI21_X1 U23060 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20751), .A(n20098), 
        .ZN(P1_U2804) );
  NAND2_X1 U23061 ( .A1(n20672), .A2(n20751), .ZN(n20664) );
  INV_X1 U23062 ( .A(n20664), .ZN(n20728) );
  OAI21_X1 U23063 ( .B1(BS16), .B2(n20099), .A(n20728), .ZN(n20726) );
  OAI21_X1 U23064 ( .B1(n20728), .B2(n20453), .A(n20726), .ZN(P1_U2805) );
  OAI21_X1 U23065 ( .B1(n20102), .B2(n20101), .A(n20100), .ZN(P1_U2806) );
  NOR4_X1 U23066 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20106) );
  NOR4_X1 U23067 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20105) );
  NOR4_X1 U23068 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20104) );
  NOR4_X1 U23069 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20103) );
  NAND4_X1 U23070 ( .A1(n20106), .A2(n20105), .A3(n20104), .A4(n20103), .ZN(
        n20112) );
  NOR4_X1 U23071 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20110) );
  AOI211_X1 U23072 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20109) );
  NOR4_X1 U23073 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20108) );
  NOR4_X1 U23074 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20107) );
  NAND4_X1 U23075 ( .A1(n20110), .A2(n20109), .A3(n20108), .A4(n20107), .ZN(
        n20111) );
  NOR2_X1 U23076 ( .A1(n20112), .A2(n20111), .ZN(n20735) );
  INV_X1 U23077 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20114) );
  NOR3_X1 U23078 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20115) );
  OAI21_X1 U23079 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20115), .A(n20735), .ZN(
        n20113) );
  OAI21_X1 U23080 ( .B1(n20735), .B2(n20114), .A(n20113), .ZN(P1_U2807) );
  INV_X1 U23081 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20727) );
  AOI21_X1 U23082 ( .B1(n20116), .B2(n20727), .A(n20115), .ZN(n20118) );
  INV_X1 U23083 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20117) );
  INV_X1 U23084 ( .A(n20735), .ZN(n20732) );
  AOI22_X1 U23085 ( .A1(n20735), .A2(n20118), .B1(n20117), .B2(n20732), .ZN(
        P1_U2808) );
  INV_X1 U23086 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20130) );
  NOR2_X1 U23087 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20119), .ZN(n20124) );
  INV_X1 U23088 ( .A(n20188), .ZN(n20120) );
  AOI22_X1 U23089 ( .A1(n20120), .A2(n20159), .B1(n20170), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n20121) );
  OAI211_X1 U23090 ( .C1(n20162), .C2(n20122), .A(n20121), .B(n9736), .ZN(
        n20123) );
  AOI21_X1 U23091 ( .B1(n20124), .B2(n20133), .A(n20123), .ZN(n20129) );
  INV_X1 U23092 ( .A(n20189), .ZN(n20127) );
  AOI22_X1 U23093 ( .A1(n20127), .A2(n20154), .B1(n20126), .B2(n20125), .ZN(
        n20128) );
  OAI211_X1 U23094 ( .C1(n20131), .C2(n20130), .A(n20129), .B(n20128), .ZN(
        P1_U2831) );
  INV_X1 U23095 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20132) );
  AOI22_X1 U23096 ( .A1(n20159), .A2(n20134), .B1(n20133), .B2(n20132), .ZN(
        n20144) );
  INV_X1 U23097 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20138) );
  INV_X1 U23098 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20135) );
  OR2_X1 U23099 ( .A1(n20136), .A2(n20135), .ZN(n20137) );
  OAI211_X1 U23100 ( .C1(n20138), .C2(n20162), .A(n20137), .B(n9736), .ZN(
        n20139) );
  AOI21_X1 U23101 ( .B1(n20150), .B2(P1_REIP_REG_7__SCAN_IN), .A(n20139), .ZN(
        n20140) );
  OAI21_X1 U23102 ( .B1(n20195), .B2(n20141), .A(n20140), .ZN(n20142) );
  INV_X1 U23103 ( .A(n20142), .ZN(n20143) );
  OAI211_X1 U23104 ( .C1(n20145), .C2(n20186), .A(n20144), .B(n20143), .ZN(
        P1_U2833) );
  AOI22_X1 U23105 ( .A1(n20146), .A2(n20159), .B1(n20170), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20147) );
  OAI211_X1 U23106 ( .C1(n20162), .C2(n20148), .A(n20147), .B(n9736), .ZN(
        n20149) );
  AOI21_X1 U23107 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20150), .A(n20149), .ZN(
        n20157) );
  NAND3_X1 U23108 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n20151) );
  OR2_X1 U23109 ( .A1(n20152), .A2(n20151), .ZN(n20179) );
  NOR2_X1 U23110 ( .A1(n20179), .A2(n20683), .ZN(n20165) );
  INV_X1 U23111 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20164) );
  NOR2_X1 U23112 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20164), .ZN(n20153) );
  AOI22_X1 U23113 ( .A1(n20155), .A2(n20154), .B1(n20165), .B2(n20153), .ZN(
        n20156) );
  OAI211_X1 U23114 ( .C1(n20158), .C2(n20186), .A(n20157), .B(n20156), .ZN(
        P1_U2834) );
  AOI22_X1 U23115 ( .A1(n20159), .A2(n20198), .B1(n20170), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20160) );
  OAI211_X1 U23116 ( .C1(n20162), .C2(n20161), .A(n20160), .B(n9736), .ZN(
        n20163) );
  AOI221_X1 U23117 ( .B1(n20181), .B2(P1_REIP_REG_5__SCAN_IN), .C1(n20165), 
        .C2(n20164), .A(n20163), .ZN(n20167) );
  NAND2_X1 U23118 ( .A1(n20201), .A2(n20182), .ZN(n20166) );
  OAI211_X1 U23119 ( .C1(n20186), .C2(n20168), .A(n20167), .B(n20166), .ZN(
        P1_U2835) );
  INV_X1 U23120 ( .A(n20169), .ZN(n20171) );
  AOI22_X1 U23121 ( .A1(n20172), .A2(n20171), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n20170), .ZN(n20173) );
  OAI21_X1 U23122 ( .B1(n20175), .B2(n20174), .A(n20173), .ZN(n20176) );
  AOI211_X1 U23123 ( .C1(n20178), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20177), .B(n20176), .ZN(n20185) );
  NAND2_X1 U23124 ( .A1(n20179), .A2(n20683), .ZN(n20180) );
  AOI22_X1 U23125 ( .A1(n20183), .A2(n20182), .B1(n20181), .B2(n20180), .ZN(
        n20184) );
  OAI211_X1 U23126 ( .C1(n20187), .C2(n20186), .A(n20185), .B(n20184), .ZN(
        P1_U2836) );
  INV_X1 U23127 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20192) );
  OAI22_X1 U23128 ( .A1(n20189), .A2(n14624), .B1(n20194), .B2(n20188), .ZN(
        n20190) );
  INV_X1 U23129 ( .A(n20190), .ZN(n20191) );
  OAI21_X1 U23130 ( .B1(n20204), .B2(n20192), .A(n20191), .ZN(P1_U2863) );
  OAI22_X1 U23131 ( .A1(n20195), .A2(n14624), .B1(n20194), .B2(n20193), .ZN(
        n20196) );
  INV_X1 U23132 ( .A(n20196), .ZN(n20197) );
  OAI21_X1 U23133 ( .B1(n20204), .B2(n20135), .A(n20197), .ZN(P1_U2865) );
  INV_X1 U23134 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20203) );
  AOI22_X1 U23135 ( .A1(n20201), .A2(n20200), .B1(n20199), .B2(n20198), .ZN(
        n20202) );
  OAI21_X1 U23136 ( .B1(n20204), .B2(n20203), .A(n20202), .ZN(P1_U2867) );
  AOI22_X1 U23137 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20206) );
  OAI21_X1 U23138 ( .B1(n12978), .B2(n20229), .A(n20206), .ZN(P1_U2921) );
  INV_X1 U23139 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20208) );
  AOI22_X1 U23140 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20207) );
  OAI21_X1 U23141 ( .B1(n20208), .B2(n20229), .A(n20207), .ZN(P1_U2922) );
  INV_X1 U23142 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20210) );
  AOI22_X1 U23143 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20209) );
  OAI21_X1 U23144 ( .B1(n20210), .B2(n20229), .A(n20209), .ZN(P1_U2923) );
  AOI22_X1 U23145 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20211) );
  OAI21_X1 U23146 ( .B1(n13952), .B2(n20229), .A(n20211), .ZN(P1_U2924) );
  AOI22_X1 U23147 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20212) );
  OAI21_X1 U23148 ( .B1(n13986), .B2(n20229), .A(n20212), .ZN(P1_U2925) );
  INV_X1 U23149 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20214) );
  AOI22_X1 U23150 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20213) );
  OAI21_X1 U23151 ( .B1(n20214), .B2(n20229), .A(n20213), .ZN(P1_U2926) );
  INV_X1 U23152 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20216) );
  AOI22_X1 U23153 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20215) );
  OAI21_X1 U23154 ( .B1(n20216), .B2(n20229), .A(n20215), .ZN(P1_U2927) );
  INV_X1 U23155 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20218) );
  AOI22_X1 U23156 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20748), .B1(n20226), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20217) );
  OAI21_X1 U23157 ( .B1(n20218), .B2(n20229), .A(n20217), .ZN(P1_U2928) );
  AOI22_X1 U23158 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20219) );
  OAI21_X1 U23159 ( .B1(n13525), .B2(n20229), .A(n20219), .ZN(P1_U2929) );
  AOI22_X1 U23160 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20220) );
  OAI21_X1 U23161 ( .B1(n13511), .B2(n20229), .A(n20220), .ZN(P1_U2930) );
  AOI22_X1 U23162 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20221) );
  OAI21_X1 U23163 ( .B1(n13258), .B2(n20229), .A(n20221), .ZN(P1_U2931) );
  AOI22_X1 U23164 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20222) );
  OAI21_X1 U23165 ( .B1(n13101), .B2(n20229), .A(n20222), .ZN(P1_U2932) );
  AOI22_X1 U23166 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20223) );
  OAI21_X1 U23167 ( .B1(n13085), .B2(n20229), .A(n20223), .ZN(P1_U2933) );
  AOI22_X1 U23168 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20224) );
  OAI21_X1 U23169 ( .B1(n13024), .B2(n20229), .A(n20224), .ZN(P1_U2934) );
  AOI22_X1 U23170 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20225) );
  OAI21_X1 U23171 ( .B1(n12913), .B2(n20229), .A(n20225), .ZN(P1_U2935) );
  AOI22_X1 U23172 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20227), .B1(n20226), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20228) );
  OAI21_X1 U23173 ( .B1(n20230), .B2(n20229), .A(n20228), .ZN(P1_U2936) );
  AOI22_X1 U23174 ( .A1(n20254), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20259), .ZN(n20232) );
  NAND2_X1 U23175 ( .A1(n20244), .A2(n20231), .ZN(n20246) );
  NAND2_X1 U23176 ( .A1(n20232), .A2(n20246), .ZN(P1_U2945) );
  AOI22_X1 U23177 ( .A1(n20254), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20234) );
  NAND2_X1 U23178 ( .A1(n20244), .A2(n20233), .ZN(n20248) );
  NAND2_X1 U23179 ( .A1(n20234), .A2(n20248), .ZN(P1_U2946) );
  AOI22_X1 U23180 ( .A1(n20254), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20236) );
  NAND2_X1 U23181 ( .A1(n20244), .A2(n20235), .ZN(n20250) );
  NAND2_X1 U23182 ( .A1(n20236), .A2(n20250), .ZN(P1_U2947) );
  AOI22_X1 U23183 ( .A1(n20254), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20238) );
  NAND2_X1 U23184 ( .A1(n20244), .A2(n20237), .ZN(n20252) );
  NAND2_X1 U23185 ( .A1(n20238), .A2(n20252), .ZN(P1_U2948) );
  AOI22_X1 U23186 ( .A1(n20254), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20240) );
  NAND2_X1 U23187 ( .A1(n20244), .A2(n20239), .ZN(n20255) );
  NAND2_X1 U23188 ( .A1(n20240), .A2(n20255), .ZN(P1_U2949) );
  AOI22_X1 U23189 ( .A1(n20254), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20242) );
  NAND2_X1 U23190 ( .A1(n20244), .A2(n20241), .ZN(n20257) );
  NAND2_X1 U23191 ( .A1(n20242), .A2(n20257), .ZN(P1_U2950) );
  AOI22_X1 U23192 ( .A1(n20254), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20259), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20245) );
  NAND2_X1 U23193 ( .A1(n20244), .A2(n20243), .ZN(n20260) );
  NAND2_X1 U23194 ( .A1(n20245), .A2(n20260), .ZN(P1_U2951) );
  AOI22_X1 U23195 ( .A1(n20254), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20247) );
  NAND2_X1 U23196 ( .A1(n20247), .A2(n20246), .ZN(P1_U2960) );
  AOI22_X1 U23197 ( .A1(n20254), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20259), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20249) );
  NAND2_X1 U23198 ( .A1(n20249), .A2(n20248), .ZN(P1_U2961) );
  AOI22_X1 U23199 ( .A1(n20254), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20259), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20251) );
  NAND2_X1 U23200 ( .A1(n20251), .A2(n20250), .ZN(P1_U2962) );
  AOI22_X1 U23201 ( .A1(n20254), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20259), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20253) );
  NAND2_X1 U23202 ( .A1(n20253), .A2(n20252), .ZN(P1_U2963) );
  AOI22_X1 U23203 ( .A1(n20254), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20259), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20256) );
  NAND2_X1 U23204 ( .A1(n20256), .A2(n20255), .ZN(P1_U2964) );
  AOI22_X1 U23205 ( .A1(n20254), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20259), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20258) );
  NAND2_X1 U23206 ( .A1(n20258), .A2(n20257), .ZN(P1_U2965) );
  AOI22_X1 U23207 ( .A1(n20254), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20259), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20261) );
  NAND2_X1 U23208 ( .A1(n20261), .A2(n20260), .ZN(P1_U2966) );
  NOR2_X1 U23209 ( .A1(n20263), .A2(n20262), .ZN(P1_U3032) );
  OR2_X1 U23210 ( .A1(n20265), .A2(n20264), .ZN(n20391) );
  INV_X1 U23211 ( .A(n9769), .ZN(n20267) );
  OAI21_X1 U23212 ( .B1(n20316), .B2(n20295), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20269) );
  NAND2_X1 U23213 ( .A1(n20269), .A2(n20548), .ZN(n20277) );
  OR2_X1 U23214 ( .A1(n20271), .A2(n20270), .ZN(n20361) );
  OR2_X1 U23215 ( .A1(n20361), .A2(n11887), .ZN(n20276) );
  INV_X1 U23216 ( .A(n20276), .ZN(n20274) );
  NAND2_X1 U23217 ( .A1(n20273), .A2(n20272), .ZN(n20359) );
  NOR2_X1 U23218 ( .A1(n20545), .A2(n20359), .ZN(n20296) );
  OAI22_X1 U23219 ( .A1(n20277), .A2(n20274), .B1(n20554), .B2(n20296), .ZN(
        n20275) );
  AOI211_X1 U23220 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20391), .A(n20329), 
        .B(n20275), .ZN(n20292) );
  AOI22_X1 U23221 ( .A1(n20603), .A2(n20296), .B1(n20295), .B2(n20610), .ZN(
        n20279) );
  OAI22_X1 U23222 ( .A1(n20277), .A2(n20276), .B1(n20485), .B2(n20391), .ZN(
        n20297) );
  AOI22_X1 U23223 ( .A1(n20604), .A2(n20297), .B1(n20316), .B2(n20546), .ZN(
        n20278) );
  OAI211_X1 U23224 ( .C1(n20292), .C2(n21006), .A(n20279), .B(n20278), .ZN(
        P1_U3033) );
  AOI22_X1 U23225 ( .A1(n20614), .A2(n20296), .B1(n20295), .B2(n20616), .ZN(
        n20281) );
  AOI22_X1 U23226 ( .A1(n20615), .A2(n20297), .B1(n20316), .B2(n20563), .ZN(
        n20280) );
  OAI211_X1 U23227 ( .C1(n20292), .C2(n20282), .A(n20281), .B(n20280), .ZN(
        P1_U3034) );
  AOI22_X1 U23228 ( .A1(n20620), .A2(n20296), .B1(n20295), .B2(n20622), .ZN(
        n20284) );
  INV_X1 U23229 ( .A(n20292), .ZN(n20298) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20298), .B1(
        n20621), .B2(n20297), .ZN(n20283) );
  OAI211_X1 U23231 ( .C1(n20625), .C2(n20326), .A(n20284), .B(n20283), .ZN(
        P1_U3035) );
  AOI22_X1 U23232 ( .A1(n20626), .A2(n20296), .B1(n20295), .B2(n20628), .ZN(
        n20286) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20298), .B1(
        n20627), .B2(n20297), .ZN(n20285) );
  OAI211_X1 U23234 ( .C1(n20631), .C2(n20326), .A(n20286), .B(n20285), .ZN(
        P1_U3036) );
  AOI22_X1 U23235 ( .A1(n20632), .A2(n20296), .B1(n20295), .B2(n20634), .ZN(
        n20288) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20298), .B1(
        n20633), .B2(n20297), .ZN(n20287) );
  OAI211_X1 U23237 ( .C1(n20637), .C2(n20326), .A(n20288), .B(n20287), .ZN(
        P1_U3037) );
  INV_X1 U23238 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20291) );
  AOI22_X1 U23239 ( .A1(n20638), .A2(n20296), .B1(n20295), .B2(n20640), .ZN(
        n20290) );
  AOI22_X1 U23240 ( .A1(n20639), .A2(n20297), .B1(n20316), .B2(n20579), .ZN(
        n20289) );
  OAI211_X1 U23241 ( .C1(n20292), .C2(n20291), .A(n20290), .B(n20289), .ZN(
        P1_U3038) );
  AOI22_X1 U23242 ( .A1(n20644), .A2(n20296), .B1(n20295), .B2(n20646), .ZN(
        n20294) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20298), .B1(
        n20645), .B2(n20297), .ZN(n20293) );
  OAI211_X1 U23244 ( .C1(n20649), .C2(n20326), .A(n20294), .B(n20293), .ZN(
        P1_U3039) );
  AOI22_X1 U23245 ( .A1(n20651), .A2(n20296), .B1(n20295), .B2(n20654), .ZN(
        n20300) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20298), .B1(
        n20653), .B2(n20297), .ZN(n20299) );
  OAI211_X1 U23247 ( .C1(n20660), .C2(n20326), .A(n20300), .B(n20299), .ZN(
        P1_U3040) );
  INV_X1 U23248 ( .A(n20361), .ZN(n20301) );
  NOR2_X1 U23249 ( .A1(n20359), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20305) );
  INV_X1 U23250 ( .A(n20305), .ZN(n20302) );
  NOR2_X1 U23251 ( .A1(n20449), .A2(n20302), .ZN(n20321) );
  AOI21_X1 U23252 ( .B1(n20301), .B2(n20450), .A(n20321), .ZN(n20303) );
  OAI22_X1 U23253 ( .A1(n20303), .A2(n20601), .B1(n20302), .B2(n12842), .ZN(
        n20322) );
  AOI22_X1 U23254 ( .A1(n20604), .A2(n20322), .B1(n20603), .B2(n20321), .ZN(
        n20307) );
  OAI211_X1 U23255 ( .C1(n20360), .C2(n20453), .A(n20518), .B(n20303), .ZN(
        n20304) );
  OAI211_X1 U23256 ( .C1(n20548), .C2(n20305), .A(n20607), .B(n20304), .ZN(
        n20323) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20323), .B1(
        n20316), .B2(n20610), .ZN(n20306) );
  OAI211_X1 U23258 ( .C1(n20613), .C2(n20358), .A(n20307), .B(n20306), .ZN(
        P1_U3041) );
  AOI22_X1 U23259 ( .A1(n20615), .A2(n20322), .B1(n20614), .B2(n20321), .ZN(
        n20309) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20323), .B1(
        n20350), .B2(n20563), .ZN(n20308) );
  OAI211_X1 U23261 ( .C1(n20566), .C2(n20326), .A(n20309), .B(n20308), .ZN(
        P1_U3042) );
  AOI22_X1 U23262 ( .A1(n20621), .A2(n20322), .B1(n20620), .B2(n20321), .ZN(
        n20311) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20323), .B1(
        n20350), .B2(n20567), .ZN(n20310) );
  OAI211_X1 U23264 ( .C1(n20570), .C2(n20326), .A(n20311), .B(n20310), .ZN(
        P1_U3043) );
  AOI22_X1 U23265 ( .A1(n20627), .A2(n20322), .B1(n20626), .B2(n20321), .ZN(
        n20313) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20323), .B1(
        n20350), .B2(n20571), .ZN(n20312) );
  OAI211_X1 U23267 ( .C1(n20574), .C2(n20326), .A(n20313), .B(n20312), .ZN(
        P1_U3044) );
  AOI22_X1 U23268 ( .A1(n20633), .A2(n20322), .B1(n20632), .B2(n20321), .ZN(
        n20315) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20323), .B1(
        n20350), .B2(n20575), .ZN(n20314) );
  OAI211_X1 U23270 ( .C1(n20578), .C2(n20326), .A(n20315), .B(n20314), .ZN(
        P1_U3045) );
  AOI22_X1 U23271 ( .A1(n20639), .A2(n20322), .B1(n20638), .B2(n20321), .ZN(
        n20318) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20323), .B1(
        n20316), .B2(n20640), .ZN(n20317) );
  OAI211_X1 U23273 ( .C1(n20643), .C2(n20358), .A(n20318), .B(n20317), .ZN(
        P1_U3046) );
  AOI22_X1 U23274 ( .A1(n20645), .A2(n20322), .B1(n20644), .B2(n20321), .ZN(
        n20320) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20323), .B1(
        n20350), .B2(n20583), .ZN(n20319) );
  OAI211_X1 U23276 ( .C1(n20586), .C2(n20326), .A(n20320), .B(n20319), .ZN(
        P1_U3047) );
  AOI22_X1 U23277 ( .A1(n20653), .A2(n20322), .B1(n20651), .B2(n20321), .ZN(
        n20325) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20323), .B1(
        n20350), .B2(n20587), .ZN(n20324) );
  OAI211_X1 U23279 ( .C1(n20594), .C2(n20326), .A(n20325), .B(n20324), .ZN(
        P1_U3048) );
  INV_X1 U23280 ( .A(n20359), .ZN(n20327) );
  NAND2_X1 U23281 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20327), .ZN(
        n20367) );
  NOR2_X1 U23282 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20367), .ZN(
        n20353) );
  AOI22_X1 U23283 ( .A1(n20603), .A2(n20353), .B1(n20380), .B2(n20546), .ZN(
        n20339) );
  NOR2_X1 U23284 ( .A1(n20361), .A2(n20551), .ZN(n20333) );
  OAI21_X1 U23285 ( .B1(n20380), .B2(n20350), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20328) );
  NAND2_X1 U23286 ( .A1(n20328), .A2(n20548), .ZN(n20337) );
  INV_X1 U23287 ( .A(n20353), .ZN(n20331) );
  AOI211_X1 U23288 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20331), .A(n20330), 
        .B(n20329), .ZN(n20332) );
  INV_X1 U23289 ( .A(n20333), .ZN(n20336) );
  INV_X1 U23290 ( .A(n20334), .ZN(n20335) );
  OAI22_X1 U23291 ( .A1(n20337), .A2(n20336), .B1(n20335), .B2(n20485), .ZN(
        n20354) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20355), .B1(
        n20604), .B2(n20354), .ZN(n20338) );
  OAI211_X1 U23293 ( .C1(n20562), .C2(n20358), .A(n20339), .B(n20338), .ZN(
        P1_U3049) );
  AOI22_X1 U23294 ( .A1(n20614), .A2(n20353), .B1(n20380), .B2(n20563), .ZN(
        n20341) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20355), .B1(
        n20615), .B2(n20354), .ZN(n20340) );
  OAI211_X1 U23296 ( .C1(n20566), .C2(n20358), .A(n20341), .B(n20340), .ZN(
        P1_U3050) );
  AOI22_X1 U23297 ( .A1(n20620), .A2(n20353), .B1(n20350), .B2(n20622), .ZN(
        n20343) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20355), .B1(
        n20621), .B2(n20354), .ZN(n20342) );
  OAI211_X1 U23299 ( .C1(n20625), .C2(n20390), .A(n20343), .B(n20342), .ZN(
        P1_U3051) );
  AOI22_X1 U23300 ( .A1(n20626), .A2(n20353), .B1(n20350), .B2(n20628), .ZN(
        n20345) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20355), .B1(
        n20627), .B2(n20354), .ZN(n20344) );
  OAI211_X1 U23302 ( .C1(n20631), .C2(n20390), .A(n20345), .B(n20344), .ZN(
        P1_U3052) );
  AOI22_X1 U23303 ( .A1(n20632), .A2(n20353), .B1(n20350), .B2(n20634), .ZN(
        n20347) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20355), .B1(
        n20633), .B2(n20354), .ZN(n20346) );
  OAI211_X1 U23305 ( .C1(n20637), .C2(n20390), .A(n20347), .B(n20346), .ZN(
        P1_U3053) );
  AOI22_X1 U23306 ( .A1(n20638), .A2(n20353), .B1(n20380), .B2(n20579), .ZN(
        n20349) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20355), .B1(
        n20639), .B2(n20354), .ZN(n20348) );
  OAI211_X1 U23308 ( .C1(n20582), .C2(n20358), .A(n20349), .B(n20348), .ZN(
        P1_U3054) );
  AOI22_X1 U23309 ( .A1(n20644), .A2(n20353), .B1(n20350), .B2(n20646), .ZN(
        n20352) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20355), .B1(
        n20645), .B2(n20354), .ZN(n20351) );
  OAI211_X1 U23311 ( .C1(n20649), .C2(n20390), .A(n20352), .B(n20351), .ZN(
        P1_U3055) );
  AOI22_X1 U23312 ( .A1(n20651), .A2(n20353), .B1(n20380), .B2(n20587), .ZN(
        n20357) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20355), .B1(
        n20653), .B2(n20354), .ZN(n20356) );
  OAI211_X1 U23314 ( .C1(n20594), .C2(n20358), .A(n20357), .B(n20356), .ZN(
        P1_U3056) );
  NOR2_X1 U23315 ( .A1(n20595), .A2(n20359), .ZN(n20385) );
  AOI22_X1 U23316 ( .A1(n20603), .A2(n20385), .B1(n20410), .B2(n20546), .ZN(
        n20371) );
  OAI21_X1 U23317 ( .B1(n20360), .B2(n20519), .A(n20518), .ZN(n20368) );
  OR2_X1 U23318 ( .A1(n20361), .A2(n20513), .ZN(n20363) );
  INV_X1 U23319 ( .A(n20385), .ZN(n20362) );
  AND2_X1 U23320 ( .A1(n20363), .A2(n20362), .ZN(n20369) );
  INV_X1 U23321 ( .A(n20369), .ZN(n20366) );
  AOI21_X1 U23322 ( .B1(n20601), .B2(n20367), .A(n20364), .ZN(n20365) );
  OAI21_X1 U23323 ( .B1(n20368), .B2(n20366), .A(n20365), .ZN(n20387) );
  OAI22_X1 U23324 ( .A1(n20369), .A2(n20368), .B1(n12842), .B2(n20367), .ZN(
        n20386) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20387), .B1(
        n20604), .B2(n20386), .ZN(n20370) );
  OAI211_X1 U23326 ( .C1(n20562), .C2(n20390), .A(n20371), .B(n20370), .ZN(
        P1_U3057) );
  AOI22_X1 U23327 ( .A1(n20614), .A2(n20385), .B1(n20380), .B2(n20616), .ZN(
        n20373) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20387), .B1(
        n20615), .B2(n20386), .ZN(n20372) );
  OAI211_X1 U23329 ( .C1(n20619), .C2(n20418), .A(n20373), .B(n20372), .ZN(
        P1_U3058) );
  AOI22_X1 U23330 ( .A1(n20620), .A2(n20385), .B1(n20380), .B2(n20622), .ZN(
        n20375) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20387), .B1(
        n20621), .B2(n20386), .ZN(n20374) );
  OAI211_X1 U23332 ( .C1(n20625), .C2(n20418), .A(n20375), .B(n20374), .ZN(
        P1_U3059) );
  AOI22_X1 U23333 ( .A1(n20626), .A2(n20385), .B1(n20410), .B2(n20571), .ZN(
        n20377) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20387), .B1(
        n20627), .B2(n20386), .ZN(n20376) );
  OAI211_X1 U23335 ( .C1(n20574), .C2(n20390), .A(n20377), .B(n20376), .ZN(
        P1_U3060) );
  AOI22_X1 U23336 ( .A1(n20632), .A2(n20385), .B1(n20380), .B2(n20634), .ZN(
        n20379) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20387), .B1(
        n20633), .B2(n20386), .ZN(n20378) );
  OAI211_X1 U23338 ( .C1(n20637), .C2(n20418), .A(n20379), .B(n20378), .ZN(
        P1_U3061) );
  AOI22_X1 U23339 ( .A1(n20638), .A2(n20385), .B1(n20380), .B2(n20640), .ZN(
        n20382) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20387), .B1(
        n20639), .B2(n20386), .ZN(n20381) );
  OAI211_X1 U23341 ( .C1(n20643), .C2(n20418), .A(n20382), .B(n20381), .ZN(
        P1_U3062) );
  AOI22_X1 U23342 ( .A1(n20644), .A2(n20385), .B1(n20410), .B2(n20583), .ZN(
        n20384) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20387), .B1(
        n20645), .B2(n20386), .ZN(n20383) );
  OAI211_X1 U23344 ( .C1(n20586), .C2(n20390), .A(n20384), .B(n20383), .ZN(
        P1_U3063) );
  AOI22_X1 U23345 ( .A1(n20651), .A2(n20385), .B1(n20410), .B2(n20587), .ZN(
        n20389) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20387), .B1(
        n20653), .B2(n20386), .ZN(n20388) );
  OAI211_X1 U23347 ( .C1(n20594), .C2(n20390), .A(n20389), .B(n20388), .ZN(
        P1_U3064) );
  NAND2_X1 U23348 ( .A1(n20551), .A2(n20518), .ZN(n20392) );
  OAI22_X1 U23349 ( .A1(n20393), .A2(n20392), .B1(n20557), .B2(n20391), .ZN(
        n20413) );
  AOI22_X1 U23350 ( .A1(n20604), .A2(n20413), .B1(n20603), .B2(n9874), .ZN(
        n20399) );
  INV_X1 U23351 ( .A(n20393), .ZN(n20420) );
  AOI21_X1 U23352 ( .B1(n20418), .B2(n20446), .A(n20453), .ZN(n20395) );
  AOI21_X1 U23353 ( .B1(n20420), .B2(n20551), .A(n20395), .ZN(n20396) );
  NOR2_X1 U23354 ( .A1(n20396), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20397) );
  INV_X1 U23355 ( .A(n20446), .ZN(n20414) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20546), .ZN(n20398) );
  OAI211_X1 U23357 ( .C1(n20562), .C2(n20418), .A(n20399), .B(n20398), .ZN(
        P1_U3065) );
  AOI22_X1 U23358 ( .A1(n20615), .A2(n20413), .B1(n20614), .B2(n9874), .ZN(
        n20401) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20563), .ZN(n20400) );
  OAI211_X1 U23360 ( .C1(n20566), .C2(n20418), .A(n20401), .B(n20400), .ZN(
        P1_U3066) );
  AOI22_X1 U23361 ( .A1(n20621), .A2(n20413), .B1(n20620), .B2(n9874), .ZN(
        n20403) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20415), .B1(
        n20410), .B2(n20622), .ZN(n20402) );
  OAI211_X1 U23363 ( .C1(n20625), .C2(n20446), .A(n20403), .B(n20402), .ZN(
        P1_U3067) );
  AOI22_X1 U23364 ( .A1(n20627), .A2(n20413), .B1(n20626), .B2(n9874), .ZN(
        n20405) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20415), .B1(
        n20410), .B2(n20628), .ZN(n20404) );
  OAI211_X1 U23366 ( .C1(n20631), .C2(n20446), .A(n20405), .B(n20404), .ZN(
        P1_U3068) );
  AOI22_X1 U23367 ( .A1(n20633), .A2(n20413), .B1(n20632), .B2(n9874), .ZN(
        n20407) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20415), .B1(
        n20410), .B2(n20634), .ZN(n20406) );
  OAI211_X1 U23369 ( .C1(n20637), .C2(n20446), .A(n20407), .B(n20406), .ZN(
        P1_U3069) );
  AOI22_X1 U23370 ( .A1(n20639), .A2(n20413), .B1(n20638), .B2(n9874), .ZN(
        n20409) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20579), .ZN(n20408) );
  OAI211_X1 U23372 ( .C1(n20582), .C2(n20418), .A(n20409), .B(n20408), .ZN(
        P1_U3070) );
  AOI22_X1 U23373 ( .A1(n20645), .A2(n20413), .B1(n20644), .B2(n9874), .ZN(
        n20412) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20415), .B1(
        n20410), .B2(n20646), .ZN(n20411) );
  OAI211_X1 U23375 ( .C1(n20649), .C2(n20446), .A(n20412), .B(n20411), .ZN(
        P1_U3071) );
  AOI22_X1 U23376 ( .A1(n20653), .A2(n20413), .B1(n20651), .B2(n9874), .ZN(
        n20417) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20587), .ZN(n20416) );
  OAI211_X1 U23378 ( .C1(n20594), .C2(n20418), .A(n20417), .B(n20416), .ZN(
        P1_U3072) );
  NOR2_X1 U23379 ( .A1(n20419), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20425) );
  INV_X1 U23380 ( .A(n20425), .ZN(n20421) );
  NOR2_X1 U23381 ( .A1(n20449), .A2(n20421), .ZN(n20440) );
  AOI21_X1 U23382 ( .B1(n20420), .B2(n20450), .A(n20440), .ZN(n20422) );
  OAI22_X1 U23383 ( .A1(n20422), .A2(n20601), .B1(n20421), .B2(n12842), .ZN(
        n20441) );
  AOI22_X1 U23384 ( .A1(n20604), .A2(n20441), .B1(n20603), .B2(n20440), .ZN(
        n20427) );
  OAI211_X1 U23385 ( .C1(n20423), .C2(n20453), .A(n20518), .B(n20422), .ZN(
        n20424) );
  OAI211_X1 U23386 ( .C1(n20548), .C2(n20425), .A(n20607), .B(n20424), .ZN(
        n20443) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20546), .ZN(n20426) );
  OAI211_X1 U23388 ( .C1(n20562), .C2(n20446), .A(n20427), .B(n20426), .ZN(
        P1_U3073) );
  AOI22_X1 U23389 ( .A1(n20615), .A2(n20441), .B1(n20614), .B2(n20440), .ZN(
        n20429) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20563), .ZN(n20428) );
  OAI211_X1 U23391 ( .C1(n20566), .C2(n20446), .A(n20429), .B(n20428), .ZN(
        P1_U3074) );
  AOI22_X1 U23392 ( .A1(n20621), .A2(n20441), .B1(n20620), .B2(n20440), .ZN(
        n20431) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20567), .ZN(n20430) );
  OAI211_X1 U23394 ( .C1(n20570), .C2(n20446), .A(n20431), .B(n20430), .ZN(
        P1_U3075) );
  AOI22_X1 U23395 ( .A1(n20627), .A2(n20441), .B1(n20626), .B2(n20440), .ZN(
        n20433) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20571), .ZN(n20432) );
  OAI211_X1 U23397 ( .C1(n20574), .C2(n20446), .A(n20433), .B(n20432), .ZN(
        P1_U3076) );
  AOI22_X1 U23398 ( .A1(n20633), .A2(n20441), .B1(n20632), .B2(n20440), .ZN(
        n20435) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20575), .ZN(n20434) );
  OAI211_X1 U23400 ( .C1(n20578), .C2(n20446), .A(n20435), .B(n20434), .ZN(
        P1_U3077) );
  AOI22_X1 U23401 ( .A1(n20639), .A2(n20441), .B1(n20638), .B2(n20440), .ZN(
        n20437) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20579), .ZN(n20436) );
  OAI211_X1 U23403 ( .C1(n20582), .C2(n20446), .A(n20437), .B(n20436), .ZN(
        P1_U3078) );
  AOI22_X1 U23404 ( .A1(n20645), .A2(n20441), .B1(n20644), .B2(n20440), .ZN(
        n20439) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20583), .ZN(n20438) );
  OAI211_X1 U23406 ( .C1(n20586), .C2(n20446), .A(n20439), .B(n20438), .ZN(
        P1_U3079) );
  AOI22_X1 U23407 ( .A1(n20653), .A2(n20441), .B1(n20651), .B2(n20440), .ZN(
        n20445) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20443), .B1(
        n20442), .B2(n20587), .ZN(n20444) );
  OAI211_X1 U23409 ( .C1(n20594), .C2(n20446), .A(n20445), .B(n20444), .ZN(
        P1_U3080) );
  INV_X1 U23410 ( .A(n20447), .ZN(n20448) );
  NOR2_X1 U23411 ( .A1(n20514), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20455) );
  INV_X1 U23412 ( .A(n20455), .ZN(n20451) );
  NOR2_X1 U23413 ( .A1(n20449), .A2(n20451), .ZN(n20471) );
  AOI21_X1 U23414 ( .B1(n20515), .B2(n20450), .A(n20471), .ZN(n20452) );
  OAI22_X1 U23415 ( .A1(n20452), .A2(n20601), .B1(n20451), .B2(n12842), .ZN(
        n20472) );
  AOI22_X1 U23416 ( .A1(n20604), .A2(n20472), .B1(n20603), .B2(n20471), .ZN(
        n20457) );
  OAI211_X1 U23417 ( .C1(n20520), .C2(n20453), .A(n20518), .B(n20452), .ZN(
        n20454) );
  OAI211_X1 U23418 ( .C1(n20548), .C2(n20455), .A(n20607), .B(n20454), .ZN(
        n20474) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(n20610), .ZN(n20456) );
  OAI211_X1 U23420 ( .C1(n20613), .C2(n20509), .A(n20457), .B(n20456), .ZN(
        P1_U3105) );
  AOI22_X1 U23421 ( .A1(n20615), .A2(n20472), .B1(n20614), .B2(n20471), .ZN(
        n20459) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(n20616), .ZN(n20458) );
  OAI211_X1 U23423 ( .C1(n20619), .C2(n20509), .A(n20459), .B(n20458), .ZN(
        P1_U3106) );
  AOI22_X1 U23424 ( .A1(n20621), .A2(n20472), .B1(n20620), .B2(n20471), .ZN(
        n20461) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(n20622), .ZN(n20460) );
  OAI211_X1 U23426 ( .C1(n20625), .C2(n20509), .A(n20461), .B(n20460), .ZN(
        P1_U3107) );
  INV_X1 U23427 ( .A(n20473), .ZN(n20470) );
  AOI22_X1 U23428 ( .A1(n20627), .A2(n20472), .B1(n20626), .B2(n20471), .ZN(
        n20463) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20474), .B1(
        n20501), .B2(n20571), .ZN(n20462) );
  OAI211_X1 U23430 ( .C1(n20574), .C2(n20470), .A(n20463), .B(n20462), .ZN(
        P1_U3108) );
  AOI22_X1 U23431 ( .A1(n20633), .A2(n20472), .B1(n20632), .B2(n20471), .ZN(
        n20465) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20474), .B1(
        n20501), .B2(n20575), .ZN(n20464) );
  OAI211_X1 U23433 ( .C1(n20578), .C2(n20470), .A(n20465), .B(n20464), .ZN(
        P1_U3109) );
  AOI22_X1 U23434 ( .A1(n20639), .A2(n20472), .B1(n20638), .B2(n20471), .ZN(
        n20467) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20474), .B1(
        n20501), .B2(n20579), .ZN(n20466) );
  OAI211_X1 U23436 ( .C1(n20582), .C2(n20470), .A(n20467), .B(n20466), .ZN(
        P1_U3110) );
  AOI22_X1 U23437 ( .A1(n20645), .A2(n20472), .B1(n20644), .B2(n20471), .ZN(
        n20469) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20474), .B1(
        n20501), .B2(n20583), .ZN(n20468) );
  OAI211_X1 U23439 ( .C1(n20586), .C2(n20470), .A(n20469), .B(n20468), .ZN(
        P1_U3111) );
  AOI22_X1 U23440 ( .A1(n20653), .A2(n20472), .B1(n20651), .B2(n20471), .ZN(
        n20476) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20474), .B1(
        n20473), .B2(n20654), .ZN(n20475) );
  OAI211_X1 U23442 ( .C1(n20660), .C2(n20509), .A(n20476), .B(n20475), .ZN(
        P1_U3112) );
  NOR2_X1 U23443 ( .A1(n20599), .A2(n20514), .ZN(n20522) );
  INV_X1 U23444 ( .A(n20522), .ZN(n20516) );
  NOR2_X1 U23445 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20516), .ZN(
        n20504) );
  INV_X1 U23446 ( .A(n20477), .ZN(n20478) );
  NAND2_X1 U23447 ( .A1(n20512), .A2(n20478), .ZN(n20530) );
  AOI22_X1 U23448 ( .A1(n20603), .A2(n20504), .B1(n20541), .B2(n20546), .ZN(
        n20490) );
  OAI21_X1 U23449 ( .B1(n20541), .B2(n20501), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20479) );
  NAND2_X1 U23450 ( .A1(n20479), .A2(n20548), .ZN(n20488) );
  AND2_X1 U23451 ( .A1(n20515), .A2(n11887), .ZN(n20484) );
  OAI211_X1 U23452 ( .C1(n20554), .C2(n20504), .A(n20481), .B(n20480), .ZN(
        n20482) );
  INV_X1 U23453 ( .A(n20482), .ZN(n20483) );
  INV_X1 U23454 ( .A(n20484), .ZN(n20487) );
  OAI22_X1 U23455 ( .A1(n20488), .A2(n20487), .B1(n20486), .B2(n20485), .ZN(
        n20505) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20506), .B1(
        n20604), .B2(n20505), .ZN(n20489) );
  OAI211_X1 U23457 ( .C1(n20562), .C2(n20509), .A(n20490), .B(n20489), .ZN(
        P1_U3113) );
  AOI22_X1 U23458 ( .A1(n20614), .A2(n20504), .B1(n20541), .B2(n20563), .ZN(
        n20492) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20506), .B1(
        n20615), .B2(n20505), .ZN(n20491) );
  OAI211_X1 U23460 ( .C1(n20566), .C2(n20509), .A(n20492), .B(n20491), .ZN(
        P1_U3114) );
  AOI22_X1 U23461 ( .A1(n20620), .A2(n20504), .B1(n20541), .B2(n20567), .ZN(
        n20494) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20506), .B1(
        n20621), .B2(n20505), .ZN(n20493) );
  OAI211_X1 U23463 ( .C1(n20570), .C2(n20509), .A(n20494), .B(n20493), .ZN(
        P1_U3115) );
  AOI22_X1 U23464 ( .A1(n20626), .A2(n20504), .B1(n20501), .B2(n20628), .ZN(
        n20496) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20506), .B1(
        n20627), .B2(n20505), .ZN(n20495) );
  OAI211_X1 U23466 ( .C1(n20631), .C2(n20530), .A(n20496), .B(n20495), .ZN(
        P1_U3116) );
  AOI22_X1 U23467 ( .A1(n20632), .A2(n20504), .B1(n20541), .B2(n20575), .ZN(
        n20498) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20506), .B1(
        n20633), .B2(n20505), .ZN(n20497) );
  OAI211_X1 U23469 ( .C1(n20578), .C2(n20509), .A(n20498), .B(n20497), .ZN(
        P1_U3117) );
  AOI22_X1 U23470 ( .A1(n20638), .A2(n20504), .B1(n20541), .B2(n20579), .ZN(
        n20500) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20506), .B1(
        n20639), .B2(n20505), .ZN(n20499) );
  OAI211_X1 U23472 ( .C1(n20582), .C2(n20509), .A(n20500), .B(n20499), .ZN(
        P1_U3118) );
  AOI22_X1 U23473 ( .A1(n20644), .A2(n20504), .B1(n20501), .B2(n20646), .ZN(
        n20503) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20506), .B1(
        n20645), .B2(n20505), .ZN(n20502) );
  OAI211_X1 U23475 ( .C1(n20649), .C2(n20530), .A(n20503), .B(n20502), .ZN(
        P1_U3119) );
  AOI22_X1 U23476 ( .A1(n20651), .A2(n20504), .B1(n20541), .B2(n20587), .ZN(
        n20508) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20506), .B1(
        n20653), .B2(n20505), .ZN(n20507) );
  OAI211_X1 U23478 ( .C1(n20594), .C2(n20509), .A(n20508), .B(n20507), .ZN(
        P1_U3120) );
  INV_X1 U23479 ( .A(n20510), .ZN(n20511) );
  INV_X1 U23480 ( .A(n20513), .ZN(n20596) );
  NOR2_X1 U23481 ( .A1(n20595), .A2(n20514), .ZN(n20539) );
  AOI21_X1 U23482 ( .B1(n20515), .B2(n20596), .A(n20539), .ZN(n20517) );
  OAI22_X1 U23483 ( .A1(n20517), .A2(n20601), .B1(n20516), .B2(n12842), .ZN(
        n20540) );
  AOI22_X1 U23484 ( .A1(n20604), .A2(n20540), .B1(n20603), .B2(n20539), .ZN(
        n20524) );
  OAI211_X1 U23485 ( .C1(n20520), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        n20521) );
  OAI211_X1 U23486 ( .C1(n20548), .C2(n20522), .A(n20607), .B(n20521), .ZN(
        n20542) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20610), .ZN(n20523) );
  OAI211_X1 U23488 ( .C1(n20613), .C2(n20593), .A(n20524), .B(n20523), .ZN(
        P1_U3121) );
  AOI22_X1 U23489 ( .A1(n20615), .A2(n20540), .B1(n20614), .B2(n20539), .ZN(
        n20526) );
  INV_X1 U23490 ( .A(n20593), .ZN(n20527) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20542), .B1(
        n20527), .B2(n20563), .ZN(n20525) );
  OAI211_X1 U23492 ( .C1(n20566), .C2(n20530), .A(n20526), .B(n20525), .ZN(
        P1_U3122) );
  AOI22_X1 U23493 ( .A1(n20621), .A2(n20540), .B1(n20620), .B2(n20539), .ZN(
        n20529) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20542), .B1(
        n20527), .B2(n20567), .ZN(n20528) );
  OAI211_X1 U23495 ( .C1(n20570), .C2(n20530), .A(n20529), .B(n20528), .ZN(
        P1_U3123) );
  AOI22_X1 U23496 ( .A1(n20627), .A2(n20540), .B1(n20626), .B2(n20539), .ZN(
        n20532) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20628), .ZN(n20531) );
  OAI211_X1 U23498 ( .C1(n20631), .C2(n20593), .A(n20532), .B(n20531), .ZN(
        P1_U3124) );
  AOI22_X1 U23499 ( .A1(n20633), .A2(n20540), .B1(n20632), .B2(n20539), .ZN(
        n20534) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20634), .ZN(n20533) );
  OAI211_X1 U23501 ( .C1(n20637), .C2(n20593), .A(n20534), .B(n20533), .ZN(
        P1_U3125) );
  AOI22_X1 U23502 ( .A1(n20639), .A2(n20540), .B1(n20638), .B2(n20539), .ZN(
        n20536) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20640), .ZN(n20535) );
  OAI211_X1 U23504 ( .C1(n20643), .C2(n20593), .A(n20536), .B(n20535), .ZN(
        P1_U3126) );
  AOI22_X1 U23505 ( .A1(n20645), .A2(n20540), .B1(n20644), .B2(n20539), .ZN(
        n20538) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20646), .ZN(n20537) );
  OAI211_X1 U23507 ( .C1(n20649), .C2(n20593), .A(n20538), .B(n20537), .ZN(
        P1_U3127) );
  AOI22_X1 U23508 ( .A1(n20653), .A2(n20540), .B1(n20651), .B2(n20539), .ZN(
        n20544) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20654), .ZN(n20543) );
  OAI211_X1 U23510 ( .C1(n20660), .C2(n20593), .A(n20544), .B(n20543), .ZN(
        P1_U3128) );
  AOI22_X1 U23511 ( .A1(n20603), .A2(n9875), .B1(n20588), .B2(n20546), .ZN(
        n20561) );
  NAND3_X1 U23512 ( .A1(n20593), .A2(n20548), .A3(n20547), .ZN(n20550) );
  NAND2_X1 U23513 ( .A1(n20550), .A2(n20549), .ZN(n20555) );
  NAND2_X1 U23514 ( .A1(n20597), .A2(n20551), .ZN(n20558) );
  AOI22_X1 U23515 ( .A1(n20555), .A2(n20558), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20556), .ZN(n20552) );
  OAI211_X1 U23516 ( .C1(n9875), .C2(n20554), .A(n20553), .B(n20552), .ZN(
        n20590) );
  INV_X1 U23517 ( .A(n20555), .ZN(n20559) );
  OAI22_X1 U23518 ( .A1(n20559), .A2(n20558), .B1(n20557), .B2(n20556), .ZN(
        n20589) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20590), .B1(
        n20604), .B2(n20589), .ZN(n20560) );
  OAI211_X1 U23520 ( .C1(n20562), .C2(n20593), .A(n20561), .B(n20560), .ZN(
        P1_U3129) );
  AOI22_X1 U23521 ( .A1(n20614), .A2(n9875), .B1(n20588), .B2(n20563), .ZN(
        n20565) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20590), .B1(
        n20615), .B2(n20589), .ZN(n20564) );
  OAI211_X1 U23523 ( .C1(n20566), .C2(n20593), .A(n20565), .B(n20564), .ZN(
        P1_U3130) );
  AOI22_X1 U23524 ( .A1(n20620), .A2(n9875), .B1(n20567), .B2(n20588), .ZN(
        n20569) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20590), .B1(
        n20621), .B2(n20589), .ZN(n20568) );
  OAI211_X1 U23526 ( .C1(n20570), .C2(n20593), .A(n20569), .B(n20568), .ZN(
        P1_U3131) );
  AOI22_X1 U23527 ( .A1(n20626), .A2(n9875), .B1(n20588), .B2(n20571), .ZN(
        n20573) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20590), .B1(
        n20627), .B2(n20589), .ZN(n20572) );
  OAI211_X1 U23529 ( .C1(n20574), .C2(n20593), .A(n20573), .B(n20572), .ZN(
        P1_U3132) );
  AOI22_X1 U23530 ( .A1(n20632), .A2(n9875), .B1(n20588), .B2(n20575), .ZN(
        n20577) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20590), .B1(
        n20633), .B2(n20589), .ZN(n20576) );
  OAI211_X1 U23532 ( .C1(n20578), .C2(n20593), .A(n20577), .B(n20576), .ZN(
        P1_U3133) );
  AOI22_X1 U23533 ( .A1(n20638), .A2(n9875), .B1(n20588), .B2(n20579), .ZN(
        n20581) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20590), .B1(
        n20639), .B2(n20589), .ZN(n20580) );
  OAI211_X1 U23535 ( .C1(n20582), .C2(n20593), .A(n20581), .B(n20580), .ZN(
        P1_U3134) );
  AOI22_X1 U23536 ( .A1(n20644), .A2(n9875), .B1(n20588), .B2(n20583), .ZN(
        n20585) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20590), .B1(
        n20645), .B2(n20589), .ZN(n20584) );
  OAI211_X1 U23538 ( .C1(n20586), .C2(n20593), .A(n20585), .B(n20584), .ZN(
        P1_U3135) );
  AOI22_X1 U23539 ( .A1(n20651), .A2(n9875), .B1(n20588), .B2(n20587), .ZN(
        n20592) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20590), .B1(
        n20653), .B2(n20589), .ZN(n20591) );
  OAI211_X1 U23541 ( .C1(n20594), .C2(n20593), .A(n20592), .B(n20591), .ZN(
        P1_U3136) );
  NOR2_X1 U23542 ( .A1(n20595), .A2(n20598), .ZN(n20650) );
  AOI21_X1 U23543 ( .B1(n20597), .B2(n20596), .A(n20650), .ZN(n20602) );
  NOR2_X1 U23544 ( .A1(n20599), .A2(n20598), .ZN(n20608) );
  INV_X1 U23545 ( .A(n20608), .ZN(n20600) );
  OAI22_X1 U23546 ( .A1(n20602), .A2(n20601), .B1(n20600), .B2(n12842), .ZN(
        n20652) );
  AOI22_X1 U23547 ( .A1(n20604), .A2(n20652), .B1(n20603), .B2(n20650), .ZN(
        n20612) );
  NOR2_X1 U23548 ( .A1(n20606), .A2(n20605), .ZN(n20609) );
  OAI21_X1 U23549 ( .B1(n20609), .B2(n20608), .A(n20607), .ZN(n20656) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20610), .ZN(n20611) );
  OAI211_X1 U23551 ( .C1(n20613), .C2(n20659), .A(n20612), .B(n20611), .ZN(
        P1_U3153) );
  AOI22_X1 U23552 ( .A1(n20615), .A2(n20652), .B1(n20614), .B2(n20650), .ZN(
        n20618) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20616), .ZN(n20617) );
  OAI211_X1 U23554 ( .C1(n20619), .C2(n20659), .A(n20618), .B(n20617), .ZN(
        P1_U3154) );
  AOI22_X1 U23555 ( .A1(n20621), .A2(n20652), .B1(n20620), .B2(n20650), .ZN(
        n20624) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20622), .ZN(n20623) );
  OAI211_X1 U23557 ( .C1(n20625), .C2(n20659), .A(n20624), .B(n20623), .ZN(
        P1_U3155) );
  AOI22_X1 U23558 ( .A1(n20627), .A2(n20652), .B1(n20626), .B2(n20650), .ZN(
        n20630) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20628), .ZN(n20629) );
  OAI211_X1 U23560 ( .C1(n20631), .C2(n20659), .A(n20630), .B(n20629), .ZN(
        P1_U3156) );
  AOI22_X1 U23561 ( .A1(n20633), .A2(n20652), .B1(n20632), .B2(n20650), .ZN(
        n20636) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20634), .ZN(n20635) );
  OAI211_X1 U23563 ( .C1(n20637), .C2(n20659), .A(n20636), .B(n20635), .ZN(
        P1_U3157) );
  AOI22_X1 U23564 ( .A1(n20639), .A2(n20652), .B1(n20638), .B2(n20650), .ZN(
        n20642) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20640), .ZN(n20641) );
  OAI211_X1 U23566 ( .C1(n20643), .C2(n20659), .A(n20642), .B(n20641), .ZN(
        P1_U3158) );
  AOI22_X1 U23567 ( .A1(n20645), .A2(n20652), .B1(n20644), .B2(n20650), .ZN(
        n20648) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20646), .ZN(n20647) );
  OAI211_X1 U23569 ( .C1(n20649), .C2(n20659), .A(n20648), .B(n20647), .ZN(
        P1_U3159) );
  AOI22_X1 U23570 ( .A1(n20653), .A2(n20652), .B1(n20651), .B2(n20650), .ZN(
        n20658) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20656), .B1(
        n20655), .B2(n20654), .ZN(n20657) );
  OAI211_X1 U23572 ( .C1(n20660), .C2(n20659), .A(n20658), .B(n20657), .ZN(
        P1_U3160) );
  NOR2_X1 U23573 ( .A1(n11886), .A2(n20661), .ZN(n20663) );
  OAI21_X1 U23574 ( .B1(n20663), .B2(n12842), .A(n20662), .ZN(P1_U3163) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20664), .ZN(
        P1_U3164) );
  AND2_X1 U23576 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20664), .ZN(
        P1_U3165) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20664), .ZN(
        P1_U3166) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20664), .ZN(
        P1_U3167) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20664), .ZN(
        P1_U3168) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20664), .ZN(
        P1_U3169) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20664), .ZN(
        P1_U3170) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20664), .ZN(
        P1_U3171) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20664), .ZN(
        P1_U3172) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20664), .ZN(
        P1_U3173) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20664), .ZN(
        P1_U3174) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20664), .ZN(
        P1_U3175) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20664), .ZN(
        P1_U3176) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20664), .ZN(
        P1_U3177) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20664), .ZN(
        P1_U3178) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20664), .ZN(
        P1_U3179) );
  AND2_X1 U23591 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20664), .ZN(
        P1_U3180) );
  AND2_X1 U23592 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20664), .ZN(
        P1_U3181) );
  AND2_X1 U23593 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20664), .ZN(
        P1_U3182) );
  AND2_X1 U23594 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20664), .ZN(
        P1_U3183) );
  AND2_X1 U23595 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20664), .ZN(
        P1_U3184) );
  AND2_X1 U23596 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20664), .ZN(
        P1_U3185) );
  AND2_X1 U23597 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20664), .ZN(P1_U3186) );
  AND2_X1 U23598 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20664), .ZN(P1_U3187) );
  AND2_X1 U23599 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20664), .ZN(P1_U3188) );
  AND2_X1 U23600 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20664), .ZN(P1_U3189) );
  AND2_X1 U23601 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20664), .ZN(P1_U3190) );
  AND2_X1 U23602 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20664), .ZN(P1_U3191) );
  AND2_X1 U23603 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20664), .ZN(P1_U3192) );
  AND2_X1 U23604 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20664), .ZN(P1_U3193) );
  NAND2_X1 U23605 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20680), .ZN(n20670) );
  NAND2_X1 U23606 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n20665) );
  OAI211_X1 U23607 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n20906), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n20665), .ZN(n20666) );
  OAI21_X1 U23608 ( .B1(n20667), .B2(n20666), .A(n20751), .ZN(n20668) );
  OAI211_X1 U23609 ( .C1(n20670), .C2(n20747), .A(n20669), .B(n20668), .ZN(
        P1_U3194) );
  NAND2_X1 U23610 ( .A1(n20906), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20673) );
  INV_X1 U23611 ( .A(n20673), .ZN(n20671) );
  AOI21_X1 U23612 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20671), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20679) );
  INV_X1 U23613 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20675) );
  OAI21_X1 U23614 ( .B1(n20747), .B2(n20673), .A(n20672), .ZN(n20674) );
  OAI211_X1 U23615 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20675), .A(HOLD), .B(
        n20674), .ZN(n20677) );
  OAI211_X1 U23616 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20906), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n12089), .ZN(n20676) );
  OAI211_X1 U23617 ( .C1(n20679), .C2(n20678), .A(n20677), .B(n20676), .ZN(
        P1_U3196) );
  OR2_X1 U23618 ( .A1(n20751), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20717) );
  OR2_X1 U23619 ( .A1(n20680), .A2(n20751), .ZN(n20720) );
  INV_X1 U23620 ( .A(n20720), .ZN(n20715) );
  AOI222_X1 U23621 ( .A1(n9735), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20751), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20715), .ZN(n20681) );
  INV_X1 U23622 ( .A(n20681), .ZN(P1_U3197) );
  AOI222_X1 U23623 ( .A1(n20715), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n9735), .ZN(n20682) );
  INV_X1 U23624 ( .A(n20682), .ZN(P1_U3198) );
  OAI222_X1 U23625 ( .A1(n20720), .A2(n20685), .B1(n20684), .B2(n20738), .C1(
        n20683), .C2(n20717), .ZN(P1_U3199) );
  AOI222_X1 U23626 ( .A1(n9735), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20715), .ZN(n20686) );
  INV_X1 U23627 ( .A(n20686), .ZN(P1_U3200) );
  AOI222_X1 U23628 ( .A1(n20715), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n9735), .ZN(n20687) );
  INV_X1 U23629 ( .A(n20687), .ZN(P1_U3201) );
  AOI222_X1 U23630 ( .A1(n9735), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20715), .ZN(n20688) );
  INV_X1 U23631 ( .A(n20688), .ZN(P1_U3202) );
  AOI222_X1 U23632 ( .A1(n20715), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n9735), .ZN(n20689) );
  INV_X1 U23633 ( .A(n20689), .ZN(P1_U3203) );
  AOI222_X1 U23634 ( .A1(n20715), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n9735), .ZN(n20690) );
  INV_X1 U23635 ( .A(n20690), .ZN(P1_U3204) );
  AOI222_X1 U23636 ( .A1(n20715), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n9735), .ZN(n20691) );
  INV_X1 U23637 ( .A(n20691), .ZN(P1_U3205) );
  AOI222_X1 U23638 ( .A1(n20715), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n9735), .ZN(n20692) );
  INV_X1 U23639 ( .A(n20692), .ZN(P1_U3206) );
  AOI22_X1 U23640 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20751), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n9735), .ZN(n20693) );
  OAI21_X1 U23641 ( .B1(n20694), .B2(n20720), .A(n20693), .ZN(P1_U3207) );
  AOI22_X1 U23642 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20751), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20715), .ZN(n20695) );
  OAI21_X1 U23643 ( .B1(n20697), .B2(n20717), .A(n20695), .ZN(P1_U3208) );
  AOI22_X1 U23644 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20751), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n9735), .ZN(n20696) );
  OAI21_X1 U23645 ( .B1(n20697), .B2(n20720), .A(n20696), .ZN(P1_U3209) );
  AOI22_X1 U23646 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20751), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20715), .ZN(n20698) );
  OAI21_X1 U23647 ( .B1(n20699), .B2(n20717), .A(n20698), .ZN(P1_U3210) );
  AOI222_X1 U23648 ( .A1(n20715), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n9735), .ZN(n20700) );
  INV_X1 U23649 ( .A(n20700), .ZN(P1_U3211) );
  AOI222_X1 U23650 ( .A1(n20715), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n9735), .ZN(n20701) );
  INV_X1 U23651 ( .A(n20701), .ZN(P1_U3212) );
  AOI222_X1 U23652 ( .A1(n9735), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20715), .ZN(n20702) );
  INV_X1 U23653 ( .A(n20702), .ZN(P1_U3213) );
  AOI222_X1 U23654 ( .A1(n9735), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20715), .ZN(n20703) );
  INV_X1 U23655 ( .A(n20703), .ZN(P1_U3214) );
  AOI22_X1 U23656 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20751), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n9735), .ZN(n20704) );
  OAI21_X1 U23657 ( .B1(n20705), .B2(n20720), .A(n20704), .ZN(P1_U3215) );
  AOI222_X1 U23658 ( .A1(n20715), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n9735), .ZN(n20706) );
  INV_X1 U23659 ( .A(n20706), .ZN(P1_U3216) );
  AOI222_X1 U23660 ( .A1(n20715), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n9735), .ZN(n20707) );
  INV_X1 U23661 ( .A(n20707), .ZN(P1_U3217) );
  AOI222_X1 U23662 ( .A1(n20715), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n9735), .ZN(n20708) );
  INV_X1 U23663 ( .A(n20708), .ZN(P1_U3218) );
  AOI222_X1 U23664 ( .A1(n20715), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n9735), .ZN(n20709) );
  INV_X1 U23665 ( .A(n20709), .ZN(P1_U3219) );
  AOI222_X1 U23666 ( .A1(n20715), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20751), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n9735), .ZN(n20710) );
  INV_X1 U23667 ( .A(n20710), .ZN(P1_U3220) );
  AOI222_X1 U23668 ( .A1(n20715), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n9735), .ZN(n20711) );
  INV_X1 U23669 ( .A(n20711), .ZN(P1_U3221) );
  AOI222_X1 U23670 ( .A1(n20715), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n9735), .ZN(n20712) );
  INV_X1 U23671 ( .A(n20712), .ZN(P1_U3222) );
  AOI222_X1 U23672 ( .A1(n20715), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n9735), .ZN(n20713) );
  INV_X1 U23673 ( .A(n20713), .ZN(P1_U3223) );
  AOI222_X1 U23674 ( .A1(n20715), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n9735), .ZN(n20714) );
  INV_X1 U23675 ( .A(n20714), .ZN(P1_U3224) );
  AOI222_X1 U23676 ( .A1(n20715), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n9735), .ZN(n20716) );
  INV_X1 U23677 ( .A(n20716), .ZN(P1_U3225) );
  INV_X1 U23678 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20866) );
  INV_X1 U23679 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20718) );
  OAI222_X1 U23680 ( .A1(n20720), .A2(n20719), .B1(n20866), .B2(n20738), .C1(
        n20718), .C2(n20717), .ZN(P1_U3226) );
  OAI22_X1 U23681 ( .A1(n20751), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20738), .ZN(n20721) );
  INV_X1 U23682 ( .A(n20721), .ZN(P1_U3458) );
  OAI22_X1 U23683 ( .A1(n20736), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20738), .ZN(n20722) );
  INV_X1 U23684 ( .A(n20722), .ZN(P1_U3459) );
  OAI22_X1 U23685 ( .A1(n20751), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20738), .ZN(n20723) );
  INV_X1 U23686 ( .A(n20723), .ZN(P1_U3460) );
  OAI22_X1 U23687 ( .A1(n20751), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20738), .ZN(n20724) );
  INV_X1 U23688 ( .A(n20724), .ZN(P1_U3461) );
  OAI21_X1 U23689 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20728), .A(n20726), 
        .ZN(n20725) );
  INV_X1 U23690 ( .A(n20725), .ZN(P1_U3464) );
  OAI21_X1 U23691 ( .B1(n20728), .B2(n20727), .A(n20726), .ZN(P1_U3465) );
  AOI211_X1 U23692 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20729) );
  AOI21_X1 U23693 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20729), .ZN(n20731) );
  INV_X1 U23694 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20730) );
  AOI22_X1 U23695 ( .A1(n20735), .A2(n20731), .B1(n20730), .B2(n20732), .ZN(
        P1_U3481) );
  NOR2_X1 U23696 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20734) );
  INV_X1 U23697 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20733) );
  AOI22_X1 U23698 ( .A1(n20735), .A2(n20734), .B1(n20733), .B2(n20732), .ZN(
        P1_U3482) );
  AOI22_X1 U23699 ( .A1(n20738), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20737), 
        .B2(n20736), .ZN(P1_U3483) );
  OAI21_X1 U23700 ( .B1(n11818), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20742) );
  NOR2_X1 U23701 ( .A1(n20740), .A2(n20739), .ZN(n20741) );
  OAI21_X1 U23702 ( .B1(n20743), .B2(n20742), .A(n20741), .ZN(n20744) );
  INV_X1 U23703 ( .A(n20744), .ZN(n20750) );
  AOI211_X1 U23704 ( .C1(n20748), .C2(n20747), .A(n20746), .B(n20745), .ZN(
        n20749) );
  MUX2_X1 U23705 ( .A(n20750), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20749), 
        .Z(P1_U3485) );
  MUX2_X1 U23706 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20751), .Z(P1_U3486) );
  AOI22_X1 U23707 ( .A1(n20753), .A2(n20904), .B1(n20752), .B2(n20906), .ZN(
        n20754) );
  AOI21_X1 U23708 ( .B1(n20904), .B2(n20852), .A(n20754), .ZN(n20760) );
  NAND2_X1 U23709 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20757) );
  OAI21_X1 U23710 ( .B1(n20757), .B2(n20756), .A(n20755), .ZN(n20758) );
  AOI22_X1 U23711 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20760), .B1(n20759), 
        .B2(n20758), .ZN(n21087) );
  NAND4_X1 U23712 ( .A1(keyinput60), .A2(keyinput73), .A3(keyinput46), .A4(
        keyinput85), .ZN(n20767) );
  INV_X1 U23713 ( .A(keyinput50), .ZN(n20761) );
  NAND4_X1 U23714 ( .A1(keyinput107), .A2(keyinput31), .A3(keyinput48), .A4(
        n20761), .ZN(n20766) );
  INV_X1 U23715 ( .A(keyinput125), .ZN(n20762) );
  NAND4_X1 U23716 ( .A1(keyinput77), .A2(keyinput122), .A3(keyinput20), .A4(
        n20762), .ZN(n20765) );
  NOR2_X1 U23717 ( .A1(keyinput104), .A2(keyinput1), .ZN(n20763) );
  NAND3_X1 U23718 ( .A1(keyinput7), .A2(keyinput76), .A3(n20763), .ZN(n20764)
         );
  NOR4_X1 U23719 ( .A1(n20767), .A2(n20766), .A3(n20765), .A4(n20764), .ZN(
        n20820) );
  INV_X1 U23720 ( .A(keyinput110), .ZN(n20768) );
  NOR4_X1 U23721 ( .A1(keyinput43), .A2(keyinput72), .A3(keyinput9), .A4(
        n20768), .ZN(n20769) );
  NAND3_X1 U23722 ( .A1(keyinput8), .A2(keyinput69), .A3(n20769), .ZN(n20773)
         );
  NOR2_X1 U23723 ( .A1(keyinput108), .A2(keyinput116), .ZN(n20770) );
  NAND3_X1 U23724 ( .A1(keyinput26), .A2(keyinput90), .A3(n20770), .ZN(n20772)
         );
  NAND4_X1 U23725 ( .A1(keyinput82), .A2(keyinput115), .A3(keyinput54), .A4(
        keyinput91), .ZN(n20771) );
  NOR4_X1 U23726 ( .A1(keyinput99), .A2(n20773), .A3(n20772), .A4(n20771), 
        .ZN(n20819) );
  INV_X1 U23727 ( .A(keyinput30), .ZN(n20789) );
  NOR4_X1 U23728 ( .A1(keyinput64), .A2(keyinput45), .A3(keyinput12), .A4(
        keyinput124), .ZN(n20774) );
  NAND3_X1 U23729 ( .A1(keyinput86), .A2(keyinput120), .A3(n20774), .ZN(n20788) );
  INV_X1 U23730 ( .A(keyinput119), .ZN(n20775) );
  NAND4_X1 U23731 ( .A1(keyinput49), .A2(keyinput21), .A3(keyinput112), .A4(
        n20775), .ZN(n20776) );
  NOR3_X1 U23732 ( .A1(keyinput93), .A2(keyinput65), .A3(n20776), .ZN(n20786)
         );
  NOR2_X1 U23733 ( .A1(keyinput23), .A2(keyinput123), .ZN(n20777) );
  NAND3_X1 U23734 ( .A1(keyinput3), .A2(keyinput95), .A3(n20777), .ZN(n20783)
         );
  NOR2_X1 U23735 ( .A1(keyinput10), .A2(keyinput98), .ZN(n20778) );
  NAND3_X1 U23736 ( .A1(keyinput39), .A2(keyinput80), .A3(n20778), .ZN(n20782)
         );
  NOR2_X1 U23737 ( .A1(keyinput61), .A2(keyinput78), .ZN(n20779) );
  NAND3_X1 U23738 ( .A1(keyinput11), .A2(keyinput84), .A3(n20779), .ZN(n20781)
         );
  NAND4_X1 U23739 ( .A1(keyinput74), .A2(keyinput121), .A3(keyinput67), .A4(
        keyinput59), .ZN(n20780) );
  NOR4_X1 U23740 ( .A1(n20783), .A2(n20782), .A3(n20781), .A4(n20780), .ZN(
        n20785) );
  INV_X1 U23741 ( .A(keyinput4), .ZN(n20784) );
  NAND4_X1 U23742 ( .A1(keyinput41), .A2(n20786), .A3(n20785), .A4(n20784), 
        .ZN(n20787) );
  NOR4_X1 U23743 ( .A1(keyinput66), .A2(n20789), .A3(n20788), .A4(n20787), 
        .ZN(n20818) );
  NOR2_X1 U23744 ( .A1(keyinput100), .A2(keyinput103), .ZN(n20790) );
  NAND3_X1 U23745 ( .A1(keyinput36), .A2(keyinput51), .A3(n20790), .ZN(n20791)
         );
  NOR3_X1 U23746 ( .A1(keyinput75), .A2(keyinput63), .A3(n20791), .ZN(n20803)
         );
  NAND4_X1 U23747 ( .A1(keyinput94), .A2(keyinput47), .A3(keyinput42), .A4(
        keyinput96), .ZN(n20801) );
  NOR2_X1 U23748 ( .A1(keyinput18), .A2(keyinput101), .ZN(n20792) );
  NAND3_X1 U23749 ( .A1(keyinput87), .A2(keyinput97), .A3(n20792), .ZN(n20800)
         );
  NOR4_X1 U23750 ( .A1(keyinput35), .A2(keyinput34), .A3(keyinput5), .A4(
        keyinput57), .ZN(n20798) );
  NAND2_X1 U23751 ( .A1(keyinput118), .A2(keyinput105), .ZN(n20793) );
  NOR3_X1 U23752 ( .A1(keyinput38), .A2(keyinput83), .A3(n20793), .ZN(n20797)
         );
  NAND2_X1 U23753 ( .A1(keyinput27), .A2(keyinput79), .ZN(n20794) );
  NOR3_X1 U23754 ( .A1(keyinput117), .A2(keyinput32), .A3(n20794), .ZN(n20796)
         );
  NOR4_X1 U23755 ( .A1(keyinput88), .A2(keyinput15), .A3(keyinput114), .A4(
        keyinput25), .ZN(n20795) );
  NAND4_X1 U23756 ( .A1(n20798), .A2(n20797), .A3(n20796), .A4(n20795), .ZN(
        n20799) );
  NOR3_X1 U23757 ( .A1(n20801), .A2(n20800), .A3(n20799), .ZN(n20802) );
  NAND4_X1 U23758 ( .A1(keyinput17), .A2(keyinput81), .A3(n20803), .A4(n20802), 
        .ZN(n20816) );
  NOR2_X1 U23759 ( .A1(keyinput68), .A2(keyinput55), .ZN(n20804) );
  NAND3_X1 U23760 ( .A1(keyinput62), .A2(keyinput70), .A3(n20804), .ZN(n20815)
         );
  NAND4_X1 U23761 ( .A1(keyinput56), .A2(keyinput71), .A3(keyinput14), .A4(
        keyinput22), .ZN(n20814) );
  NOR4_X1 U23762 ( .A1(keyinput109), .A2(keyinput92), .A3(keyinput16), .A4(
        keyinput33), .ZN(n20812) );
  NOR4_X1 U23763 ( .A1(keyinput44), .A2(keyinput52), .A3(keyinput127), .A4(
        keyinput2), .ZN(n20811) );
  NAND4_X1 U23764 ( .A1(keyinput6), .A2(keyinput111), .A3(keyinput102), .A4(
        keyinput106), .ZN(n20809) );
  NAND4_X1 U23765 ( .A1(keyinput19), .A2(keyinput58), .A3(keyinput113), .A4(
        keyinput28), .ZN(n20808) );
  NAND4_X1 U23766 ( .A1(keyinput53), .A2(keyinput0), .A3(keyinput89), .A4(
        keyinput40), .ZN(n20807) );
  NOR2_X1 U23767 ( .A1(keyinput29), .A2(keyinput13), .ZN(n20805) );
  NAND3_X1 U23768 ( .A1(keyinput24), .A2(keyinput37), .A3(n20805), .ZN(n20806)
         );
  NOR4_X1 U23769 ( .A1(n20809), .A2(n20808), .A3(n20807), .A4(n20806), .ZN(
        n20810) );
  NAND3_X1 U23770 ( .A1(n20812), .A2(n20811), .A3(n20810), .ZN(n20813) );
  NOR4_X1 U23771 ( .A1(n20816), .A2(n20815), .A3(n20814), .A4(n20813), .ZN(
        n20817) );
  NAND4_X1 U23772 ( .A1(n20820), .A2(n20819), .A3(n20818), .A4(n20817), .ZN(
        n21084) );
  AOI22_X1 U23773 ( .A1(n13101), .A2(keyinput55), .B1(keyinput14), .B2(n20822), 
        .ZN(n20821) );
  OAI221_X1 U23774 ( .B1(n13101), .B2(keyinput55), .C1(n20822), .C2(keyinput14), .A(n20821), .ZN(n20832) );
  AOI22_X1 U23775 ( .A1(n20825), .A2(keyinput68), .B1(keyinput70), .B2(n20824), 
        .ZN(n20823) );
  OAI221_X1 U23776 ( .B1(n20825), .B2(keyinput68), .C1(n20824), .C2(keyinput70), .A(n20823), .ZN(n20831) );
  AOI22_X1 U23777 ( .A1(n14798), .A2(keyinput71), .B1(n10766), .B2(keyinput62), 
        .ZN(n20826) );
  OAI221_X1 U23778 ( .B1(n14798), .B2(keyinput71), .C1(n10766), .C2(keyinput62), .A(n20826), .ZN(n20830) );
  XOR2_X1 U23779 ( .A(n14718), .B(keyinput22), .Z(n20828) );
  XNOR2_X1 U23780 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput19), 
        .ZN(n20827) );
  NAND2_X1 U23781 ( .A1(n20828), .A2(n20827), .ZN(n20829) );
  NOR4_X1 U23782 ( .A1(n20832), .A2(n20831), .A3(n20830), .A4(n20829), .ZN(
        n20884) );
  INV_X1 U23783 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U23784 ( .A1(n20835), .A2(keyinput111), .B1(n20834), .B2(
        keyinput102), .ZN(n20833) );
  OAI221_X1 U23785 ( .B1(n20835), .B2(keyinput111), .C1(n20834), .C2(
        keyinput102), .A(n20833), .ZN(n20838) );
  INV_X1 U23786 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20836) );
  XNOR2_X1 U23787 ( .A(n20836), .B(keyinput24), .ZN(n20837) );
  NOR2_X1 U23788 ( .A1(n20838), .A2(n20837), .ZN(n20849) );
  AOI22_X1 U23789 ( .A1(n14210), .A2(keyinput58), .B1(keyinput113), .B2(n20840), .ZN(n20839) );
  OAI221_X1 U23790 ( .B1(n14210), .B2(keyinput58), .C1(n20840), .C2(
        keyinput113), .A(n20839), .ZN(n20841) );
  INV_X1 U23791 ( .A(n20841), .ZN(n20848) );
  INV_X1 U23792 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20844) );
  INV_X1 U23793 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n20843) );
  AOI22_X1 U23794 ( .A1(n20844), .A2(keyinput28), .B1(keyinput6), .B2(n20843), 
        .ZN(n20842) );
  OAI221_X1 U23795 ( .B1(n20844), .B2(keyinput28), .C1(n20843), .C2(keyinput6), 
        .A(n20842), .ZN(n20845) );
  INV_X1 U23796 ( .A(n20845), .ZN(n20847) );
  XNOR2_X1 U23797 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B(keyinput106), .ZN(
        n20846) );
  AND4_X1 U23798 ( .A1(n20849), .A2(n20848), .A3(n20847), .A4(n20846), .ZN(
        n20883) );
  AOI22_X1 U23799 ( .A1(n20852), .A2(keyinput29), .B1(n20851), .B2(keyinput53), 
        .ZN(n20850) );
  OAI221_X1 U23800 ( .B1(n20852), .B2(keyinput29), .C1(n20851), .C2(keyinput53), .A(n20850), .ZN(n20864) );
  INV_X1 U23801 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n20855) );
  INV_X1 U23802 ( .A(keyinput89), .ZN(n20854) );
  AOI22_X1 U23803 ( .A1(n20855), .A2(keyinput0), .B1(
        P2_DATAWIDTH_REG_15__SCAN_IN), .B2(n20854), .ZN(n20853) );
  OAI221_X1 U23804 ( .B1(n20855), .B2(keyinput0), .C1(n20854), .C2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A(n20853), .ZN(n20863) );
  INV_X1 U23805 ( .A(keyinput40), .ZN(n20857) );
  AOI22_X1 U23806 ( .A1(n12673), .A2(keyinput37), .B1(
        P3_DATAWIDTH_REG_7__SCAN_IN), .B2(n20857), .ZN(n20856) );
  OAI221_X1 U23807 ( .B1(n12673), .B2(keyinput37), .C1(n20857), .C2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A(n20856), .ZN(n20862) );
  AOI22_X1 U23808 ( .A1(n20860), .A2(keyinput13), .B1(keyinput44), .B2(n20859), 
        .ZN(n20858) );
  OAI221_X1 U23809 ( .B1(n20860), .B2(keyinput13), .C1(n20859), .C2(keyinput44), .A(n20858), .ZN(n20861) );
  NOR4_X1 U23810 ( .A1(n20864), .A2(n20863), .A3(n20862), .A4(n20861), .ZN(
        n20882) );
  AOI22_X1 U23811 ( .A1(n20867), .A2(keyinput52), .B1(n20866), .B2(keyinput127), .ZN(n20865) );
  OAI221_X1 U23812 ( .B1(n20867), .B2(keyinput52), .C1(n20866), .C2(
        keyinput127), .A(n20865), .ZN(n20880) );
  INV_X1 U23813 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n20869) );
  AOI22_X1 U23814 ( .A1(n20870), .A2(keyinput2), .B1(keyinput109), .B2(n20869), 
        .ZN(n20868) );
  OAI221_X1 U23815 ( .B1(n20870), .B2(keyinput2), .C1(n20869), .C2(keyinput109), .A(n20868), .ZN(n20879) );
  INV_X1 U23816 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U23817 ( .A1(n20873), .A2(keyinput92), .B1(keyinput16), .B2(n20872), 
        .ZN(n20871) );
  OAI221_X1 U23818 ( .B1(n20873), .B2(keyinput92), .C1(n20872), .C2(keyinput16), .A(n20871), .ZN(n20878) );
  INV_X1 U23819 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n20876) );
  INV_X1 U23820 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n20875) );
  AOI22_X1 U23821 ( .A1(n20876), .A2(keyinput33), .B1(n20875), .B2(keyinput66), 
        .ZN(n20874) );
  OAI221_X1 U23822 ( .B1(n20876), .B2(keyinput33), .C1(n20875), .C2(keyinput66), .A(n20874), .ZN(n20877) );
  NOR4_X1 U23823 ( .A1(n20880), .A2(n20879), .A3(n20878), .A4(n20877), .ZN(
        n20881) );
  NAND4_X1 U23824 ( .A1(n20884), .A2(n20883), .A3(n20882), .A4(n20881), .ZN(
        n21082) );
  AOI22_X1 U23825 ( .A1(n13952), .A2(keyinput30), .B1(keyinput64), .B2(n20886), 
        .ZN(n20885) );
  OAI221_X1 U23826 ( .B1(n13952), .B2(keyinput30), .C1(n20886), .C2(keyinput64), .A(n20885), .ZN(n20898) );
  INV_X1 U23827 ( .A(DATAI_23_), .ZN(n20889) );
  AOI22_X1 U23828 ( .A1(n20889), .A2(keyinput45), .B1(keyinput86), .B2(n20888), 
        .ZN(n20887) );
  OAI221_X1 U23829 ( .B1(n20889), .B2(keyinput45), .C1(n20888), .C2(keyinput86), .A(n20887), .ZN(n20897) );
  INV_X1 U23830 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U23831 ( .A1(n20892), .A2(keyinput120), .B1(n20891), .B2(keyinput12), .ZN(n20890) );
  OAI221_X1 U23832 ( .B1(n20892), .B2(keyinput120), .C1(n20891), .C2(
        keyinput12), .A(n20890), .ZN(n20896) );
  INV_X1 U23833 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n20894) );
  AOI22_X1 U23834 ( .A1(n20894), .A2(keyinput124), .B1(n13708), .B2(keyinput41), .ZN(n20893) );
  OAI221_X1 U23835 ( .B1(n20894), .B2(keyinput124), .C1(n13708), .C2(
        keyinput41), .A(n20893), .ZN(n20895) );
  NOR4_X1 U23836 ( .A1(n20898), .A2(n20897), .A3(n20896), .A4(n20895), .ZN(
        n20951) );
  AOI22_X1 U23837 ( .A1(n20901), .A2(keyinput4), .B1(keyinput49), .B2(n20900), 
        .ZN(n20899) );
  OAI221_X1 U23838 ( .B1(n20901), .B2(keyinput4), .C1(n20900), .C2(keyinput49), 
        .A(n20899), .ZN(n20913) );
  AOI22_X1 U23839 ( .A1(n20904), .A2(keyinput119), .B1(n20903), .B2(keyinput93), .ZN(n20902) );
  OAI221_X1 U23840 ( .B1(n20904), .B2(keyinput119), .C1(n20903), .C2(
        keyinput93), .A(n20902), .ZN(n20912) );
  AOI22_X1 U23841 ( .A1(n20907), .A2(keyinput65), .B1(keyinput21), .B2(n20906), 
        .ZN(n20905) );
  OAI221_X1 U23842 ( .B1(n20907), .B2(keyinput65), .C1(n20906), .C2(keyinput21), .A(n20905), .ZN(n20911) );
  INV_X1 U23843 ( .A(keyinput10), .ZN(n20909) );
  AOI22_X1 U23844 ( .A1(n15975), .A2(keyinput112), .B1(
        P2_DATAWIDTH_REG_29__SCAN_IN), .B2(n20909), .ZN(n20908) );
  OAI221_X1 U23845 ( .B1(n15975), .B2(keyinput112), .C1(n20909), .C2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A(n20908), .ZN(n20910) );
  NOR4_X1 U23846 ( .A1(n20913), .A2(n20912), .A3(n20911), .A4(n20910), .ZN(
        n20950) );
  AOI22_X1 U23847 ( .A1(n20916), .A2(keyinput80), .B1(keyinput23), .B2(n20915), 
        .ZN(n20914) );
  OAI221_X1 U23848 ( .B1(n20916), .B2(keyinput80), .C1(n20915), .C2(keyinput23), .A(n20914), .ZN(n20919) );
  XNOR2_X1 U23849 ( .A(n20917), .B(keyinput123), .ZN(n20918) );
  NOR2_X1 U23850 ( .A1(n20919), .A2(n20918), .ZN(n20931) );
  INV_X1 U23851 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20921) );
  AOI22_X1 U23852 ( .A1(n20922), .A2(keyinput39), .B1(keyinput98), .B2(n20921), 
        .ZN(n20920) );
  OAI221_X1 U23853 ( .B1(n20922), .B2(keyinput39), .C1(n20921), .C2(keyinput98), .A(n20920), .ZN(n20923) );
  INV_X1 U23854 ( .A(n20923), .ZN(n20930) );
  INV_X1 U23855 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n20926) );
  AOI22_X1 U23856 ( .A1(n20926), .A2(keyinput3), .B1(keyinput95), .B2(n20925), 
        .ZN(n20924) );
  OAI221_X1 U23857 ( .B1(n20926), .B2(keyinput3), .C1(n20925), .C2(keyinput95), 
        .A(n20924), .ZN(n20927) );
  INV_X1 U23858 ( .A(n20927), .ZN(n20929) );
  XNOR2_X1 U23859 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B(keyinput74), .ZN(
        n20928) );
  AND4_X1 U23860 ( .A1(n20931), .A2(n20930), .A3(n20929), .A4(n20928), .ZN(
        n20949) );
  AOI22_X1 U23861 ( .A1(n20934), .A2(keyinput121), .B1(keyinput61), .B2(n20933), .ZN(n20932) );
  OAI221_X1 U23862 ( .B1(n20934), .B2(keyinput121), .C1(n20933), .C2(
        keyinput61), .A(n20932), .ZN(n20947) );
  AOI22_X1 U23863 ( .A1(n20937), .A2(keyinput11), .B1(keyinput78), .B2(n20936), 
        .ZN(n20935) );
  OAI221_X1 U23864 ( .B1(n20937), .B2(keyinput11), .C1(n20936), .C2(keyinput78), .A(n20935), .ZN(n20946) );
  INV_X1 U23865 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20940) );
  INV_X1 U23866 ( .A(keyinput67), .ZN(n20939) );
  AOI22_X1 U23867 ( .A1(n20940), .A2(keyinput84), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n20939), .ZN(n20938) );
  OAI221_X1 U23868 ( .B1(n20940), .B2(keyinput84), .C1(n20939), .C2(
        P3_ADDRESS_REG_29__SCAN_IN), .A(n20938), .ZN(n20945) );
  INV_X1 U23869 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U23870 ( .A1(n20943), .A2(keyinput99), .B1(n20942), .B2(keyinput59), 
        .ZN(n20941) );
  OAI221_X1 U23871 ( .B1(n20943), .B2(keyinput99), .C1(n20942), .C2(keyinput59), .A(n20941), .ZN(n20944) );
  NOR4_X1 U23872 ( .A1(n20947), .A2(n20946), .A3(n20945), .A4(n20944), .ZN(
        n20948) );
  NAND4_X1 U23873 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n21081) );
  AOI22_X1 U23874 ( .A1(n20954), .A2(keyinput47), .B1(keyinput97), .B2(n20953), 
        .ZN(n20952) );
  OAI221_X1 U23875 ( .B1(n20954), .B2(keyinput47), .C1(n20953), .C2(keyinput97), .A(n20952), .ZN(n20967) );
  INV_X1 U23876 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20957) );
  AOI22_X1 U23877 ( .A1(n20957), .A2(keyinput18), .B1(keyinput94), .B2(n20956), 
        .ZN(n20955) );
  OAI221_X1 U23878 ( .B1(n20957), .B2(keyinput18), .C1(n20956), .C2(keyinput94), .A(n20955), .ZN(n20966) );
  INV_X1 U23879 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20960) );
  INV_X1 U23880 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n20959) );
  AOI22_X1 U23881 ( .A1(n20960), .A2(keyinput96), .B1(keyinput88), .B2(n20959), 
        .ZN(n20958) );
  OAI221_X1 U23882 ( .B1(n20960), .B2(keyinput96), .C1(n20959), .C2(keyinput88), .A(n20958), .ZN(n20965) );
  INV_X1 U23883 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20963) );
  INV_X1 U23884 ( .A(keyinput42), .ZN(n20962) );
  AOI22_X1 U23885 ( .A1(n20963), .A2(keyinput101), .B1(
        P3_BYTEENABLE_REG_0__SCAN_IN), .B2(n20962), .ZN(n20961) );
  OAI221_X1 U23886 ( .B1(n20963), .B2(keyinput101), .C1(n20962), .C2(
        P3_BYTEENABLE_REG_0__SCAN_IN), .A(n20961), .ZN(n20964) );
  NOR4_X1 U23887 ( .A1(n20967), .A2(n20966), .A3(n20965), .A4(n20964), .ZN(
        n21016) );
  AOI22_X1 U23888 ( .A1(n20970), .A2(keyinput34), .B1(n20969), .B2(keyinput5), 
        .ZN(n20968) );
  OAI221_X1 U23889 ( .B1(n20970), .B2(keyinput34), .C1(n20969), .C2(keyinput5), 
        .A(n20968), .ZN(n20982) );
  AOI22_X1 U23890 ( .A1(n20972), .A2(keyinput105), .B1(n13403), .B2(keyinput35), .ZN(n20971) );
  OAI221_X1 U23891 ( .B1(n20972), .B2(keyinput105), .C1(n13403), .C2(
        keyinput35), .A(n20971), .ZN(n20981) );
  INV_X1 U23892 ( .A(P3_UWORD_REG_13__SCAN_IN), .ZN(n20974) );
  AOI22_X1 U23893 ( .A1(n20975), .A2(keyinput118), .B1(keyinput87), .B2(n20974), .ZN(n20973) );
  OAI221_X1 U23894 ( .B1(n20975), .B2(keyinput118), .C1(n20974), .C2(
        keyinput87), .A(n20973), .ZN(n20980) );
  INV_X1 U23895 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n20978) );
  AOI22_X1 U23896 ( .A1(n20978), .A2(keyinput57), .B1(keyinput83), .B2(n20977), 
        .ZN(n20976) );
  OAI221_X1 U23897 ( .B1(n20978), .B2(keyinput57), .C1(n20977), .C2(keyinput83), .A(n20976), .ZN(n20979) );
  NOR4_X1 U23898 ( .A1(n20982), .A2(n20981), .A3(n20980), .A4(n20979), .ZN(
        n21015) );
  AOI22_X1 U23899 ( .A1(n20985), .A2(keyinput63), .B1(n20984), .B2(keyinput103), .ZN(n20983) );
  OAI221_X1 U23900 ( .B1(n20985), .B2(keyinput63), .C1(n20984), .C2(
        keyinput103), .A(n20983), .ZN(n20997) );
  AOI22_X1 U23901 ( .A1(n20987), .A2(keyinput36), .B1(keyinput75), .B2(n12709), 
        .ZN(n20986) );
  OAI221_X1 U23902 ( .B1(n20987), .B2(keyinput36), .C1(n12709), .C2(keyinput75), .A(n20986), .ZN(n20996) );
  AOI22_X1 U23903 ( .A1(n20990), .A2(keyinput81), .B1(n20989), .B2(keyinput56), 
        .ZN(n20988) );
  OAI221_X1 U23904 ( .B1(n20990), .B2(keyinput81), .C1(n20989), .C2(keyinput56), .A(n20988), .ZN(n20995) );
  INV_X1 U23905 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20993) );
  INV_X1 U23906 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U23907 ( .A1(n20993), .A2(keyinput51), .B1(n20992), .B2(keyinput17), 
        .ZN(n20991) );
  OAI221_X1 U23908 ( .B1(n20993), .B2(keyinput51), .C1(n20992), .C2(keyinput17), .A(n20991), .ZN(n20994) );
  NOR4_X1 U23909 ( .A1(n20997), .A2(n20996), .A3(n20995), .A4(n20994), .ZN(
        n21014) );
  AOI22_X1 U23910 ( .A1(n21000), .A2(keyinput79), .B1(keyinput114), .B2(n20999), .ZN(n20998) );
  OAI221_X1 U23911 ( .B1(n21000), .B2(keyinput79), .C1(n20999), .C2(
        keyinput114), .A(n20998), .ZN(n21012) );
  AOI22_X1 U23912 ( .A1(n21003), .A2(keyinput15), .B1(keyinput117), .B2(n21002), .ZN(n21001) );
  OAI221_X1 U23913 ( .B1(n21003), .B2(keyinput15), .C1(n21002), .C2(
        keyinput117), .A(n21001), .ZN(n21011) );
  INV_X1 U23914 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n21005) );
  AOI22_X1 U23915 ( .A1(n21006), .A2(keyinput27), .B1(keyinput100), .B2(n21005), .ZN(n21004) );
  OAI221_X1 U23916 ( .B1(n21006), .B2(keyinput27), .C1(n21005), .C2(
        keyinput100), .A(n21004), .ZN(n21010) );
  INV_X1 U23917 ( .A(P3_LWORD_REG_7__SCAN_IN), .ZN(n21008) );
  AOI22_X1 U23918 ( .A1(n14628), .A2(keyinput25), .B1(keyinput32), .B2(n21008), 
        .ZN(n21007) );
  OAI221_X1 U23919 ( .B1(n14628), .B2(keyinput25), .C1(n21008), .C2(keyinput32), .A(n21007), .ZN(n21009) );
  NOR4_X1 U23920 ( .A1(n21012), .A2(n21011), .A3(n21010), .A4(n21009), .ZN(
        n21013) );
  NAND4_X1 U23921 ( .A1(n21016), .A2(n21015), .A3(n21014), .A4(n21013), .ZN(
        n21080) );
  INV_X1 U23922 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21019) );
  AOI22_X1 U23923 ( .A1(n21019), .A2(keyinput116), .B1(keyinput54), .B2(n21018), .ZN(n21017) );
  OAI221_X1 U23924 ( .B1(n21019), .B2(keyinput116), .C1(n21018), .C2(
        keyinput54), .A(n21017), .ZN(n21032) );
  AOI22_X1 U23925 ( .A1(n21022), .A2(keyinput115), .B1(keyinput26), .B2(n21021), .ZN(n21020) );
  OAI221_X1 U23926 ( .B1(n21022), .B2(keyinput115), .C1(n21021), .C2(
        keyinput26), .A(n21020), .ZN(n21031) );
  INV_X1 U23927 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n21025) );
  INV_X1 U23928 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n21024) );
  AOI22_X1 U23929 ( .A1(n21025), .A2(keyinput90), .B1(n21024), .B2(keyinput31), 
        .ZN(n21023) );
  OAI221_X1 U23930 ( .B1(n21025), .B2(keyinput90), .C1(n21024), .C2(keyinput31), .A(n21023), .ZN(n21030) );
  AOI22_X1 U23931 ( .A1(n21028), .A2(keyinput91), .B1(n21027), .B2(keyinput108), .ZN(n21026) );
  OAI221_X1 U23932 ( .B1(n21028), .B2(keyinput91), .C1(n21027), .C2(
        keyinput108), .A(n21026), .ZN(n21029) );
  NOR4_X1 U23933 ( .A1(n21032), .A2(n21031), .A3(n21030), .A4(n21029), .ZN(
        n21078) );
  XOR2_X1 U23934 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput8), .Z(
        n21033) );
  AOI21_X1 U23935 ( .B1(n21085), .B2(keyinput126), .A(n21033), .ZN(n21036) );
  XNOR2_X1 U23936 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput110), 
        .ZN(n21035) );
  XNOR2_X1 U23937 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(keyinput69), 
        .ZN(n21034) );
  NAND3_X1 U23938 ( .A1(n21036), .A2(n21035), .A3(n21034), .ZN(n21045) );
  INV_X1 U23939 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n21039) );
  AOI22_X1 U23940 ( .A1(n21039), .A2(keyinput9), .B1(n21038), .B2(keyinput82), 
        .ZN(n21037) );
  OAI221_X1 U23941 ( .B1(n21039), .B2(keyinput9), .C1(n21038), .C2(keyinput82), 
        .A(n21037), .ZN(n21044) );
  INV_X1 U23942 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n21041) );
  AOI22_X1 U23943 ( .A1(n21042), .A2(keyinput43), .B1(keyinput72), .B2(n21041), 
        .ZN(n21040) );
  OAI221_X1 U23944 ( .B1(n21042), .B2(keyinput43), .C1(n21041), .C2(keyinput72), .A(n21040), .ZN(n21043) );
  NOR3_X1 U23945 ( .A1(n21045), .A2(n21044), .A3(n21043), .ZN(n21077) );
  INV_X1 U23946 ( .A(DATAI_17_), .ZN(n21048) );
  INV_X1 U23947 ( .A(keyinput76), .ZN(n21047) );
  AOI22_X1 U23948 ( .A1(n21048), .A2(keyinput122), .B1(P2_D_C_N_REG_SCAN_IN), 
        .B2(n21047), .ZN(n21046) );
  OAI221_X1 U23949 ( .B1(n21048), .B2(keyinput122), .C1(n21047), .C2(
        P2_D_C_N_REG_SCAN_IN), .A(n21046), .ZN(n21060) );
  INV_X1 U23950 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n21051) );
  AOI22_X1 U23951 ( .A1(n21051), .A2(keyinput1), .B1(keyinput104), .B2(n21050), 
        .ZN(n21049) );
  OAI221_X1 U23952 ( .B1(n21051), .B2(keyinput1), .C1(n21050), .C2(keyinput104), .A(n21049), .ZN(n21059) );
  INV_X1 U23953 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21053) );
  AOI22_X1 U23954 ( .A1(n13728), .A2(keyinput125), .B1(n21053), .B2(keyinput38), .ZN(n21052) );
  OAI221_X1 U23955 ( .B1(n13728), .B2(keyinput125), .C1(n21053), .C2(
        keyinput38), .A(n21052), .ZN(n21058) );
  INV_X1 U23956 ( .A(keyinput77), .ZN(n21055) );
  AOI22_X1 U23957 ( .A1(n21056), .A2(keyinput20), .B1(
        P2_DATAWIDTH_REG_19__SCAN_IN), .B2(n21055), .ZN(n21054) );
  OAI221_X1 U23958 ( .B1(n21056), .B2(keyinput20), .C1(n21055), .C2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A(n21054), .ZN(n21057) );
  NOR4_X1 U23959 ( .A1(n21060), .A2(n21059), .A3(n21058), .A4(n21057), .ZN(
        n21076) );
  AOI22_X1 U23960 ( .A1(n21063), .A2(keyinput48), .B1(keyinput60), .B2(n21062), 
        .ZN(n21061) );
  OAI221_X1 U23961 ( .B1(n21063), .B2(keyinput48), .C1(n21062), .C2(keyinput60), .A(n21061), .ZN(n21074) );
  INV_X1 U23962 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n21065) );
  AOI22_X1 U23963 ( .A1(n21065), .A2(keyinput107), .B1(n12721), .B2(keyinput50), .ZN(n21064) );
  OAI221_X1 U23964 ( .B1(n21065), .B2(keyinput107), .C1(n12721), .C2(
        keyinput50), .A(n21064), .ZN(n21073) );
  INV_X1 U23965 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21067) );
  AOI22_X1 U23966 ( .A1(n21068), .A2(keyinput85), .B1(keyinput7), .B2(n21067), 
        .ZN(n21066) );
  OAI221_X1 U23967 ( .B1(n21068), .B2(keyinput85), .C1(n21067), .C2(keyinput7), 
        .A(n21066), .ZN(n21072) );
  AOI22_X1 U23968 ( .A1(n21070), .A2(keyinput73), .B1(keyinput46), .B2(n10344), 
        .ZN(n21069) );
  OAI221_X1 U23969 ( .B1(n21070), .B2(keyinput73), .C1(n10344), .C2(keyinput46), .A(n21069), .ZN(n21071) );
  NOR4_X1 U23970 ( .A1(n21074), .A2(n21073), .A3(n21072), .A4(n21071), .ZN(
        n21075) );
  NAND4_X1 U23971 ( .A1(n21078), .A2(n21077), .A3(n21076), .A4(n21075), .ZN(
        n21079) );
  NOR4_X1 U23972 ( .A1(n21082), .A2(n21081), .A3(n21080), .A4(n21079), .ZN(
        n21083) );
  OAI221_X1 U23973 ( .B1(n21085), .B2(keyinput126), .C1(n21085), .C2(n21084), 
        .A(n21083), .ZN(n21086) );
  XOR2_X1 U23974 ( .A(n21087), .B(n21086), .Z(P2_U3211) );
  AND2_X1 U11876 ( .A1(n13217), .A2(n11673), .ZN(n11759) );
  INV_X2 U11189 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18933) );
  NAND2_X2 U13156 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10244), .ZN(
        n17275) );
  AND2_X1 U13723 ( .A1(n10756), .A2(n10747), .ZN(n10749) );
  INV_X2 U11311 ( .A(n19206), .ZN(n19190) );
  NOR2_X1 U12872 ( .A1(n11666), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11673) );
  AND2_X2 U11287 ( .A1(n11672), .A2(n13217), .ZN(n11845) );
  CLKBUF_X1 U11224 ( .A(n11630), .Z(n9764) );
  CLKBUF_X1 U11235 ( .A(n18803), .Z(n9773) );
  CLKBUF_X1 U11241 ( .A(n17619), .Z(n17626) );
  CLKBUF_X1 U11272 ( .A(n18917), .Z(n18910) );
  CLKBUF_X1 U11273 ( .A(n16630), .Z(n16638) );
  AND3_X1 U11290 ( .A1(n10276), .A2(n10275), .A3(n10274), .ZN(n21088) );
  CLKBUF_X1 U11572 ( .A(n11845), .Z(n14283) );
endmodule

