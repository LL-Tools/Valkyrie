

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356;

  NOR2_X1 U2523 ( .A1(n4578), .A2(n4579), .ZN(n4577) );
  CLKBUF_X2 U2525 ( .A(n3043), .Z(n2493) );
  NAND2_X1 U2526 ( .A1(n2934), .A2(n2933), .ZN(n3099) );
  NAND2_X1 U2527 ( .A1(n2788), .A2(n2787), .ZN(n5183) );
  AND2_X1 U2528 ( .A1(n4952), .A2(n4959), .ZN(n2579) );
  INV_X1 U2529 ( .A(IR_REG_18__SCAN_IN), .ZN(n4981) );
  BUF_X1 U2530 ( .A(n3128), .Z(n3875) );
  INV_X1 U2531 ( .A(n3810), .ZN(n3873) );
  BUF_X1 U2532 ( .A(n2957), .Z(n2956) );
  INV_X1 U2533 ( .A(n3240), .ZN(n3216) );
  INV_X1 U2534 ( .A(n3099), .ZN(n2980) );
  AND2_X1 U2535 ( .A1(n2738), .A2(n2737), .ZN(n2758) );
  INV_X2 U2536 ( .A(n3128), .ZN(n2499) );
  NAND2_X1 U2537 ( .A1(n4488), .A2(n4489), .ZN(n4491) );
  INV_X1 U2538 ( .A(IR_REG_20__SCAN_IN), .ZN(n4985) );
  MUX2_X1 U2539 ( .A(n5167), .B(DATAI_0_), .S(n4162), .Z(n3094) );
  AND2_X1 U2540 ( .A1(n2777), .A2(n2864), .ZN(n4671) );
  CLKBUF_X3 U2541 ( .A(n4162), .Z(n2488) );
  NAND2_X2 U2542 ( .A1(n2794), .A2(n5183), .ZN(n4162) );
  AOI21_X2 U2543 ( .B1(n3937), .B2(n4501), .A(n3936), .ZN(n4588) );
  OAI21_X2 U2544 ( .B1(n5202), .B2(n2626), .A(n2625), .ZN(n5119) );
  NAND2_X2 U2545 ( .A1(n2692), .A2(n2693), .ZN(n5202) );
  XNOR2_X2 U2546 ( .A(n2725), .B(n2724), .ZN(n3409) );
  INV_X1 U2547 ( .A(n3872), .ZN(n2489) );
  AND2_X2 U2548 ( .A1(n2959), .A2(n2956), .ZN(n3044) );
  INV_X1 U2549 ( .A(n2976), .ZN(n2490) );
  INV_X1 U2550 ( .A(n2976), .ZN(n2491) );
  AND2_X2 U2551 ( .A1(n2959), .A2(n2958), .ZN(n2976) );
  OR2_X2 U2553 ( .A1(n3035), .A2(n3036), .ZN(n3117) );
  NOR2_X2 U2555 ( .A1(n5160), .A2(n2745), .ZN(n2847) );
  XNOR2_X2 U2556 ( .A(n2901), .B(n4985), .ZN(n2923) );
  NAND2_X2 U2557 ( .A1(n2900), .A2(n2899), .ZN(n2901) );
  INV_X1 U2558 ( .A(n2896), .ZN(n2898) );
  AND2_X1 U2559 ( .A1(n2896), .A2(n4669), .ZN(n3006) );
  XNOR2_X2 U2560 ( .A(n2867), .B(n4804), .ZN(n2896) );
  AOI21_X2 U2561 ( .B1(REG2_REG_15__SCAN_IN), .B2(n5150), .A(n5146), .ZN(n2741) );
  OAI21_X1 U2562 ( .B1(n2642), .B2(n2640), .A(n3857), .ZN(n2639) );
  INV_X1 U2563 ( .A(n2642), .ZN(n2641) );
  NOR2_X1 U2564 ( .A1(n3493), .A2(n2607), .ZN(n2730) );
  OR2_X1 U2565 ( .A1(n3577), .A2(n3576), .ZN(n3581) );
  AND2_X1 U2566 ( .A1(n2657), .A2(n3575), .ZN(n3576) );
  OR2_X1 U2567 ( .A1(n3547), .A2(n3546), .ZN(n3575) );
  NAND2_X2 U2568 ( .A1(n3221), .A2(n3222), .ZN(n3058) );
  OR2_X1 U2569 ( .A1(n3543), .A2(n5290), .ZN(n3544) );
  NAND2_X2 U2570 ( .A1(n3016), .A2(n5307), .ZN(n5282) );
  NAND2_X1 U2571 ( .A1(n3104), .A2(n4158), .ZN(n3248) );
  AND2_X2 U2572 ( .A1(n3005), .A2(n3004), .ZN(n5296) );
  NOR2_X1 U2573 ( .A1(n3368), .A2(n3363), .ZN(n3254) );
  INV_X1 U2574 ( .A(n2493), .ZN(n3831) );
  INV_X1 U2575 ( .A(n4251), .ZN(n3206) );
  NAND2_X1 U2576 ( .A1(n4079), .A2(n4082), .ZN(n3024) );
  NAND4_X1 U2577 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n4248)
         );
  NAND4_X1 U2578 ( .A1(n3011), .A2(n3010), .A3(n3009), .A4(n3008), .ZN(n4251)
         );
  NAND4_X1 U2579 ( .A1(n3050), .A2(n3049), .A3(n3048), .A4(n3047), .ZN(n4250)
         );
  INV_X1 U2580 ( .A(n2495), .ZN(n2496) );
  INV_X2 U2581 ( .A(n2495), .ZN(n2497) );
  INV_X1 U2582 ( .A(n5211), .ZN(n4674) );
  INV_X1 U2583 ( .A(n3006), .ZN(n2495) );
  NAND2_X1 U2584 ( .A1(n2754), .A2(n2900), .ZN(n5211) );
  INV_X4 U2585 ( .A(n3156), .ZN(n3353) );
  MUX2_X1 U2586 ( .A(n2899), .B(n2769), .S(IR_REG_25__SCAN_IN), .Z(n2771) );
  NAND2_X1 U2587 ( .A1(n2895), .A2(n2894), .ZN(n2897) );
  NAND2_X1 U2588 ( .A1(n2762), .A2(n2899), .ZN(n2739) );
  NOR2_X2 U2589 ( .A1(n2647), .A2(n2646), .ZN(n2645) );
  NAND4_X2 U2590 ( .A1(n2579), .A2(n2659), .A3(n2658), .A4(n2677), .ZN(n2703)
         );
  INV_X2 U2591 ( .A(n2663), .ZN(n2899) );
  INV_X1 U2592 ( .A(IR_REG_8__SCAN_IN), .ZN(n4963) );
  INV_X1 U2593 ( .A(IR_REG_19__SCAN_IN), .ZN(n2759) );
  INV_X1 U2594 ( .A(IR_REG_5__SCAN_IN), .ZN(n4959) );
  INV_X1 U2595 ( .A(IR_REG_7__SCAN_IN), .ZN(n2709) );
  INV_X1 U2596 ( .A(IR_REG_2__SCAN_IN), .ZN(n4952) );
  NOR2_X2 U2597 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2677)
         );
  CLKBUF_X1 U2598 ( .A(IR_REG_0__SCAN_IN), .Z(n5167) );
  CLKBUF_X1 U2599 ( .A(n3043), .Z(n2492) );
  NAND2_X1 U2600 ( .A1(n3044), .A2(n3292), .ZN(n3043) );
  NAND2_X1 U2601 ( .A1(n4443), .A2(n3939), .ZN(n4446) );
  NOR2_X4 U2602 ( .A1(n3422), .A2(n4111), .ZN(n3532) );
  AOI21_X1 U2603 ( .B1(n2494), .B2(n4252), .A(n2963), .ZN(n2966) );
  NAND4_X2 U2604 ( .A1(n2946), .A2(n2945), .A3(n2944), .A4(n2943), .ZN(n4252)
         );
  AOI21_X2 U2605 ( .B1(n3628), .B2(n3627), .A(n3626), .ZN(n3707) );
  INV_X1 U2606 ( .A(n2492), .ZN(n2494) );
  NOR2_X2 U2607 ( .A1(n4446), .A2(n4418), .ZN(n4403) );
  NOR2_X2 U2608 ( .A1(n4526), .A2(n3938), .ZN(n4509) );
  INV_X1 U2610 ( .A(n3128), .ZN(n2498) );
  INV_X2 U2611 ( .A(n2976), .ZN(n3128) );
  NOR2_X2 U2612 ( .A1(n3833), .A2(n3832), .ZN(n4002) );
  AND2_X1 U2613 ( .A1(n2670), .A2(n2513), .ZN(n2570) );
  AOI21_X1 U2614 ( .B1(n2549), .B2(n2547), .A(n2517), .ZN(n2546) );
  INV_X1 U2615 ( .A(n2551), .ZN(n2547) );
  AND2_X1 U2616 ( .A1(n2541), .A2(n2528), .ZN(n2533) );
  NAND2_X1 U2617 ( .A1(n2628), .A2(n2631), .ZN(n3984) );
  AND2_X1 U2618 ( .A1(n2632), .A2(n4023), .ZN(n2631) );
  NAND2_X1 U2619 ( .A1(n4024), .A2(n2633), .ZN(n2632) );
  INV_X1 U2620 ( .A(n4034), .ZN(n3796) );
  INV_X1 U2621 ( .A(n3007), .ZN(n3836) );
  XNOR2_X1 U2622 ( .A(n2805), .B(n5206), .ZN(n5199) );
  NAND2_X1 U2623 ( .A1(n2622), .A2(n2621), .ZN(n2620) );
  AND2_X1 U2624 ( .A1(n2624), .A2(REG2_REG_8__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U2625 ( .A1(n3903), .A2(n3902), .ZN(n3904) );
  OAI22_X1 U2626 ( .A1(n4376), .A2(n2558), .B1(n4399), .B2(n4378), .ZN(n2557)
         );
  NAND2_X1 U2627 ( .A1(n4181), .A2(n4180), .ZN(n2558) );
  INV_X1 U2628 ( .A(n2541), .ZN(n2538) );
  MUX2_X1 U2629 ( .A(n2899), .B(n2893), .S(IR_REG_29__SCAN_IN), .Z(n2895) );
  OR2_X1 U2630 ( .A1(n3585), .A2(n3584), .ZN(n3586) );
  INV_X1 U2631 ( .A(n2679), .ZN(n2616) );
  NOR2_X1 U2632 ( .A1(n3232), .A2(n2814), .ZN(n2815) );
  NOR2_X1 U2633 ( .A1(n2720), .A2(n2813), .ZN(n2814) );
  AND2_X1 U2634 ( .A1(n4676), .A2(REG2_REG_11__SCAN_IN), .ZN(n2607) );
  AND2_X1 U2635 ( .A1(n4324), .A2(n3909), .ZN(n4206) );
  OR2_X1 U2636 ( .A1(n4433), .A2(n4425), .ZN(n4395) );
  INV_X1 U2637 ( .A(n3243), .ZN(n2529) );
  OAI22_X1 U2638 ( .A1(n2536), .A2(n2506), .B1(n3276), .B2(n3275), .ZN(n2532)
         );
  AND2_X1 U2639 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n3061) );
  AND2_X1 U2640 ( .A1(n4114), .A2(n4103), .ZN(n4159) );
  NAND2_X1 U2641 ( .A1(n3022), .A2(n3036), .ZN(n4079) );
  AND4_X1 U2642 ( .A1(n2775), .A2(n2774), .A3(n2763), .A4(n2779), .ZN(n2776)
         );
  INV_X1 U2643 ( .A(IR_REG_23__SCAN_IN), .ZN(n2779) );
  INV_X1 U2644 ( .A(IR_REG_6__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U2645 ( .A1(n3855), .A2(n2643), .ZN(n2642) );
  OR2_X1 U2646 ( .A1(n4066), .A2(n3856), .ZN(n3855) );
  NAND2_X1 U2647 ( .A1(n3150), .A2(REG3_REG_22__SCAN_IN), .ZN(n3801) );
  AND4_X2 U2648 ( .A1(n2910), .A2(n2909), .A3(n2908), .A4(n2907), .ZN(n2971)
         );
  NOR2_X1 U2649 ( .A1(n2874), .A2(n2870), .ZN(n2778) );
  NAND2_X1 U2650 ( .A1(n2864), .A2(n2899), .ZN(n2786) );
  NAND2_X1 U2651 ( .A1(n2786), .A2(n2785), .ZN(n2788) );
  NOR2_X1 U2652 ( .A1(n5112), .A2(n5111), .ZN(n5110) );
  AOI22_X1 U2653 ( .A1(n2800), .A2(n5227), .B1(REG2_REG_2__SCAN_IN), .B2(n5180), .ZN(n5171) );
  NOR2_X1 U2654 ( .A1(n5174), .A2(n2648), .ZN(n2803) );
  NAND2_X1 U2655 ( .A1(n5075), .A2(n2616), .ZN(n2615) );
  OR2_X1 U2656 ( .A1(n2680), .A2(n2617), .ZN(n2613) );
  NAND2_X1 U2657 ( .A1(n2680), .A2(n2614), .ZN(n2610) );
  NOR2_X1 U2658 ( .A1(n5075), .A2(n2616), .ZN(n2614) );
  NAND2_X1 U2659 ( .A1(n2627), .A2(REG2_REG_4__SCAN_IN), .ZN(n2626) );
  INV_X1 U2660 ( .A(n5120), .ZN(n2627) );
  AND2_X1 U2661 ( .A1(n5126), .A2(REG1_REG_5__SCAN_IN), .ZN(n2807) );
  NOR2_X1 U2662 ( .A1(n5119), .A2(n2701), .ZN(n2705) );
  AND2_X1 U2663 ( .A1(n5126), .A2(REG2_REG_5__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U2664 ( .A1(n5138), .A2(n2650), .ZN(n2812) );
  NAND2_X1 U2665 ( .A1(n2620), .A2(n2619), .ZN(n2725) );
  AND2_X1 U2666 ( .A1(n2623), .A2(n2519), .ZN(n2619) );
  NOR2_X1 U2667 ( .A1(n3487), .A2(n2582), .ZN(n2817) );
  AND2_X1 U2668 ( .A1(n4676), .A2(REG1_REG_11__SCAN_IN), .ZN(n2582) );
  NOR2_X1 U2669 ( .A1(n3673), .A2(n3674), .ZN(n3672) );
  INV_X1 U2670 ( .A(n2834), .ZN(n2592) );
  OAI21_X1 U2671 ( .B1(n5153), .B2(n2589), .A(n2586), .ZN(n2585) );
  INV_X1 U2672 ( .A(n2587), .ZN(n2586) );
  OAI21_X1 U2673 ( .B1(n2589), .B2(n2591), .A(n2588), .ZN(n2587) );
  NAND2_X1 U2674 ( .A1(n2592), .A2(n2590), .ZN(n2588) );
  NOR2_X1 U2675 ( .A1(n4376), .A2(n2560), .ZN(n2559) );
  INV_X1 U2676 ( .A(n4373), .ZN(n4376) );
  OR2_X1 U2677 ( .A1(n3801), .A2(n3800), .ZN(n3818) );
  AOI21_X1 U2678 ( .B1(n2546), .B2(n2548), .A(n2518), .ZN(n2544) );
  AND2_X1 U2679 ( .A1(n2514), .A2(n3900), .ZN(n2551) );
  NAND2_X1 U2680 ( .A1(n2550), .A2(n2514), .ZN(n2549) );
  OR2_X1 U2681 ( .A1(n4465), .A2(n4481), .ZN(n3900) );
  NAND2_X1 U2682 ( .A1(n3148), .A2(REG3_REG_19__SCAN_IN), .ZN(n3752) );
  NOR2_X1 U2683 ( .A1(n3638), .A2(n3719), .ZN(n3714) );
  INV_X1 U2684 ( .A(n4465), .ZN(n4508) );
  NAND2_X1 U2685 ( .A1(n3898), .A2(n3897), .ZN(n3899) );
  INV_X1 U2686 ( .A(n4505), .ZN(n3898) );
  INV_X1 U2687 ( .A(n5295), .ZN(n4549) );
  AOI21_X1 U2688 ( .B1(n2567), .B2(n2565), .A(n2503), .ZN(n2563) );
  INV_X1 U2689 ( .A(n3242), .ZN(n2537) );
  AND2_X1 U2690 ( .A1(n3243), .A2(n2506), .ZN(n2539) );
  INV_X1 U2691 ( .A(n4249), .ZN(n4058) );
  NOR2_X1 U2692 ( .A1(n3244), .A2(n2542), .ZN(n2541) );
  INV_X1 U2693 ( .A(n3241), .ZN(n2542) );
  OR2_X1 U2694 ( .A1(n5338), .A2(n5211), .ZN(n3013) );
  INV_X1 U2695 ( .A(n3947), .ZN(n4330) );
  OR2_X1 U2696 ( .A1(n3810), .A2(n2904), .ZN(n5272) );
  AND2_X1 U2697 ( .A1(n3021), .A2(n3020), .ZN(n3025) );
  AND2_X1 U2698 ( .A1(n2891), .A2(n4167), .ZN(n2947) );
  OAI21_X1 U2699 ( .B1(n2993), .B2(D_REG_0__SCAN_IN), .A(n2926), .ZN(n3201) );
  XNOR2_X1 U2700 ( .A(n2784), .B(n5001), .ZN(n2794) );
  NAND2_X1 U2701 ( .A1(n2788), .A2(n2899), .ZN(n2784) );
  OR2_X1 U2702 ( .A1(n2733), .A2(IR_REG_14__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U2703 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2674)
         );
  INV_X1 U2704 ( .A(n3986), .ZN(n3779) );
  NAND2_X1 U2705 ( .A1(n3825), .A2(n3824), .ZN(n4399) );
  OR2_X1 U2706 ( .A1(n4385), .A2(n3836), .ZN(n3825) );
  XNOR2_X1 U2707 ( .A(n2812), .B(n4678), .ZN(n3084) );
  XNOR2_X1 U2708 ( .A(n2824), .B(n2823), .ZN(n4280) );
  NAND2_X1 U2709 ( .A1(n5153), .A2(n2591), .ZN(n2844) );
  OAI21_X1 U2710 ( .B1(n4312), .B2(n4210), .A(n4578), .ZN(n4586) );
  XNOR2_X1 U2711 ( .A(n3910), .B(n4138), .ZN(n4589) );
  NAND2_X1 U2712 ( .A1(n2574), .A2(n2572), .ZN(n3910) );
  INV_X1 U2713 ( .A(n2573), .ZN(n2572) );
  AND3_X1 U2714 ( .A1(n4434), .A2(n4395), .A3(n4176), .ZN(n4202) );
  AND3_X1 U2715 ( .A1(n4461), .A2(n3912), .A3(n3916), .ZN(n4197) );
  INV_X1 U2716 ( .A(n3975), .ZN(n3379) );
  INV_X1 U2717 ( .A(n3751), .ZN(n2633) );
  NOR2_X1 U2718 ( .A1(n2634), .A2(n2630), .ZN(n2629) );
  INV_X1 U2719 ( .A(n4024), .ZN(n2634) );
  INV_X1 U2720 ( .A(n3964), .ZN(n2630) );
  INV_X1 U2721 ( .A(n3230), .ZN(n2624) );
  NOR2_X1 U2722 ( .A1(n4265), .A2(n2603), .ZN(n2734) );
  AND2_X1 U2723 ( .A1(n4675), .A2(REG2_REG_13__SCAN_IN), .ZN(n2603) );
  INV_X1 U2724 ( .A(n2833), .ZN(n2590) );
  OR2_X1 U2725 ( .A1(n2592), .A2(n2590), .ZN(n2589) );
  OR2_X1 U2726 ( .A1(n4399), .A2(n4386), .ZN(n3924) );
  INV_X1 U2727 ( .A(n2549), .ZN(n2548) );
  AND2_X1 U2728 ( .A1(n2502), .A2(n2565), .ZN(n2564) );
  NAND2_X1 U2729 ( .A1(n2568), .A2(n2515), .ZN(n2567) );
  NAND2_X1 U2730 ( .A1(n2569), .A2(n3651), .ZN(n2568) );
  INV_X1 U2731 ( .A(n3611), .ZN(n2569) );
  INV_X1 U2732 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3481) );
  INV_X1 U2733 ( .A(n4378), .ZN(n4386) );
  NOR2_X2 U2734 ( .A1(n4491), .A2(n4464), .ZN(n4443) );
  INV_X1 U2735 ( .A(n4481), .ZN(n4489) );
  INV_X1 U2736 ( .A(n4503), .ZN(n4510) );
  BUF_X1 U2737 ( .A(n4509), .Z(n4527) );
  AOI21_X1 U2738 ( .B1(n3609), .B2(n2502), .A(n2567), .ZN(n3680) );
  NOR2_X2 U2739 ( .A1(n3605), .A2(n5281), .ZN(n3648) );
  INV_X1 U2740 ( .A(n3094), .ZN(n2953) );
  AND4_X1 U2741 ( .A1(n2938), .A2(n2935), .A3(n2936), .A4(n2937), .ZN(n2981)
         );
  INV_X1 U2742 ( .A(IR_REG_21__SCAN_IN), .ZN(n4989) );
  INV_X1 U2743 ( .A(n2662), .ZN(n2646) );
  AND2_X1 U2744 ( .A1(n2488), .A2(DATAI_27_), .ZN(n3947) );
  NAND2_X1 U2745 ( .A1(n4066), .A2(n3856), .ZN(n3857) );
  OR2_X1 U2746 ( .A1(n2492), .A2(n2971), .ZN(n2969) );
  NAND2_X1 U2747 ( .A1(n3963), .A2(n3964), .ZN(n3962) );
  OR2_X1 U2748 ( .A1(n3449), .A2(n3481), .ZN(n3474) );
  INV_X1 U2749 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4268) );
  INV_X1 U2750 ( .A(n3448), .ZN(n3446) );
  AND2_X1 U2751 ( .A1(n3038), .A2(n2985), .ZN(n2635) );
  NAND2_X1 U2752 ( .A1(n3171), .A2(n3170), .ZN(n2644) );
  INV_X1 U2753 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3136) );
  NOR2_X1 U2754 ( .A1(n3137), .A2(n3136), .ZN(n3176) );
  AND2_X1 U2755 ( .A1(n3848), .A2(n3847), .ZN(n3849) );
  INV_X1 U2756 ( .A(n4241), .ZN(n3682) );
  INV_X1 U2757 ( .A(n4559), .ZN(n4561) );
  AND2_X1 U2758 ( .A1(n4234), .A2(n4673), .ZN(n2996) );
  NAND2_X1 U2759 ( .A1(n3007), .A2(REG3_REG_1__SCAN_IN), .ZN(n2937) );
  OR2_X1 U2760 ( .A1(n3156), .A2(n5223), .ZN(n2936) );
  AND2_X1 U2761 ( .A1(n5219), .A2(REG1_REG_1__SCAN_IN), .ZN(n2799) );
  NOR2_X1 U2762 ( .A1(n5173), .A2(n5175), .ZN(n5174) );
  NOR2_X1 U2763 ( .A1(n2618), .A2(n2612), .ZN(n2611) );
  INV_X1 U2764 ( .A(n2615), .ZN(n2612) );
  NOR2_X1 U2765 ( .A1(n5199), .A2(n5236), .ZN(n5198) );
  NOR2_X1 U2766 ( .A1(n2880), .A2(n2706), .ZN(n5132) );
  OR2_X1 U2767 ( .A1(n5132), .A2(n5131), .ZN(n5129) );
  OR2_X1 U2768 ( .A1(n2884), .A2(n2809), .ZN(n2581) );
  NAND2_X1 U2769 ( .A1(n5129), .A2(n2708), .ZN(n2714) );
  NAND2_X1 U2770 ( .A1(n2716), .A2(n2624), .ZN(n2623) );
  INV_X1 U2771 ( .A(n2715), .ZN(n2716) );
  NAND2_X1 U2772 ( .A1(n2602), .A2(REG1_REG_8__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U2773 ( .A1(n2649), .A2(n2602), .ZN(n2600) );
  INV_X1 U2774 ( .A(n3233), .ZN(n2602) );
  NAND3_X1 U2775 ( .A1(n2709), .A2(n2660), .A3(n4963), .ZN(n2661) );
  INV_X1 U2776 ( .A(IR_REG_9__SCAN_IN), .ZN(n2660) );
  OR2_X1 U2777 ( .A1(n3408), .A2(n2726), .ZN(n2609) );
  OR2_X1 U2778 ( .A1(n3672), .A2(n2731), .ZN(n2605) );
  OAI21_X1 U2779 ( .B1(n2751), .B2(IR_REG_18__SCAN_IN), .A(n2899), .ZN(n2753)
         );
  NAND2_X1 U2780 ( .A1(n2753), .A2(n2759), .ZN(n2900) );
  NOR2_X1 U2781 ( .A1(n2843), .A2(n2831), .ZN(n2591) );
  NOR2_X1 U2782 ( .A1(n4303), .A2(n2577), .ZN(n2575) );
  OAI22_X1 U2783 ( .A1(n4303), .A2(n2578), .B1(n4314), .B2(n4324), .ZN(n2573)
         );
  NAND2_X1 U2784 ( .A1(n3928), .A2(n4342), .ZN(n3905) );
  OR2_X1 U2785 ( .A1(n4134), .A2(n4205), .ZN(n4322) );
  OAI22_X1 U2786 ( .A1(n2553), .A2(n2552), .B1(n2555), .B2(n2656), .ZN(n4337)
         );
  NAND2_X1 U2787 ( .A1(n2559), .A2(n2561), .ZN(n2552) );
  NOR2_X1 U2788 ( .A1(n2557), .A2(n2516), .ZN(n2555) );
  AND2_X1 U2789 ( .A1(n2488), .A2(DATAI_25_), .ZN(n4360) );
  NAND2_X1 U2790 ( .A1(n3151), .A2(REG3_REG_24__SCAN_IN), .ZN(n3834) );
  AND2_X1 U2791 ( .A1(n2488), .A2(DATAI_23_), .ZN(n4398) );
  NAND2_X1 U2792 ( .A1(n3149), .A2(REG3_REG_20__SCAN_IN), .ZN(n3768) );
  INV_X1 U2793 ( .A(n3752), .ZN(n3149) );
  NOR2_X1 U2794 ( .A1(n3561), .A2(n3600), .ZN(n3594) );
  NAND2_X1 U2795 ( .A1(n3594), .A2(REG3_REG_16__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U2796 ( .A1(n4553), .A2(n3683), .ZN(n4550) );
  OR2_X1 U2797 ( .A1(n4454), .A2(n4198), .ZN(n3685) );
  NOR2_X1 U2798 ( .A1(n3474), .A2(n4268), .ZN(n3549) );
  NAND2_X1 U2799 ( .A1(n3549), .A2(REG3_REG_14__SCAN_IN), .ZN(n3561) );
  INV_X1 U2800 ( .A(n4243), .ZN(n3513) );
  CLKBUF_X1 U2801 ( .A(n3506), .Z(n3530) );
  AND2_X1 U2802 ( .A1(n3334), .A2(REG3_REG_10__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U2803 ( .A1(n3351), .A2(REG3_REG_11__SCAN_IN), .ZN(n3449) );
  AND2_X1 U2804 ( .A1(n3528), .A2(n3526), .ZN(n3503) );
  OR2_X1 U2805 ( .A1(n3189), .A2(n4921), .ZN(n3280) );
  INV_X1 U2806 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4943) );
  NOR2_X1 U2807 ( .A1(n3280), .A2(n4943), .ZN(n3334) );
  NAND2_X1 U2808 ( .A1(n2533), .A2(n3242), .ZN(n2530) );
  NAND2_X1 U2809 ( .A1(n2529), .A2(n2528), .ZN(n2527) );
  INV_X1 U2810 ( .A(n4247), .ZN(n3976) );
  INV_X1 U2811 ( .A(n4581), .ZN(n4560) );
  INV_X1 U2812 ( .A(n4398), .ZN(n4406) );
  INV_X1 U2814 ( .A(n4443), .ZN(n4472) );
  INV_X1 U2815 ( .A(n3893), .ZN(n3690) );
  OR2_X2 U2816 ( .A1(n3689), .A2(n3893), .ZN(n4526) );
  INV_X1 U2817 ( .A(n3679), .ZN(n3657) );
  NAND2_X1 U2818 ( .A1(n3609), .A2(n3608), .ZN(n2566) );
  CLKBUF_X1 U2819 ( .A(n3648), .Z(n3649) );
  CLKBUF_X1 U2820 ( .A(n3388), .Z(n3420) );
  NOR2_X2 U2821 ( .A1(n3117), .A2(n3223), .ZN(n3217) );
  NAND2_X1 U2822 ( .A1(n5212), .A2(n2947), .ZN(n4581) );
  NAND2_X1 U2823 ( .A1(n2953), .A2(n2980), .ZN(n3035) );
  INV_X1 U2824 ( .A(n4501), .ZN(n4554) );
  NAND2_X1 U2825 ( .A1(n2873), .A2(n4671), .ZN(n2993) );
  NOR2_X1 U2826 ( .A1(n2767), .A2(n2766), .ZN(n2770) );
  NAND2_X1 U2827 ( .A1(n2770), .A2(n4996), .ZN(n2772) );
  NAND2_X1 U2828 ( .A1(n2747), .A2(n4980), .ZN(n2751) );
  INV_X1 U2829 ( .A(n2746), .ZN(n2747) );
  NAND2_X1 U2830 ( .A1(n4162), .A2(DATAI_1_), .ZN(n2933) );
  CLKBUF_X1 U2831 ( .A(n3984), .Z(n3985) );
  NAND2_X1 U2832 ( .A1(n2636), .A2(n3038), .ZN(n2988) );
  CLKBUF_X1 U2833 ( .A(n3724), .Z(n3711) );
  AND2_X1 U2834 ( .A1(n3005), .A2(n5184), .ZN(n5284) );
  INV_X1 U2835 ( .A(n5284), .ZN(n4071) );
  INV_X1 U2836 ( .A(n5300), .ZN(n4068) );
  NAND2_X1 U2837 ( .A1(n3866), .A2(n3865), .ZN(n4341) );
  NAND2_X1 U2838 ( .A1(n3841), .A2(n3840), .ZN(n4344) );
  OR2_X1 U2839 ( .A1(n4366), .A2(n3836), .ZN(n3841) );
  NAND2_X1 U2840 ( .A1(n3807), .A2(n3806), .ZN(n4379) );
  NAND2_X1 U2841 ( .A1(n3791), .A2(n3790), .ZN(n4433) );
  NAND2_X1 U2842 ( .A1(n3774), .A2(n3773), .ZN(n4419) );
  NAND2_X1 U2843 ( .A1(n3743), .A2(n3742), .ZN(n4465) );
  OAI211_X1 U2844 ( .C1(n4513), .C2(n3836), .A(n3718), .B(n3717), .ZN(n4524)
         );
  NAND4_X1 U2845 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n4505)
         );
  NAND4_X1 U2846 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n5295)
         );
  NAND4_X1 U2847 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n4244)
         );
  INV_X1 U2848 ( .A(n2971), .ZN(n4254) );
  OR2_X1 U2849 ( .A1(n2786), .A2(n2785), .ZN(n2787) );
  XNOR2_X1 U2850 ( .A(n2803), .B(n5075), .ZN(n4261) );
  NAND2_X1 U2851 ( .A1(n4261), .A2(REG1_REG_3__SCAN_IN), .ZN(n4260) );
  NOR2_X1 U2852 ( .A1(n5202), .A2(n5203), .ZN(n5201) );
  NAND2_X1 U2853 ( .A1(n2599), .A2(REG1_REG_4__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U2854 ( .A1(n2655), .A2(n2599), .ZN(n2597) );
  INV_X1 U2855 ( .A(n5124), .ZN(n2599) );
  NOR2_X1 U2856 ( .A1(n2881), .A2(n2882), .ZN(n2880) );
  NAND2_X1 U2857 ( .A1(n2581), .A2(n2580), .ZN(n5138) );
  INV_X1 U2858 ( .A(n5135), .ZN(n2580) );
  NOR2_X1 U2859 ( .A1(n3084), .A2(n3083), .ZN(n3082) );
  NOR2_X1 U2860 ( .A1(n3080), .A2(n3081), .ZN(n3079) );
  NAND2_X1 U2861 ( .A1(n2620), .A2(n2623), .ZN(n3229) );
  NOR2_X1 U2862 ( .A1(n3409), .A2(n3410), .ZN(n3408) );
  AND2_X1 U2863 ( .A1(n2609), .A2(n2608), .ZN(n3493) );
  INV_X1 U2864 ( .A(n3494), .ZN(n2608) );
  INV_X1 U2865 ( .A(n2609), .ZN(n3495) );
  XNOR2_X1 U2866 ( .A(n2817), .B(n3671), .ZN(n3668) );
  NOR2_X1 U2867 ( .A1(n3668), .A2(n5278), .ZN(n3667) );
  AND2_X1 U2868 ( .A1(n2605), .A2(n2604), .ZN(n4265) );
  INV_X1 U2869 ( .A(n4267), .ZN(n2604) );
  INV_X1 U2870 ( .A(n2605), .ZN(n4266) );
  NOR2_X1 U2871 ( .A1(n4280), .A2(n4281), .ZN(n4279) );
  OAI21_X1 U2872 ( .B1(n4280), .B2(n2595), .A(n2594), .ZN(n5142) );
  NAND2_X1 U2873 ( .A1(n2596), .A2(REG1_REG_14__SCAN_IN), .ZN(n2595) );
  INV_X1 U2874 ( .A(n5143), .ZN(n2596) );
  OR2_X1 U2875 ( .A1(n5106), .A2(n5184), .ZN(n5181) );
  NAND2_X1 U2876 ( .A1(n2584), .A2(n2583), .ZN(n2840) );
  INV_X1 U2877 ( .A(n2557), .ZN(n2554) );
  NAND2_X1 U2878 ( .A1(n4393), .A2(n2559), .ZN(n2556) );
  NAND2_X1 U2879 ( .A1(n2545), .A2(n2549), .ZN(n4432) );
  NAND2_X1 U2880 ( .A1(n3901), .A2(n2551), .ZN(n2545) );
  AOI21_X1 U2881 ( .B1(n2539), .B2(n2538), .A(n2507), .ZN(n2534) );
  NAND2_X1 U2882 ( .A1(n2537), .A2(n2539), .ZN(n2535) );
  NAND2_X1 U2883 ( .A1(n2540), .A2(n3243), .ZN(n3260) );
  NAND2_X1 U2884 ( .A1(n4545), .A2(n5340), .ZN(n4518) );
  NAND2_X1 U2885 ( .A1(n3015), .A2(n3014), .ZN(n5307) );
  OR2_X1 U2886 ( .A1(n4586), .A2(n5338), .ZN(n4587) );
  OAI21_X1 U2887 ( .B1(n4331), .B2(n4330), .A(n4329), .ZN(n4640) );
  AND2_X2 U2888 ( .A1(n2928), .A2(n3201), .ZN(n5348) );
  INV_X1 U2889 ( .A(n5091), .ZN(n5101) );
  NAND2_X1 U2890 ( .A1(n2894), .A2(n2899), .ZN(n2867) );
  BUF_X1 U2891 ( .A(n2794), .Z(n3004) );
  AND2_X1 U2892 ( .A1(n3068), .A2(STATE_REG_SCAN_IN), .ZN(n2879) );
  INV_X1 U2893 ( .A(n4167), .ZN(n4673) );
  AND2_X1 U2894 ( .A1(n2669), .A2(n2668), .ZN(n5150) );
  AND2_X1 U2895 ( .A1(n2673), .A2(n2727), .ZN(n4676) );
  AND2_X1 U2896 ( .A1(n2713), .A2(n2717), .ZN(n4678) );
  OR2_X1 U2897 ( .A1(n2677), .A2(n2663), .ZN(n2678) );
  CLKBUF_X1 U2898 ( .A(n2797), .Z(n5219) );
  OAI211_X1 U2899 ( .C1(n2505), .C2(n2593), .A(n2844), .B(n5177), .ZN(n2851)
         );
  AOI21_X1 U2900 ( .B1(n4412), .B2(n4394), .A(n2652), .ZN(n4393) );
  AND2_X1 U2901 ( .A1(n3446), .A2(n3443), .ZN(n2500) );
  AND2_X1 U2902 ( .A1(n2531), .A2(n2527), .ZN(n2501) );
  AND2_X1 U2903 ( .A1(n3608), .A2(n3651), .ZN(n2502) );
  INV_X1 U2904 ( .A(n4462), .ZN(n2550) );
  NOR2_X1 U2905 ( .A1(n5295), .A2(n3679), .ZN(n2503) );
  OR2_X1 U2906 ( .A1(n4524), .A2(n4503), .ZN(n2504) );
  AND2_X1 U2907 ( .A1(n5153), .A2(n2832), .ZN(n2505) );
  OR2_X1 U2908 ( .A1(n4248), .A2(n4057), .ZN(n2506) );
  INV_X2 U2909 ( .A(IR_REG_31__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U2910 ( .A1(n2556), .A2(n2554), .ZN(n4355) );
  AND2_X1 U2911 ( .A1(n4248), .A2(n4057), .ZN(n2507) );
  NOR2_X1 U2912 ( .A1(n3995), .A2(n3849), .ZN(n2508) );
  NAND2_X1 U2913 ( .A1(n2714), .A2(n4678), .ZN(n2715) );
  AND2_X1 U2914 ( .A1(n2677), .A2(n4952), .ZN(n2681) );
  AND2_X1 U2915 ( .A1(n2681), .A2(n2658), .ZN(n2695) );
  NAND2_X1 U2916 ( .A1(n3989), .A2(n3983), .ZN(n4031) );
  NOR2_X1 U2917 ( .A1(n4279), .A2(n2826), .ZN(n2509) );
  NAND2_X1 U2918 ( .A1(n5075), .A2(n2686), .ZN(n2510) );
  NAND2_X1 U2919 ( .A1(n2670), .A2(n2645), .ZN(n2511) );
  OR2_X1 U2920 ( .A1(n3275), .A2(n2507), .ZN(n2536) );
  INV_X1 U2921 ( .A(n2536), .ZN(n2528) );
  AND2_X1 U2922 ( .A1(n2645), .A2(n4989), .ZN(n2512) );
  AND2_X1 U2923 ( .A1(n2785), .A2(n5001), .ZN(n2513) );
  OR2_X1 U2924 ( .A1(n4439), .A2(n4464), .ZN(n2514) );
  OAI21_X1 U2925 ( .B1(n4393), .B2(n4181), .A(n4180), .ZN(n4372) );
  NAND2_X1 U2926 ( .A1(n3962), .A2(n3751), .ZN(n4022) );
  INV_X1 U2927 ( .A(n4180), .ZN(n2560) );
  OR2_X1 U2928 ( .A1(n4242), .A2(n5281), .ZN(n2515) );
  AND2_X1 U2929 ( .A1(n4381), .A2(n4364), .ZN(n2516) );
  NOR2_X1 U2930 ( .A1(n4419), .A2(n4444), .ZN(n2517) );
  NOR2_X1 U2931 ( .A1(n4467), .A2(n3939), .ZN(n2518) );
  INV_X1 U2932 ( .A(n2653), .ZN(n2578) );
  INV_X1 U2933 ( .A(n2656), .ZN(n2561) );
  INV_X1 U2934 ( .A(n2577), .ZN(n2576) );
  NAND2_X1 U2935 ( .A1(n3908), .A2(n3905), .ZN(n2577) );
  NAND2_X1 U2936 ( .A1(n3901), .A2(n3900), .ZN(n4452) );
  OR2_X1 U2937 ( .A1(n2720), .A2(n2719), .ZN(n2519) );
  AND2_X1 U2938 ( .A1(n3796), .A2(n3983), .ZN(n2520) );
  OR2_X1 U2939 ( .A1(n4508), .A2(n4489), .ZN(n2521) );
  NAND2_X1 U2940 ( .A1(n2644), .A2(n3172), .ZN(n3186) );
  NAND2_X1 U2941 ( .A1(n3242), .A2(n3241), .ZN(n3376) );
  NAND2_X1 U2942 ( .A1(n2566), .A2(n3611), .ZN(n3652) );
  NAND2_X1 U2943 ( .A1(n2535), .A2(n2534), .ZN(n3277) );
  NAND2_X1 U2944 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  NAND2_X1 U2945 ( .A1(n3348), .A2(n3347), .ZN(n3444) );
  NOR2_X1 U2946 ( .A1(n3079), .A2(n2716), .ZN(n2522) );
  NOR2_X1 U2947 ( .A1(n3082), .A2(n2649), .ZN(n2523) );
  AND2_X1 U2948 ( .A1(n4552), .A2(n4100), .ZN(n4155) );
  INV_X1 U2949 ( .A(n4155), .ZN(n2565) );
  NAND2_X1 U2950 ( .A1(n2637), .A2(n2985), .ZN(n2986) );
  NOR2_X1 U2951 ( .A1(n5201), .A2(n2694), .ZN(n2524) );
  NOR2_X1 U2952 ( .A1(n5198), .A2(n2655), .ZN(n2525) );
  AND2_X1 U2953 ( .A1(n2591), .A2(n2592), .ZN(n2526) );
  INV_X1 U2954 ( .A(n2843), .ZN(n2593) );
  XNOR2_X1 U2955 ( .A(n2674), .B(IR_REG_1__SCAN_IN), .ZN(n2797) );
  OR2_X4 U2956 ( .A1(n3369), .A2(n4057), .ZN(n3267) );
  NAND2_X2 U2957 ( .A1(n3383), .A2(n4146), .ZN(n3509) );
  OR2_X1 U2958 ( .A1(n2941), .A2(n4075), .ZN(n3027) );
  AOI21_X2 U2959 ( .B1(n4340), .B2(n4130), .A(n4139), .ZN(n4323) );
  AOI21_X2 U2960 ( .B1(n3262), .B2(n4087), .A(n4091), .ZN(n3278) );
  NOR2_X2 U2961 ( .A1(n4321), .A2(n4205), .ZN(n4308) );
  NAND2_X1 U2962 ( .A1(n3684), .A2(n4156), .ZN(n4453) );
  AND2_X2 U2963 ( .A1(n2645), .A2(n2776), .ZN(n2571) );
  NAND2_X1 U2964 ( .A1(n2530), .A2(n2501), .ZN(n3392) );
  INV_X1 U2965 ( .A(n2532), .ZN(n2531) );
  NAND2_X1 U2966 ( .A1(n3242), .A2(n2541), .ZN(n2540) );
  NAND2_X1 U2967 ( .A1(n3901), .A2(n2546), .ZN(n2543) );
  NAND2_X1 U2968 ( .A1(n2543), .A2(n2544), .ZN(n4412) );
  INV_X1 U2969 ( .A(n4393), .ZN(n2553) );
  NAND2_X1 U2970 ( .A1(n3609), .A2(n2564), .ZN(n2562) );
  NAND2_X1 U2971 ( .A1(n2562), .A2(n2563), .ZN(n4540) );
  NAND2_X1 U2972 ( .A1(n2571), .A2(n2670), .ZN(n2864) );
  NAND2_X1 U2973 ( .A1(n2571), .A2(n2570), .ZN(n2892) );
  AOI21_X1 U2974 ( .B1(n3906), .B2(n2576), .A(n2653), .ZN(n4304) );
  NAND2_X1 U2975 ( .A1(n3906), .A2(n2575), .ZN(n2574) );
  NAND2_X1 U2976 ( .A1(n3906), .A2(n3905), .ZN(n4320) );
  NAND3_X1 U2977 ( .A1(n2579), .A2(n2658), .A3(n2677), .ZN(n2698) );
  NOR2_X2 U2978 ( .A1(n2703), .A2(n2661), .ZN(n2721) );
  INV_X1 U2979 ( .A(n2581), .ZN(n5136) );
  NOR2_X1 U2980 ( .A1(n2885), .A2(n2886), .ZN(n2884) );
  XNOR2_X1 U2981 ( .A(n2808), .B(n3164), .ZN(n2885) );
  NOR2_X1 U2982 ( .A1(n3488), .A2(n3489), .ZN(n3487) );
  NAND2_X1 U2983 ( .A1(n5153), .A2(n2526), .ZN(n2583) );
  INV_X1 U2984 ( .A(n2585), .ZN(n2584) );
  NAND2_X1 U2985 ( .A1(n2826), .A2(n2596), .ZN(n2594) );
  OAI21_X1 U2986 ( .B1(n5199), .B2(n2598), .A(n2597), .ZN(n5123) );
  OAI21_X1 U2987 ( .B1(n3084), .B2(n2601), .A(n2600), .ZN(n3232) );
  NOR2_X1 U2988 ( .A1(n5108), .A2(n5186), .ZN(n5107) );
  OAI21_X1 U2989 ( .B1(n2797), .B2(REG2_REG_1__SCAN_IN), .A(n2606), .ZN(n5108)
         );
  NAND2_X1 U2990 ( .A1(n2797), .A2(REG2_REG_1__SCAN_IN), .ZN(n2606) );
  INV_X1 U2991 ( .A(n5219), .ZN(n2675) );
  NOR2_X1 U2992 ( .A1(n5107), .A2(n2676), .ZN(n5170) );
  INV_X1 U2993 ( .A(n5075), .ZN(n2617) );
  NAND2_X1 U2994 ( .A1(n2680), .A2(n2679), .ZN(n2686) );
  NAND3_X1 U2995 ( .A1(n2613), .A2(n2615), .A3(n2610), .ZN(n4257) );
  NAND3_X1 U2996 ( .A1(n2613), .A2(n2611), .A3(n2610), .ZN(n4255) );
  INV_X1 U2997 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2618) );
  INV_X1 U2998 ( .A(n3080), .ZN(n2622) );
  NAND2_X1 U2999 ( .A1(n2694), .A2(n2627), .ZN(n2625) );
  NAND2_X1 U3000 ( .A1(n3963), .A2(n2629), .ZN(n2628) );
  NAND3_X1 U3001 ( .A1(n2637), .A2(n2635), .A3(n2636), .ZN(n3039) );
  NAND2_X1 U3002 ( .A1(n2964), .A2(n2965), .ZN(n2636) );
  NAND2_X1 U3003 ( .A1(n2966), .A2(n2967), .ZN(n3038) );
  NAND2_X1 U3004 ( .A1(n3097), .A2(n3098), .ZN(n2637) );
  NOR2_X1 U3005 ( .A1(n3994), .A2(n3996), .ZN(n3995) );
  INV_X1 U3006 ( .A(n2638), .ZN(n3945) );
  AOI21_X1 U3007 ( .B1(n3994), .B2(n2641), .A(n2639), .ZN(n2638) );
  INV_X1 U3008 ( .A(n3996), .ZN(n2640) );
  INV_X1 U3009 ( .A(n3849), .ZN(n2643) );
  NAND2_X1 U3010 ( .A1(n3444), .A2(n2500), .ZN(n3580) );
  NAND2_X1 U3011 ( .A1(n3989), .A2(n2520), .ZN(n4032) );
  NAND2_X2 U3012 ( .A1(n3780), .A2(n3779), .ZN(n3989) );
  NAND3_X1 U3013 ( .A1(n2644), .A2(n2651), .A3(n3172), .ZN(n3320) );
  NAND2_X1 U3014 ( .A1(n2670), .A2(n2662), .ZN(n2762) );
  NAND2_X1 U3015 ( .A1(n2670), .A2(n2512), .ZN(n2789) );
  AOI211_X2 U3016 ( .C1(n4504), .C2(n4341), .A(n4311), .B(n4310), .ZN(n4591)
         );
  NAND2_X1 U3017 ( .A1(n3353), .A2(REG2_REG_0__SCAN_IN), .ZN(n2908) );
  AOI22_X1 U3018 ( .A1(n2976), .A2(n3094), .B1(n2968), .B2(n5167), .ZN(n2970)
         );
  XNOR2_X1 U3019 ( .A(n2765), .B(IR_REG_24__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U3020 ( .A1(n2782), .A2(n2899), .ZN(n2765) );
  OR2_X2 U3021 ( .A1(n2761), .A2(n2760), .ZN(n2647) );
  AND2_X1 U3022 ( .A1(n2800), .A2(REG1_REG_2__SCAN_IN), .ZN(n2648) );
  AND2_X1 U3023 ( .A1(n2812), .A2(n4678), .ZN(n2649) );
  OR2_X1 U3024 ( .A1(n2811), .A2(n2810), .ZN(n2650) );
  OR2_X1 U3025 ( .A1(n5106), .A2(n4231), .ZN(n5200) );
  INV_X1 U3026 ( .A(n5200), .ZN(n2795) );
  OR2_X1 U3027 ( .A1(n5106), .A2(n4670), .ZN(n5197) );
  INV_X1 U3028 ( .A(IR_REG_27__SCAN_IN), .ZN(n2785) );
  AND2_X1 U3029 ( .A1(n3188), .A2(n3187), .ZN(n2651) );
  AND2_X1 U3030 ( .A1(n4433), .A2(n4418), .ZN(n2652) );
  INV_X1 U3031 ( .A(n3024), .ZN(n3023) );
  NAND2_X1 U3032 ( .A1(n3758), .A2(n3757), .ZN(n4439) );
  AOI21_X1 U3033 ( .B1(n4349), .B2(n3007), .A(n3853), .ZN(n3928) );
  INV_X1 U3034 ( .A(n3928), .ZN(n3903) );
  INV_X1 U3035 ( .A(n4677), .ZN(n2720) );
  AND2_X1 U3036 ( .A1(n4341), .A2(n3947), .ZN(n2653) );
  AND2_X1 U3037 ( .A1(n3871), .A2(n3870), .ZN(n2654) );
  AND2_X1 U3038 ( .A1(n2805), .A2(n5206), .ZN(n2655) );
  AND2_X1 U3039 ( .A1(n4344), .A2(n4360), .ZN(n2656) );
  NAND2_X1 U3040 ( .A1(n3574), .A2(n3573), .ZN(n2657) );
  INV_X1 U3041 ( .A(n4464), .ZN(n4473) );
  AND2_X1 U3042 ( .A1(n2488), .A2(DATAI_20_), .ZN(n4464) );
  OR4_X1 U3043 ( .A1(n5011), .A2(n5010), .A3(n5009), .A4(n5008), .ZN(n5026) );
  INV_X1 U3044 ( .A(n2758), .ZN(n2761) );
  INV_X1 U3045 ( .A(n4342), .ZN(n3902) );
  AND2_X1 U3046 ( .A1(n5219), .A2(REG2_REG_1__SCAN_IN), .ZN(n2676) );
  INV_X1 U3047 ( .A(n3044), .ZN(n3872) );
  INV_X1 U3048 ( .A(n3785), .ZN(n3150) );
  INV_X1 U3049 ( .A(n5206), .ZN(n2689) );
  INV_X1 U3050 ( .A(n2824), .ZN(n2825) );
  INV_X1 U3051 ( .A(n3818), .ZN(n3151) );
  INV_X1 U3052 ( .A(n3737), .ZN(n3148) );
  NAND2_X1 U3053 ( .A1(n2923), .A2(n4673), .ZN(n2957) );
  INV_X1 U3054 ( .A(n3938), .ZN(n3897) );
  INV_X1 U3055 ( .A(n4245), .ZN(n3394) );
  INV_X1 U3056 ( .A(n3956), .ZN(n3813) );
  INV_X1 U3057 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4921) );
  OR2_X1 U3058 ( .A1(n3859), .A2(n3152), .ZN(n3861) );
  OR2_X1 U3059 ( .A1(n3834), .A2(n4741), .ZN(n3859) );
  INV_X1 U3060 ( .A(n3046), .ZN(n3884) );
  INV_X1 U3061 ( .A(n3413), .ZN(n2724) );
  INV_X1 U3062 ( .A(n4284), .ZN(n2823) );
  INV_X1 U3063 ( .A(n2749), .ZN(n2750) );
  NOR2_X1 U3064 ( .A1(n4455), .A2(n4454), .ZN(n4520) );
  NAND2_X1 U3065 ( .A1(n3061), .A2(REG3_REG_5__SCAN_IN), .ZN(n3137) );
  OR2_X1 U3066 ( .A1(n4240), .A2(n3893), .ZN(n3894) );
  INV_X1 U3067 ( .A(n3500), .ZN(n3531) );
  OR2_X1 U3068 ( .A1(n3768), .A2(n4928), .ZN(n3785) );
  OR2_X1 U3069 ( .A1(n2490), .A2(n2971), .ZN(n2972) );
  INV_X1 U3070 ( .A(n4419), .ZN(n4467) );
  INV_X1 U3071 ( .A(n4344), .ZN(n4381) );
  AND2_X1 U3072 ( .A1(n3861), .A2(n3860), .ZN(n4332) );
  NAND2_X1 U3073 ( .A1(n3714), .A2(REG3_REG_18__SCAN_IN), .ZN(n3737) );
  NOR2_X1 U3074 ( .A1(n3667), .A2(n2818), .ZN(n4274) );
  NAND2_X1 U3075 ( .A1(n3907), .A2(n4330), .ZN(n3908) );
  INV_X1 U3076 ( .A(n4439), .ZN(n4483) );
  INV_X1 U3077 ( .A(n3685), .ZN(n4156) );
  INV_X1 U3078 ( .A(n4548), .ZN(n4504) );
  INV_X1 U3079 ( .A(n4360), .ZN(n4364) );
  INV_X1 U3080 ( .A(n4444), .ZN(n3939) );
  OAI21_X1 U3081 ( .B1(n3895), .B2(n4156), .A(n3894), .ZN(n4537) );
  INV_X1 U3082 ( .A(n3036), .ZN(n3106) );
  AND2_X1 U3083 ( .A1(n3015), .A2(n3069), .ZN(n3202) );
  INV_X1 U3084 ( .A(IR_REG_10__SCAN_IN), .ZN(n4772) );
  AND2_X1 U3085 ( .A1(n2488), .A2(DATAI_21_), .ZN(n4444) );
  AND2_X1 U3086 ( .A1(n2488), .A2(DATAI_24_), .ZN(n4378) );
  AND2_X1 U3087 ( .A1(n2488), .A2(DATAI_22_), .ZN(n4418) );
  OR2_X1 U3088 ( .A1(n4315), .A2(n3836), .ZN(n3162) );
  OR2_X1 U3089 ( .A1(n4035), .A2(n3836), .ZN(n3791) );
  NOR2_X1 U3090 ( .A1(n4131), .A2(n4206), .ZN(n4303) );
  NAND2_X1 U3091 ( .A1(n4545), .A2(n3293), .ZN(n5309) );
  INV_X1 U3092 ( .A(n4546), .ZN(n4525) );
  INV_X1 U3093 ( .A(n5309), .ZN(n5352) );
  NAND2_X1 U3094 ( .A1(n2906), .A2(n2905), .ZN(n4501) );
  INV_X1 U3095 ( .A(n5272), .ZN(n5340) );
  AND4_X1 U3096 ( .A1(n3202), .A2(n2925), .A3(n3013), .A4(n2924), .ZN(n2928)
         );
  AND2_X1 U3097 ( .A1(n2959), .A2(n2879), .ZN(n3015) );
  AND2_X1 U3098 ( .A1(n2837), .A2(n2836), .ZN(n5196) );
  NAND2_X1 U3099 ( .A1(n3072), .A2(STATE_REG_SCAN_IN), .ZN(n5300) );
  OR2_X1 U3100 ( .A1(n3012), .A2(n2998), .ZN(n5291) );
  AND2_X1 U3101 ( .A1(n3162), .A2(n3161), .ZN(n4324) );
  NAND4_X1 U3102 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n4241)
         );
  OR2_X1 U3103 ( .A1(n2959), .A2(n2852), .ZN(n4253) );
  AOI21_X1 U3104 ( .B1(n5196), .B2(ADDR_REG_18__SCAN_IN), .A(n4048), .ZN(n2849) );
  AND2_X2 U3105 ( .A1(n2928), .A2(n2995), .ZN(n5344) );
  INV_X1 U3106 ( .A(n5344), .ZN(n5342) );
  INV_X1 U3107 ( .A(n5348), .ZN(n5345) );
  AND2_X1 U3108 ( .A1(n2685), .A2(n2687), .ZN(n5075) );
  NOR2_X2 U3109 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2658)
         );
  AND2_X2 U3110 ( .A1(n2721), .A2(n4772), .ZN(n2670) );
  NOR2_X1 U3111 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2662)
         );
  NAND2_X1 U3112 ( .A1(n2899), .A2(IR_REG_13__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3113 ( .A1(n2739), .A2(n2664), .ZN(n2733) );
  NAND2_X1 U3114 ( .A1(n2665), .A2(n2899), .ZN(n2667) );
  INV_X1 U3115 ( .A(IR_REG_15__SCAN_IN), .ZN(n4783) );
  NAND2_X1 U3116 ( .A1(n2667), .A2(n4783), .ZN(n2669) );
  NAND2_X1 U3117 ( .A1(n2669), .A2(n2899), .ZN(n2666) );
  INV_X1 U3118 ( .A(IR_REG_16__SCAN_IN), .ZN(n4782) );
  XNOR2_X1 U3119 ( .A(n2666), .B(n4782), .ZN(n4299) );
  INV_X1 U3120 ( .A(n4299), .ZN(n3629) );
  OR2_X1 U3121 ( .A1(n2667), .A2(n4783), .ZN(n2668) );
  XNOR2_X1 U3122 ( .A(n2739), .B(IR_REG_13__SCAN_IN), .ZN(n4675) );
  OR2_X1 U3123 ( .A1(n2670), .A2(n2663), .ZN(n2672) );
  INV_X1 U3124 ( .A(n2672), .ZN(n2671) );
  NAND2_X1 U3125 ( .A1(n2671), .A2(IR_REG_11__SCAN_IN), .ZN(n2673) );
  INV_X1 U3126 ( .A(IR_REG_11__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U3127 ( .A1(n2672), .A2(n4967), .ZN(n2727) );
  INV_X1 U3128 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3081) );
  NAND2_X1 U3129 ( .A1(n5167), .A2(REG2_REG_0__SCAN_IN), .ZN(n5186) );
  INV_X1 U3130 ( .A(REG2_REG_1__SCAN_IN), .ZN(n5223) );
  XNOR2_X2 U3131 ( .A(n2678), .B(IR_REG_2__SCAN_IN), .ZN(n2800) );
  INV_X1 U3132 ( .A(REG2_REG_2__SCAN_IN), .ZN(n5227) );
  INV_X1 U3133 ( .A(n2800), .ZN(n5180) );
  NOR2_X1 U3134 ( .A1(n5170), .A2(n5171), .ZN(n5169) );
  INV_X1 U3135 ( .A(n5169), .ZN(n2680) );
  NAND2_X1 U3136 ( .A1(n2800), .A2(REG2_REG_2__SCAN_IN), .ZN(n2679) );
  NOR2_X1 U3137 ( .A1(n2681), .A2(n2663), .ZN(n2682) );
  NAND2_X1 U3138 ( .A1(n2682), .A2(IR_REG_3__SCAN_IN), .ZN(n2685) );
  INV_X1 U3139 ( .A(n2682), .ZN(n2684) );
  INV_X1 U3140 ( .A(IR_REG_3__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3141 ( .A1(n2684), .A2(n2683), .ZN(n2687) );
  NAND2_X1 U3142 ( .A1(n4255), .A2(n2510), .ZN(n2691) );
  INV_X1 U3143 ( .A(n2691), .ZN(n2690) );
  NAND2_X1 U3144 ( .A1(n2687), .A2(n2899), .ZN(n2688) );
  XNOR2_X1 U3145 ( .A(n2688), .B(IR_REG_4__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U3146 ( .A1(n2690), .A2(n2689), .ZN(n2692) );
  NAND2_X1 U3147 ( .A1(n2691), .A2(n5206), .ZN(n2693) );
  INV_X1 U31480 ( .A(REG2_REG_4__SCAN_IN), .ZN(n5203) );
  INV_X1 U31490 ( .A(n2693), .ZN(n2694) );
  NOR2_X1 U3150 ( .A1(n2695), .A2(n2663), .ZN(n2696) );
  MUX2_X1 U3151 ( .A(n2663), .B(n2696), .S(IR_REG_5__SCAN_IN), .Z(n2697) );
  INV_X1 U3152 ( .A(n2697), .ZN(n2699) );
  AND2_X1 U3153 ( .A1(n2699), .A2(n2698), .ZN(n5126) );
  NAND2_X1 U3154 ( .A1(n5126), .A2(REG2_REG_5__SCAN_IN), .ZN(n2700) );
  OAI21_X1 U3155 ( .B1(n5126), .B2(REG2_REG_5__SCAN_IN), .A(n2700), .ZN(n5120)
         );
  NAND2_X1 U3156 ( .A1(n2698), .A2(n2899), .ZN(n2702) );
  MUX2_X1 U3157 ( .A(n2899), .B(n2702), .S(IR_REG_6__SCAN_IN), .Z(n2704) );
  NAND2_X1 U3158 ( .A1(n2704), .A2(n2703), .ZN(n3164) );
  XNOR2_X1 U3159 ( .A(n2705), .B(n3164), .ZN(n2881) );
  INV_X1 U3160 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2882) );
  NOR2_X1 U3161 ( .A1(n2705), .A2(n3164), .ZN(n2706) );
  NAND2_X1 U3162 ( .A1(n2703), .A2(n2899), .ZN(n2710) );
  XNOR2_X1 U3163 ( .A(n2710), .B(IR_REG_7__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U3164 ( .A1(n5137), .A2(REG2_REG_7__SCAN_IN), .ZN(n2708) );
  OR2_X1 U3165 ( .A1(n5137), .A2(REG2_REG_7__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U3166 ( .A1(n2708), .A2(n2707), .ZN(n5131) );
  NAND2_X1 U3167 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  NAND2_X1 U3168 ( .A1(n2711), .A2(n2899), .ZN(n2712) );
  OR2_X1 U3169 ( .A1(n2712), .A2(n4963), .ZN(n2713) );
  NAND2_X1 U3170 ( .A1(n2712), .A2(n4963), .ZN(n2717) );
  OAI21_X1 U3171 ( .B1(n2714), .B2(n4678), .A(n2715), .ZN(n3080) );
  INV_X1 U3172 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U3173 ( .A1(n2717), .A2(n2899), .ZN(n2718) );
  XNOR2_X1 U3174 ( .A(n2718), .B(IR_REG_9__SCAN_IN), .ZN(n4677) );
  MUX2_X1 U3175 ( .A(n2719), .B(REG2_REG_9__SCAN_IN), .S(n4677), .Z(n3230) );
  INV_X1 U3176 ( .A(n2725), .ZN(n2723) );
  OR2_X1 U3177 ( .A1(n2721), .A2(n2663), .ZN(n2722) );
  XNOR2_X1 U3178 ( .A(n2722), .B(n4772), .ZN(n3413) );
  NOR2_X1 U3179 ( .A1(n2723), .A2(n3413), .ZN(n2726) );
  INV_X1 U3180 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3410) );
  INV_X1 U3181 ( .A(n4676), .ZN(n3492) );
  AOI22_X1 U3182 ( .A1(n4676), .A2(n3533), .B1(REG2_REG_11__SCAN_IN), .B2(
        n3492), .ZN(n3494) );
  NAND2_X1 U3183 ( .A1(n2727), .A2(n2899), .ZN(n2729) );
  INV_X1 U3184 ( .A(IR_REG_12__SCAN_IN), .ZN(n2728) );
  XNOR2_X1 U3185 ( .A(n2729), .B(n2728), .ZN(n3671) );
  NOR2_X1 U3186 ( .A1(n2730), .A2(n3671), .ZN(n2731) );
  INV_X1 U3187 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3674) );
  XNOR2_X1 U3188 ( .A(n2730), .B(n3671), .ZN(n3673) );
  INV_X1 U3189 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2732) );
  MUX2_X1 U3190 ( .A(n2732), .B(REG2_REG_13__SCAN_IN), .S(n4675), .Z(n4267) );
  XNOR2_X1 U3191 ( .A(n2733), .B(IR_REG_14__SCAN_IN), .ZN(n4284) );
  NOR2_X1 U3192 ( .A1(n2734), .A2(n4284), .ZN(n2735) );
  INV_X1 U3193 ( .A(REG2_REG_14__SCAN_IN), .ZN(n5313) );
  XNOR2_X1 U3194 ( .A(n2734), .B(n4284), .ZN(n4286) );
  NOR2_X1 U3195 ( .A1(n5313), .A2(n4286), .ZN(n4285) );
  NOR2_X1 U3196 ( .A1(n2735), .A2(n4285), .ZN(n5148) );
  NAND2_X1 U3197 ( .A1(n5150), .A2(REG2_REG_15__SCAN_IN), .ZN(n2736) );
  OAI21_X1 U3198 ( .B1(n5150), .B2(REG2_REG_15__SCAN_IN), .A(n2736), .ZN(n5147) );
  NOR2_X1 U3199 ( .A1(n5148), .A2(n5147), .ZN(n5146) );
  XNOR2_X1 U3200 ( .A(n3629), .B(n2741), .ZN(n4294) );
  INV_X1 U3201 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4293) );
  NOR2_X2 U3203 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2737)
         );
  NAND2_X1 U3204 ( .A1(n2739), .A2(n2758), .ZN(n2746) );
  NAND2_X1 U3205 ( .A1(n2746), .A2(n2899), .ZN(n2740) );
  XNOR2_X1 U3206 ( .A(n2740), .B(IR_REG_17__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U3207 ( .A1(n5156), .A2(REG2_REG_17__SCAN_IN), .ZN(n2744) );
  OAI21_X1 U3208 ( .B1(n5156), .B2(REG2_REG_17__SCAN_IN), .A(n2744), .ZN(n5162) );
  INV_X1 U3209 ( .A(n5162), .ZN(n2742) );
  NAND2_X1 U32100 ( .A1(n2741), .A2(n4299), .ZN(n5159) );
  NAND2_X1 U32110 ( .A1(n2742), .A2(n5159), .ZN(n2743) );
  AOI21_X1 U32120 ( .B1(n4294), .B2(n4293), .A(n2743), .ZN(n5160) );
  INV_X1 U32130 ( .A(n2744), .ZN(n2745) );
  NAND2_X1 U32140 ( .A1(n2751), .A2(n2899), .ZN(n2748) );
  XNOR2_X1 U32150 ( .A(n2748), .B(IR_REG_18__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U32160 ( .A1(n5327), .A2(REG2_REG_18__SCAN_IN), .ZN(n2749) );
  OAI21_X1 U32170 ( .B1(n5327), .B2(REG2_REG_18__SCAN_IN), .A(n2749), .ZN(
        n2846) );
  NOR2_X1 U32180 ( .A1(n2847), .A2(n2846), .ZN(n2845) );
  NOR2_X1 U32190 ( .A1(n2845), .A2(n2750), .ZN(n2757) );
  INV_X1 U32200 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2755) );
  INV_X1 U32210 ( .A(n2753), .ZN(n2752) );
  NAND2_X1 U32220 ( .A1(n2752), .A2(IR_REG_19__SCAN_IN), .ZN(n2754) );
  MUX2_X1 U32230 ( .A(n2755), .B(REG2_REG_19__SCAN_IN), .S(n5211), .Z(n2756)
         );
  XNOR2_X1 U32240 ( .A(n2757), .B(n2756), .ZN(n2796) );
  INV_X2 U32250 ( .A(IR_REG_17__SCAN_IN), .ZN(n4980) );
  NAND4_X1 U32260 ( .A1(n4985), .A2(n2759), .A3(n4981), .A4(n4980), .ZN(n2760)
         );
  INV_X1 U32270 ( .A(n2789), .ZN(n2764) );
  INV_X1 U32280 ( .A(IR_REG_22__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U32290 ( .A1(n2764), .A2(n2763), .ZN(n2767) );
  NAND2_X1 U32300 ( .A1(n2767), .A2(n2899), .ZN(n2780) );
  NAND2_X1 U32310 ( .A1(n2780), .A2(n2779), .ZN(n2782) );
  INV_X1 U32320 ( .A(n2871), .ZN(n2874) );
  INV_X1 U32330 ( .A(IR_REG_24__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U32340 ( .A1(n2779), .A2(n4796), .ZN(n2766) );
  INV_X1 U32350 ( .A(n2770), .ZN(n2768) );
  NAND2_X1 U32360 ( .A1(n2768), .A2(IR_REG_31__SCAN_IN), .ZN(n2769) );
  INV_X1 U32370 ( .A(IR_REG_25__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U32380 ( .A1(n2771), .A2(n2772), .ZN(n2870) );
  NAND2_X1 U32390 ( .A1(n2772), .A2(n2899), .ZN(n2773) );
  MUX2_X1 U32400 ( .A(n2899), .B(n2773), .S(IR_REG_26__SCAN_IN), .Z(n2777) );
  NOR2_X1 U32410 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2775) );
  NOR2_X1 U32420 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2774) );
  NAND2_X1 U32430 ( .A1(n2778), .A2(n4671), .ZN(n2959) );
  OR2_X1 U32440 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  NAND2_X1 U32450 ( .A1(n2782), .A2(n2781), .ZN(n3068) );
  INV_X1 U32460 ( .A(n3015), .ZN(n3000) );
  INV_X1 U32470 ( .A(n3068), .ZN(n2783) );
  NAND2_X1 U32480 ( .A1(n2783), .A2(STATE_REG_SCAN_IN), .ZN(n4236) );
  NAND2_X1 U32490 ( .A1(n3000), .A2(n4236), .ZN(n2837) );
  INV_X1 U32500 ( .A(IR_REG_28__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U32510 ( .A1(n2789), .A2(n2899), .ZN(n2790) );
  XNOR2_X1 U32520 ( .A(n2790), .B(n2763), .ZN(n2891) );
  INV_X1 U32530 ( .A(n2891), .ZN(n4234) );
  NAND2_X1 U32540 ( .A1(n2511), .A2(n2899), .ZN(n2791) );
  MUX2_X1 U32550 ( .A(n2899), .B(n2791), .S(IR_REG_21__SCAN_IN), .Z(n2792) );
  NAND2_X1 U32560 ( .A1(n2792), .A2(n2789), .ZN(n4167) );
  NAND2_X1 U32570 ( .A1(n2996), .A2(n3068), .ZN(n2793) );
  AND2_X1 U32580 ( .A1(n2488), .A2(n2793), .ZN(n2835) );
  NAND2_X1 U32590 ( .A1(n2837), .A2(n2835), .ZN(n5106) );
  OR2_X1 U32600 ( .A1(n3004), .A2(n5183), .ZN(n4231) );
  NAND2_X1 U32610 ( .A1(n2796), .A2(n2795), .ZN(n2842) );
  INV_X1 U32620 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5278) );
  INV_X1 U32630 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2798) );
  MUX2_X1 U32640 ( .A(n2798), .B(REG1_REG_1__SCAN_IN), .S(n2797), .Z(n5112) );
  NAND2_X1 U32650 ( .A1(n5167), .A2(REG1_REG_0__SCAN_IN), .ZN(n5111) );
  NOR2_X1 U32660 ( .A1(n5110), .A2(n2799), .ZN(n5173) );
  INV_X1 U32670 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2801) );
  MUX2_X1 U32680 ( .A(n2801), .B(REG1_REG_2__SCAN_IN), .S(n2800), .Z(n5175) );
  INV_X1 U32690 ( .A(n2803), .ZN(n2802) );
  NAND2_X1 U32700 ( .A1(n5075), .A2(n2802), .ZN(n2804) );
  NAND2_X1 U32710 ( .A1(n2804), .A2(n4260), .ZN(n2805) );
  INV_X1 U32720 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U32730 ( .A1(n5126), .A2(REG1_REG_5__SCAN_IN), .ZN(n2806) );
  OAI21_X1 U32740 ( .B1(n5126), .B2(REG1_REG_5__SCAN_IN), .A(n2806), .ZN(n5124) );
  NOR2_X1 U32750 ( .A1(n5123), .A2(n2807), .ZN(n2808) );
  INV_X1 U32760 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2886) );
  NOR2_X1 U32770 ( .A1(n2808), .A2(n3164), .ZN(n2809) );
  XNOR2_X1 U32780 ( .A(n5137), .B(REG1_REG_7__SCAN_IN), .ZN(n5135) );
  INV_X1 U32790 ( .A(n5137), .ZN(n2811) );
  INV_X1 U32800 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2810) );
  INV_X1 U32810 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3083) );
  INV_X1 U32820 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2813) );
  MUX2_X1 U32830 ( .A(n2813), .B(REG1_REG_9__SCAN_IN), .S(n4677), .Z(n3233) );
  NOR2_X1 U32840 ( .A1(n2815), .A2(n3413), .ZN(n2816) );
  INV_X1 U32850 ( .A(REG1_REG_10__SCAN_IN), .ZN(n5262) );
  XNOR2_X1 U32860 ( .A(n2815), .B(n3413), .ZN(n3415) );
  NOR2_X1 U32870 ( .A1(n5262), .A2(n3415), .ZN(n3414) );
  NOR2_X1 U32880 ( .A1(n2816), .A2(n3414), .ZN(n3488) );
  INV_X1 U32890 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5269) );
  AOI22_X1 U32900 ( .A1(n4676), .A2(n5269), .B1(REG1_REG_11__SCAN_IN), .B2(
        n3492), .ZN(n3489) );
  NOR2_X1 U32910 ( .A1(n2817), .A2(n3671), .ZN(n2818) );
  INV_X1 U32920 ( .A(n4274), .ZN(n2821) );
  INV_X1 U32930 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2819) );
  MUX2_X1 U32940 ( .A(n2819), .B(REG1_REG_13__SCAN_IN), .S(n4675), .Z(n4273)
         );
  INV_X1 U32950 ( .A(n4273), .ZN(n2820) );
  NAND2_X1 U32960 ( .A1(n2821), .A2(n2820), .ZN(n4271) );
  NAND2_X1 U32970 ( .A1(n4675), .A2(REG1_REG_13__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U32980 ( .A1(n4271), .A2(n2822), .ZN(n2824) );
  INV_X1 U32990 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4281) );
  NOR2_X1 U33000 ( .A1(n2825), .A2(n4284), .ZN(n2826) );
  NAND2_X1 U33010 ( .A1(n5150), .A2(REG1_REG_15__SCAN_IN), .ZN(n2827) );
  OAI21_X1 U33020 ( .B1(n5150), .B2(REG1_REG_15__SCAN_IN), .A(n2827), .ZN(
        n5143) );
  AND2_X1 U33030 ( .A1(n5150), .A2(REG1_REG_15__SCAN_IN), .ZN(n2828) );
  NOR2_X1 U33040 ( .A1(n5142), .A2(n2828), .ZN(n2829) );
  XNOR2_X1 U33050 ( .A(n2829), .B(n3629), .ZN(n4292) );
  INV_X1 U33060 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U33070 ( .A1(n4292), .A2(n4626), .ZN(n4291) );
  NAND2_X1 U33080 ( .A1(n2829), .A2(n4299), .ZN(n2830) );
  NAND2_X1 U33090 ( .A1(n4291), .A2(n2830), .ZN(n5154) );
  NOR2_X1 U33100 ( .A1(n5156), .A2(REG1_REG_17__SCAN_IN), .ZN(n2831) );
  AOI21_X1 U33110 ( .B1(REG1_REG_17__SCAN_IN), .B2(n5156), .A(n2831), .ZN(
        n5155) );
  NAND2_X1 U33120 ( .A1(n5154), .A2(n5155), .ZN(n5153) );
  INV_X1 U33130 ( .A(n2831), .ZN(n2832) );
  NAND2_X1 U33140 ( .A1(n5327), .A2(REG1_REG_18__SCAN_IN), .ZN(n2833) );
  OAI21_X1 U33150 ( .B1(n5327), .B2(REG1_REG_18__SCAN_IN), .A(n2833), .ZN(
        n2843) );
  INV_X1 U33160 ( .A(REG1_REG_19__SCAN_IN), .ZN(n5343) );
  MUX2_X1 U33170 ( .A(n5343), .B(REG1_REG_19__SCAN_IN), .S(n5211), .Z(n2834)
         );
  INV_X1 U33180 ( .A(n5183), .ZN(n4670) );
  INV_X1 U33190 ( .A(n5197), .ZN(n5177) );
  INV_X1 U33200 ( .A(n3004), .ZN(n5184) );
  INV_X1 U33210 ( .A(n2835), .ZN(n2836) );
  INV_X1 U33220 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3736) );
  NOR2_X1 U33230 ( .A1(STATE_REG_SCAN_IN), .A2(n3736), .ZN(n3967) );
  AOI21_X1 U33240 ( .B1(n5196), .B2(ADDR_REG_19__SCAN_IN), .A(n3967), .ZN(
        n2838) );
  OAI21_X1 U33250 ( .B1(n5211), .B2(n5181), .A(n2838), .ZN(n2839) );
  AOI21_X1 U33260 ( .B1(n2840), .B2(n5177), .A(n2839), .ZN(n2841) );
  NAND2_X1 U33270 ( .A1(n2842), .A2(n2841), .ZN(U3259) );
  AOI21_X1 U33280 ( .B1(n2847), .B2(n2846), .A(n2845), .ZN(n2848) );
  INV_X1 U33290 ( .A(n5181), .ZN(n5207) );
  AOI22_X1 U33300 ( .A1(n2848), .A2(n2795), .B1(n5327), .B2(n5207), .ZN(n2850)
         );
  AND2_X1 U33310 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4048) );
  NAND3_X1 U33320 ( .A1(n2851), .A2(n2850), .A3(n2849), .ZN(U3258) );
  INV_X1 U33330 ( .A(n2879), .ZN(n2852) );
  INV_X2 U33340 ( .A(n4253), .ZN(U4043) );
  INV_X1 U33350 ( .A(DATAI_12_), .ZN(n2853) );
  MUX2_X1 U33360 ( .A(n3671), .B(n2853), .S(U3149), .Z(n2854) );
  INV_X1 U33370 ( .A(n2854), .ZN(U3340) );
  INV_X1 U33380 ( .A(DATAI_14_), .ZN(n2855) );
  MUX2_X1 U33390 ( .A(n2855), .B(n4284), .S(STATE_REG_SCAN_IN), .Z(n2856) );
  INV_X1 U33400 ( .A(n2856), .ZN(U3338) );
  INV_X1 U33410 ( .A(DATAI_22_), .ZN(n2857) );
  MUX2_X1 U33420 ( .A(n2857), .B(n2891), .S(STATE_REG_SCAN_IN), .Z(n2858) );
  INV_X1 U33430 ( .A(n2858), .ZN(U3330) );
  INV_X1 U33440 ( .A(DATAI_28_), .ZN(n2859) );
  MUX2_X1 U33450 ( .A(n2859), .B(n3004), .S(STATE_REG_SCAN_IN), .Z(n2860) );
  INV_X1 U33460 ( .A(n2860), .ZN(U3324) );
  INV_X1 U33470 ( .A(DATAI_23_), .ZN(n2861) );
  AOI21_X1 U33480 ( .B1(n2861), .B2(U3149), .A(n2879), .ZN(U3329) );
  INV_X1 U33490 ( .A(DATAI_16_), .ZN(n2862) );
  MUX2_X1 U33500 ( .A(n2862), .B(n4299), .S(STATE_REG_SCAN_IN), .Z(n2863) );
  INV_X1 U33510 ( .A(n2863), .ZN(U3336) );
  INV_X1 U33520 ( .A(n2892), .ZN(n2866) );
  INV_X1 U3353 ( .A(IR_REG_29__SCAN_IN), .ZN(n2865) );
  NAND2_X1 U33540 ( .A1(n2866), .A2(n2865), .ZN(n2894) );
  INV_X1 U3355 ( .A(IR_REG_30__SCAN_IN), .ZN(n4804) );
  INV_X1 U3356 ( .A(DATAI_30_), .ZN(n2868) );
  MUX2_X1 U3357 ( .A(n2896), .B(n2868), .S(U3149), .Z(n2869) );
  INV_X1 U3358 ( .A(n2869), .ZN(U3322) );
  NAND2_X1 U3359 ( .A1(n2870), .A2(B_REG_SCAN_IN), .ZN(n2872) );
  MUX2_X1 U3360 ( .A(n2872), .B(B_REG_SCAN_IN), .S(n2871), .Z(n2873) );
  NAND2_X1 U3361 ( .A1(n2993), .A2(n3015), .ZN(n5091) );
  INV_X1 U3362 ( .A(D_REG_0__SCAN_IN), .ZN(n2876) );
  INV_X1 U3363 ( .A(n4671), .ZN(n2877) );
  NAND2_X1 U3364 ( .A1(n2877), .A2(n2874), .ZN(n2926) );
  INV_X1 U3365 ( .A(n2926), .ZN(n2875) );
  AOI22_X1 U3366 ( .A1(n5091), .A2(n2876), .B1(n2879), .B2(n2875), .ZN(U3458)
         );
  INV_X1 U3367 ( .A(D_REG_1__SCAN_IN), .ZN(n2989) );
  NAND2_X1 U3368 ( .A1(n2877), .A2(n2870), .ZN(n2991) );
  INV_X1 U3369 ( .A(n2991), .ZN(n2878) );
  AOI22_X1 U3370 ( .A1(n5091), .A2(n2989), .B1(n2879), .B2(n2878), .ZN(U3459)
         );
  NOR2_X1 U3371 ( .A1(n5196), .A2(U4043), .ZN(U3148) );
  AOI21_X1 U3372 ( .B1(n2882), .B2(n2881), .A(n2880), .ZN(n2889) );
  AND2_X1 U3373 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n4060) );
  AOI21_X1 U3374 ( .B1(n5196), .B2(ADDR_REG_6__SCAN_IN), .A(n4060), .ZN(n2883)
         );
  OAI21_X1 U3375 ( .B1(n5181), .B2(n3164), .A(n2883), .ZN(n2888) );
  AOI211_X1 U3376 ( .C1(n2886), .C2(n2885), .A(n2884), .B(n5197), .ZN(n2887)
         );
  AOI211_X1 U3377 ( .C1(n2889), .C2(n2795), .A(n2888), .B(n2887), .ZN(n2890)
         );
  INV_X1 U3378 ( .A(n2890), .ZN(U3246) );
  NAND2_X1 U3379 ( .A1(n2892), .A2(n2899), .ZN(n2893) );
  INV_X1 U3380 ( .A(n2897), .ZN(n4669) );
  NAND2_X1 U3381 ( .A1(n3006), .A2(REG1_REG_1__SCAN_IN), .ZN(n2938) );
  AND2_X4 U3382 ( .A1(n2896), .A2(n2897), .ZN(n3046) );
  NAND2_X1 U3383 ( .A1(n3046), .A2(REG0_REG_1__SCAN_IN), .ZN(n2935) );
  NAND2_X2 U3384 ( .A1(n2898), .A2(n2897), .ZN(n3156) );
  AND2_X4 U3385 ( .A1(n2898), .A2(n4669), .ZN(n3007) );
  NAND2_X1 U3386 ( .A1(n3004), .A2(n2996), .ZN(n4546) );
  NAND2_X1 U3387 ( .A1(n5211), .A2(n4234), .ZN(n2902) );
  AND2_X4 U3388 ( .A1(n2956), .A2(n2902), .ZN(n3810) );
  AND2_X1 U3389 ( .A1(n2996), .A2(n5211), .ZN(n2903) );
  NAND2_X1 U3390 ( .A1(n2923), .A2(n2903), .ZN(n2999) );
  INV_X1 U3391 ( .A(n2999), .ZN(n2904) );
  INV_X1 U3392 ( .A(n2923), .ZN(n5212) );
  NAND2_X1 U3393 ( .A1(n5212), .A2(n4673), .ZN(n2906) );
  NAND2_X1 U3394 ( .A1(n4674), .A2(n4234), .ZN(n2905) );
  NAND2_X1 U3395 ( .A1(n3006), .A2(REG1_REG_0__SCAN_IN), .ZN(n2910) );
  NAND2_X1 U3396 ( .A1(n3007), .A2(REG3_REG_0__SCAN_IN), .ZN(n2909) );
  NAND2_X1 U3397 ( .A1(n3046), .A2(REG0_REG_0__SCAN_IN), .ZN(n2907) );
  OR2_X1 U3398 ( .A1(n2971), .A2(n3094), .ZN(n4077) );
  NAND2_X1 U3399 ( .A1(n2971), .A2(n3094), .ZN(n4075) );
  NAND2_X1 U3400 ( .A1(n4077), .A2(n4075), .ZN(n4157) );
  OAI21_X1 U3401 ( .B1(n5340), .B2(n4501), .A(n4157), .ZN(n2911) );
  OAI21_X1 U3402 ( .B1(n2981), .B2(n4546), .A(n2911), .ZN(n5213) );
  AOI21_X1 U3403 ( .B1(n2947), .B2(n3094), .A(n5213), .ZN(n5215) );
  NAND2_X1 U3404 ( .A1(n4501), .A2(n2996), .ZN(n3069) );
  INV_X1 U3405 ( .A(n2993), .ZN(n2922) );
  NOR2_X1 U3406 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_27__SCAN_IN), .ZN(n2915) );
  NOR4_X1 U3407 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2914) );
  NOR4_X1 U3408 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2913) );
  NOR4_X1 U3409 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2912) );
  AND4_X1 U3410 ( .A1(n2915), .A2(n2914), .A3(n2913), .A4(n2912), .ZN(n2921)
         );
  NOR4_X1 U3411 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2919) );
  NOR4_X1 U3412 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2918) );
  NOR4_X1 U3413 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2917) );
  NOR4_X1 U3414 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2916) );
  AND4_X1 U3415 ( .A1(n2919), .A2(n2918), .A3(n2917), .A4(n2916), .ZN(n2920)
         );
  NAND2_X1 U3416 ( .A1(n2921), .A2(n2920), .ZN(n2990) );
  NAND2_X1 U3417 ( .A1(n2922), .A2(n2990), .ZN(n2925) );
  NAND2_X2 U3418 ( .A1(n2947), .A2(n2923), .ZN(n5338) );
  OAI21_X1 U3419 ( .B1(n2993), .B2(D_REG_1__SCAN_IN), .A(n2991), .ZN(n2924) );
  INV_X1 U3420 ( .A(n3201), .ZN(n2995) );
  NAND2_X1 U3421 ( .A1(n5342), .A2(REG1_REG_0__SCAN_IN), .ZN(n2927) );
  OAI21_X1 U3422 ( .B1(n5215), .B2(n5342), .A(n2927), .ZN(U3518) );
  INV_X1 U3423 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2931) );
  INV_X1 U3424 ( .A(n5215), .ZN(n2929) );
  NAND2_X1 U3425 ( .A1(n2929), .A2(n5348), .ZN(n2930) );
  OAI21_X1 U3426 ( .B1(n5348), .B2(n2931), .A(n2930), .ZN(U3467) );
  INV_X1 U3427 ( .A(n4162), .ZN(n2932) );
  NAND2_X1 U3428 ( .A1(n2932), .A2(n5219), .ZN(n2934) );
  NAND2_X1 U3429 ( .A1(n2981), .A2(n3099), .ZN(n3026) );
  NAND4_X2 U3430 ( .A1(n2938), .A2(n2937), .A3(n2936), .A4(n2935), .ZN(n3002)
         );
  NAND2_X1 U3431 ( .A1(n3002), .A2(n2980), .ZN(n4076) );
  NAND2_X1 U3432 ( .A1(n3026), .A2(n4076), .ZN(n2941) );
  INV_X1 U3433 ( .A(n2941), .ZN(n4161) );
  INV_X1 U3434 ( .A(n3094), .ZN(n2939) );
  NOR2_X1 U3435 ( .A1(n2971), .A2(n2939), .ZN(n2940) );
  NAND2_X1 U3436 ( .A1(n2941), .A2(n2940), .ZN(n3021) );
  NAND3_X1 U3437 ( .A1(n3021), .A2(n3094), .A3(n5340), .ZN(n2942) );
  NAND2_X1 U3438 ( .A1(n5184), .A2(n2996), .ZN(n4548) );
  OAI211_X1 U3439 ( .C1(n4161), .C2(n4554), .A(n2942), .B(n4548), .ZN(n2952)
         );
  NAND2_X1 U3440 ( .A1(n3046), .A2(REG0_REG_2__SCAN_IN), .ZN(n2946) );
  NAND2_X1 U3441 ( .A1(n3006), .A2(REG1_REG_2__SCAN_IN), .ZN(n2945) );
  OR2_X1 U3442 ( .A1(n3156), .A2(n5227), .ZN(n2944) );
  NAND2_X1 U3443 ( .A1(n3007), .A2(REG3_REG_2__SCAN_IN), .ZN(n2943) );
  AOI22_X1 U3444 ( .A1(n4252), .A2(n4525), .B1(n3099), .B2(n4560), .ZN(n2948)
         );
  OAI21_X1 U3445 ( .B1(n3027), .B2(n4554), .A(n2948), .ZN(n2951) );
  AOI22_X1 U3446 ( .A1(n3021), .A2(n5340), .B1(n2953), .B2(n4501), .ZN(n2949)
         );
  NOR2_X1 U3447 ( .A1(n2949), .A2(n4161), .ZN(n2950) );
  AOI211_X1 U3448 ( .C1(n4254), .C2(n2952), .A(n2951), .B(n2950), .ZN(n5224)
         );
  INV_X1 U3449 ( .A(n5338), .ZN(n5277) );
  NAND2_X1 U3450 ( .A1(n5344), .A2(n5277), .ZN(n4628) );
  INV_X1 U3451 ( .A(n4628), .ZN(n3308) );
  INV_X1 U3452 ( .A(n3035), .ZN(n2954) );
  AOI21_X1 U3453 ( .B1(n3099), .B2(n3094), .A(n2954), .ZN(n5221) );
  AOI22_X1 U3454 ( .A1(n3308), .A2(n5221), .B1(n5342), .B2(REG1_REG_1__SCAN_IN), .ZN(n2955) );
  OAI21_X1 U3455 ( .B1(n5224), .B2(n5342), .A(n2955), .ZN(U3519) );
  MUX2_X1 U3456 ( .A(n2800), .B(DATAI_2_), .S(n4162), .Z(n3036) );
  NAND2_X1 U3457 ( .A1(n3044), .A2(n3036), .ZN(n2961) );
  INV_X1 U34580 ( .A(n2957), .ZN(n2958) );
  NAND2_X1 U34590 ( .A1(n2976), .A2(n4252), .ZN(n2960) );
  NAND2_X1 U3460 ( .A1(n2961), .A2(n2960), .ZN(n2962) );
  XNOR2_X1 U3461 ( .A(n2962), .B(n3810), .ZN(n2967) );
  INV_X1 U3462 ( .A(n2967), .ZN(n2965) );
  OR2_X2 U3463 ( .A1(n5338), .A2(n4674), .ZN(n3292) );
  NOR2_X1 U3464 ( .A1(n3128), .A2(n3106), .ZN(n2963) );
  INV_X1 U3465 ( .A(n2966), .ZN(n2964) );
  INV_X1 U3466 ( .A(n2959), .ZN(n2968) );
  NAND2_X1 U34670 ( .A1(n2970), .A2(n2969), .ZN(n3093) );
  INV_X1 U3468 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U34690 ( .A1(n3044), .A2(n3094), .ZN(n2973) );
  OAI211_X1 U3470 ( .C1(n2959), .C2(n5102), .A(n2973), .B(n2972), .ZN(n3092)
         );
  NAND2_X1 U34710 ( .A1(n3093), .A2(n3092), .ZN(n2975) );
  NAND2_X1 U3472 ( .A1(n2973), .A2(n3810), .ZN(n2974) );
  NAND2_X1 U34730 ( .A1(n2975), .A2(n2974), .ZN(n3097) );
  NAND2_X1 U3474 ( .A1(n2976), .A2(n3002), .ZN(n2978) );
  NAND2_X1 U34750 ( .A1(n3044), .A2(n3099), .ZN(n2977) );
  NAND2_X1 U3476 ( .A1(n2978), .A2(n2977), .ZN(n2979) );
  XNOR2_X1 U34770 ( .A(n2979), .B(n3810), .ZN(n2982) );
  OAI22_X1 U3478 ( .A1(n2492), .A2(n2981), .B1(n2491), .B2(n2980), .ZN(n2983)
         );
  XNOR2_X1 U34790 ( .A(n2982), .B(n2983), .ZN(n3098) );
  INV_X1 U3480 ( .A(n2982), .ZN(n2984) );
  NAND2_X1 U34810 ( .A1(n2984), .A2(n2983), .ZN(n2985) );
  INV_X1 U3482 ( .A(n3039), .ZN(n2987) );
  AOI21_X1 U34830 ( .B1(n2988), .B2(n2986), .A(n2987), .ZN(n3019) );
  NOR2_X1 U3484 ( .A1(n2990), .A2(n2989), .ZN(n2992) );
  OAI21_X1 U34850 ( .B1(n2993), .B2(n2992), .A(n2991), .ZN(n2994) );
  INV_X1 U3486 ( .A(n2994), .ZN(n3203) );
  NAND2_X1 U34870 ( .A1(n2995), .A2(n3203), .ZN(n3003) );
  INV_X1 U3488 ( .A(n3003), .ZN(n3001) );
  NAND2_X1 U34890 ( .A1(n3001), .A2(n3015), .ZN(n3012) );
  INV_X1 U3490 ( .A(n2996), .ZN(n2997) );
  NAND3_X1 U34910 ( .A1(n3013), .A2(n2997), .A3(n4581), .ZN(n2998) );
  NOR2_X1 U3492 ( .A1(n3000), .A2(n2999), .ZN(n4232) );
  AND2_X1 U34930 ( .A1(n3001), .A2(n4232), .ZN(n3005) );
  NAND2_X1 U3494 ( .A1(n3003), .A2(n3013), .ZN(n3071) );
  NAND2_X1 U34950 ( .A1(n3071), .A2(n3202), .ZN(n3100) );
  AOI22_X1 U3496 ( .A1(n5284), .A2(n3002), .B1(REG3_REG_2__SCAN_IN), .B2(n3100), .ZN(n3018) );
  NAND2_X1 U34970 ( .A1(n3006), .A2(REG1_REG_3__SCAN_IN), .ZN(n3011) );
  INV_X1 U3498 ( .A(REG3_REG_3__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U34990 ( .A1(n3007), .A2(n5229), .ZN(n3010) );
  NAND2_X1 U3500 ( .A1(n3353), .A2(REG2_REG_3__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U35010 ( .A1(n3046), .A2(REG0_REG_3__SCAN_IN), .ZN(n3008) );
  OR2_X1 U3502 ( .A1(n3012), .A2(n4581), .ZN(n3016) );
  INV_X1 U35030 ( .A(n3013), .ZN(n3014) );
  AOI22_X1 U3504 ( .A1(n5296), .A2(n4251), .B1(n5282), .B2(n3036), .ZN(n3017)
         );
  OAI211_X1 U35050 ( .C1(n3019), .C2(n5291), .A(n3018), .B(n3017), .ZN(U3234)
         );
  NAND2_X1 U35060 ( .A1(n3002), .A2(n3099), .ZN(n3020) );
  INV_X1 U35070 ( .A(n4252), .ZN(n3022) );
  NAND2_X1 U35080 ( .A1(n3106), .A2(n4252), .ZN(n4082) );
  NAND2_X1 U35090 ( .A1(n3025), .A2(n3024), .ZN(n3108) );
  OAI21_X1 U35100 ( .B1(n3025), .B2(n3024), .A(n3108), .ZN(n3033) );
  NAND2_X1 U35110 ( .A1(n3027), .A2(n3026), .ZN(n3028) );
  NAND2_X1 U35120 ( .A1(n3028), .A2(n3023), .ZN(n3109) );
  OAI21_X1 U35130 ( .B1(n3023), .B2(n3028), .A(n3109), .ZN(n3029) );
  NAND2_X1 U35140 ( .A1(n3029), .A2(n4501), .ZN(n3031) );
  AOI22_X1 U35150 ( .A1(n4525), .A2(n4251), .B1(n3002), .B2(n4504), .ZN(n3030)
         );
  OAI211_X1 U35160 ( .C1(n4581), .C2(n3106), .A(n3031), .B(n3030), .ZN(n3032)
         );
  AOI21_X1 U35170 ( .B1(n5340), .B2(n3033), .A(n3032), .ZN(n5228) );
  INV_X1 U35180 ( .A(n3117), .ZN(n3034) );
  AOI21_X1 U35190 ( .B1(n3036), .B2(n3035), .A(n3034), .ZN(n5225) );
  AOI22_X1 U35200 ( .A1(n3308), .A2(n5225), .B1(n5342), .B2(
        REG1_REG_2__SCAN_IN), .ZN(n3037) );
  OAI21_X1 U35210 ( .B1(n5228), .B2(n5342), .A(n3037), .ZN(U3520) );
  NAND2_X1 U35220 ( .A1(n3039), .A2(n3038), .ZN(n3221) );
  NAND2_X1 U35230 ( .A1(n2976), .A2(n4251), .ZN(n3041) );
  INV_X2 U35240 ( .A(n3872), .ZN(n3826) );
  MUX2_X1 U35250 ( .A(n5075), .B(DATAI_3_), .S(n2488), .Z(n3223) );
  NAND2_X1 U35260 ( .A1(n3044), .A2(n3223), .ZN(n3040) );
  NAND2_X1 U35270 ( .A1(n3041), .A2(n3040), .ZN(n3042) );
  XNOR2_X1 U35280 ( .A(n3042), .B(n3810), .ZN(n3056) );
  INV_X1 U35290 ( .A(n3223), .ZN(n3205) );
  OAI22_X1 U35300 ( .A1(n2493), .A2(n3206), .B1(n3128), .B2(n3205), .ZN(n3054)
         );
  XNOR2_X1 U35310 ( .A(n3056), .B(n3054), .ZN(n3222) );
  MUX2_X1 U35320 ( .A(n5206), .B(DATAI_4_), .S(n2488), .Z(n3240) );
  NAND2_X1 U35330 ( .A1(n2489), .A2(n3240), .ZN(n3052) );
  NAND2_X1 U35340 ( .A1(n2497), .A2(REG1_REG_4__SCAN_IN), .ZN(n3050) );
  NOR2_X1 U35350 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n3045) );
  NOR2_X1 U35360 ( .A1(n3061), .A2(n3045), .ZN(n3073) );
  NAND2_X1 U35370 ( .A1(n3007), .A2(n3073), .ZN(n3049) );
  NAND2_X1 U35380 ( .A1(n3353), .A2(REG2_REG_4__SCAN_IN), .ZN(n3048) );
  NAND2_X1 U35390 ( .A1(n3046), .A2(REG0_REG_4__SCAN_IN), .ZN(n3047) );
  NAND2_X1 U35400 ( .A1(n2976), .A2(n4250), .ZN(n3051) );
  NAND2_X1 U35410 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  XNOR2_X1 U35420 ( .A(n3053), .B(n3810), .ZN(n3122) );
  INV_X1 U35430 ( .A(n4250), .ZN(n3209) );
  OAI22_X1 U35440 ( .A1(n2493), .A2(n3209), .B1(n3875), .B2(n3216), .ZN(n3123)
         );
  XNOR2_X1 U35450 ( .A(n3122), .B(n3123), .ZN(n3059) );
  INV_X1 U35460 ( .A(n3054), .ZN(n3055) );
  NAND2_X1 U35470 ( .A1(n3056), .A2(n3055), .ZN(n3060) );
  AND2_X1 U35480 ( .A1(n3059), .A2(n3060), .ZN(n3057) );
  NAND2_X1 U35490 ( .A1(n3058), .A2(n3057), .ZN(n3171) );
  INV_X1 U35500 ( .A(n5291), .ZN(n4055) );
  NAND2_X1 U35510 ( .A1(n3171), .A2(n4055), .ZN(n3078) );
  AOI21_X1 U35520 ( .B1(n3058), .B2(n3060), .A(n3059), .ZN(n3077) );
  OAI21_X1 U35530 ( .B1(n3061), .B2(REG3_REG_5__SCAN_IN), .A(n3137), .ZN(n3372) );
  INV_X1 U35540 ( .A(n3372), .ZN(n3062) );
  NAND2_X1 U35550 ( .A1(n3007), .A2(n3062), .ZN(n3066) );
  NAND2_X1 U35560 ( .A1(n2496), .A2(REG1_REG_5__SCAN_IN), .ZN(n3065) );
  NAND2_X1 U35570 ( .A1(n3353), .A2(REG2_REG_5__SCAN_IN), .ZN(n3064) );
  NAND2_X1 U35580 ( .A1(n3046), .A2(REG0_REG_5__SCAN_IN), .ZN(n3063) );
  NAND4_X1 U35590 ( .A1(n3066), .A2(n3065), .A3(n3064), .A4(n3063), .ZN(n4249)
         );
  AOI22_X1 U35600 ( .A1(n5296), .A2(n4249), .B1(n5282), .B2(n3240), .ZN(n3076)
         );
  INV_X1 U35610 ( .A(REG3_REG_4__SCAN_IN), .ZN(n3067) );
  NOR2_X1 U35620 ( .A1(STATE_REG_SCAN_IN), .A2(n3067), .ZN(n5195) );
  AND3_X1 U35630 ( .A1(n3069), .A2(n2959), .A3(n3068), .ZN(n3070) );
  NAND2_X1 U35640 ( .A1(n3071), .A2(n3070), .ZN(n3072) );
  INV_X1 U35650 ( .A(n3073), .ZN(n3218) );
  NOR2_X1 U35660 ( .A1(n5300), .A2(n3218), .ZN(n3074) );
  AOI211_X1 U35670 ( .C1(n5284), .C2(n4251), .A(n5195), .B(n3074), .ZN(n3075)
         );
  OAI211_X1 U35680 ( .C1(n3078), .C2(n3077), .A(n3076), .B(n3075), .ZN(U3227)
         );
  AOI211_X1 U35690 ( .C1(n3081), .C2(n3080), .A(n3079), .B(n5200), .ZN(n3089)
         );
  AOI211_X1 U35700 ( .C1(n3084), .C2(n3083), .A(n3082), .B(n5197), .ZN(n3088)
         );
  INV_X1 U35710 ( .A(n4678), .ZN(n3086) );
  AND2_X1 U35720 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n3978) );
  AOI21_X1 U35730 ( .B1(n5196), .B2(ADDR_REG_8__SCAN_IN), .A(n3978), .ZN(n3085) );
  OAI21_X1 U35740 ( .B1(n5181), .B2(n3086), .A(n3085), .ZN(n3087) );
  OR3_X1 U35750 ( .A1(n3089), .A2(n3088), .A3(n3087), .ZN(U3248) );
  NAND2_X1 U35760 ( .A1(n5348), .A2(n5277), .ZN(n4666) );
  INV_X1 U35770 ( .A(n4666), .ZN(n3312) );
  AOI22_X1 U35780 ( .A1(n3312), .A2(n5225), .B1(REG0_REG_2__SCAN_IN), .B2(
        n5345), .ZN(n3090) );
  OAI21_X1 U35790 ( .B1(n5228), .B2(n5345), .A(n3090), .ZN(U3471) );
  AOI22_X1 U35800 ( .A1(n3312), .A2(n5221), .B1(REG0_REG_1__SCAN_IN), .B2(
        n5345), .ZN(n3091) );
  OAI21_X1 U35810 ( .B1(n5224), .B2(n5345), .A(n3091), .ZN(U3469) );
  XNOR2_X1 U3582 ( .A(n3093), .B(n3092), .ZN(n5185) );
  AOI22_X1 U3583 ( .A1(n5296), .A2(n3002), .B1(REG3_REG_0__SCAN_IN), .B2(n3100), .ZN(n3096) );
  NAND2_X1 U3584 ( .A1(n5282), .A2(n3094), .ZN(n3095) );
  OAI211_X1 U3585 ( .C1(n5185), .C2(n5291), .A(n3096), .B(n3095), .ZN(U3229)
         );
  XNOR2_X1 U3586 ( .A(n3098), .B(n3097), .ZN(n3103) );
  AOI22_X1 U3587 ( .A1(n5296), .A2(n4252), .B1(n5282), .B2(n3099), .ZN(n3102)
         );
  AOI22_X1 U3588 ( .A1(n5284), .A2(n4254), .B1(REG3_REG_1__SCAN_IN), .B2(n3100), .ZN(n3101) );
  OAI211_X1 U3589 ( .C1(n3103), .C2(n5291), .A(n3102), .B(n3101), .ZN(U3219)
         );
  NAND2_X1 U3590 ( .A1(n3109), .A2(n4079), .ZN(n3104) );
  NAND2_X1 U3591 ( .A1(n3206), .A2(n3223), .ZN(n3247) );
  NAND2_X1 U3592 ( .A1(n3205), .A2(n4251), .ZN(n4081) );
  AND2_X1 U3593 ( .A1(n3247), .A2(n4081), .ZN(n4158) );
  INV_X1 U3594 ( .A(n3248), .ZN(n3116) );
  AOI22_X1 U3595 ( .A1(n4525), .A2(n4250), .B1(n4252), .B2(n4504), .ZN(n3105)
         );
  OAI21_X1 U3596 ( .B1(n3205), .B2(n4581), .A(n3105), .ZN(n3115) );
  NAND2_X1 U3597 ( .A1(n3022), .A2(n3106), .ZN(n3107) );
  NAND2_X1 U3598 ( .A1(n3108), .A2(n3107), .ZN(n3208) );
  INV_X1 U3599 ( .A(n3208), .ZN(n3111) );
  NAND3_X1 U3600 ( .A1(n3109), .A2(n4501), .A3(n4079), .ZN(n3110) );
  OAI21_X1 U3601 ( .B1(n3111), .B2(n5272), .A(n3110), .ZN(n3113) );
  NOR2_X1 U3602 ( .A1(n3208), .A2(n5272), .ZN(n3112) );
  MUX2_X1 U3603 ( .A(n3113), .B(n3112), .S(n4158), .Z(n3114) );
  AOI211_X1 U3604 ( .C1(n3116), .C2(n4501), .A(n3115), .B(n3114), .ZN(n5232)
         );
  AOI21_X1 U3605 ( .B1(n3223), .B2(n3117), .A(n3217), .ZN(n5230) );
  INV_X1 U3606 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3118) );
  NOR2_X1 U3607 ( .A1(n5348), .A2(n3118), .ZN(n3119) );
  AOI21_X1 U3608 ( .B1(n3312), .B2(n5230), .A(n3119), .ZN(n3120) );
  OAI21_X1 U3609 ( .B1(n5232), .B2(n5345), .A(n3120), .ZN(U3473) );
  AOI22_X1 U3610 ( .A1(n3308), .A2(n5230), .B1(n5342), .B2(REG1_REG_3__SCAN_IN), .ZN(n3121) );
  OAI21_X1 U3611 ( .B1(n5232), .B2(n5342), .A(n3121), .ZN(U3521) );
  INV_X1 U3612 ( .A(n3122), .ZN(n3124) );
  NAND2_X1 U3613 ( .A1(n3124), .A2(n3123), .ZN(n3169) );
  NAND2_X1 U3614 ( .A1(n3171), .A2(n3169), .ZN(n3135) );
  MUX2_X1 U3615 ( .A(n5126), .B(DATAI_5_), .S(n2488), .Z(n3363) );
  NAND2_X1 U3616 ( .A1(n3826), .A2(n3363), .ZN(n3126) );
  NAND2_X1 U3617 ( .A1(n2498), .A2(n4249), .ZN(n3125) );
  NAND2_X1 U3618 ( .A1(n3126), .A2(n3125), .ZN(n3127) );
  XNOR2_X1 U3619 ( .A(n3127), .B(n3873), .ZN(n3132) );
  INV_X1 U3620 ( .A(n3132), .ZN(n3130) );
  INV_X1 U3621 ( .A(n3363), .ZN(n3370) );
  OAI22_X1 U3622 ( .A1(n2493), .A2(n4058), .B1(n3875), .B2(n3370), .ZN(n3131)
         );
  INV_X1 U3623 ( .A(n3131), .ZN(n3129) );
  AND2_X1 U3624 ( .A1(n3130), .A2(n3129), .ZN(n4052) );
  INV_X1 U3625 ( .A(n4052), .ZN(n3133) );
  NAND2_X1 U3626 ( .A1(n3132), .A2(n3131), .ZN(n3168) );
  NAND2_X1 U3627 ( .A1(n3133), .A2(n3168), .ZN(n3134) );
  NOR2_X1 U3628 ( .A1(n3135), .A2(n3134), .ZN(n4054) );
  AOI21_X1 U3629 ( .B1(n3135), .B2(n3134), .A(n4054), .ZN(n3147) );
  NAND2_X1 U3630 ( .A1(n2497), .A2(REG1_REG_6__SCAN_IN), .ZN(n3142) );
  AND2_X1 U3631 ( .A1(n3137), .A2(n3136), .ZN(n3138) );
  NOR2_X1 U3632 ( .A1(n3176), .A2(n3138), .ZN(n4061) );
  NAND2_X1 U3633 ( .A1(n3007), .A2(n4061), .ZN(n3141) );
  NAND2_X1 U3634 ( .A1(n3353), .A2(REG2_REG_6__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U3635 ( .A1(n3046), .A2(REG0_REG_6__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U3636 ( .A1(n5296), .A2(n4248), .B1(n5282), .B2(n3363), .ZN(n3146)
         );
  INV_X1 U3637 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3143) );
  NOR2_X1 U3638 ( .A1(STATE_REG_SCAN_IN), .A2(n3143), .ZN(n5121) );
  NOR2_X1 U3639 ( .A1(n5300), .A2(n3372), .ZN(n3144) );
  AOI211_X1 U3640 ( .C1(n5284), .C2(n4250), .A(n5121), .B(n3144), .ZN(n3145)
         );
  OAI211_X1 U3641 ( .C1(n3147), .C2(n5291), .A(n3146), .B(n3145), .ZN(U3224)
         );
  NAND2_X1 U3642 ( .A1(n3176), .A2(REG3_REG_7__SCAN_IN), .ZN(n3189) );
  INV_X1 U3643 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3600) );
  INV_X1 U3644 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3719) );
  INV_X1 U3645 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4928) );
  INV_X1 U3646 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3800) );
  INV_X1 U3647 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U3648 ( .A1(REG3_REG_26__SCAN_IN), .A2(REG3_REG_27__SCAN_IN), .ZN(
        n3152) );
  INV_X1 U3649 ( .A(n3861), .ZN(n3153) );
  NAND2_X1 U3650 ( .A1(n3153), .A2(REG3_REG_28__SCAN_IN), .ZN(n3880) );
  INV_X1 U3651 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3154) );
  NAND2_X1 U3652 ( .A1(n3861), .A2(n3154), .ZN(n3155) );
  NAND2_X1 U3653 ( .A1(n3880), .A2(n3155), .ZN(n4315) );
  INV_X1 U3654 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U3655 ( .A1(n3006), .A2(REG1_REG_28__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U3656 ( .A1(n3353), .A2(REG2_REG_28__SCAN_IN), .ZN(n3157) );
  OAI211_X1 U3657 ( .C1(n3159), .C2(n3884), .A(n3158), .B(n3157), .ZN(n3160)
         );
  INV_X1 U3658 ( .A(n3160), .ZN(n3161) );
  NAND2_X1 U3659 ( .A1(n4253), .A2(DATAO_REG_28__SCAN_IN), .ZN(n3163) );
  OAI21_X1 U3660 ( .B1(n4324), .B2(n4253), .A(n3163), .ZN(U3578) );
  NAND2_X1 U3661 ( .A1(n2976), .A2(n4248), .ZN(n3166) );
  INV_X1 U3662 ( .A(n3164), .ZN(n5074) );
  MUX2_X1 U3663 ( .A(n5074), .B(DATAI_6_), .S(n2488), .Z(n4057) );
  NAND2_X1 U3664 ( .A1(n2489), .A2(n4057), .ZN(n3165) );
  NAND2_X1 U3665 ( .A1(n3166), .A2(n3165), .ZN(n3167) );
  XNOR2_X1 U3666 ( .A(n3167), .B(n3810), .ZN(n3175) );
  INV_X1 U3667 ( .A(n4248), .ZN(n3263) );
  INV_X1 U3668 ( .A(n4057), .ZN(n3245) );
  OAI22_X1 U3669 ( .A1(n2493), .A2(n3263), .B1(n3875), .B2(n3245), .ZN(n3173)
         );
  XNOR2_X1 U3670 ( .A(n3175), .B(n3173), .ZN(n4053) );
  AND3_X1 U3671 ( .A1(n4053), .A2(n3169), .A3(n3168), .ZN(n3170) );
  NAND2_X1 U3672 ( .A1(n4053), .A2(n4052), .ZN(n3172) );
  INV_X1 U3673 ( .A(n3186), .ZN(n3185) );
  INV_X1 U3674 ( .A(n3173), .ZN(n3174) );
  NAND2_X1 U3675 ( .A1(n3175), .A2(n3174), .ZN(n3187) );
  NAND2_X1 U3676 ( .A1(n2497), .A2(REG1_REG_7__SCAN_IN), .ZN(n3181) );
  OR2_X1 U3677 ( .A1(n3176), .A2(REG3_REG_7__SCAN_IN), .ZN(n3177) );
  AND2_X1 U3678 ( .A1(n3189), .A2(n3177), .ZN(n3268) );
  NAND2_X1 U3679 ( .A1(n3007), .A2(n3268), .ZN(n3180) );
  NAND2_X1 U3680 ( .A1(n3353), .A2(REG2_REG_7__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U3681 ( .A1(n3046), .A2(REG0_REG_7__SCAN_IN), .ZN(n3178) );
  NAND4_X1 U3682 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n4247)
         );
  NAND2_X1 U3683 ( .A1(n2498), .A2(n4247), .ZN(n3183) );
  MUX2_X1 U3684 ( .A(n5137), .B(DATAI_7_), .S(n2488), .Z(n3274) );
  NAND2_X1 U3685 ( .A1(n3826), .A2(n3274), .ZN(n3182) );
  NAND2_X1 U3686 ( .A1(n3183), .A2(n3182), .ZN(n3184) );
  XNOR2_X1 U3687 ( .A(n3184), .B(n3810), .ZN(n3316) );
  INV_X1 U3688 ( .A(n3274), .ZN(n3261) );
  OAI22_X1 U3689 ( .A1(n2493), .A2(n3976), .B1(n3875), .B2(n3261), .ZN(n3317)
         );
  XNOR2_X1 U3690 ( .A(n3316), .B(n3317), .ZN(n3188) );
  AOI21_X1 U3691 ( .B1(n3185), .B2(n3187), .A(n3188), .ZN(n3200) );
  NAND2_X1 U3692 ( .A1(n3320), .A2(n4055), .ZN(n3199) );
  NAND2_X1 U3693 ( .A1(n2496), .A2(REG1_REG_8__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U3694 ( .A1(n3189), .A2(n4921), .ZN(n3190) );
  AND2_X1 U3695 ( .A1(n3280), .A2(n3190), .ZN(n3979) );
  NAND2_X1 U3696 ( .A1(n3007), .A2(n3979), .ZN(n3193) );
  NAND2_X1 U3697 ( .A1(n3353), .A2(REG2_REG_8__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U3698 ( .A1(n3046), .A2(REG0_REG_8__SCAN_IN), .ZN(n3191) );
  NAND4_X1 U3699 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n4246)
         );
  AOI22_X1 U3700 ( .A1(n5296), .A2(n4246), .B1(n5282), .B2(n3274), .ZN(n3198)
         );
  INV_X1 U3701 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3195) );
  NOR2_X1 U3702 ( .A1(STATE_REG_SCAN_IN), .A2(n3195), .ZN(n5133) );
  NOR2_X1 U3703 ( .A1(n4071), .A2(n3263), .ZN(n3196) );
  AOI211_X1 U3704 ( .C1(n4068), .C2(n3268), .A(n5133), .B(n3196), .ZN(n3197)
         );
  OAI211_X1 U3705 ( .C1(n3200), .C2(n3199), .A(n3198), .B(n3197), .ZN(U3210)
         );
  NAND3_X1 U3706 ( .A1(n3203), .A2(n3202), .A3(n3201), .ZN(n3204) );
  NAND2_X2 U3707 ( .A1(n3204), .A2(n5307), .ZN(n4545) );
  NOR2_X1 U3708 ( .A1(n4251), .A2(n3223), .ZN(n3207) );
  OAI22_X1 U3709 ( .A1(n3208), .A2(n3207), .B1(n3206), .B2(n3205), .ZN(n3239)
         );
  NAND2_X1 U3710 ( .A1(n3209), .A2(n3240), .ZN(n3246) );
  NAND2_X1 U3711 ( .A1(n3216), .A2(n4250), .ZN(n4089) );
  NAND2_X1 U3712 ( .A1(n3246), .A2(n4089), .ZN(n3238) );
  XNOR2_X1 U3713 ( .A(n3239), .B(n3238), .ZN(n3215) );
  NAND2_X1 U3714 ( .A1(n3248), .A2(n3247), .ZN(n3210) );
  INV_X1 U3715 ( .A(n3238), .ZN(n4145) );
  XNOR2_X1 U3716 ( .A(n3210), .B(n4145), .ZN(n3213) );
  AOI22_X1 U3717 ( .A1(n4504), .A2(n4251), .B1(n4249), .B2(n4525), .ZN(n3211)
         );
  OAI21_X1 U3718 ( .B1(n3216), .B2(n4581), .A(n3211), .ZN(n3212) );
  AOI21_X1 U3719 ( .B1(n3213), .B2(n4501), .A(n3212), .ZN(n3214) );
  OAI21_X1 U3720 ( .B1(n3215), .B2(n5272), .A(n3214), .ZN(n5235) );
  NAND2_X1 U3721 ( .A1(n3217), .A2(n3216), .ZN(n3368) );
  OAI211_X1 U3722 ( .C1(n3217), .C2(n3216), .A(n3368), .B(n5277), .ZN(n5233)
         );
  OAI22_X1 U3723 ( .A1(n5233), .A2(n4674), .B1(n5307), .B2(n3218), .ZN(n3219)
         );
  OAI21_X1 U3724 ( .B1(n5235), .B2(n3219), .A(n4545), .ZN(n3220) );
  OAI21_X1 U3725 ( .B1(n5203), .B2(n4545), .A(n3220), .ZN(U3286) );
  OAI21_X1 U3726 ( .B1(n3222), .B2(n3221), .A(n3058), .ZN(n3227) );
  AOI22_X1 U3727 ( .A1(n5296), .A2(n4250), .B1(n5282), .B2(n3223), .ZN(n3225)
         );
  NOR2_X1 U3728 ( .A1(STATE_REG_SCAN_IN), .A2(n5229), .ZN(n4259) );
  AOI21_X1 U3729 ( .B1(n5284), .B2(n4252), .A(n4259), .ZN(n3224) );
  OAI211_X1 U3730 ( .C1(REG3_REG_3__SCAN_IN), .C2(n5300), .A(n3225), .B(n3224), 
        .ZN(n3226) );
  AOI21_X1 U3731 ( .B1(n3227), .B2(n4055), .A(n3226), .ZN(n3228) );
  INV_X1 U3732 ( .A(n3228), .ZN(U3215) );
  AOI21_X1 U3733 ( .B1(n3230), .B2(n2522), .A(n3229), .ZN(n3236) );
  NOR2_X1 U3734 ( .A1(STATE_REG_SCAN_IN), .A2(n4943), .ZN(n4018) );
  AOI21_X1 U3735 ( .B1(n5196), .B2(ADDR_REG_9__SCAN_IN), .A(n4018), .ZN(n3231)
         );
  OAI21_X1 U3736 ( .B1(n5181), .B2(n2720), .A(n3231), .ZN(n3235) );
  AOI211_X1 U3737 ( .C1(n2523), .C2(n3233), .A(n5197), .B(n3232), .ZN(n3234)
         );
  AOI211_X1 U3738 ( .C1(n2795), .C2(n3236), .A(n3235), .B(n3234), .ZN(n3237)
         );
  INV_X1 U3739 ( .A(n3237), .ZN(U3249) );
  NAND2_X1 U3740 ( .A1(n3239), .A2(n3238), .ZN(n3242) );
  NAND2_X1 U3741 ( .A1(n4250), .A2(n3240), .ZN(n3241) );
  AND2_X1 U3742 ( .A1(n4249), .A2(n3363), .ZN(n3244) );
  NAND2_X1 U3743 ( .A1(n4058), .A2(n3370), .ZN(n3243) );
  NAND2_X1 U3744 ( .A1(n3245), .A2(n4248), .ZN(n4087) );
  INV_X1 U3745 ( .A(n4087), .ZN(n4109) );
  NOR2_X1 U3746 ( .A1(n3245), .A2(n4248), .ZN(n4091) );
  OR2_X1 U3747 ( .A1(n4109), .A2(n4091), .ZN(n4144) );
  XNOR2_X1 U3748 ( .A(n3260), .B(n4144), .ZN(n3299) );
  AND2_X1 U3749 ( .A1(n3247), .A2(n3246), .ZN(n4084) );
  NAND2_X1 U3750 ( .A1(n3248), .A2(n4084), .ZN(n3249) );
  NAND2_X1 U3751 ( .A1(n3249), .A2(n4089), .ZN(n3364) );
  AND2_X1 U3752 ( .A1(n3370), .A2(n4249), .ZN(n4086) );
  OR2_X1 U3753 ( .A1(n3364), .A2(n4086), .ZN(n3250) );
  NAND2_X1 U3754 ( .A1(n4058), .A2(n3363), .ZN(n4107) );
  NAND2_X1 U3755 ( .A1(n3250), .A2(n4107), .ZN(n3262) );
  XNOR2_X1 U3756 ( .A(n3262), .B(n4144), .ZN(n3253) );
  OAI22_X1 U3757 ( .A1(n4058), .A2(n4548), .B1(n3976), .B2(n4546), .ZN(n3251)
         );
  AOI21_X1 U3758 ( .B1(n4057), .B2(n4560), .A(n3251), .ZN(n3252) );
  OAI21_X1 U3759 ( .B1(n3253), .B2(n4554), .A(n3252), .ZN(n3303) );
  AOI21_X1 U3760 ( .B1(n5340), .B2(n3299), .A(n3303), .ZN(n3259) );
  INV_X1 U3761 ( .A(n3254), .ZN(n3369) );
  NAND2_X1 U3762 ( .A1(n3369), .A2(n4057), .ZN(n3255) );
  NAND2_X1 U3763 ( .A1(n3267), .A2(n3255), .ZN(n3301) );
  INV_X1 U3764 ( .A(n3301), .ZN(n3257) );
  AOI22_X1 U3765 ( .A1(n3257), .A2(n3312), .B1(REG0_REG_6__SCAN_IN), .B2(n5345), .ZN(n3256) );
  OAI21_X1 U3766 ( .B1(n3259), .B2(n5345), .A(n3256), .ZN(U3479) );
  AOI22_X1 U3767 ( .A1(n3257), .A2(n3308), .B1(n5342), .B2(REG1_REG_6__SCAN_IN), .ZN(n3258) );
  OAI21_X1 U3768 ( .B1(n3259), .B2(n5342), .A(n3258), .ZN(U3524) );
  NAND2_X1 U3769 ( .A1(n3976), .A2(n3274), .ZN(n4093) );
  NAND2_X1 U3770 ( .A1(n3261), .A2(n4247), .ZN(n3381) );
  NAND2_X1 U3771 ( .A1(n4093), .A2(n3381), .ZN(n3276) );
  INV_X1 U3772 ( .A(n3276), .ZN(n4148) );
  XNOR2_X1 U3773 ( .A(n3277), .B(n4148), .ZN(n5248) );
  INV_X1 U3774 ( .A(n5248), .ZN(n3273) );
  XNOR2_X1 U3775 ( .A(n3278), .B(n4148), .ZN(n3266) );
  INV_X1 U3776 ( .A(n4246), .ZN(n4016) );
  OAI22_X1 U3777 ( .A1(n3263), .A2(n4548), .B1(n4016), .B2(n4546), .ZN(n3264)
         );
  AOI21_X1 U3778 ( .B1(n3274), .B2(n4560), .A(n3264), .ZN(n3265) );
  OAI21_X1 U3779 ( .B1(n3266), .B2(n4554), .A(n3265), .ZN(n5246) );
  NOR2_X4 U3780 ( .A1(n3267), .A2(n3274), .ZN(n3289) );
  AOI211_X1 U3781 ( .C1(n3274), .C2(n3267), .A(n5338), .B(n3289), .ZN(n5247)
         );
  INV_X1 U3782 ( .A(n5247), .ZN(n3270) );
  NAND2_X1 U3783 ( .A1(n4545), .A2(n5211), .ZN(n4512) );
  INV_X2 U3784 ( .A(n4545), .ZN(n5356) );
  INV_X1 U3785 ( .A(n5307), .ZN(n5302) );
  AOI22_X1 U3786 ( .A1(n5356), .A2(REG2_REG_7__SCAN_IN), .B1(n3268), .B2(n5302), .ZN(n3269) );
  OAI21_X1 U3787 ( .B1(n3270), .B2(n4512), .A(n3269), .ZN(n3271) );
  AOI21_X1 U3788 ( .B1(n5246), .B2(n4545), .A(n3271), .ZN(n3272) );
  OAI21_X1 U3789 ( .B1(n4518), .B2(n3273), .A(n3272), .ZN(U3283) );
  AND2_X1 U3790 ( .A1(n4247), .A2(n3274), .ZN(n3275) );
  MUX2_X1 U3791 ( .A(n4678), .B(DATAI_8_), .S(n2488), .Z(n3975) );
  NAND2_X1 U3792 ( .A1(n4016), .A2(n3379), .ZN(n3423) );
  NAND2_X1 U3793 ( .A1(n4246), .A2(n3975), .ZN(n3391) );
  NAND2_X1 U3794 ( .A1(n3423), .A2(n3391), .ZN(n4168) );
  XOR2_X1 U3795 ( .A(n3392), .B(n4168), .Z(n3307) );
  INV_X1 U3796 ( .A(n3307), .ZN(n3298) );
  NAND2_X1 U3797 ( .A1(n3278), .A2(n4093), .ZN(n3382) );
  NAND2_X1 U3798 ( .A1(n3382), .A2(n3381), .ZN(n3279) );
  XNOR2_X1 U3799 ( .A(n3279), .B(n4168), .ZN(n3288) );
  NAND2_X1 U3800 ( .A1(n2497), .A2(REG1_REG_9__SCAN_IN), .ZN(n3285) );
  AND2_X1 U3801 ( .A1(n3280), .A2(n4943), .ZN(n3281) );
  NOR2_X1 U3802 ( .A1(n3334), .A2(n3281), .ZN(n5251) );
  NAND2_X1 U3803 ( .A1(n3007), .A2(n5251), .ZN(n3284) );
  NAND2_X1 U3804 ( .A1(n3353), .A2(REG2_REG_9__SCAN_IN), .ZN(n3283) );
  NAND2_X1 U3805 ( .A1(n3046), .A2(REG0_REG_9__SCAN_IN), .ZN(n3282) );
  NAND4_X1 U3806 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n4245)
         );
  OAI22_X1 U3807 ( .A1(n3394), .A2(n4546), .B1(n3976), .B2(n4548), .ZN(n3286)
         );
  AOI21_X1 U3808 ( .B1(n3975), .B2(n4560), .A(n3286), .ZN(n3287) );
  OAI21_X1 U3809 ( .B1(n3288), .B2(n4554), .A(n3287), .ZN(n3306) );
  INV_X1 U3810 ( .A(n3289), .ZN(n3291) );
  NAND2_X1 U3811 ( .A1(n3289), .A2(n3379), .ZN(n3388) );
  INV_X1 U3812 ( .A(n3420), .ZN(n3290) );
  AOI21_X1 U3813 ( .B1(n3975), .B2(n3291), .A(n3290), .ZN(n3313) );
  INV_X1 U3814 ( .A(n3313), .ZN(n3295) );
  INV_X1 U3815 ( .A(n3292), .ZN(n3293) );
  AOI22_X1 U3816 ( .A1(n5356), .A2(REG2_REG_8__SCAN_IN), .B1(n3979), .B2(n5302), .ZN(n3294) );
  OAI21_X1 U3817 ( .B1(n3295), .B2(n5309), .A(n3294), .ZN(n3296) );
  AOI21_X1 U3818 ( .B1(n3306), .B2(n4545), .A(n3296), .ZN(n3297) );
  OAI21_X1 U3819 ( .B1(n3298), .B2(n4518), .A(n3297), .ZN(U3282) );
  INV_X1 U3820 ( .A(n3299), .ZN(n3305) );
  AOI22_X1 U3821 ( .A1(n5356), .A2(REG2_REG_6__SCAN_IN), .B1(n4061), .B2(n5302), .ZN(n3300) );
  OAI21_X1 U3822 ( .B1(n3301), .B2(n5309), .A(n3300), .ZN(n3302) );
  AOI21_X1 U3823 ( .B1(n3303), .B2(n4545), .A(n3302), .ZN(n3304) );
  OAI21_X1 U3824 ( .B1(n3305), .B2(n4518), .A(n3304), .ZN(U3284) );
  AOI21_X1 U3825 ( .B1(n3307), .B2(n5340), .A(n3306), .ZN(n3315) );
  AOI22_X1 U3826 ( .A1(n3313), .A2(n3308), .B1(n5342), .B2(REG1_REG_8__SCAN_IN), .ZN(n3309) );
  OAI21_X1 U3827 ( .B1(n3315), .B2(n5342), .A(n3309), .ZN(U3526) );
  INV_X1 U3828 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3310) );
  NOR2_X1 U3829 ( .A1(n5348), .A2(n3310), .ZN(n3311) );
  AOI21_X1 U3830 ( .B1(n3313), .B2(n3312), .A(n3311), .ZN(n3314) );
  OAI21_X1 U3831 ( .B1(n3315), .B2(n5345), .A(n3314), .ZN(U3483) );
  INV_X1 U3832 ( .A(n3316), .ZN(n3318) );
  NAND2_X1 U3833 ( .A1(n3318), .A2(n3317), .ZN(n3319) );
  AND2_X2 U3834 ( .A1(n3320), .A2(n3319), .ZN(n3973) );
  NAND2_X1 U3835 ( .A1(n3826), .A2(n3975), .ZN(n3322) );
  NAND2_X1 U3836 ( .A1(n2499), .A2(n4246), .ZN(n3321) );
  NAND2_X1 U3837 ( .A1(n3322), .A2(n3321), .ZN(n3323) );
  XNOR2_X1 U3838 ( .A(n3323), .B(n3810), .ZN(n3325) );
  NOR2_X1 U3839 ( .A1(n3875), .A2(n3379), .ZN(n3324) );
  AOI21_X1 U3840 ( .B1(n3831), .B2(n4246), .A(n3324), .ZN(n3326) );
  NAND2_X1 U3841 ( .A1(n3325), .A2(n3326), .ZN(n3330) );
  INV_X1 U3842 ( .A(n3325), .ZN(n3328) );
  INV_X1 U3843 ( .A(n3326), .ZN(n3327) );
  NAND2_X1 U3844 ( .A1(n3328), .A2(n3327), .ZN(n3329) );
  AND2_X1 U3845 ( .A1(n3330), .A2(n3329), .ZN(n3972) );
  NAND2_X1 U3846 ( .A1(n3973), .A2(n3972), .ZN(n3971) );
  NAND2_X1 U3847 ( .A1(n3971), .A2(n3330), .ZN(n4012) );
  MUX2_X1 U3848 ( .A(n4677), .B(DATAI_9_), .S(n2488), .Z(n4015) );
  NAND2_X1 U3849 ( .A1(n3826), .A2(n4015), .ZN(n3332) );
  NAND2_X1 U3850 ( .A1(n2499), .A2(n4245), .ZN(n3331) );
  NAND2_X1 U3851 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  XNOR2_X1 U3852 ( .A(n3333), .B(n3810), .ZN(n3346) );
  INV_X1 U3853 ( .A(n4015), .ZN(n3393) );
  OAI22_X1 U3854 ( .A1(n2493), .A2(n3394), .B1(n3128), .B2(n3393), .ZN(n3344)
         );
  XNOR2_X1 U3855 ( .A(n3346), .B(n3344), .ZN(n4013) );
  NAND2_X1 U3856 ( .A1(n4012), .A2(n4013), .ZN(n3348) );
  MUX2_X1 U3857 ( .A(n2724), .B(DATAI_10_), .S(n2488), .Z(n4111) );
  NAND2_X1 U3858 ( .A1(n3826), .A2(n4111), .ZN(n3342) );
  NAND2_X1 U3859 ( .A1(n2496), .A2(REG1_REG_10__SCAN_IN), .ZN(n3340) );
  NOR2_X1 U3860 ( .A1(n3334), .A2(REG3_REG_10__SCAN_IN), .ZN(n3335) );
  OR2_X1 U3861 ( .A1(n3351), .A2(n3335), .ZN(n3389) );
  INV_X1 U3862 ( .A(n3389), .ZN(n3336) );
  NAND2_X1 U3863 ( .A1(n3007), .A2(n3336), .ZN(n3339) );
  NAND2_X1 U3864 ( .A1(n3353), .A2(REG2_REG_10__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U3865 ( .A1(n3046), .A2(REG0_REG_10__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U3866 ( .A1(n2499), .A2(n4244), .ZN(n3341) );
  NAND2_X1 U3867 ( .A1(n3342), .A2(n3341), .ZN(n3343) );
  XNOR2_X1 U3868 ( .A(n3343), .B(n3810), .ZN(n3440) );
  INV_X1 U3869 ( .A(n4244), .ZN(n4110) );
  INV_X1 U3870 ( .A(n4111), .ZN(n3510) );
  OAI22_X1 U3871 ( .A1(n2493), .A2(n4110), .B1(n3128), .B2(n3510), .ZN(n3441)
         );
  XNOR2_X1 U3872 ( .A(n3440), .B(n3441), .ZN(n3349) );
  INV_X1 U3873 ( .A(n3344), .ZN(n3345) );
  NAND2_X1 U3874 ( .A1(n3346), .A2(n3345), .ZN(n3350) );
  AND2_X1 U3875 ( .A1(n3349), .A2(n3350), .ZN(n3347) );
  NAND2_X1 U3876 ( .A1(n3444), .A2(n4055), .ZN(n3362) );
  AOI21_X1 U3877 ( .B1(n3348), .B2(n3350), .A(n3349), .ZN(n3361) );
  NAND2_X1 U3878 ( .A1(n2496), .A2(REG1_REG_11__SCAN_IN), .ZN(n3357) );
  OR2_X1 U3879 ( .A1(n3351), .A2(REG3_REG_11__SCAN_IN), .ZN(n3352) );
  AND2_X1 U3880 ( .A1(n3449), .A2(n3352), .ZN(n3525) );
  NAND2_X1 U3881 ( .A1(n3007), .A2(n3525), .ZN(n3356) );
  NAND2_X1 U3882 ( .A1(n3353), .A2(REG2_REG_11__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U3883 ( .A1(n3046), .A2(REG0_REG_11__SCAN_IN), .ZN(n3354) );
  NAND4_X1 U3884 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n4243)
         );
  AOI22_X1 U3885 ( .A1(n5296), .A2(n4243), .B1(n5282), .B2(n4111), .ZN(n3360)
         );
  AND2_X1 U3886 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3411) );
  NOR2_X1 U3887 ( .A1(n5300), .A2(n3389), .ZN(n3358) );
  AOI211_X1 U3888 ( .C1(n5284), .C2(n4245), .A(n3411), .B(n3358), .ZN(n3359)
         );
  OAI211_X1 U3889 ( .C1(n3362), .C2(n3361), .A(n3360), .B(n3359), .ZN(U3214)
         );
  XNOR2_X1 U3890 ( .A(n4249), .B(n3363), .ZN(n4177) );
  XOR2_X1 U3891 ( .A(n4177), .B(n3364), .Z(n3367) );
  AOI22_X1 U3892 ( .A1(n4504), .A2(n4250), .B1(n4248), .B2(n4525), .ZN(n3365)
         );
  OAI21_X1 U3893 ( .B1(n3370), .B2(n4581), .A(n3365), .ZN(n3366) );
  AOI21_X1 U3894 ( .B1(n3367), .B2(n4501), .A(n3366), .ZN(n5239) );
  INV_X1 U3895 ( .A(n3368), .ZN(n3371) );
  OAI21_X1 U3896 ( .B1(n3371), .B2(n3370), .A(n3369), .ZN(n5240) );
  INV_X1 U3897 ( .A(n5240), .ZN(n3375) );
  INV_X1 U3898 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3373) );
  OAI22_X1 U3899 ( .A1(n4545), .A2(n3373), .B1(n3372), .B2(n5307), .ZN(n3374)
         );
  AOI21_X1 U3900 ( .B1(n3375), .B2(n5352), .A(n3374), .ZN(n3378) );
  XNOR2_X1 U3901 ( .A(n3376), .B(n4177), .ZN(n5242) );
  INV_X1 U3902 ( .A(n4518), .ZN(n4568) );
  NAND2_X1 U3903 ( .A1(n5242), .A2(n4568), .ZN(n3377) );
  OAI211_X1 U3904 ( .C1(n5239), .C2(n5356), .A(n3378), .B(n3377), .ZN(U3285)
         );
  NAND2_X1 U3905 ( .A1(n3379), .A2(n4246), .ZN(n3380) );
  AND2_X1 U3906 ( .A1(n3381), .A2(n3380), .ZN(n4112) );
  NAND2_X1 U3907 ( .A1(n3382), .A2(n4112), .ZN(n3424) );
  NAND2_X1 U3908 ( .A1(n4016), .A2(n3975), .ZN(n4096) );
  NAND2_X1 U3909 ( .A1(n3424), .A2(n4096), .ZN(n3383) );
  NAND2_X1 U3910 ( .A1(n3394), .A2(n4015), .ZN(n4095) );
  NAND2_X1 U3911 ( .A1(n3393), .A2(n4245), .ZN(n4106) );
  NAND2_X1 U3912 ( .A1(n4095), .A2(n4106), .ZN(n3398) );
  INV_X1 U3913 ( .A(n3398), .ZN(n4146) );
  NAND2_X1 U3914 ( .A1(n3509), .A2(n4095), .ZN(n3384) );
  XNOR2_X1 U3915 ( .A(n4244), .B(n4111), .ZN(n4174) );
  XNOR2_X1 U3916 ( .A(n3384), .B(n4174), .ZN(n3385) );
  NAND2_X1 U3917 ( .A1(n3385), .A2(n4501), .ZN(n3387) );
  AOI22_X1 U3918 ( .A1(n4504), .A2(n4245), .B1(n4243), .B2(n4525), .ZN(n3386)
         );
  OAI211_X1 U3919 ( .C1(n4581), .C2(n3510), .A(n3387), .B(n3386), .ZN(n5260)
         );
  INV_X1 U3920 ( .A(n5260), .ZN(n3407) );
  OR2_X2 U3921 ( .A1(n3388), .A2(n4015), .ZN(n3422) );
  AOI21_X1 U3922 ( .B1(n4111), .B2(n3422), .A(n3532), .ZN(n5261) );
  OAI22_X1 U3923 ( .A1(n4545), .A2(n3410), .B1(n3389), .B2(n5307), .ZN(n3390)
         );
  AOI21_X1 U3924 ( .B1(n5261), .B2(n5352), .A(n3390), .ZN(n3406) );
  NAND2_X1 U3925 ( .A1(n3392), .A2(n3391), .ZN(n3400) );
  NAND2_X1 U3926 ( .A1(n3394), .A2(n3393), .ZN(n3397) );
  AND2_X1 U3927 ( .A1(n3423), .A2(n3397), .ZN(n3401) );
  INV_X1 U3928 ( .A(n4174), .ZN(n3395) );
  AND2_X1 U3929 ( .A1(n3401), .A2(n3395), .ZN(n3396) );
  NAND2_X1 U3930 ( .A1(n3400), .A2(n3396), .ZN(n3504) );
  INV_X1 U3931 ( .A(n3397), .ZN(n3399) );
  OR2_X1 U3932 ( .A1(n3399), .A2(n3398), .ZN(n3402) );
  OR2_X1 U3933 ( .A1(n4174), .A2(n3402), .ZN(n3501) );
  AND2_X1 U3934 ( .A1(n3504), .A2(n3501), .ZN(n5258) );
  NAND2_X1 U3935 ( .A1(n3400), .A2(n3401), .ZN(n3403) );
  AND2_X1 U3936 ( .A1(n3403), .A2(n3402), .ZN(n3404) );
  NAND2_X1 U3937 ( .A1(n3404), .A2(n4174), .ZN(n5257) );
  NAND3_X1 U3938 ( .A1(n5258), .A2(n5257), .A3(n4568), .ZN(n3405) );
  OAI211_X1 U3939 ( .C1(n3407), .C2(n5356), .A(n3406), .B(n3405), .ZN(U3280)
         );
  AOI21_X1 U3940 ( .B1(n3410), .B2(n3409), .A(n3408), .ZN(n3418) );
  AOI21_X1 U3941 ( .B1(n5196), .B2(ADDR_REG_10__SCAN_IN), .A(n3411), .ZN(n3412) );
  OAI21_X1 U3942 ( .B1(n5181), .B2(n3413), .A(n3412), .ZN(n3417) );
  AOI211_X1 U3943 ( .C1(n3415), .C2(n5262), .A(n3414), .B(n5197), .ZN(n3416)
         );
  AOI211_X1 U3944 ( .C1(n3418), .C2(n2795), .A(n3417), .B(n3416), .ZN(n3419)
         );
  INV_X1 U3945 ( .A(n3419), .ZN(U3250) );
  NAND2_X1 U3946 ( .A1(n3420), .A2(n4015), .ZN(n3421) );
  NAND2_X1 U3947 ( .A1(n3422), .A2(n3421), .ZN(n5253) );
  NAND2_X1 U3948 ( .A1(n3400), .A2(n3423), .ZN(n3427) );
  INV_X1 U3949 ( .A(n3427), .ZN(n3426) );
  NAND3_X1 U3950 ( .A1(n3424), .A2(n4501), .A3(n4096), .ZN(n3425) );
  OAI21_X1 U3951 ( .B1(n3426), .B2(n5272), .A(n3425), .ZN(n3429) );
  NOR2_X1 U3952 ( .A1(n3427), .A2(n5272), .ZN(n3428) );
  MUX2_X1 U3953 ( .A(n3429), .B(n3428), .S(n4146), .Z(n3433) );
  AOI22_X1 U3954 ( .A1(n4504), .A2(n4246), .B1(n4244), .B2(n4525), .ZN(n3431)
         );
  NAND2_X1 U3955 ( .A1(n4015), .A2(n4560), .ZN(n3430) );
  OAI211_X1 U3956 ( .C1(n3509), .C2(n4554), .A(n3431), .B(n3430), .ZN(n3432)
         );
  NOR2_X1 U3957 ( .A1(n3433), .A2(n3432), .ZN(n5256) );
  MUX2_X1 U3958 ( .A(n2813), .B(n5256), .S(n5344), .Z(n3434) );
  OAI21_X1 U3959 ( .B1(n5253), .B2(n4628), .A(n3434), .ZN(U3527) );
  INV_X1 U3960 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3435) );
  MUX2_X1 U3961 ( .A(n3435), .B(n5256), .S(n5348), .Z(n3436) );
  OAI21_X1 U3962 ( .B1(n5253), .B2(n4666), .A(n3436), .ZN(U3485) );
  MUX2_X1 U3963 ( .A(n4676), .B(DATAI_11_), .S(n2488), .Z(n3500) );
  NAND2_X1 U3964 ( .A1(n3826), .A2(n3500), .ZN(n3438) );
  NAND2_X1 U3965 ( .A1(n2499), .A2(n4243), .ZN(n3437) );
  NAND2_X1 U3966 ( .A1(n3438), .A2(n3437), .ZN(n3439) );
  XNOR2_X1 U3967 ( .A(n3439), .B(n3873), .ZN(n3460) );
  OAI22_X1 U3968 ( .A1(n2493), .A2(n3513), .B1(n3128), .B2(n3531), .ZN(n3461)
         );
  XNOR2_X1 U3969 ( .A(n3460), .B(n3461), .ZN(n3448) );
  INV_X1 U3970 ( .A(n3440), .ZN(n3442) );
  NAND2_X1 U3971 ( .A1(n3442), .A2(n3441), .ZN(n3443) );
  INV_X1 U3972 ( .A(n3580), .ZN(n3447) );
  AOI21_X1 U3973 ( .B1(n3448), .B2(n3445), .A(n3447), .ZN(n3459) );
  NAND2_X1 U3974 ( .A1(n2496), .A2(REG1_REG_12__SCAN_IN), .ZN(n3454) );
  NAND2_X1 U3975 ( .A1(n3449), .A2(n3481), .ZN(n3450) );
  AND2_X1 U3976 ( .A1(n3474), .A2(n3450), .ZN(n3473) );
  NAND2_X1 U3977 ( .A1(n3007), .A2(n3473), .ZN(n3453) );
  NAND2_X1 U3978 ( .A1(n3353), .A2(REG2_REG_12__SCAN_IN), .ZN(n3452) );
  NAND2_X1 U3979 ( .A1(n3046), .A2(REG0_REG_12__SCAN_IN), .ZN(n3451) );
  NAND4_X1 U3980 ( .A1(n3454), .A2(n3453), .A3(n3452), .A4(n3451), .ZN(n5283)
         );
  AOI22_X1 U3981 ( .A1(n5296), .A2(n5283), .B1(n5282), .B2(n3500), .ZN(n3458)
         );
  INV_X1 U3982 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3455) );
  NOR2_X1 U3983 ( .A1(STATE_REG_SCAN_IN), .A2(n3455), .ZN(n3490) );
  NOR2_X1 U3984 ( .A1(n4071), .A2(n4110), .ZN(n3456) );
  AOI211_X1 U3985 ( .C1(n4068), .C2(n3525), .A(n3490), .B(n3456), .ZN(n3457)
         );
  OAI211_X1 U3986 ( .C1(n3459), .C2(n5291), .A(n3458), .B(n3457), .ZN(U3233)
         );
  INV_X1 U3987 ( .A(n3460), .ZN(n3463) );
  INV_X1 U3988 ( .A(n3461), .ZN(n3462) );
  NAND2_X1 U3989 ( .A1(n3463), .A2(n3462), .ZN(n3578) );
  NAND2_X1 U3990 ( .A1(n3580), .A2(n3578), .ZN(n5286) );
  INV_X1 U3991 ( .A(n3671), .ZN(n3464) );
  MUX2_X1 U3992 ( .A(n3464), .B(DATAI_12_), .S(n2488), .Z(n3515) );
  NAND2_X1 U3993 ( .A1(n3826), .A2(n3515), .ZN(n3466) );
  NAND2_X1 U3994 ( .A1(n2499), .A2(n5283), .ZN(n3465) );
  NAND2_X1 U3995 ( .A1(n3466), .A2(n3465), .ZN(n3467) );
  XNOR2_X1 U3996 ( .A(n3467), .B(n3873), .ZN(n3471) );
  INV_X1 U3997 ( .A(n3471), .ZN(n3469) );
  INV_X1 U3998 ( .A(n5283), .ZN(n3616) );
  INV_X1 U3999 ( .A(n3515), .ZN(n3610) );
  OAI22_X1 U4000 ( .A1(n2493), .A2(n3616), .B1(n3875), .B2(n3610), .ZN(n3470)
         );
  INV_X1 U4001 ( .A(n3470), .ZN(n3468) );
  NAND2_X1 U4002 ( .A1(n3469), .A2(n3468), .ZN(n5287) );
  NAND2_X1 U4003 ( .A1(n3471), .A2(n3470), .ZN(n5285) );
  NAND2_X1 U4004 ( .A1(n5287), .A2(n5285), .ZN(n3472) );
  XNOR2_X1 U4005 ( .A(n5286), .B(n3472), .ZN(n3486) );
  INV_X1 U4006 ( .A(n3473), .ZN(n3507) );
  NAND2_X1 U4007 ( .A1(n2497), .A2(REG1_REG_13__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4008 ( .A1(n3474), .A2(n4268), .ZN(n3476) );
  INV_X1 U4009 ( .A(n3549), .ZN(n3475) );
  NAND2_X1 U4010 ( .A1(n3476), .A2(n3475), .ZN(n5299) );
  INV_X1 U4011 ( .A(n5299), .ZN(n5303) );
  NAND2_X1 U4012 ( .A1(n3007), .A2(n5303), .ZN(n3479) );
  NAND2_X1 U4013 ( .A1(n3353), .A2(REG2_REG_13__SCAN_IN), .ZN(n3478) );
  NAND2_X1 U4014 ( .A1(n3046), .A2(REG0_REG_13__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4015 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n4242)
         );
  AOI22_X1 U4016 ( .A1(n5296), .A2(n4242), .B1(n5282), .B2(n3515), .ZN(n3483)
         );
  NOR2_X1 U4017 ( .A1(STATE_REG_SCAN_IN), .A2(n3481), .ZN(n3669) );
  AOI21_X1 U4018 ( .B1(n5284), .B2(n4243), .A(n3669), .ZN(n3482) );
  OAI211_X1 U4019 ( .C1(n3507), .C2(n5300), .A(n3483), .B(n3482), .ZN(n3484)
         );
  INV_X1 U4020 ( .A(n3484), .ZN(n3485) );
  OAI21_X1 U4021 ( .B1(n3486), .B2(n5291), .A(n3485), .ZN(U3221) );
  AOI21_X1 U4022 ( .B1(n3489), .B2(n3488), .A(n3487), .ZN(n3498) );
  AOI21_X1 U4023 ( .B1(n5196), .B2(ADDR_REG_11__SCAN_IN), .A(n3490), .ZN(n3491) );
  OAI21_X1 U4024 ( .B1(n5181), .B2(n3492), .A(n3491), .ZN(n3497) );
  AOI211_X1 U4025 ( .C1(n3495), .C2(n3494), .A(n3493), .B(n5200), .ZN(n3496)
         );
  AOI211_X1 U4026 ( .C1(n5177), .C2(n3498), .A(n3497), .B(n3496), .ZN(n3499)
         );
  INV_X1 U4027 ( .A(n3499), .ZN(U3251) );
  NAND2_X1 U4028 ( .A1(n3513), .A2(n3500), .ZN(n4114) );
  NAND2_X1 U4029 ( .A1(n3531), .A2(n4243), .ZN(n4103) );
  INV_X1 U4030 ( .A(n4159), .ZN(n3528) );
  NAND2_X1 U4031 ( .A1(n4244), .A2(n4111), .ZN(n3502) );
  AND2_X1 U4032 ( .A1(n3502), .A2(n3501), .ZN(n3526) );
  NAND2_X1 U4033 ( .A1(n3504), .A2(n3503), .ZN(n3527) );
  NAND2_X1 U4034 ( .A1(n3513), .A2(n3531), .ZN(n3505) );
  NAND2_X1 U4035 ( .A1(n3527), .A2(n3505), .ZN(n3609) );
  NAND2_X1 U4036 ( .A1(n3616), .A2(n3515), .ZN(n4115) );
  NAND2_X1 U4037 ( .A1(n3610), .A2(n5283), .ZN(n3654) );
  NAND2_X1 U4038 ( .A1(n4115), .A2(n3654), .ZN(n3608) );
  INV_X1 U4039 ( .A(n3608), .ZN(n4149) );
  XNOR2_X1 U4040 ( .A(n3609), .B(n4149), .ZN(n5273) );
  NAND2_X1 U4041 ( .A1(n3532), .A2(n3531), .ZN(n3506) );
  OR2_X2 U4042 ( .A1(n3506), .A2(n3515), .ZN(n3605) );
  INV_X1 U40430 ( .A(n3605), .ZN(n3607) );
  AOI21_X1 U4044 ( .B1(n3515), .B2(n3530), .A(n3607), .ZN(n5276) );
  OAI22_X1 U4045 ( .A1(n4545), .A2(n3674), .B1(n3507), .B2(n5307), .ZN(n3508)
         );
  AOI21_X1 U4046 ( .B1(n5276), .B2(n5352), .A(n3508), .ZN(n3519) );
  NAND3_X1 U4047 ( .A1(n3509), .A2(n4174), .A3(n4095), .ZN(n3511) );
  NAND2_X1 U4048 ( .A1(n3510), .A2(n4244), .ZN(n4102) );
  NAND2_X1 U4049 ( .A1(n3511), .A2(n4102), .ZN(n3520) );
  NAND2_X1 U4050 ( .A1(n3520), .A2(n4159), .ZN(n3512) );
  NAND2_X1 U4051 ( .A1(n3512), .A2(n4103), .ZN(n3614) );
  XNOR2_X1 U4052 ( .A(n3614), .B(n4149), .ZN(n3517) );
  INV_X1 U4053 ( .A(n4242), .ZN(n3612) );
  OAI22_X1 U4054 ( .A1(n3612), .A2(n4546), .B1(n3513), .B2(n4548), .ZN(n3514)
         );
  AOI21_X1 U4055 ( .B1(n3515), .B2(n4560), .A(n3514), .ZN(n3516) );
  OAI21_X1 U4056 ( .B1(n3517), .B2(n4554), .A(n3516), .ZN(n5275) );
  NAND2_X1 U4057 ( .A1(n5275), .A2(n4545), .ZN(n3518) );
  OAI211_X1 U4058 ( .C1(n5273), .C2(n4518), .A(n3519), .B(n3518), .ZN(U3278)
         );
  XOR2_X1 U4059 ( .A(n4159), .B(n3520), .Z(n3523) );
  AOI22_X1 U4060 ( .A1(n4504), .A2(n4244), .B1(n5283), .B2(n4525), .ZN(n3521)
         );
  OAI21_X1 U4061 ( .B1(n3531), .B2(n4581), .A(n3521), .ZN(n3522) );
  AOI21_X1 U4062 ( .B1(n3523), .B2(n4501), .A(n3522), .ZN(n5265) );
  INV_X1 U4063 ( .A(n5265), .ZN(n3524) );
  AOI21_X1 U4064 ( .B1(n3525), .B2(n5302), .A(n3524), .ZN(n3536) );
  AND2_X1 U4065 ( .A1(n3504), .A2(n3526), .ZN(n3529) );
  OAI21_X1 U4066 ( .B1(n3529), .B2(n3528), .A(n3527), .ZN(n5268) );
  OAI21_X1 U4067 ( .B1(n3532), .B2(n3531), .A(n3530), .ZN(n5266) );
  INV_X1 U4068 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3533) );
  OAI22_X1 U4069 ( .A1(n5266), .A2(n5309), .B1(n3533), .B2(n4545), .ZN(n3534)
         );
  AOI21_X1 U4070 ( .B1(n5268), .B2(n4568), .A(n3534), .ZN(n3535) );
  OAI21_X1 U4071 ( .B1(n3536), .B2(n5356), .A(n3535), .ZN(U3279) );
  MUX2_X1 U4072 ( .A(n4675), .B(DATAI_13_), .S(n2488), .Z(n5281) );
  NAND2_X1 U4073 ( .A1(n3826), .A2(n5281), .ZN(n3538) );
  NAND2_X1 U4074 ( .A1(n2498), .A2(n4242), .ZN(n3537) );
  NAND2_X1 U4075 ( .A1(n3538), .A2(n3537), .ZN(n3539) );
  XNOR2_X1 U4076 ( .A(n3539), .B(n3810), .ZN(n3542) );
  INV_X1 U4077 ( .A(n5281), .ZN(n3613) );
  OAI22_X1 U4078 ( .A1(n2493), .A2(n3612), .B1(n3875), .B2(n3613), .ZN(n3541)
         );
  INV_X1 U4079 ( .A(n3541), .ZN(n3540) );
  NAND2_X1 U4080 ( .A1(n3542), .A2(n3540), .ZN(n3545) );
  INV_X1 U4081 ( .A(n3545), .ZN(n3543) );
  XNOR2_X1 U4082 ( .A(n3542), .B(n3541), .ZN(n5290) );
  AND2_X1 U4083 ( .A1(n5285), .A2(n3544), .ZN(n3583) );
  NAND2_X1 U4084 ( .A1(n5286), .A2(n3583), .ZN(n3548) );
  INV_X1 U4085 ( .A(n3544), .ZN(n3547) );
  AND2_X1 U4086 ( .A1(n5287), .A2(n3545), .ZN(n3546) );
  NAND2_X1 U4087 ( .A1(n3548), .A2(n3575), .ZN(n3560) );
  MUX2_X1 U4088 ( .A(n2823), .B(DATAI_14_), .S(n2488), .Z(n3679) );
  NAND2_X1 U4089 ( .A1(n3826), .A2(n3679), .ZN(n3556) );
  NAND2_X1 U4090 ( .A1(n2496), .A2(REG1_REG_14__SCAN_IN), .ZN(n3554) );
  OAI21_X1 U4091 ( .B1(REG3_REG_14__SCAN_IN), .B2(n3549), .A(n3561), .ZN(n5308) );
  INV_X1 U4092 ( .A(n5308), .ZN(n3550) );
  NAND2_X1 U4093 ( .A1(n3007), .A2(n3550), .ZN(n3553) );
  NAND2_X1 U4094 ( .A1(n3353), .A2(REG2_REG_14__SCAN_IN), .ZN(n3552) );
  NAND2_X1 U4095 ( .A1(n3046), .A2(REG0_REG_14__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4096 ( .A1(n2499), .A2(n5295), .ZN(n3555) );
  NAND2_X1 U4097 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  XNOR2_X1 U4098 ( .A(n3557), .B(n3810), .ZN(n3574) );
  NOR2_X1 U4099 ( .A1(n3875), .A2(n3657), .ZN(n3558) );
  AOI21_X1 U4100 ( .B1(n3831), .B2(n5295), .A(n3558), .ZN(n3573) );
  XNOR2_X1 U4101 ( .A(n3574), .B(n3573), .ZN(n3559) );
  XNOR2_X1 U4102 ( .A(n3560), .B(n3559), .ZN(n3570) );
  NAND2_X1 U4103 ( .A1(n2497), .A2(REG1_REG_15__SCAN_IN), .ZN(n3565) );
  AOI21_X1 U4104 ( .B1(n3561), .B2(n3600), .A(n3594), .ZN(n4542) );
  NAND2_X1 U4105 ( .A1(n3007), .A2(n4542), .ZN(n3564) );
  NAND2_X1 U4106 ( .A1(n3353), .A2(REG2_REG_15__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U4107 ( .A1(n3046), .A2(REG0_REG_15__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4108 ( .A1(n5296), .A2(n4241), .B1(n5282), .B2(n3679), .ZN(n3569)
         );
  INV_X1 U4109 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3566) );
  NOR2_X1 U4110 ( .A1(STATE_REG_SCAN_IN), .A2(n3566), .ZN(n4282) );
  NOR2_X1 U4111 ( .A1(n5300), .A2(n5308), .ZN(n3567) );
  AOI211_X1 U4112 ( .C1(n5284), .C2(n4242), .A(n4282), .B(n3567), .ZN(n3568)
         );
  OAI211_X1 U4113 ( .C1(n3570), .C2(n5291), .A(n3569), .B(n3568), .ZN(U3212)
         );
  MUX2_X1 U4114 ( .A(n5150), .B(DATAI_15_), .S(n2488), .Z(n4559) );
  OAI22_X1 U4115 ( .A1(n2493), .A2(n3682), .B1(n3128), .B2(n4561), .ZN(n3627)
         );
  INV_X1 U4116 ( .A(n3574), .ZN(n3572) );
  INV_X1 U4117 ( .A(n3573), .ZN(n3571) );
  NAND2_X1 U4118 ( .A1(n3572), .A2(n3571), .ZN(n3582) );
  INV_X1 U4119 ( .A(n3582), .ZN(n3577) );
  AND2_X1 U4120 ( .A1(n3578), .A2(n3581), .ZN(n3579) );
  NAND2_X1 U4121 ( .A1(n3580), .A2(n3579), .ZN(n3587) );
  INV_X1 U4122 ( .A(n3581), .ZN(n3585) );
  AND2_X1 U4123 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  NAND2_X1 U4124 ( .A1(n3587), .A2(n3586), .ZN(n3592) );
  NAND2_X1 U4125 ( .A1(n3826), .A2(n4559), .ZN(n3589) );
  NAND2_X1 U4126 ( .A1(n2499), .A2(n4241), .ZN(n3588) );
  NAND2_X1 U4127 ( .A1(n3589), .A2(n3588), .ZN(n3590) );
  XNOR2_X1 U4128 ( .A(n3590), .B(n3873), .ZN(n3591) );
  OR2_X2 U4129 ( .A1(n3592), .A2(n3591), .ZN(n3628) );
  NAND2_X1 U4130 ( .A1(n3592), .A2(n3591), .ZN(n3625) );
  NAND2_X1 U4131 ( .A1(n3628), .A2(n3625), .ZN(n3593) );
  XOR2_X1 U4132 ( .A(n3627), .B(n3593), .Z(n3604) );
  NAND2_X1 U4133 ( .A1(n2497), .A2(REG1_REG_16__SCAN_IN), .ZN(n3599) );
  OAI21_X1 U4134 ( .B1(n3594), .B2(REG3_REG_16__SCAN_IN), .A(n3638), .ZN(n3692) );
  INV_X1 U4135 ( .A(n3692), .ZN(n3595) );
  NAND2_X1 U4136 ( .A1(n3007), .A2(n3595), .ZN(n3598) );
  NAND2_X1 U4137 ( .A1(n3353), .A2(REG2_REG_16__SCAN_IN), .ZN(n3597) );
  NAND2_X1 U4138 ( .A1(n3046), .A2(REG0_REG_16__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4139 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n4240)
         );
  AOI22_X1 U4140 ( .A1(n5296), .A2(n4240), .B1(n5282), .B2(n4559), .ZN(n3603)
         );
  NOR2_X1 U4141 ( .A1(STATE_REG_SCAN_IN), .A2(n3600), .ZN(n5144) );
  NOR2_X1 U4142 ( .A1(n4071), .A2(n4549), .ZN(n3601) );
  AOI211_X1 U4143 ( .C1(n4068), .C2(n4542), .A(n5144), .B(n3601), .ZN(n3602)
         );
  OAI211_X1 U4144 ( .C1(n3604), .C2(n5291), .A(n3603), .B(n3602), .ZN(U3238)
         );
  INV_X1 U4145 ( .A(n3649), .ZN(n3606) );
  OAI21_X1 U4146 ( .B1(n3607), .B2(n3613), .A(n3606), .ZN(n5301) );
  INV_X1 U4147 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3622) );
  NAND2_X1 U4148 ( .A1(n3616), .A2(n3610), .ZN(n3611) );
  NAND2_X1 U4149 ( .A1(n3612), .A2(n5281), .ZN(n4118) );
  NAND2_X1 U4150 ( .A1(n3613), .A2(n4242), .ZN(n3653) );
  NAND2_X1 U4151 ( .A1(n4118), .A2(n3653), .ZN(n3651) );
  XNOR2_X1 U4152 ( .A(n3652), .B(n3651), .ZN(n3621) );
  NAND2_X1 U4153 ( .A1(n3614), .A2(n4115), .ZN(n3655) );
  NAND2_X1 U4154 ( .A1(n3655), .A2(n3654), .ZN(n3615) );
  INV_X1 U4155 ( .A(n3651), .ZN(n4150) );
  XNOR2_X1 U4156 ( .A(n3615), .B(n4150), .ZN(n3619) );
  OAI22_X1 U4157 ( .A1(n3616), .A2(n4548), .B1(n4549), .B2(n4546), .ZN(n3617)
         );
  AOI21_X1 U4158 ( .B1(n5281), .B2(n4560), .A(n3617), .ZN(n3618) );
  OAI21_X1 U4159 ( .B1(n3619), .B2(n4554), .A(n3618), .ZN(n3620) );
  AOI21_X1 U4160 ( .B1(n3621), .B2(n5340), .A(n3620), .ZN(n5306) );
  MUX2_X1 U4161 ( .A(n3622), .B(n5306), .S(n5348), .Z(n3623) );
  OAI21_X1 U4162 ( .B1(n5301), .B2(n4666), .A(n3623), .ZN(U3493) );
  MUX2_X1 U4163 ( .A(n2819), .B(n5306), .S(n5344), .Z(n3624) );
  OAI21_X1 U4164 ( .B1(n5301), .B2(n4628), .A(n3624), .ZN(U3531) );
  INV_X1 U4165 ( .A(n3625), .ZN(n3626) );
  MUX2_X1 U4166 ( .A(n3629), .B(DATAI_16_), .S(n2488), .Z(n3893) );
  NAND2_X1 U4167 ( .A1(n3826), .A2(n3893), .ZN(n3631) );
  NAND2_X1 U4168 ( .A1(n2499), .A2(n4240), .ZN(n3630) );
  NAND2_X1 U4169 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  XNOR2_X1 U4170 ( .A(n3632), .B(n3873), .ZN(n3636) );
  INV_X1 U4171 ( .A(n3636), .ZN(n3634) );
  INV_X1 U4172 ( .A(n4240), .ZN(n4547) );
  OAI22_X1 U4173 ( .A1(n2493), .A2(n4547), .B1(n2491), .B2(n3690), .ZN(n3635)
         );
  INV_X1 U4174 ( .A(n3635), .ZN(n3633) );
  NAND2_X1 U4175 ( .A1(n3634), .A2(n3633), .ZN(n3708) );
  NAND2_X1 U4176 ( .A1(n3636), .A2(n3635), .ZN(n3706) );
  NAND2_X1 U4177 ( .A1(n3708), .A2(n3706), .ZN(n3637) );
  XNOR2_X1 U4178 ( .A(n3707), .B(n3637), .ZN(n3647) );
  AOI22_X1 U4179 ( .A1(n5284), .A2(n4241), .B1(n5282), .B2(n3893), .ZN(n3644)
         );
  AOI21_X1 U4180 ( .B1(n3638), .B2(n3719), .A(n3714), .ZN(n4530) );
  NAND2_X1 U4181 ( .A1(n3007), .A2(n4530), .ZN(n3642) );
  NAND2_X1 U4182 ( .A1(n2496), .A2(REG1_REG_17__SCAN_IN), .ZN(n3641) );
  NAND2_X1 U4183 ( .A1(n3353), .A2(REG2_REG_17__SCAN_IN), .ZN(n3640) );
  NAND2_X1 U4184 ( .A1(n3046), .A2(REG0_REG_17__SCAN_IN), .ZN(n3639) );
  INV_X1 U4185 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4935) );
  NOR2_X1 U4186 ( .A1(STATE_REG_SCAN_IN), .A2(n4935), .ZN(n4296) );
  AOI21_X1 U4187 ( .B1(n5296), .B2(n4505), .A(n4296), .ZN(n3643) );
  OAI211_X1 U4188 ( .C1(n3692), .C2(n5300), .A(n3644), .B(n3643), .ZN(n3645)
         );
  INV_X1 U4189 ( .A(n3645), .ZN(n3646) );
  OAI21_X1 U4190 ( .B1(n3647), .B2(n5291), .A(n3646), .ZN(U3223) );
  AND2_X2 U4191 ( .A1(n3648), .A2(n3657), .ZN(n4562) );
  NOR2_X1 U4192 ( .A1(n3649), .A2(n3657), .ZN(n3650) );
  OR2_X1 U4193 ( .A1(n4562), .A2(n3650), .ZN(n5310) );
  AND2_X1 U4194 ( .A1(n3680), .A2(n5340), .ZN(n3659) );
  AND2_X1 U4195 ( .A1(n3654), .A2(n3653), .ZN(n4120) );
  NAND2_X1 U4196 ( .A1(n3655), .A2(n4120), .ZN(n3656) );
  NAND2_X1 U4197 ( .A1(n3656), .A2(n4118), .ZN(n4194) );
  OAI22_X1 U4198 ( .A1(n3680), .A2(n5272), .B1(n4554), .B2(n4194), .ZN(n3658)
         );
  NAND2_X1 U4199 ( .A1(n4549), .A2(n3679), .ZN(n4552) );
  NAND2_X1 U4200 ( .A1(n3657), .A2(n5295), .ZN(n4100) );
  MUX2_X1 U4201 ( .A(n3659), .B(n3658), .S(n2565), .Z(n3663) );
  NAND2_X2 U4202 ( .A1(n4194), .A2(n4155), .ZN(n4553) );
  AOI22_X1 U4203 ( .A1(n4525), .A2(n4241), .B1(n4242), .B2(n4504), .ZN(n3661)
         );
  NAND2_X1 U4204 ( .A1(n3679), .A2(n4560), .ZN(n3660) );
  OAI211_X1 U4205 ( .C1(n4553), .C2(n4554), .A(n3661), .B(n3660), .ZN(n3662)
         );
  NOR2_X1 U4206 ( .A1(n3663), .A2(n3662), .ZN(n5314) );
  INV_X1 U4207 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3664) );
  MUX2_X1 U4208 ( .A(n5314), .B(n3664), .S(n5345), .Z(n3665) );
  OAI21_X1 U4209 ( .B1(n5310), .B2(n4666), .A(n3665), .ZN(U3495) );
  MUX2_X1 U4210 ( .A(n5314), .B(n4281), .S(n5342), .Z(n3666) );
  OAI21_X1 U4211 ( .B1(n5310), .B2(n4628), .A(n3666), .ZN(U3532) );
  AOI21_X1 U4212 ( .B1(n5278), .B2(n3668), .A(n3667), .ZN(n3677) );
  AOI21_X1 U4213 ( .B1(n5196), .B2(ADDR_REG_12__SCAN_IN), .A(n3669), .ZN(n3670) );
  OAI21_X1 U4214 ( .B1(n5181), .B2(n3671), .A(n3670), .ZN(n3676) );
  AOI211_X1 U4215 ( .C1(n3674), .C2(n3673), .A(n3672), .B(n5200), .ZN(n3675)
         );
  AOI211_X1 U4216 ( .C1(n5177), .C2(n3677), .A(n3676), .B(n3675), .ZN(n3678)
         );
  INV_X1 U4217 ( .A(n3678), .ZN(U3252) );
  NOR2_X1 U4218 ( .A1(n4241), .A2(n4559), .ZN(n3681) );
  OAI22_X1 U4219 ( .A1(n4540), .A2(n3681), .B1(n3682), .B2(n4561), .ZN(n3895)
         );
  NAND2_X1 U4220 ( .A1(n3690), .A2(n4240), .ZN(n3911) );
  INV_X1 U4221 ( .A(n3911), .ZN(n4454) );
  NOR2_X1 U4222 ( .A1(n3690), .A2(n4240), .ZN(n4198) );
  XNOR2_X1 U4223 ( .A(n3895), .B(n4156), .ZN(n4625) );
  INV_X1 U4224 ( .A(n4625), .ZN(n3696) );
  NAND2_X1 U4225 ( .A1(n3682), .A2(n4559), .ZN(n4191) );
  NAND2_X1 U4226 ( .A1(n4561), .A2(n4241), .ZN(n4101) );
  NAND2_X1 U4227 ( .A1(n4191), .A2(n4101), .ZN(n4541) );
  INV_X1 U4228 ( .A(n4552), .ZN(n4193) );
  NOR2_X1 U4229 ( .A1(n4541), .A2(n4193), .ZN(n3683) );
  NAND2_X1 U4230 ( .A1(n4550), .A2(n4101), .ZN(n3684) );
  NAND3_X1 U4231 ( .A1(n4550), .A2(n3685), .A3(n4101), .ZN(n3686) );
  NAND3_X1 U4232 ( .A1(n4453), .A2(n4501), .A3(n3686), .ZN(n3688) );
  AOI22_X1 U4233 ( .A1(n4504), .A2(n4241), .B1(n4505), .B2(n4525), .ZN(n3687)
         );
  OAI211_X1 U4234 ( .C1(n4581), .C2(n3690), .A(n3688), .B(n3687), .ZN(n4624)
         );
  NAND2_X1 U4235 ( .A1(n4562), .A2(n4561), .ZN(n3689) );
  INV_X1 U4236 ( .A(n3689), .ZN(n3691) );
  OAI21_X1 U4237 ( .B1(n3691), .B2(n3690), .A(n4526), .ZN(n4667) );
  NOR2_X1 U4238 ( .A1(n4667), .A2(n5309), .ZN(n3694) );
  OAI22_X1 U4239 ( .A1(n4545), .A2(n4293), .B1(n3692), .B2(n5307), .ZN(n3693)
         );
  AOI211_X1 U4240 ( .C1(n4624), .C2(n4545), .A(n3694), .B(n3693), .ZN(n3695)
         );
  OAI21_X1 U4241 ( .B1(n3696), .B2(n4518), .A(n3695), .ZN(U3274) );
  NAND2_X1 U4242 ( .A1(n2499), .A2(n4505), .ZN(n3698) );
  MUX2_X1 U4243 ( .A(n5156), .B(DATAI_17_), .S(n2488), .Z(n3938) );
  NAND2_X1 U4244 ( .A1(n3826), .A2(n3938), .ZN(n3697) );
  NAND2_X1 U4245 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  XNOR2_X1 U4246 ( .A(n3699), .B(n3810), .ZN(n3701) );
  NOR2_X1 U4247 ( .A1(n3128), .A2(n3897), .ZN(n3700) );
  AOI21_X1 U4248 ( .B1(n3831), .B2(n4505), .A(n3700), .ZN(n3702) );
  NAND2_X1 U4249 ( .A1(n3701), .A2(n3702), .ZN(n4041) );
  INV_X1 U4250 ( .A(n3701), .ZN(n3704) );
  INV_X1 U4251 ( .A(n3702), .ZN(n3703) );
  NAND2_X1 U4252 ( .A1(n3704), .A2(n3703), .ZN(n3705) );
  AND2_X1 U4253 ( .A1(n4041), .A2(n3705), .ZN(n3712) );
  NAND2_X1 U4254 ( .A1(n3707), .A2(n3706), .ZN(n3709) );
  NAND2_X1 U4255 ( .A1(n3709), .A2(n3708), .ZN(n3710) );
  NAND2_X1 U4256 ( .A1(n3710), .A2(n3712), .ZN(n3724) );
  OAI21_X1 U4257 ( .B1(n3712), .B2(n3710), .A(n3711), .ZN(n3713) );
  INV_X1 U4258 ( .A(n3713), .ZN(n3723) );
  OAI21_X1 U4259 ( .B1(n3714), .B2(REG3_REG_18__SCAN_IN), .A(n3737), .ZN(n4513) );
  NAND2_X1 U4260 ( .A1(n3353), .A2(REG2_REG_18__SCAN_IN), .ZN(n3716) );
  NAND2_X1 U4261 ( .A1(n3046), .A2(REG0_REG_18__SCAN_IN), .ZN(n3715) );
  AND2_X1 U4262 ( .A1(n3716), .A2(n3715), .ZN(n3718) );
  NAND2_X1 U4263 ( .A1(n2497), .A2(REG1_REG_18__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4264 ( .A1(n5296), .A2(n4524), .B1(n5282), .B2(n3938), .ZN(n3722)
         );
  NOR2_X1 U4265 ( .A1(STATE_REG_SCAN_IN), .A2(n3719), .ZN(n5163) );
  NOR2_X1 U4266 ( .A1(n4071), .A2(n4547), .ZN(n3720) );
  AOI211_X1 U4267 ( .C1(n4068), .C2(n4530), .A(n5163), .B(n3720), .ZN(n3721)
         );
  OAI211_X1 U4268 ( .C1(n3723), .C2(n5291), .A(n3722), .B(n3721), .ZN(U3225)
         );
  NAND2_X1 U4269 ( .A1(n3724), .A2(n4041), .ZN(n3734) );
  NAND2_X1 U4270 ( .A1(n4524), .A2(n2499), .ZN(n3726) );
  MUX2_X1 U4271 ( .A(n5327), .B(DATAI_18_), .S(n2488), .Z(n4503) );
  NAND2_X1 U4272 ( .A1(n3826), .A2(n4503), .ZN(n3725) );
  NAND2_X1 U4273 ( .A1(n3726), .A2(n3725), .ZN(n3727) );
  XNOR2_X1 U4274 ( .A(n3727), .B(n3810), .ZN(n3729) );
  NOR2_X1 U4275 ( .A1(n3128), .A2(n4510), .ZN(n3728) );
  AOI21_X1 U4276 ( .B1(n3831), .B2(n4524), .A(n3728), .ZN(n3730) );
  NAND2_X1 U4277 ( .A1(n3729), .A2(n3730), .ZN(n3735) );
  INV_X1 U4278 ( .A(n3729), .ZN(n3732) );
  INV_X1 U4279 ( .A(n3730), .ZN(n3731) );
  NAND2_X1 U4280 ( .A1(n3732), .A2(n3731), .ZN(n3733) );
  AND2_X1 U4281 ( .A1(n3735), .A2(n3733), .ZN(n4043) );
  NAND2_X1 U4282 ( .A1(n3734), .A2(n4043), .ZN(n4044) );
  NAND2_X1 U4283 ( .A1(n4044), .A2(n3735), .ZN(n3963) );
  NAND2_X1 U4284 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  NAND2_X1 U4285 ( .A1(n3752), .A2(n3738), .ZN(n4492) );
  OR2_X1 U4286 ( .A1(n4492), .A2(n3836), .ZN(n3743) );
  NAND2_X1 U4287 ( .A1(n2496), .A2(REG1_REG_19__SCAN_IN), .ZN(n3740) );
  NAND2_X1 U4288 ( .A1(n3046), .A2(REG0_REG_19__SCAN_IN), .ZN(n3739) );
  OAI211_X1 U4289 ( .C1(n3156), .C2(n2755), .A(n3740), .B(n3739), .ZN(n3741)
         );
  INV_X1 U4290 ( .A(n3741), .ZN(n3742) );
  NAND2_X1 U4291 ( .A1(n4465), .A2(n2499), .ZN(n3745) );
  MUX2_X1 U4292 ( .A(n4674), .B(DATAI_19_), .S(n2488), .Z(n4481) );
  NAND2_X1 U4293 ( .A1(n3826), .A2(n4481), .ZN(n3744) );
  NAND2_X1 U4294 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  XNOR2_X1 U4295 ( .A(n3746), .B(n3873), .ZN(n3748) );
  NOR2_X1 U4296 ( .A1(n3128), .A2(n4489), .ZN(n3747) );
  AOI21_X1 U4297 ( .B1(n3831), .B2(n4465), .A(n3747), .ZN(n3749) );
  XNOR2_X1 U4298 ( .A(n3748), .B(n3749), .ZN(n3964) );
  INV_X1 U4299 ( .A(n3748), .ZN(n3750) );
  NAND2_X1 U4300 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  INV_X1 U4301 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U4302 ( .A1(n3752), .A2(n4755), .ZN(n3753) );
  NAND2_X1 U4303 ( .A1(n3768), .A2(n3753), .ZN(n4475) );
  OR2_X1 U4304 ( .A1(n4475), .A2(n3836), .ZN(n3758) );
  INV_X1 U4305 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U4306 ( .A1(n2497), .A2(REG1_REG_20__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4307 ( .A1(n3353), .A2(REG2_REG_20__SCAN_IN), .ZN(n3754) );
  OAI211_X1 U4308 ( .C1(n4660), .C2(n3884), .A(n3755), .B(n3754), .ZN(n3756)
         );
  INV_X1 U4309 ( .A(n3756), .ZN(n3757) );
  NAND2_X1 U4310 ( .A1(n4439), .A2(n2499), .ZN(n3760) );
  NAND2_X1 U4311 ( .A1(n3826), .A2(n4464), .ZN(n3759) );
  NAND2_X1 U4312 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  XNOR2_X1 U4313 ( .A(n3761), .B(n3873), .ZN(n3764) );
  NAND2_X1 U4314 ( .A1(n4439), .A2(n3831), .ZN(n3763) );
  NAND2_X1 U4315 ( .A1(n2499), .A2(n4464), .ZN(n3762) );
  NAND2_X1 U4316 ( .A1(n3763), .A2(n3762), .ZN(n3765) );
  NAND2_X1 U4317 ( .A1(n3764), .A2(n3765), .ZN(n4024) );
  INV_X1 U4318 ( .A(n3764), .ZN(n3767) );
  INV_X1 U4319 ( .A(n3765), .ZN(n3766) );
  NAND2_X1 U4320 ( .A1(n3767), .A2(n3766), .ZN(n4023) );
  INV_X1 U4321 ( .A(n3984), .ZN(n3780) );
  NAND2_X1 U4322 ( .A1(n3768), .A2(n4928), .ZN(n3769) );
  AND2_X1 U4323 ( .A1(n3785), .A2(n3769), .ZN(n4447) );
  NAND2_X1 U4324 ( .A1(n4447), .A2(n3007), .ZN(n3774) );
  INV_X1 U4325 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4656) );
  NAND2_X1 U4326 ( .A1(n2497), .A2(REG1_REG_21__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4327 ( .A1(n3353), .A2(REG2_REG_21__SCAN_IN), .ZN(n3770) );
  OAI211_X1 U4328 ( .C1(n4656), .C2(n3884), .A(n3771), .B(n3770), .ZN(n3772)
         );
  INV_X1 U4329 ( .A(n3772), .ZN(n3773) );
  NAND2_X1 U4330 ( .A1(n4419), .A2(n2499), .ZN(n3776) );
  NAND2_X1 U4331 ( .A1(n3826), .A2(n4444), .ZN(n3775) );
  NAND2_X1 U4332 ( .A1(n3776), .A2(n3775), .ZN(n3777) );
  XNOR2_X1 U4333 ( .A(n3777), .B(n3810), .ZN(n3781) );
  NOR2_X1 U4334 ( .A1(n3128), .A2(n3939), .ZN(n3778) );
  AOI21_X1 U4335 ( .B1(n4419), .B2(n3831), .A(n3778), .ZN(n3782) );
  AND2_X1 U4336 ( .A1(n3781), .A2(n3782), .ZN(n3986) );
  INV_X1 U4337 ( .A(n3781), .ZN(n3784) );
  INV_X1 U4338 ( .A(n3782), .ZN(n3783) );
  NAND2_X1 U4339 ( .A1(n3784), .A2(n3783), .ZN(n3983) );
  INV_X1 U4340 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4036) );
  NAND2_X1 U4341 ( .A1(n3785), .A2(n4036), .ZN(n3786) );
  NAND2_X1 U4342 ( .A1(n3801), .A2(n3786), .ZN(n4035) );
  INV_X1 U4343 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U4344 ( .A1(n2496), .A2(REG1_REG_22__SCAN_IN), .ZN(n3788) );
  NAND2_X1 U4345 ( .A1(n3353), .A2(REG2_REG_22__SCAN_IN), .ZN(n3787) );
  OAI211_X1 U4346 ( .C1(n4652), .C2(n3884), .A(n3788), .B(n3787), .ZN(n3789)
         );
  INV_X1 U4347 ( .A(n3789), .ZN(n3790) );
  NAND2_X1 U4348 ( .A1(n4433), .A2(n2499), .ZN(n3793) );
  NAND2_X1 U4349 ( .A1(n3826), .A2(n4418), .ZN(n3792) );
  NAND2_X1 U4350 ( .A1(n3793), .A2(n3792), .ZN(n3794) );
  XNOR2_X1 U4351 ( .A(n3794), .B(n3810), .ZN(n3798) );
  INV_X1 U4352 ( .A(n4418), .ZN(n4425) );
  NOR2_X1 U4353 ( .A1(n2491), .A2(n4425), .ZN(n3795) );
  AOI21_X1 U4354 ( .B1(n4433), .B2(n3831), .A(n3795), .ZN(n3797) );
  XNOR2_X1 U4355 ( .A(n3798), .B(n3797), .ZN(n4034) );
  NAND2_X1 U4356 ( .A1(n3798), .A2(n3797), .ZN(n3799) );
  NAND2_X1 U4357 ( .A1(n4032), .A2(n3799), .ZN(n3955) );
  INV_X1 U4358 ( .A(n3955), .ZN(n3814) );
  NAND2_X1 U4359 ( .A1(n3801), .A2(n3800), .ZN(n3802) );
  AND2_X1 U4360 ( .A1(n3818), .A2(n3802), .ZN(n4407) );
  NAND2_X1 U4361 ( .A1(n4407), .A2(n3007), .ZN(n3807) );
  INV_X1 U4362 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U4363 ( .A1(n2496), .A2(REG1_REG_23__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4364 ( .A1(n3353), .A2(REG2_REG_23__SCAN_IN), .ZN(n3803) );
  OAI211_X1 U4365 ( .C1(n4648), .C2(n3884), .A(n3804), .B(n3803), .ZN(n3805)
         );
  INV_X1 U4366 ( .A(n3805), .ZN(n3806) );
  NAND2_X1 U4367 ( .A1(n4379), .A2(n2499), .ZN(n3809) );
  NAND2_X1 U4368 ( .A1(n3826), .A2(n4398), .ZN(n3808) );
  NAND2_X1 U4369 ( .A1(n3809), .A2(n3808), .ZN(n3811) );
  XNOR2_X1 U4370 ( .A(n3811), .B(n3810), .ZN(n3816) );
  NOR2_X1 U4371 ( .A1(n3128), .A2(n4406), .ZN(n3812) );
  AOI21_X1 U4372 ( .B1(n4379), .B2(n3831), .A(n3812), .ZN(n3815) );
  XNOR2_X1 U4373 ( .A(n3816), .B(n3815), .ZN(n3956) );
  NAND2_X1 U4374 ( .A1(n3814), .A2(n3813), .ZN(n3953) );
  OR2_X1 U4375 ( .A1(n3816), .A2(n3815), .ZN(n3817) );
  NAND2_X1 U4376 ( .A1(n3953), .A2(n3817), .ZN(n3833) );
  INV_X1 U4377 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U4378 ( .A1(n3818), .A2(n4939), .ZN(n3819) );
  NAND2_X1 U4379 ( .A1(n3834), .A2(n3819), .ZN(n4385) );
  INV_X1 U4380 ( .A(REG0_REG_24__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4381 ( .A1(n2497), .A2(REG1_REG_24__SCAN_IN), .ZN(n3821) );
  NAND2_X1 U4382 ( .A1(n3353), .A2(REG2_REG_24__SCAN_IN), .ZN(n3820) );
  OAI211_X1 U4383 ( .C1(n3822), .C2(n3884), .A(n3821), .B(n3820), .ZN(n3823)
         );
  INV_X1 U4384 ( .A(n3823), .ZN(n3824) );
  NAND2_X1 U4385 ( .A1(n4399), .A2(n2498), .ZN(n3828) );
  NAND2_X1 U4386 ( .A1(n3826), .A2(n4378), .ZN(n3827) );
  NAND2_X1 U4387 ( .A1(n3828), .A2(n3827), .ZN(n3829) );
  XNOR2_X1 U4388 ( .A(n3829), .B(n3873), .ZN(n3832) );
  AOI22_X1 U4389 ( .A1(n4399), .A2(n3831), .B1(n2499), .B2(n4378), .ZN(n4005)
         );
  NAND2_X1 U4390 ( .A1(n3833), .A2(n3832), .ZN(n4003) );
  OAI21_X1 U4391 ( .B1(n4002), .B2(n4005), .A(n4003), .ZN(n3994) );
  NAND2_X1 U4392 ( .A1(n3834), .A2(n4741), .ZN(n3835) );
  NAND2_X1 U4393 ( .A1(n3859), .A2(n3835), .ZN(n4366) );
  INV_X1 U4394 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4643) );
  NAND2_X1 U4395 ( .A1(n2497), .A2(REG1_REG_25__SCAN_IN), .ZN(n3838) );
  NAND2_X1 U4396 ( .A1(n3353), .A2(REG2_REG_25__SCAN_IN), .ZN(n3837) );
  OAI211_X1 U4397 ( .C1(n3884), .C2(n4643), .A(n3838), .B(n3837), .ZN(n3839)
         );
  INV_X1 U4398 ( .A(n3839), .ZN(n3840) );
  NAND2_X1 U4399 ( .A1(n4344), .A2(n2499), .ZN(n3843) );
  NAND2_X1 U4400 ( .A1(n3826), .A2(n4360), .ZN(n3842) );
  NAND2_X1 U4401 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  XNOR2_X1 U4402 ( .A(n3844), .B(n3873), .ZN(n3845) );
  OAI22_X1 U4403 ( .A1(n4381), .A2(n2493), .B1(n2490), .B2(n4364), .ZN(n3846)
         );
  XNOR2_X1 U4404 ( .A(n3845), .B(n3846), .ZN(n3996) );
  INV_X1 U4405 ( .A(n3845), .ZN(n3848) );
  INV_X1 U4406 ( .A(n3846), .ZN(n3847) );
  XNOR2_X1 U4407 ( .A(n3859), .B(REG3_REG_26__SCAN_IN), .ZN(n4349) );
  INV_X1 U4408 ( .A(REG0_REG_26__SCAN_IN), .ZN(n3852) );
  NAND2_X1 U4409 ( .A1(n2496), .A2(REG1_REG_26__SCAN_IN), .ZN(n3851) );
  NAND2_X1 U4410 ( .A1(n3353), .A2(REG2_REG_26__SCAN_IN), .ZN(n3850) );
  OAI211_X1 U4411 ( .C1(n3852), .C2(n3884), .A(n3851), .B(n3850), .ZN(n3853)
         );
  NAND2_X1 U4412 ( .A1(n2488), .A2(DATAI_26_), .ZN(n4342) );
  OAI22_X1 U4413 ( .A1(n3928), .A2(n2491), .B1(n3872), .B2(n4342), .ZN(n3854)
         );
  XNOR2_X1 U4414 ( .A(n3854), .B(n3873), .ZN(n4066) );
  OAI22_X1 U4415 ( .A1(n3928), .A2(n2493), .B1(n4342), .B2(n3128), .ZN(n3856)
         );
  INV_X1 U4416 ( .A(n3856), .ZN(n4065) );
  INV_X1 U4417 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3858) );
  INV_X1 U4418 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4914) );
  OAI21_X1 U4419 ( .B1(n3859), .B2(n3858), .A(n4914), .ZN(n3860) );
  NAND2_X1 U4420 ( .A1(n4332), .A2(n3007), .ZN(n3866) );
  INV_X1 U4421 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U4422 ( .A1(n3006), .A2(REG1_REG_27__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4423 ( .A1(n3353), .A2(REG2_REG_27__SCAN_IN), .ZN(n3862) );
  OAI211_X1 U4424 ( .C1(n4638), .C2(n3884), .A(n3863), .B(n3862), .ZN(n3864)
         );
  INV_X1 U4425 ( .A(n3864), .ZN(n3865) );
  INV_X1 U4426 ( .A(n4341), .ZN(n3907) );
  OAI22_X1 U4427 ( .A1(n3907), .A2(n2493), .B1(n2491), .B2(n4330), .ZN(n3870)
         );
  NAND2_X1 U4428 ( .A1(n4341), .A2(n2499), .ZN(n3868) );
  NAND2_X1 U4429 ( .A1(n3826), .A2(n3947), .ZN(n3867) );
  NAND2_X1 U4430 ( .A1(n3868), .A2(n3867), .ZN(n3869) );
  XNOR2_X1 U4431 ( .A(n3869), .B(n3873), .ZN(n3871) );
  XOR2_X1 U4432 ( .A(n3870), .B(n3871), .Z(n3946) );
  AOI21_X2 U4433 ( .B1(n3945), .B2(n3946), .A(n2654), .ZN(n3879) );
  NAND2_X1 U4434 ( .A1(n2488), .A2(DATAI_28_), .ZN(n4314) );
  OAI22_X1 U4435 ( .A1(n4324), .A2(n3128), .B1(n3872), .B2(n4314), .ZN(n3874)
         );
  XNOR2_X1 U4436 ( .A(n3874), .B(n3873), .ZN(n3877) );
  OAI22_X1 U4437 ( .A1(n4324), .A2(n2493), .B1(n3128), .B2(n4314), .ZN(n3876)
         );
  XNOR2_X1 U4438 ( .A(n3877), .B(n3876), .ZN(n3878) );
  XNOR2_X1 U4439 ( .A(n3879), .B(n3878), .ZN(n3892) );
  INV_X1 U4440 ( .A(n3880), .ZN(n3940) );
  NAND2_X1 U4441 ( .A1(n3940), .A2(n3007), .ZN(n3887) );
  INV_X1 U4442 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3883) );
  NAND2_X1 U4443 ( .A1(n3006), .A2(REG1_REG_29__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4444 ( .A1(n3353), .A2(REG2_REG_29__SCAN_IN), .ZN(n3881) );
  OAI211_X1 U4445 ( .C1(n3884), .C2(n3883), .A(n3882), .B(n3881), .ZN(n3885)
         );
  INV_X1 U4446 ( .A(n3885), .ZN(n3886) );
  NAND2_X1 U4447 ( .A1(n3887), .A2(n3886), .ZN(n4239) );
  NAND2_X1 U4448 ( .A1(n4239), .A2(n5296), .ZN(n3889) );
  INV_X1 U4449 ( .A(n4314), .ZN(n3909) );
  AOI22_X1 U4450 ( .A1(n5282), .A2(n3909), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3888) );
  OAI211_X1 U4451 ( .C1(n4315), .C2(n5300), .A(n3889), .B(n3888), .ZN(n3890)
         );
  AOI21_X1 U4452 ( .B1(n5284), .B2(n4341), .A(n3890), .ZN(n3891) );
  OAI21_X1 U4453 ( .B1(n3892), .B2(n5291), .A(n3891), .ZN(U3217) );
  NOR2_X1 U4454 ( .A1(n3897), .A2(n4505), .ZN(n4456) );
  INV_X1 U4455 ( .A(n4456), .ZN(n3896) );
  NAND2_X1 U4456 ( .A1(n3897), .A2(n4505), .ZN(n4457) );
  NAND2_X1 U4457 ( .A1(n3896), .A2(n4457), .ZN(n4536) );
  NAND2_X1 U4458 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U4459 ( .A1(n4535), .A2(n3899), .ZN(n4498) );
  NOR2_X1 U4460 ( .A1(n4524), .A2(n4510), .ZN(n3913) );
  INV_X1 U4461 ( .A(n3913), .ZN(n4458) );
  NAND2_X1 U4462 ( .A1(n4524), .A2(n4510), .ZN(n4478) );
  NAND2_X1 U4463 ( .A1(n4458), .A2(n4478), .ZN(n4499) );
  NAND2_X1 U4464 ( .A1(n4498), .A2(n4499), .ZN(n4497) );
  NAND2_X1 U4465 ( .A1(n4497), .A2(n2504), .ZN(n4486) );
  NAND2_X1 U4466 ( .A1(n4486), .A2(n2521), .ZN(n3901) );
  OR2_X1 U4467 ( .A1(n4439), .A2(n4473), .ZN(n3914) );
  NAND2_X1 U4468 ( .A1(n4439), .A2(n4473), .ZN(n3916) );
  NAND2_X1 U4469 ( .A1(n3914), .A2(n3916), .ZN(n4462) );
  NAND2_X1 U4470 ( .A1(n4433), .A2(n4425), .ZN(n3918) );
  NAND2_X1 U4471 ( .A1(n4395), .A2(n3918), .ZN(n4394) );
  NOR2_X1 U4472 ( .A1(n4379), .A2(n4398), .ZN(n4181) );
  NAND2_X1 U4473 ( .A1(n4379), .A2(n4398), .ZN(n4180) );
  NAND2_X1 U4474 ( .A1(n4399), .A2(n4386), .ZN(n4356) );
  NAND2_X1 U4475 ( .A1(n3924), .A2(n4356), .ZN(n4373) );
  NAND2_X1 U4476 ( .A1(n4337), .A2(n3904), .ZN(n3906) );
  NOR2_X1 U4477 ( .A1(n4324), .A2(n3909), .ZN(n4131) );
  NAND2_X1 U4478 ( .A1(n2488), .A2(DATAI_29_), .ZN(n4210) );
  XNOR2_X1 U4479 ( .A(n4239), .B(n4210), .ZN(n4138) );
  NAND2_X1 U4480 ( .A1(n4465), .A2(n4489), .ZN(n4154) );
  AND2_X1 U4481 ( .A1(n4478), .A2(n4154), .ZN(n4461) );
  AND2_X1 U4482 ( .A1(n4457), .A2(n3911), .ZN(n3912) );
  NAND2_X1 U4483 ( .A1(n4453), .A2(n4197), .ZN(n4435) );
  OAI21_X1 U4484 ( .B1(n3913), .B2(n4456), .A(n4461), .ZN(n3915) );
  NAND2_X1 U4485 ( .A1(n4508), .A2(n4481), .ZN(n4459) );
  NAND3_X1 U4486 ( .A1(n3915), .A2(n3914), .A3(n4459), .ZN(n3917) );
  NAND2_X1 U4487 ( .A1(n3917), .A2(n3916), .ZN(n4434) );
  OR2_X1 U4488 ( .A1(n4419), .A2(n3939), .ZN(n4176) );
  NAND2_X1 U4489 ( .A1(n4435), .A2(n4202), .ZN(n3923) );
  NAND2_X1 U4490 ( .A1(n4419), .A2(n3939), .ZN(n4415) );
  NAND2_X1 U4491 ( .A1(n3918), .A2(n4415), .ZN(n3919) );
  NAND2_X1 U4492 ( .A1(n3919), .A2(n4395), .ZN(n3921) );
  NAND2_X1 U4493 ( .A1(n4379), .A2(n4406), .ZN(n3920) );
  NAND2_X1 U4494 ( .A1(n3921), .A2(n3920), .ZN(n4200) );
  INV_X1 U4495 ( .A(n4200), .ZN(n3922) );
  NAND2_X1 U4496 ( .A1(n3923), .A2(n3922), .ZN(n4375) );
  OR2_X1 U4497 ( .A1(n4379), .A2(n4406), .ZN(n4374) );
  NAND2_X1 U4498 ( .A1(n3924), .A2(n4374), .ZN(n4203) );
  INV_X1 U4499 ( .A(n4203), .ZN(n3925) );
  NAND2_X1 U4500 ( .A1(n4375), .A2(n3925), .ZN(n4357) );
  NAND2_X1 U4501 ( .A1(n4344), .A2(n4364), .ZN(n4141) );
  NAND2_X1 U4502 ( .A1(n4141), .A2(n4356), .ZN(n4208) );
  INV_X1 U4503 ( .A(n4208), .ZN(n4128) );
  NAND2_X1 U4504 ( .A1(n4357), .A2(n4128), .ZN(n3927) );
  NOR2_X1 U4505 ( .A1(n4344), .A2(n4364), .ZN(n4143) );
  INV_X1 U4506 ( .A(n4143), .ZN(n3926) );
  NAND2_X1 U4507 ( .A1(n3927), .A2(n3926), .ZN(n4340) );
  OR2_X1 U4508 ( .A1(n3928), .A2(n3902), .ZN(n4130) );
  AND2_X1 U4509 ( .A1(n3928), .A2(n3902), .ZN(n4139) );
  AND2_X1 U4510 ( .A1(n4341), .A2(n4330), .ZN(n4134) );
  NOR2_X1 U4511 ( .A1(n4341), .A2(n4330), .ZN(n4205) );
  NOR2_X1 U4512 ( .A1(n4323), .A2(n4322), .ZN(n4321) );
  INV_X1 U4513 ( .A(n4303), .ZN(n4307) );
  NOR2_X1 U4514 ( .A1(n4308), .A2(n4307), .ZN(n4306) );
  NOR2_X1 U4515 ( .A1(n4306), .A2(n4206), .ZN(n3929) );
  XNOR2_X1 U4516 ( .A(n3929), .B(n4138), .ZN(n3937) );
  NAND2_X1 U4517 ( .A1(n3006), .A2(REG1_REG_30__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U4518 ( .A1(n3353), .A2(REG2_REG_30__SCAN_IN), .ZN(n3931) );
  NAND2_X1 U4519 ( .A1(n3046), .A2(REG0_REG_30__SCAN_IN), .ZN(n3930) );
  NAND3_X1 U4520 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n4238) );
  INV_X1 U4521 ( .A(B_REG_SCAN_IN), .ZN(n3933) );
  NOR2_X1 U4522 ( .A1(n5183), .A2(n3933), .ZN(n3934) );
  NOR2_X1 U4523 ( .A1(n4546), .A2(n3934), .ZN(n4571) );
  INV_X1 U4524 ( .A(n4210), .ZN(n4133) );
  AOI22_X1 U4525 ( .A1(n4238), .A2(n4571), .B1(n4560), .B2(n4133), .ZN(n3935)
         );
  OAI21_X1 U4526 ( .B1(n4324), .B2(n4548), .A(n3935), .ZN(n3936) );
  INV_X1 U4527 ( .A(n4588), .ZN(n3943) );
  AND2_X2 U4528 ( .A1(n4509), .A2(n4510), .ZN(n4488) );
  AND2_X2 U4529 ( .A1(n4403), .A2(n4406), .ZN(n4404) );
  AND2_X2 U4530 ( .A1(n4404), .A2(n4386), .ZN(n4388) );
  NAND2_X1 U4531 ( .A1(n4388), .A2(n4364), .ZN(n4350) );
  OR2_X2 U4532 ( .A1(n4350), .A2(n3902), .ZN(n4598) );
  NOR2_X4 U4533 ( .A1(n4598), .A2(n3947), .ZN(n4328) );
  AOI22_X1 U4534 ( .A1(n3940), .A2(n5302), .B1(REG2_REG_29__SCAN_IN), .B2(
        n5356), .ZN(n3941) );
  OAI21_X1 U4535 ( .B1(n4586), .B2(n5309), .A(n3941), .ZN(n3942) );
  AOI21_X1 U4536 ( .B1(n3943), .B2(n4545), .A(n3942), .ZN(n3944) );
  OAI21_X1 U4537 ( .B1(n4589), .B2(n4518), .A(n3944), .ZN(U3354) );
  XNOR2_X1 U4538 ( .A(n3945), .B(n3946), .ZN(n3952) );
  INV_X1 U4539 ( .A(n5296), .ZN(n4007) );
  AOI22_X1 U4540 ( .A1(n5282), .A2(n3947), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3949) );
  NAND2_X1 U4541 ( .A1(n4332), .A2(n4068), .ZN(n3948) );
  OAI211_X1 U4542 ( .C1(n4324), .C2(n4007), .A(n3949), .B(n3948), .ZN(n3950)
         );
  AOI21_X1 U4543 ( .B1(n5284), .B2(n3903), .A(n3950), .ZN(n3951) );
  OAI21_X1 U4544 ( .B1(n3952), .B2(n5291), .A(n3951), .ZN(U3211) );
  INV_X1 U4545 ( .A(n3953), .ZN(n3954) );
  AOI211_X1 U4546 ( .C1(n3956), .C2(n3955), .A(n5291), .B(n3954), .ZN(n3961)
         );
  INV_X1 U4547 ( .A(n4407), .ZN(n3959) );
  AOI22_X1 U4548 ( .A1(n4399), .A2(n5296), .B1(n5282), .B2(n4398), .ZN(n3958)
         );
  AOI22_X1 U4549 ( .A1(n5284), .A2(n4433), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3957) );
  OAI211_X1 U4550 ( .C1(n3959), .C2(n5300), .A(n3958), .B(n3957), .ZN(n3960)
         );
  OR2_X1 U4551 ( .A1(n3961), .A2(n3960), .ZN(U3213) );
  OAI21_X1 U4552 ( .B1(n3964), .B2(n3963), .A(n3962), .ZN(n3965) );
  INV_X1 U4553 ( .A(n3965), .ZN(n3970) );
  AOI22_X1 U4554 ( .A1(n5296), .A2(n4439), .B1(n5282), .B2(n4481), .ZN(n3969)
         );
  NOR2_X1 U4555 ( .A1(n5300), .A2(n4492), .ZN(n3966) );
  AOI211_X1 U4556 ( .C1(n5284), .C2(n4524), .A(n3967), .B(n3966), .ZN(n3968)
         );
  OAI211_X1 U4557 ( .C1(n3970), .C2(n5291), .A(n3969), .B(n3968), .ZN(U3216)
         );
  OAI21_X1 U4558 ( .B1(n3973), .B2(n3972), .A(n3971), .ZN(n3974) );
  NAND2_X1 U4559 ( .A1(n3974), .A2(n4055), .ZN(n3982) );
  AOI22_X1 U4560 ( .A1(n5296), .A2(n4245), .B1(n5282), .B2(n3975), .ZN(n3981)
         );
  NOR2_X1 U4561 ( .A1(n4071), .A2(n3976), .ZN(n3977) );
  AOI211_X1 U4562 ( .C1(n4068), .C2(n3979), .A(n3978), .B(n3977), .ZN(n3980)
         );
  NAND3_X1 U4563 ( .A1(n3982), .A2(n3981), .A3(n3980), .ZN(U3218) );
  INV_X1 U4564 ( .A(n3983), .ZN(n3987) );
  OAI21_X1 U4565 ( .B1(n3987), .B2(n3986), .A(n3985), .ZN(n3988) );
  AOI22_X1 U4566 ( .A1(n3989), .A2(n3988), .B1(n3780), .B2(n3987), .ZN(n3993)
         );
  AOI22_X1 U4567 ( .A1(n5296), .A2(n4433), .B1(n5282), .B2(n4444), .ZN(n3992)
         );
  OAI22_X1 U4568 ( .A1(n4071), .A2(n4483), .B1(STATE_REG_SCAN_IN), .B2(n4928), 
        .ZN(n3990) );
  AOI21_X1 U4569 ( .B1(n4447), .B2(n4068), .A(n3990), .ZN(n3991) );
  OAI211_X1 U4570 ( .C1(n3993), .C2(n5291), .A(n3992), .B(n3991), .ZN(U3220)
         );
  AOI21_X1 U4571 ( .B1(n3996), .B2(n3994), .A(n3995), .ZN(n4001) );
  AOI22_X1 U4572 ( .A1(n4399), .A2(n5284), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3998) );
  NAND2_X1 U4573 ( .A1(n5282), .A2(n4360), .ZN(n3997) );
  OAI211_X1 U4574 ( .C1(n5300), .C2(n4366), .A(n3998), .B(n3997), .ZN(n3999)
         );
  AOI21_X1 U4575 ( .B1(n3903), .B2(n5296), .A(n3999), .ZN(n4000) );
  OAI21_X1 U4576 ( .B1(n4001), .B2(n5291), .A(n4000), .ZN(U3222) );
  INV_X1 U4577 ( .A(n4002), .ZN(n4004) );
  NAND2_X1 U4578 ( .A1(n4004), .A2(n4003), .ZN(n4006) );
  XNOR2_X1 U4579 ( .A(n4006), .B(n4005), .ZN(n4011) );
  INV_X1 U4580 ( .A(n4379), .ZN(n4422) );
  OAI22_X1 U4581 ( .A1(n4071), .A2(n4422), .B1(STATE_REG_SCAN_IN), .B2(n4939), 
        .ZN(n4009) );
  OAI22_X1 U4582 ( .A1(n4381), .A2(n4007), .B1(n5300), .B2(n4385), .ZN(n4008)
         );
  AOI211_X1 U4583 ( .C1(n4378), .C2(n5282), .A(n4009), .B(n4008), .ZN(n4010)
         );
  OAI21_X1 U4584 ( .B1(n4011), .B2(n5291), .A(n4010), .ZN(U3226) );
  OAI21_X1 U4585 ( .B1(n4013), .B2(n4012), .A(n3348), .ZN(n4014) );
  NAND2_X1 U4586 ( .A1(n4014), .A2(n4055), .ZN(n4021) );
  AOI22_X1 U4587 ( .A1(n5296), .A2(n4244), .B1(n5282), .B2(n4015), .ZN(n4020)
         );
  NOR2_X1 U4588 ( .A1(n4071), .A2(n4016), .ZN(n4017) );
  AOI211_X1 U4589 ( .C1(n4068), .C2(n5251), .A(n4018), .B(n4017), .ZN(n4019)
         );
  NAND3_X1 U4590 ( .A1(n4021), .A2(n4020), .A3(n4019), .ZN(U3228) );
  NAND2_X1 U4591 ( .A1(n4024), .A2(n4023), .ZN(n4025) );
  XNOR2_X1 U4592 ( .A(n4022), .B(n4025), .ZN(n4030) );
  AOI22_X1 U4593 ( .A1(n5296), .A2(n4419), .B1(n5282), .B2(n4464), .ZN(n4027)
         );
  AOI22_X1 U4594 ( .A1(n5284), .A2(n4465), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4026) );
  OAI211_X1 U4595 ( .C1(n4475), .C2(n5300), .A(n4027), .B(n4026), .ZN(n4028)
         );
  INV_X1 U4596 ( .A(n4028), .ZN(n4029) );
  OAI21_X1 U4597 ( .B1(n4030), .B2(n5291), .A(n4029), .ZN(U3230) );
  INV_X1 U4598 ( .A(n4032), .ZN(n4033) );
  AOI21_X1 U4599 ( .B1(n4034), .B2(n4031), .A(n4033), .ZN(n4040) );
  AOI22_X1 U4600 ( .A1(n5296), .A2(n4379), .B1(n5282), .B2(n4418), .ZN(n4039)
         );
  INV_X1 U4601 ( .A(n4035), .ZN(n4427) );
  OAI22_X1 U4602 ( .A1(n4071), .A2(n4467), .B1(STATE_REG_SCAN_IN), .B2(n4036), 
        .ZN(n4037) );
  AOI21_X1 U4603 ( .B1(n4427), .B2(n4068), .A(n4037), .ZN(n4038) );
  OAI211_X1 U4604 ( .C1(n4040), .C2(n5291), .A(n4039), .B(n4038), .ZN(U3232)
         );
  INV_X1 U4605 ( .A(n4041), .ZN(n4042) );
  NOR2_X1 U4606 ( .A1(n4043), .A2(n4042), .ZN(n4046) );
  INV_X1 U4607 ( .A(n4044), .ZN(n4045) );
  AOI21_X1 U4608 ( .B1(n4046), .B2(n3711), .A(n4045), .ZN(n4051) );
  AOI22_X1 U4609 ( .A1(n5296), .A2(n4465), .B1(n5282), .B2(n4503), .ZN(n4050)
         );
  NOR2_X1 U4610 ( .A1(n5300), .A2(n4513), .ZN(n4047) );
  AOI211_X1 U4611 ( .C1(n5284), .C2(n4505), .A(n4048), .B(n4047), .ZN(n4049)
         );
  OAI211_X1 U4612 ( .C1(n4051), .C2(n5291), .A(n4050), .B(n4049), .ZN(U3235)
         );
  NOR3_X1 U4613 ( .A1(n4054), .A2(n4053), .A3(n4052), .ZN(n4056) );
  OAI21_X1 U4614 ( .B1(n4056), .B2(n3186), .A(n4055), .ZN(n4064) );
  AOI22_X1 U4615 ( .A1(n5296), .A2(n4247), .B1(n5282), .B2(n4057), .ZN(n4063)
         );
  NOR2_X1 U4616 ( .A1(n4071), .A2(n4058), .ZN(n4059) );
  AOI211_X1 U4617 ( .C1(n4068), .C2(n4061), .A(n4060), .B(n4059), .ZN(n4062)
         );
  NAND3_X1 U4618 ( .A1(n4064), .A2(n4063), .A3(n4062), .ZN(U3236) );
  XNOR2_X1 U4619 ( .A(n4066), .B(n4065), .ZN(n4067) );
  XNOR2_X1 U4620 ( .A(n2508), .B(n4067), .ZN(n4074) );
  AOI22_X1 U4621 ( .A1(n5282), .A2(n3902), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4070) );
  NAND2_X1 U4622 ( .A1(n4349), .A2(n4068), .ZN(n4069) );
  OAI211_X1 U4623 ( .C1(n4381), .C2(n4071), .A(n4070), .B(n4069), .ZN(n4072)
         );
  AOI21_X1 U4624 ( .B1(n5296), .B2(n4341), .A(n4072), .ZN(n4073) );
  OAI21_X1 U4625 ( .B1(n4074), .B2(n5291), .A(n4073), .ZN(U3237) );
  NOR2_X1 U4626 ( .A1(n4139), .A2(n4143), .ZN(n4207) );
  INV_X1 U4627 ( .A(n4075), .ZN(n4078) );
  OAI211_X1 U4628 ( .C1(n4078), .C2(n4673), .A(n4077), .B(n4076), .ZN(n4080)
         );
  NAND3_X1 U4629 ( .A1(n4080), .A2(n4079), .A3(n3026), .ZN(n4083) );
  NAND3_X1 U4630 ( .A1(n4083), .A2(n4082), .A3(n4081), .ZN(n4085) );
  NAND2_X1 U4631 ( .A1(n4085), .A2(n4084), .ZN(n4090) );
  INV_X1 U4632 ( .A(n4086), .ZN(n4088) );
  NAND4_X1 U4633 ( .A1(n4090), .A2(n4089), .A3(n4088), .A4(n4087), .ZN(n4094)
         );
  INV_X1 U4634 ( .A(n4091), .ZN(n4092) );
  NAND3_X1 U4635 ( .A1(n4094), .A2(n4093), .A3(n4092), .ZN(n4099) );
  INV_X1 U4636 ( .A(n4095), .ZN(n4098) );
  INV_X1 U4637 ( .A(n4096), .ZN(n4097) );
  AOI211_X1 U4638 ( .C1(n4099), .C2(n4112), .A(n4098), .B(n4097), .ZN(n4125)
         );
  NAND2_X1 U4639 ( .A1(n4101), .A2(n4100), .ZN(n4122) );
  INV_X1 U4640 ( .A(n4122), .ZN(n4105) );
  NAND2_X1 U4641 ( .A1(n4103), .A2(n4102), .ZN(n4116) );
  INV_X1 U4642 ( .A(n4116), .ZN(n4104) );
  NAND4_X1 U4643 ( .A1(n4105), .A2(n4120), .A3(n4104), .A4(n4106), .ZN(n4124)
         );
  INV_X1 U4644 ( .A(n4106), .ZN(n4108) );
  NOR3_X1 U4645 ( .A1(n4109), .A2(n4108), .A3(n4107), .ZN(n4113) );
  AOI22_X1 U4646 ( .A1(n4113), .A2(n4112), .B1(n4111), .B2(n4110), .ZN(n4117)
         );
  OAI211_X1 U4647 ( .C1(n4117), .C2(n4116), .A(n4115), .B(n4114), .ZN(n4121)
         );
  NAND3_X1 U4648 ( .A1(n4552), .A2(n4191), .A3(n4118), .ZN(n4119) );
  AOI21_X1 U4649 ( .B1(n4121), .B2(n4120), .A(n4119), .ZN(n4123) );
  AND2_X1 U4650 ( .A1(n4122), .A2(n4191), .ZN(n4195) );
  OAI22_X1 U4651 ( .A1(n4125), .A2(n4124), .B1(n4123), .B2(n4195), .ZN(n4126)
         );
  OAI21_X1 U4652 ( .B1(n4198), .B2(n4126), .A(n4197), .ZN(n4127) );
  AOI21_X1 U4653 ( .B1(n4202), .B2(n4127), .A(n4200), .ZN(n4129) );
  OAI21_X1 U4654 ( .B1(n4129), .B2(n4203), .A(n4128), .ZN(n4136) );
  INV_X1 U4655 ( .A(n4130), .ZN(n4140) );
  INV_X1 U4656 ( .A(n4239), .ZN(n4305) );
  INV_X1 U4657 ( .A(n4131), .ZN(n4132) );
  OAI21_X1 U4658 ( .B1(n4305), .B2(n4133), .A(n4132), .ZN(n4214) );
  NOR3_X1 U4659 ( .A1(n4134), .A2(n4140), .A3(n4214), .ZN(n4216) );
  INV_X1 U4660 ( .A(n4216), .ZN(n4135) );
  AOI21_X1 U4661 ( .B1(n4207), .B2(n4136), .A(n4135), .ZN(n4137) );
  INV_X1 U4662 ( .A(n4137), .ZN(n4187) );
  INV_X1 U4663 ( .A(n4138), .ZN(n4185) );
  OR2_X1 U4664 ( .A1(n4140), .A2(n4139), .ZN(n4338) );
  INV_X1 U4665 ( .A(n4338), .ZN(n4339) );
  INV_X1 U4666 ( .A(n4141), .ZN(n4142) );
  NOR2_X1 U4667 ( .A1(n4143), .A2(n4142), .ZN(n4358) );
  INV_X1 U4668 ( .A(n4144), .ZN(n4147) );
  NAND4_X1 U4669 ( .A1(n4147), .A2(n4146), .A3(n4145), .A4(n3023), .ZN(n4153)
         );
  INV_X1 U4670 ( .A(n4536), .ZN(n4151) );
  NAND4_X1 U4671 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4152)
         );
  NOR2_X1 U4672 ( .A1(n4153), .A2(n4152), .ZN(n4175) );
  AND2_X1 U4673 ( .A1(n4459), .A2(n4154), .ZN(n4487) );
  INV_X1 U4674 ( .A(n4541), .ZN(n4551) );
  AND4_X1 U4675 ( .A1(n4156), .A2(n4155), .A3(n4487), .A4(n4551), .ZN(n4173)
         );
  INV_X1 U4676 ( .A(n4157), .ZN(n4160) );
  NAND4_X1 U4677 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4171)
         );
  NAND2_X1 U4678 ( .A1(n2488), .A2(DATAI_30_), .ZN(n4580) );
  NAND2_X1 U4679 ( .A1(n2496), .A2(REG1_REG_31__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U4680 ( .A1(n3353), .A2(REG2_REG_31__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U4681 ( .A1(n3046), .A2(REG0_REG_31__SCAN_IN), .ZN(n4163) );
  NAND3_X1 U4682 ( .A1(n4165), .A2(n4164), .A3(n4163), .ZN(n4572) );
  NAND2_X1 U4683 ( .A1(n2488), .A2(DATAI_31_), .ZN(n4573) );
  NAND2_X1 U4684 ( .A1(n4572), .A2(n4573), .ZN(n4221) );
  OAI21_X1 U4685 ( .B1(n4238), .B2(n4580), .A(n4221), .ZN(n4166) );
  INV_X1 U4686 ( .A(n4166), .ZN(n4211) );
  NAND3_X1 U4687 ( .A1(n4211), .A2(n4168), .A3(n4167), .ZN(n4169) );
  OR2_X1 U4688 ( .A1(n4169), .A2(n4499), .ZN(n4170) );
  NOR2_X1 U4689 ( .A1(n4171), .A2(n4170), .ZN(n4172) );
  NAND4_X1 U4690 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4179)
         );
  AND2_X1 U4691 ( .A1(n4176), .A2(n4415), .ZN(n4437) );
  NAND3_X1 U4692 ( .A1(n4437), .A2(n2550), .A3(n4177), .ZN(n4178) );
  NOR3_X1 U4693 ( .A1(n4179), .A2(n4394), .A3(n4178), .ZN(n4182) );
  OR2_X1 U4694 ( .A1(n4181), .A2(n2560), .ZN(n4397) );
  NAND4_X1 U4695 ( .A1(n4358), .A2(n4376), .A3(n4182), .A4(n4397), .ZN(n4183)
         );
  NOR2_X1 U4696 ( .A1(n4322), .A2(n4183), .ZN(n4184) );
  NAND4_X1 U4697 ( .A1(n4303), .A2(n4185), .A3(n4339), .A4(n4184), .ZN(n4186)
         );
  MUX2_X1 U4698 ( .A(n4187), .B(n4186), .S(n5212), .Z(n4229) );
  INV_X1 U4699 ( .A(n4572), .ZN(n4188) );
  INV_X1 U4700 ( .A(n4573), .ZN(n4570) );
  NAND2_X1 U4701 ( .A1(n4188), .A2(n4570), .ZN(n4190) );
  NAND2_X1 U4702 ( .A1(n4238), .A2(n4580), .ZN(n4189) );
  AND2_X1 U4703 ( .A1(n4190), .A2(n4189), .ZN(n4223) );
  INV_X1 U4704 ( .A(n4223), .ZN(n4228) );
  INV_X1 U4705 ( .A(n4191), .ZN(n4192) );
  NOR3_X1 U4706 ( .A1(n4194), .A2(n4193), .A3(n4192), .ZN(n4196) );
  NOR2_X1 U4707 ( .A1(n4196), .A2(n4195), .ZN(n4199) );
  OAI21_X1 U4708 ( .B1(n4199), .B2(n4198), .A(n4197), .ZN(n4201) );
  AOI21_X1 U4709 ( .B1(n4202), .B2(n4201), .A(n4200), .ZN(n4204) );
  NOR2_X1 U4710 ( .A1(n4204), .A2(n4203), .ZN(n4209) );
  NOR2_X1 U4711 ( .A1(n4206), .A2(n4205), .ZN(n4215) );
  OAI211_X1 U4712 ( .C1(n4209), .C2(n4208), .A(n4207), .B(n4215), .ZN(n4218)
         );
  OR2_X1 U4713 ( .A1(n4239), .A2(n4210), .ZN(n4212) );
  AND2_X1 U4714 ( .A1(n4212), .A2(n4211), .ZN(n4213) );
  INV_X1 U4715 ( .A(n4213), .ZN(n4217) );
  OAI21_X1 U4716 ( .B1(n4215), .B2(n4214), .A(n4213), .ZN(n4222) );
  OAI22_X1 U4717 ( .A1(n4218), .A2(n4217), .B1(n4222), .B2(n4216), .ZN(n4219)
         );
  OAI21_X1 U4718 ( .B1(n4580), .B2(n4572), .A(n4219), .ZN(n4220) );
  OAI211_X1 U4719 ( .C1(n4223), .C2(n4573), .A(n4220), .B(n4673), .ZN(n4226)
         );
  INV_X1 U4720 ( .A(n4221), .ZN(n4224) );
  OAI21_X1 U4721 ( .B1(n4224), .B2(n4223), .A(n4222), .ZN(n4225) );
  MUX2_X1 U4722 ( .A(n4226), .B(n4225), .S(n2923), .Z(n4227) );
  OAI21_X1 U4723 ( .B1(n4229), .B2(n4228), .A(n4227), .ZN(n4230) );
  XNOR2_X1 U4724 ( .A(n4230), .B(n4674), .ZN(n4237) );
  INV_X1 U4725 ( .A(n4231), .ZN(n5188) );
  NAND2_X1 U4726 ( .A1(n4232), .A2(n5188), .ZN(n4233) );
  OAI211_X1 U4727 ( .C1(n4234), .C2(n4236), .A(n4233), .B(B_REG_SCAN_IN), .ZN(
        n4235) );
  OAI21_X1 U4728 ( .B1(n4237), .B2(n4236), .A(n4235), .ZN(U3239) );
  MUX2_X1 U4729 ( .A(DATAO_REG_31__SCAN_IN), .B(n4572), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4730 ( .A(DATAO_REG_30__SCAN_IN), .B(n4238), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4731 ( .A(n4239), .B(DATAO_REG_29__SCAN_IN), .S(n4253), .Z(U3579)
         );
  MUX2_X1 U4732 ( .A(n4341), .B(DATAO_REG_27__SCAN_IN), .S(n4253), .Z(U3577)
         );
  MUX2_X1 U4733 ( .A(DATAO_REG_26__SCAN_IN), .B(n3903), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4734 ( .A(n4344), .B(DATAO_REG_25__SCAN_IN), .S(n4253), .Z(U3575)
         );
  MUX2_X1 U4735 ( .A(n4399), .B(DATAO_REG_24__SCAN_IN), .S(n4253), .Z(U3574)
         );
  MUX2_X1 U4736 ( .A(DATAO_REG_23__SCAN_IN), .B(n4379), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4737 ( .A(DATAO_REG_22__SCAN_IN), .B(n4433), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4738 ( .A(DATAO_REG_21__SCAN_IN), .B(n4419), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4739 ( .A(DATAO_REG_20__SCAN_IN), .B(n4439), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4740 ( .A(DATAO_REG_19__SCAN_IN), .B(n4465), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4741 ( .A(DATAO_REG_18__SCAN_IN), .B(n4524), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4742 ( .A(DATAO_REG_17__SCAN_IN), .B(n4505), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4743 ( .A(DATAO_REG_16__SCAN_IN), .B(n4240), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4744 ( .A(DATAO_REG_15__SCAN_IN), .B(n4241), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4745 ( .A(DATAO_REG_14__SCAN_IN), .B(n5295), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4746 ( .A(DATAO_REG_13__SCAN_IN), .B(n4242), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4747 ( .A(DATAO_REG_12__SCAN_IN), .B(n5283), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4748 ( .A(DATAO_REG_11__SCAN_IN), .B(n4243), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4749 ( .A(DATAO_REG_10__SCAN_IN), .B(n4244), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4750 ( .A(DATAO_REG_9__SCAN_IN), .B(n4245), .S(U4043), .Z(U3559) );
  MUX2_X1 U4751 ( .A(DATAO_REG_8__SCAN_IN), .B(n4246), .S(U4043), .Z(U3558) );
  MUX2_X1 U4752 ( .A(DATAO_REG_7__SCAN_IN), .B(n4247), .S(U4043), .Z(U3557) );
  MUX2_X1 U4753 ( .A(DATAO_REG_6__SCAN_IN), .B(n4248), .S(U4043), .Z(U3556) );
  MUX2_X1 U4754 ( .A(DATAO_REG_5__SCAN_IN), .B(n4249), .S(U4043), .Z(U3555) );
  MUX2_X1 U4755 ( .A(DATAO_REG_4__SCAN_IN), .B(n4250), .S(U4043), .Z(U3554) );
  MUX2_X1 U4756 ( .A(DATAO_REG_3__SCAN_IN), .B(n4251), .S(U4043), .Z(U3553) );
  MUX2_X1 U4757 ( .A(DATAO_REG_2__SCAN_IN), .B(n4252), .S(U4043), .Z(U3552) );
  MUX2_X1 U4758 ( .A(DATAO_REG_1__SCAN_IN), .B(n3002), .S(U4043), .Z(U3551) );
  MUX2_X1 U4759 ( .A(n4254), .B(DATAO_REG_0__SCAN_IN), .S(n4253), .Z(U3550) );
  INV_X1 U4760 ( .A(n4255), .ZN(n4256) );
  AOI21_X1 U4761 ( .B1(n2618), .B2(n4257), .A(n4256), .ZN(n4258) );
  AOI22_X1 U4762 ( .A1(n2795), .A2(n4258), .B1(n5207), .B2(n5075), .ZN(n4264)
         );
  AOI21_X1 U4763 ( .B1(n5196), .B2(ADDR_REG_3__SCAN_IN), .A(n4259), .ZN(n4263)
         );
  OAI211_X1 U4764 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4261), .A(n5177), .B(n4260), 
        .ZN(n4262) );
  NAND3_X1 U4765 ( .A1(n4264), .A2(n4263), .A3(n4262), .ZN(U3243) );
  AOI21_X1 U4766 ( .B1(n4267), .B2(n4266), .A(n4265), .ZN(n4277) );
  INV_X1 U4767 ( .A(n4675), .ZN(n4270) );
  NOR2_X1 U4768 ( .A1(STATE_REG_SCAN_IN), .A2(n4268), .ZN(n5294) );
  AOI21_X1 U4769 ( .B1(n5196), .B2(ADDR_REG_13__SCAN_IN), .A(n5294), .ZN(n4269) );
  OAI21_X1 U4770 ( .B1(n5181), .B2(n4270), .A(n4269), .ZN(n4276) );
  INV_X1 U4771 ( .A(n4271), .ZN(n4272) );
  AOI211_X1 U4772 ( .C1(n4274), .C2(n4273), .A(n5197), .B(n4272), .ZN(n4275)
         );
  AOI211_X1 U4773 ( .C1(n2795), .C2(n4277), .A(n4276), .B(n4275), .ZN(n4278)
         );
  INV_X1 U4774 ( .A(n4278), .ZN(U3253) );
  AOI21_X1 U4775 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(n4289) );
  AOI21_X1 U4776 ( .B1(n5196), .B2(ADDR_REG_14__SCAN_IN), .A(n4282), .ZN(n4283) );
  OAI21_X1 U4777 ( .B1(n5181), .B2(n4284), .A(n4283), .ZN(n4288) );
  AOI211_X1 U4778 ( .C1(n5313), .C2(n4286), .A(n4285), .B(n5200), .ZN(n4287)
         );
  AOI211_X1 U4779 ( .C1(n5177), .C2(n4289), .A(n4288), .B(n4287), .ZN(n4290)
         );
  INV_X1 U4780 ( .A(n4290), .ZN(U3254) );
  OAI21_X1 U4781 ( .B1(n4292), .B2(n4626), .A(n4291), .ZN(n4301) );
  NAND2_X1 U4782 ( .A1(n4294), .A2(n4293), .ZN(n5158) );
  OAI21_X1 U4783 ( .B1(n4294), .B2(n4293), .A(n5158), .ZN(n4295) );
  NAND2_X1 U4784 ( .A1(n4295), .A2(n2795), .ZN(n4298) );
  AOI21_X1 U4785 ( .B1(n5196), .B2(ADDR_REG_16__SCAN_IN), .A(n4296), .ZN(n4297) );
  OAI211_X1 U4786 ( .C1(n5181), .C2(n4299), .A(n4298), .B(n4297), .ZN(n4300)
         );
  AOI21_X1 U4787 ( .B1(n5177), .B2(n4301), .A(n4300), .ZN(n4302) );
  INV_X1 U4788 ( .A(n4302), .ZN(U3256) );
  XNOR2_X1 U4789 ( .A(n4304), .B(n4303), .ZN(n4592) );
  OAI22_X1 U4790 ( .A1(n4305), .A2(n4546), .B1(n4314), .B2(n4581), .ZN(n4311)
         );
  AOI21_X1 U4791 ( .B1(n4308), .B2(n4307), .A(n4306), .ZN(n4309) );
  NOR2_X1 U4792 ( .A1(n4309), .A2(n4554), .ZN(n4310) );
  INV_X1 U4793 ( .A(n4591), .ZN(n4317) );
  INV_X1 U4794 ( .A(n4312), .ZN(n4313) );
  OAI211_X1 U4795 ( .C1(n4328), .C2(n4314), .A(n4313), .B(n5277), .ZN(n4590)
         );
  OAI22_X1 U4796 ( .A1(n4590), .A2(n4674), .B1(n5307), .B2(n4315), .ZN(n4316)
         );
  OAI21_X1 U4797 ( .B1(n4317), .B2(n4316), .A(n4545), .ZN(n4319) );
  NAND2_X1 U4798 ( .A1(n5356), .A2(REG2_REG_28__SCAN_IN), .ZN(n4318) );
  OAI211_X1 U4799 ( .C1(n4592), .C2(n4518), .A(n4319), .B(n4318), .ZN(U3262)
         );
  XNOR2_X1 U4800 ( .A(n4320), .B(n4322), .ZN(n4594) );
  INV_X1 U4801 ( .A(n4594), .ZN(n4336) );
  AOI21_X1 U4802 ( .B1(n4323), .B2(n4322), .A(n4321), .ZN(n4327) );
  OAI22_X1 U4803 ( .A1(n4324), .A2(n4546), .B1(n4330), .B2(n4581), .ZN(n4325)
         );
  AOI21_X1 U4804 ( .B1(n4504), .B2(n3903), .A(n4325), .ZN(n4326) );
  OAI21_X1 U4805 ( .B1(n4327), .B2(n4554), .A(n4326), .ZN(n4593) );
  INV_X1 U4806 ( .A(n4598), .ZN(n4331) );
  INV_X1 U4807 ( .A(n4328), .ZN(n4329) );
  AOI22_X1 U4808 ( .A1(n4332), .A2(n5302), .B1(REG2_REG_27__SCAN_IN), .B2(
        n5356), .ZN(n4333) );
  OAI21_X1 U4809 ( .B1(n4640), .B2(n5309), .A(n4333), .ZN(n4334) );
  AOI21_X1 U4810 ( .B1(n4593), .B2(n4545), .A(n4334), .ZN(n4335) );
  OAI21_X1 U4811 ( .B1(n4336), .B2(n4518), .A(n4335), .ZN(U3263) );
  XOR2_X1 U4812 ( .A(n4338), .B(n4337), .Z(n4601) );
  XNOR2_X1 U4813 ( .A(n4340), .B(n4339), .ZN(n4348) );
  NAND2_X1 U4814 ( .A1(n4341), .A2(n4525), .ZN(n4346) );
  NOR2_X1 U4815 ( .A1(n4581), .A2(n4342), .ZN(n4343) );
  AOI21_X1 U4816 ( .B1(n4344), .B2(n4504), .A(n4343), .ZN(n4345) );
  NAND2_X1 U4817 ( .A1(n4346), .A2(n4345), .ZN(n4347) );
  AOI21_X1 U4818 ( .B1(n4348), .B2(n4501), .A(n4347), .ZN(n4600) );
  AOI22_X1 U4819 ( .A1(n4349), .A2(n5302), .B1(REG2_REG_26__SCAN_IN), .B2(
        n5356), .ZN(n4352) );
  NAND2_X1 U4820 ( .A1(n4350), .A2(n3902), .ZN(n4597) );
  NAND3_X1 U4821 ( .A1(n4598), .A2(n5352), .A3(n4597), .ZN(n4351) );
  OAI211_X1 U4822 ( .C1(n4600), .C2(n5356), .A(n4352), .B(n4351), .ZN(n4353)
         );
  INV_X1 U4823 ( .A(n4353), .ZN(n4354) );
  OAI21_X1 U4824 ( .B1(n4601), .B2(n4518), .A(n4354), .ZN(U3264) );
  XOR2_X1 U4825 ( .A(n4358), .B(n4355), .Z(n4603) );
  INV_X1 U4826 ( .A(n4603), .ZN(n4371) );
  NAND2_X1 U4827 ( .A1(n4357), .A2(n4356), .ZN(n4359) );
  XNOR2_X1 U4828 ( .A(n4359), .B(n4358), .ZN(n4363) );
  AOI22_X1 U4829 ( .A1(n4399), .A2(n4504), .B1(n4360), .B2(n4560), .ZN(n4362)
         );
  NAND2_X1 U4830 ( .A1(n3903), .A2(n4525), .ZN(n4361) );
  OAI211_X1 U4831 ( .C1(n4363), .C2(n4554), .A(n4362), .B(n4361), .ZN(n4602)
         );
  OR2_X1 U4832 ( .A1(n4388), .A2(n4364), .ZN(n4365) );
  NAND2_X1 U4833 ( .A1(n4350), .A2(n4365), .ZN(n4645) );
  INV_X1 U4834 ( .A(n4366), .ZN(n4367) );
  AOI22_X1 U4835 ( .A1(n4367), .A2(n5302), .B1(REG2_REG_25__SCAN_IN), .B2(
        n5356), .ZN(n4368) );
  OAI21_X1 U4836 ( .B1(n4645), .B2(n5309), .A(n4368), .ZN(n4369) );
  AOI21_X1 U4837 ( .B1(n4545), .B2(n4602), .A(n4369), .ZN(n4370) );
  OAI21_X1 U4838 ( .B1(n4371), .B2(n4518), .A(n4370), .ZN(U3265) );
  XNOR2_X1 U4839 ( .A(n4372), .B(n4373), .ZN(n4608) );
  NAND2_X1 U4840 ( .A1(n4375), .A2(n4374), .ZN(n4377) );
  XNOR2_X1 U4841 ( .A(n4377), .B(n4376), .ZN(n4383) );
  AOI22_X1 U4842 ( .A1(n4379), .A2(n4504), .B1(n4378), .B2(n4560), .ZN(n4380)
         );
  OAI21_X1 U4843 ( .B1(n4381), .B2(n4546), .A(n4380), .ZN(n4382) );
  AOI21_X1 U4844 ( .B1(n4383), .B2(n4501), .A(n4382), .ZN(n4607) );
  INV_X1 U4845 ( .A(n4607), .ZN(n4391) );
  INV_X1 U4846 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4384) );
  OAI22_X1 U4847 ( .A1(n4385), .A2(n5307), .B1(n4384), .B2(n4545), .ZN(n4390)
         );
  OAI21_X1 U4848 ( .B1(n4404), .B2(n4386), .A(n5277), .ZN(n4387) );
  OR2_X1 U4849 ( .A1(n4388), .A2(n4387), .ZN(n4606) );
  NOR2_X1 U4850 ( .A1(n4606), .A2(n4512), .ZN(n4389) );
  AOI211_X1 U4851 ( .C1(n4545), .C2(n4391), .A(n4390), .B(n4389), .ZN(n4392)
         );
  OAI21_X1 U4852 ( .B1(n4608), .B2(n4518), .A(n4392), .ZN(U3266) );
  XOR2_X1 U4853 ( .A(n4397), .B(n4393), .Z(n4610) );
  INV_X1 U4854 ( .A(n4610), .ZN(n4411) );
  NAND3_X1 U4855 ( .A1(n4435), .A2(n4437), .A3(n4434), .ZN(n4436) );
  INV_X1 U4856 ( .A(n4394), .ZN(n4414) );
  NAND3_X1 U4857 ( .A1(n4436), .A2(n4414), .A3(n4415), .ZN(n4413) );
  NAND2_X1 U4858 ( .A1(n4413), .A2(n4395), .ZN(n4396) );
  XOR2_X1 U4859 ( .A(n4397), .B(n4396), .Z(n4402) );
  AOI22_X1 U4860 ( .A1(n4433), .A2(n4504), .B1(n4398), .B2(n4560), .ZN(n4401)
         );
  NAND2_X1 U4861 ( .A1(n4399), .A2(n4525), .ZN(n4400) );
  OAI211_X1 U4862 ( .C1(n4402), .C2(n4554), .A(n4401), .B(n4400), .ZN(n4609)
         );
  INV_X1 U4863 ( .A(n4404), .ZN(n4405) );
  OAI21_X1 U4864 ( .B1(n4423), .B2(n4406), .A(n4405), .ZN(n4650) );
  AOI22_X1 U4865 ( .A1(n5356), .A2(REG2_REG_23__SCAN_IN), .B1(n4407), .B2(
        n5302), .ZN(n4408) );
  OAI21_X1 U4866 ( .B1(n4650), .B2(n5309), .A(n4408), .ZN(n4409) );
  AOI21_X1 U4867 ( .B1(n4609), .B2(n4545), .A(n4409), .ZN(n4410) );
  OAI21_X1 U4868 ( .B1(n4411), .B2(n4518), .A(n4410), .ZN(U3267) );
  XNOR2_X1 U4869 ( .A(n4412), .B(n4414), .ZN(n4614) );
  INV_X1 U4870 ( .A(n4614), .ZN(n4431) );
  INV_X1 U4871 ( .A(n4413), .ZN(n4417) );
  AOI21_X1 U4872 ( .B1(n4436), .B2(n4415), .A(n4414), .ZN(n4416) );
  OAI21_X1 U4873 ( .B1(n4417), .B2(n4416), .A(n4501), .ZN(n4421) );
  AOI22_X1 U4874 ( .A1(n4419), .A2(n4504), .B1(n4418), .B2(n4560), .ZN(n4420)
         );
  OAI211_X1 U4875 ( .C1(n4422), .C2(n4546), .A(n4421), .B(n4420), .ZN(n4613)
         );
  INV_X1 U4876 ( .A(n4446), .ZN(n4426) );
  INV_X1 U4877 ( .A(n4423), .ZN(n4424) );
  OAI21_X1 U4878 ( .B1(n4426), .B2(n4425), .A(n4424), .ZN(n4654) );
  AOI22_X1 U4879 ( .A1(n5356), .A2(REG2_REG_22__SCAN_IN), .B1(n4427), .B2(
        n5302), .ZN(n4428) );
  OAI21_X1 U4880 ( .B1(n4654), .B2(n5309), .A(n4428), .ZN(n4429) );
  AOI21_X1 U4881 ( .B1(n4613), .B2(n4545), .A(n4429), .ZN(n4430) );
  OAI21_X1 U4882 ( .B1(n4431), .B2(n4518), .A(n4430), .ZN(U3268) );
  XNOR2_X1 U4883 ( .A(n4432), .B(n4437), .ZN(n4618) );
  INV_X1 U4884 ( .A(n4618), .ZN(n4451) );
  INV_X1 U4885 ( .A(n4433), .ZN(n4442) );
  AND2_X1 U4886 ( .A1(n4435), .A2(n4434), .ZN(n4438) );
  OAI211_X1 U4887 ( .C1(n4438), .C2(n4437), .A(n4501), .B(n4436), .ZN(n4441)
         );
  AOI22_X1 U4888 ( .A1(n4439), .A2(n4504), .B1(n4444), .B2(n4560), .ZN(n4440)
         );
  OAI211_X1 U4889 ( .C1(n4442), .C2(n4546), .A(n4441), .B(n4440), .ZN(n4617)
         );
  NAND2_X1 U4890 ( .A1(n4472), .A2(n4444), .ZN(n4445) );
  NAND2_X1 U4891 ( .A1(n4446), .A2(n4445), .ZN(n4658) );
  AOI22_X1 U4892 ( .A1(n5356), .A2(REG2_REG_21__SCAN_IN), .B1(n4447), .B2(
        n5302), .ZN(n4448) );
  OAI21_X1 U4893 ( .B1(n4658), .B2(n5309), .A(n4448), .ZN(n4449) );
  AOI21_X1 U4894 ( .B1(n4617), .B2(n4545), .A(n4449), .ZN(n4450) );
  OAI21_X1 U4895 ( .B1(n4451), .B2(n4518), .A(n4450), .ZN(U3269) );
  XNOR2_X1 U4896 ( .A(n4452), .B(n2550), .ZN(n4471) );
  INV_X1 U4897 ( .A(n4453), .ZN(n4455) );
  AOI21_X1 U4898 ( .B1(n4520), .B2(n4457), .A(n4456), .ZN(n4500) );
  NAND2_X1 U4899 ( .A1(n4500), .A2(n4458), .ZN(n4479) );
  INV_X1 U4900 ( .A(n4459), .ZN(n4460) );
  AOI21_X1 U4901 ( .B1(n4479), .B2(n4461), .A(n4460), .ZN(n4463) );
  XNOR2_X1 U4902 ( .A(n4463), .B(n4462), .ZN(n4469) );
  AOI22_X1 U4903 ( .A1(n4465), .A2(n4504), .B1(n4464), .B2(n4560), .ZN(n4466)
         );
  OAI21_X1 U4904 ( .B1(n4467), .B2(n4546), .A(n4466), .ZN(n4468) );
  AOI21_X1 U4905 ( .B1(n4469), .B2(n4501), .A(n4468), .ZN(n4470) );
  OAI21_X1 U4906 ( .B1(n4471), .B2(n5272), .A(n4470), .ZN(n4621) );
  MUX2_X1 U4907 ( .A(REG2_REG_20__SCAN_IN), .B(n4621), .S(n4545), .Z(n4477) );
  INV_X1 U4908 ( .A(n4491), .ZN(n4474) );
  OAI21_X1 U4909 ( .B1(n4474), .B2(n4473), .A(n4472), .ZN(n4662) );
  OAI22_X1 U4910 ( .A1(n4662), .A2(n5309), .B1(n4475), .B2(n5307), .ZN(n4476)
         );
  OR2_X1 U4911 ( .A1(n4477), .A2(n4476), .ZN(U3270) );
  NAND2_X1 U4912 ( .A1(n4479), .A2(n4478), .ZN(n4480) );
  XOR2_X1 U4913 ( .A(n4487), .B(n4480), .Z(n4485) );
  AOI22_X1 U4914 ( .A1(n4524), .A2(n4504), .B1(n4560), .B2(n4481), .ZN(n4482)
         );
  OAI21_X1 U4915 ( .B1(n4483), .B2(n4546), .A(n4482), .ZN(n4484) );
  AOI21_X1 U4916 ( .B1(n4485), .B2(n4501), .A(n4484), .ZN(n5336) );
  XOR2_X1 U4917 ( .A(n4487), .B(n4486), .Z(n5341) );
  NAND2_X1 U4918 ( .A1(n5341), .A2(n4568), .ZN(n4496) );
  OR2_X1 U4919 ( .A1(n4488), .A2(n4489), .ZN(n4490) );
  NAND2_X1 U4920 ( .A1(n4491), .A2(n4490), .ZN(n5337) );
  INV_X1 U4921 ( .A(n5337), .ZN(n4494) );
  OAI22_X1 U4922 ( .A1(n4545), .A2(n2755), .B1(n4492), .B2(n5307), .ZN(n4493)
         );
  AOI21_X1 U4923 ( .B1(n4494), .B2(n5352), .A(n4493), .ZN(n4495) );
  OAI211_X1 U4924 ( .C1(n5356), .C2(n5336), .A(n4496), .B(n4495), .ZN(U3271)
         );
  OAI21_X1 U4925 ( .B1(n4498), .B2(n4499), .A(n4497), .ZN(n5332) );
  INV_X1 U4926 ( .A(n5332), .ZN(n4519) );
  XNOR2_X1 U4927 ( .A(n4500), .B(n4499), .ZN(n4502) );
  NAND2_X1 U4928 ( .A1(n4502), .A2(n4501), .ZN(n4507) );
  AOI22_X1 U4929 ( .A1(n4505), .A2(n4504), .B1(n4503), .B2(n4560), .ZN(n4506)
         );
  OAI211_X1 U4930 ( .C1(n4508), .C2(n4546), .A(n4507), .B(n4506), .ZN(n5330)
         );
  NOR2_X1 U4931 ( .A1(n4527), .A2(n4510), .ZN(n4511) );
  OR3_X1 U4932 ( .A1(n4488), .A2(n4511), .A3(n5338), .ZN(n5329) );
  NOR2_X1 U4933 ( .A1(n5329), .A2(n4512), .ZN(n4516) );
  INV_X1 U4934 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4514) );
  OAI22_X1 U4935 ( .A1(n4545), .A2(n4514), .B1(n4513), .B2(n5307), .ZN(n4515)
         );
  AOI211_X1 U4936 ( .C1(n5330), .C2(n4545), .A(n4516), .B(n4515), .ZN(n4517)
         );
  OAI21_X1 U4937 ( .B1(n4519), .B2(n4518), .A(n4517), .ZN(U3272) );
  OAI22_X1 U4938 ( .A1(n4547), .A2(n4548), .B1(n3897), .B2(n4581), .ZN(n4523)
         );
  XNOR2_X1 U4939 ( .A(n4520), .B(n4536), .ZN(n4521) );
  NOR2_X1 U4940 ( .A1(n4521), .A2(n4554), .ZN(n4522) );
  AOI211_X1 U4941 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4522), .ZN(n5320)
         );
  INV_X1 U4942 ( .A(n4526), .ZN(n4529) );
  INV_X1 U4943 ( .A(n4527), .ZN(n4528) );
  OAI21_X1 U4944 ( .B1(n4529), .B2(n3897), .A(n4528), .ZN(n5321) );
  INV_X1 U4945 ( .A(n5321), .ZN(n4534) );
  INV_X1 U4946 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4532) );
  INV_X1 U4947 ( .A(n4530), .ZN(n4531) );
  OAI22_X1 U4948 ( .A1(n4545), .A2(n4532), .B1(n4531), .B2(n5307), .ZN(n4533)
         );
  AOI21_X1 U4949 ( .B1(n4534), .B2(n5352), .A(n4533), .ZN(n4539) );
  OAI21_X1 U4950 ( .B1(n4537), .B2(n4536), .A(n4535), .ZN(n5323) );
  NAND2_X1 U4951 ( .A1(n5323), .A2(n4568), .ZN(n4538) );
  OAI211_X1 U4952 ( .C1(n5320), .C2(n5356), .A(n4539), .B(n4538), .ZN(U3273)
         );
  XNOR2_X1 U4953 ( .A(n4540), .B(n4541), .ZN(n5316) );
  INV_X1 U4954 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4544) );
  INV_X1 U4955 ( .A(n4542), .ZN(n4543) );
  OAI22_X1 U4956 ( .A1(n4545), .A2(n4544), .B1(n4543), .B2(n5307), .ZN(n4567)
         );
  OAI22_X1 U4957 ( .A1(n4549), .A2(n4548), .B1(n4547), .B2(n4546), .ZN(n4558)
         );
  INV_X1 U4958 ( .A(n4550), .ZN(n4556) );
  AOI21_X1 U4959 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(n4555) );
  NOR3_X1 U4960 ( .A1(n4556), .A2(n4555), .A3(n4554), .ZN(n4557) );
  AOI211_X1 U4961 ( .C1(n4560), .C2(n4559), .A(n4558), .B(n4557), .ZN(n4565)
         );
  XNOR2_X1 U4962 ( .A(n4562), .B(n4561), .ZN(n4563) );
  OAI21_X1 U4963 ( .B1(n4563), .B2(n5338), .A(n4565), .ZN(n5315) );
  INV_X1 U4964 ( .A(n5315), .ZN(n4564) );
  AOI211_X1 U4965 ( .C1(n4674), .C2(n4565), .A(n5356), .B(n4564), .ZN(n4566)
         );
  AOI211_X1 U4966 ( .C1(n4568), .C2(n5316), .A(n4567), .B(n4566), .ZN(n4569)
         );
  INV_X1 U4967 ( .A(n4569), .ZN(U3275) );
  INV_X1 U4968 ( .A(n4580), .ZN(n4579) );
  XNOR2_X1 U4969 ( .A(n4577), .B(n4570), .ZN(n5353) );
  INV_X1 U4970 ( .A(n5353), .ZN(n4631) );
  INV_X1 U4971 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U4972 ( .A1(n4572), .A2(n4571), .ZN(n4583) );
  OR2_X1 U4973 ( .A1(n4581), .A2(n4573), .ZN(n4574) );
  AND2_X1 U4974 ( .A1(n4583), .A2(n4574), .ZN(n5355) );
  MUX2_X1 U4975 ( .A(n4575), .B(n5355), .S(n5344), .Z(n4576) );
  OAI21_X1 U4976 ( .B1(n4631), .B2(n4628), .A(n4576), .ZN(U3549) );
  AOI21_X1 U4977 ( .B1(n4579), .B2(n4578), .A(n4577), .ZN(n5349) );
  INV_X1 U4978 ( .A(n5349), .ZN(n4634) );
  INV_X1 U4979 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4584) );
  OR2_X1 U4980 ( .A1(n4581), .A2(n4580), .ZN(n4582) );
  AND2_X1 U4981 ( .A1(n4583), .A2(n4582), .ZN(n5351) );
  MUX2_X1 U4982 ( .A(n4584), .B(n5351), .S(n5344), .Z(n4585) );
  OAI21_X1 U4983 ( .B1(n4634), .B2(n4628), .A(n4585), .ZN(U3548) );
  OAI211_X1 U4984 ( .C1(n4589), .C2(n5272), .A(n4588), .B(n4587), .ZN(n4635)
         );
  MUX2_X1 U4985 ( .A(REG1_REG_29__SCAN_IN), .B(n4635), .S(n5344), .Z(U3547) );
  OAI211_X1 U4986 ( .C1(n4592), .C2(n5272), .A(n4591), .B(n4590), .ZN(n4636)
         );
  MUX2_X1 U4987 ( .A(REG1_REG_28__SCAN_IN), .B(n4636), .S(n5344), .Z(U3546) );
  INV_X1 U4988 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4595) );
  AOI21_X1 U4989 ( .B1(n4594), .B2(n5340), .A(n4593), .ZN(n4637) );
  MUX2_X1 U4990 ( .A(n4595), .B(n4637), .S(n5344), .Z(n4596) );
  OAI21_X1 U4991 ( .B1(n4640), .B2(n4628), .A(n4596), .ZN(U3545) );
  NAND3_X1 U4992 ( .A1(n4598), .A2(n5277), .A3(n4597), .ZN(n4599) );
  OAI211_X1 U4993 ( .C1(n4601), .C2(n5272), .A(n4600), .B(n4599), .ZN(n4641)
         );
  MUX2_X1 U4994 ( .A(REG1_REG_26__SCAN_IN), .B(n4641), .S(n5344), .Z(U3544) );
  INV_X1 U4995 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4604) );
  AOI21_X1 U4996 ( .B1(n4603), .B2(n5340), .A(n4602), .ZN(n4642) );
  MUX2_X1 U4997 ( .A(n4604), .B(n4642), .S(n5344), .Z(n4605) );
  OAI21_X1 U4998 ( .B1(n4628), .B2(n4645), .A(n4605), .ZN(U3543) );
  OAI211_X1 U4999 ( .C1(n4608), .C2(n5272), .A(n4607), .B(n4606), .ZN(n4646)
         );
  MUX2_X1 U5000 ( .A(REG1_REG_24__SCAN_IN), .B(n4646), .S(n5344), .Z(U3542) );
  INV_X1 U5001 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4611) );
  AOI21_X1 U5002 ( .B1(n4610), .B2(n5340), .A(n4609), .ZN(n4647) );
  MUX2_X1 U5003 ( .A(n4611), .B(n4647), .S(n5344), .Z(n4612) );
  OAI21_X1 U5004 ( .B1(n4628), .B2(n4650), .A(n4612), .ZN(U3541) );
  INV_X1 U5005 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4615) );
  AOI21_X1 U5006 ( .B1(n4614), .B2(n5340), .A(n4613), .ZN(n4651) );
  MUX2_X1 U5007 ( .A(n4615), .B(n4651), .S(n5344), .Z(n4616) );
  OAI21_X1 U5008 ( .B1(n4628), .B2(n4654), .A(n4616), .ZN(U3540) );
  INV_X1 U5009 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4619) );
  AOI21_X1 U5010 ( .B1(n4618), .B2(n5340), .A(n4617), .ZN(n4655) );
  MUX2_X1 U5011 ( .A(n4619), .B(n4655), .S(n5344), .Z(n4620) );
  OAI21_X1 U5012 ( .B1(n4628), .B2(n4658), .A(n4620), .ZN(U3539) );
  INV_X1 U5013 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4622) );
  INV_X1 U5014 ( .A(n4621), .ZN(n4659) );
  MUX2_X1 U5015 ( .A(n4622), .B(n4659), .S(n5344), .Z(n4623) );
  OAI21_X1 U5016 ( .B1(n4662), .B2(n4628), .A(n4623), .ZN(U3538) );
  AOI21_X1 U5017 ( .B1(n4625), .B2(n5340), .A(n4624), .ZN(n4663) );
  MUX2_X1 U5018 ( .A(n4626), .B(n4663), .S(n5344), .Z(n4627) );
  OAI21_X1 U5019 ( .B1(n4667), .B2(n4628), .A(n4627), .ZN(U3534) );
  INV_X1 U5020 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4629) );
  MUX2_X1 U5021 ( .A(n4629), .B(n5355), .S(n5348), .Z(n4630) );
  OAI21_X1 U5022 ( .B1(n4631), .B2(n4666), .A(n4630), .ZN(U3517) );
  INV_X1 U5023 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4632) );
  MUX2_X1 U5024 ( .A(n4632), .B(n5351), .S(n5348), .Z(n4633) );
  OAI21_X1 U5025 ( .B1(n4634), .B2(n4666), .A(n4633), .ZN(U3516) );
  MUX2_X1 U5026 ( .A(REG0_REG_29__SCAN_IN), .B(n4635), .S(n5348), .Z(U3515) );
  MUX2_X1 U5027 ( .A(REG0_REG_28__SCAN_IN), .B(n4636), .S(n5348), .Z(U3514) );
  MUX2_X1 U5028 ( .A(n4638), .B(n4637), .S(n5348), .Z(n4639) );
  OAI21_X1 U5029 ( .B1(n4640), .B2(n4666), .A(n4639), .ZN(U3513) );
  MUX2_X1 U5030 ( .A(REG0_REG_26__SCAN_IN), .B(n4641), .S(n5348), .Z(U3512) );
  MUX2_X1 U5031 ( .A(n4643), .B(n4642), .S(n5348), .Z(n4644) );
  OAI21_X1 U5032 ( .B1(n4645), .B2(n4666), .A(n4644), .ZN(U3511) );
  MUX2_X1 U5033 ( .A(REG0_REG_24__SCAN_IN), .B(n4646), .S(n5348), .Z(U3510) );
  MUX2_X1 U5034 ( .A(n4648), .B(n4647), .S(n5348), .Z(n4649) );
  OAI21_X1 U5035 ( .B1(n4650), .B2(n4666), .A(n4649), .ZN(U3509) );
  MUX2_X1 U5036 ( .A(n4652), .B(n4651), .S(n5348), .Z(n4653) );
  OAI21_X1 U5037 ( .B1(n4654), .B2(n4666), .A(n4653), .ZN(U3508) );
  MUX2_X1 U5038 ( .A(n4656), .B(n4655), .S(n5348), .Z(n4657) );
  OAI21_X1 U5039 ( .B1(n4658), .B2(n4666), .A(n4657), .ZN(U3507) );
  MUX2_X1 U5040 ( .A(n4660), .B(n4659), .S(n5348), .Z(n4661) );
  OAI21_X1 U5041 ( .B1(n4662), .B2(n4666), .A(n4661), .ZN(U3506) );
  INV_X1 U5042 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4664) );
  MUX2_X1 U5043 ( .A(n4664), .B(n4663), .S(n5348), .Z(n4665) );
  OAI21_X1 U5044 ( .B1(n4667), .B2(n4666), .A(n4665), .ZN(U3499) );
  NOR3_X1 U5045 ( .A1(n2894), .A2(IR_REG_30__SCAN_IN), .A3(n2663), .ZN(n4668)
         );
  MUX2_X1 U5046 ( .A(DATAI_31_), .B(n4668), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5047 ( .A(n4669), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5048 ( .A(DATAI_27_), .B(n4670), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5049 ( .A(n4671), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  INV_X1 U5050 ( .A(n2870), .ZN(n4672) );
  MUX2_X1 U5051 ( .A(n4672), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5052 ( .A(DATAI_24_), .B(n2871), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5053 ( .A(n4673), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5054 ( .A(n5212), .B(DATAI_20_), .S(U3149), .Z(U3332) );
  MUX2_X1 U5055 ( .A(n4674), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5056 ( .A(DATAI_17_), .B(n5156), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U5057 ( .A(n5150), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5058 ( .A(DATAI_13_), .B(n4675), .S(STATE_REG_SCAN_IN), .Z(U3339)
         );
  MUX2_X1 U5059 ( .A(n4676), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5060 ( .A(n2724), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5061 ( .A(DATAI_9_), .B(n4677), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5062 ( .A(n4678), .B(DATAI_8_), .S(U3149), .Z(n5073) );
  XNOR2_X1 U5063 ( .A(DATAI_30_), .B(keyinput_1), .ZN(n4681) );
  XNOR2_X1 U5064 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n4680) );
  XNOR2_X1 U5065 ( .A(DATAI_31_), .B(keyinput_0), .ZN(n4679) );
  NOR3_X1 U5066 ( .A1(n4681), .A2(n4680), .A3(n4679), .ZN(n4685) );
  XOR2_X1 U5067 ( .A(DATAI_27_), .B(keyinput_4), .Z(n4684) );
  XNOR2_X1 U5068 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n4683) );
  XNOR2_X1 U5069 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n4682) );
  NOR4_X1 U5070 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4688)
         );
  XOR2_X1 U5071 ( .A(DATAI_25_), .B(keyinput_6), .Z(n4687) );
  XNOR2_X1 U5072 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n4686) );
  NOR3_X1 U5073 ( .A1(n4688), .A2(n4687), .A3(n4686), .ZN(n4691) );
  XOR2_X1 U5074 ( .A(DATAI_23_), .B(keyinput_8), .Z(n4690) );
  XOR2_X1 U5075 ( .A(DATAI_22_), .B(keyinput_9), .Z(n4689) );
  NOR3_X1 U5076 ( .A1(n4691), .A2(n4690), .A3(n4689), .ZN(n4694) );
  XOR2_X1 U5077 ( .A(DATAI_21_), .B(keyinput_10), .Z(n4693) );
  XOR2_X1 U5078 ( .A(DATAI_20_), .B(keyinput_11), .Z(n4692) );
  NOR3_X1 U5079 ( .A1(n4694), .A2(n4693), .A3(n4692), .ZN(n4698) );
  XNOR2_X1 U5080 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n4697) );
  XOR2_X1 U5081 ( .A(DATAI_18_), .B(keyinput_13), .Z(n4696) );
  XOR2_X1 U5082 ( .A(DATAI_17_), .B(keyinput_14), .Z(n4695) );
  OAI211_X1 U5083 ( .C1(n4698), .C2(n4697), .A(n4696), .B(n4695), .ZN(n4701)
         );
  XOR2_X1 U5084 ( .A(DATAI_16_), .B(keyinput_15), .Z(n4700) );
  XNOR2_X1 U5085 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n4699) );
  NAND3_X1 U5086 ( .A1(n4701), .A2(n4700), .A3(n4699), .ZN(n4704) );
  XNOR2_X1 U5087 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n4703) );
  XNOR2_X1 U5088 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n4702) );
  NAND3_X1 U5089 ( .A1(n4704), .A2(n4703), .A3(n4702), .ZN(n4707) );
  XOR2_X1 U5090 ( .A(DATAI_12_), .B(keyinput_19), .Z(n4706) );
  XNOR2_X1 U5091 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n4705) );
  NAND3_X1 U5092 ( .A1(n4707), .A2(n4706), .A3(n4705), .ZN(n4710) );
  XNOR2_X1 U5093 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n4709) );
  XNOR2_X1 U5094 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n4708) );
  AOI21_X1 U5095 ( .B1(n4710), .B2(n4709), .A(n4708), .ZN(n4718) );
  XNOR2_X1 U5096 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n4717) );
  XNOR2_X1 U5097 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n4716) );
  XOR2_X1 U5098 ( .A(DATAI_8_), .B(keyinput_23), .Z(n4714) );
  XOR2_X1 U5099 ( .A(DATAI_6_), .B(keyinput_25), .Z(n4713) );
  XNOR2_X1 U5100 ( .A(DATAI_5_), .B(keyinput_26), .ZN(n4712) );
  XNOR2_X1 U5101 ( .A(DATAI_3_), .B(keyinput_28), .ZN(n4711) );
  NAND4_X1 U5102 ( .A1(n4714), .A2(n4713), .A3(n4712), .A4(n4711), .ZN(n4715)
         );
  NOR4_X1 U5103 ( .A1(n4718), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4722)
         );
  XOR2_X1 U5104 ( .A(DATAI_2_), .B(keyinput_29), .Z(n4721) );
  XOR2_X1 U5105 ( .A(DATAI_1_), .B(keyinput_30), .Z(n4720) );
  XNOR2_X1 U5106 ( .A(DATAI_0_), .B(keyinput_31), .ZN(n4719) );
  OAI211_X1 U5107 ( .C1(n4722), .C2(n4721), .A(n4720), .B(n4719), .ZN(n4725)
         );
  XNOR2_X1 U5108 ( .A(STATE_REG_SCAN_IN), .B(keyinput_32), .ZN(n4724) );
  XOR2_X1 U5109 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .Z(n4723) );
  AOI21_X1 U5110 ( .B1(n4725), .B2(n4724), .A(n4723), .ZN(n4728) );
  XNOR2_X1 U5111 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_34), .ZN(n4727) );
  XNOR2_X1 U5112 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_35), .ZN(n4726) );
  NOR3_X1 U5113 ( .A1(n4728), .A2(n4727), .A3(n4726), .ZN(n4731) );
  XNOR2_X1 U5114 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_36), .ZN(n4730) );
  XNOR2_X1 U5115 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_37), .ZN(n4729) );
  NOR3_X1 U5116 ( .A1(n4731), .A2(n4730), .A3(n4729), .ZN(n4737) );
  XNOR2_X1 U5117 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_38), .ZN(n4736) );
  XNOR2_X1 U5118 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_41), .ZN(n4734) );
  XNOR2_X1 U5119 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_40), .ZN(n4733) );
  XNOR2_X1 U5120 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .ZN(n4732) );
  NOR3_X1 U5121 ( .A1(n4734), .A2(n4733), .A3(n4732), .ZN(n4735) );
  OAI21_X1 U5122 ( .B1(n4737), .B2(n4736), .A(n4735), .ZN(n4740) );
  XNOR2_X1 U5123 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n4739) );
  XNOR2_X1 U5124 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_43), .ZN(n4738) );
  AOI21_X1 U5125 ( .B1(n4740), .B2(n4739), .A(n4738), .ZN(n4744) );
  XNOR2_X1 U5126 ( .A(n4741), .B(keyinput_45), .ZN(n4743) );
  XNOR2_X1 U5127 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_44), .ZN(n4742) );
  NOR3_X1 U5128 ( .A1(n4744), .A2(n4743), .A3(n4742), .ZN(n4747) );
  XNOR2_X1 U5129 ( .A(n4935), .B(keyinput_46), .ZN(n4746) );
  XOR2_X1 U5130 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .Z(n4745) );
  NOR3_X1 U5131 ( .A1(n4747), .A2(n4746), .A3(n4745), .ZN(n4750) );
  XNOR2_X1 U5132 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_49), .ZN(n4749) );
  XNOR2_X1 U5133 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_48), .ZN(n4748) );
  NOR3_X1 U5134 ( .A1(n4750), .A2(n4749), .A3(n4748), .ZN(n4754) );
  XOR2_X1 U5135 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .Z(n4753) );
  XNOR2_X1 U5136 ( .A(n4943), .B(keyinput_51), .ZN(n4752) );
  XNOR2_X1 U5137 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .ZN(n4751) );
  NOR4_X1 U5138 ( .A1(n4754), .A2(n4753), .A3(n4752), .A4(n4751), .ZN(n4759)
         );
  XOR2_X1 U5139 ( .A(n5167), .B(keyinput_55), .Z(n4758) );
  XNOR2_X1 U5140 ( .A(n4755), .B(keyinput_53), .ZN(n4757) );
  XNOR2_X1 U5141 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .ZN(n4756) );
  NOR4_X1 U5142 ( .A1(n4759), .A2(n4758), .A3(n4757), .A4(n4756), .ZN(n4762)
         );
  XNOR2_X1 U5143 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .ZN(n4761) );
  XNOR2_X1 U5144 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n4760) );
  OAI21_X1 U5145 ( .B1(n4762), .B2(n4761), .A(n4760), .ZN(n4765) );
  XNOR2_X1 U5146 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_58), .ZN(n4764) );
  XOR2_X1 U5147 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_59), .Z(n4763) );
  AOI21_X1 U5148 ( .B1(n4765), .B2(n4764), .A(n4763), .ZN(n4768) );
  XNOR2_X1 U5149 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4767) );
  XNOR2_X1 U5150 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n4766) );
  OAI21_X1 U5151 ( .B1(n4768), .B2(n4767), .A(n4766), .ZN(n4771) );
  XNOR2_X1 U5152 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n4770) );
  XNOR2_X1 U5153 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n4769) );
  NAND3_X1 U5154 ( .A1(n4771), .A2(n4770), .A3(n4769), .ZN(n4778) );
  XNOR2_X1 U5155 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .ZN(n4777) );
  XNOR2_X1 U5156 ( .A(n4772), .B(keyinput_65), .ZN(n4775) );
  XNOR2_X1 U5157 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_66), .ZN(n4774) );
  XNOR2_X1 U5158 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_67), .ZN(n4773) );
  NAND3_X1 U5159 ( .A1(n4775), .A2(n4774), .A3(n4773), .ZN(n4776) );
  AOI21_X1 U5160 ( .B1(n4778), .B2(n4777), .A(n4776), .ZN(n4781) );
  XOR2_X1 U5161 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_68), .Z(n4780) );
  XNOR2_X1 U5162 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n4779) );
  NOR3_X1 U5163 ( .A1(n4781), .A2(n4780), .A3(n4779), .ZN(n4786) );
  XNOR2_X1 U5164 ( .A(n4782), .B(keyinput_71), .ZN(n4785) );
  XNOR2_X1 U5165 ( .A(n4783), .B(keyinput_70), .ZN(n4784) );
  NOR3_X1 U5166 ( .A1(n4786), .A2(n4785), .A3(n4784), .ZN(n4789) );
  XNOR2_X1 U5167 ( .A(n4981), .B(keyinput_73), .ZN(n4788) );
  XNOR2_X1 U5168 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_72), .ZN(n4787) );
  NOR3_X1 U5169 ( .A1(n4789), .A2(n4788), .A3(n4787), .ZN(n4792) );
  XNOR2_X1 U5170 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_74), .ZN(n4791) );
  XNOR2_X1 U5171 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_75), .ZN(n4790) );
  NOR3_X1 U5172 ( .A1(n4792), .A2(n4791), .A3(n4790), .ZN(n4795) );
  XNOR2_X1 U5173 ( .A(n4989), .B(keyinput_76), .ZN(n4794) );
  XNOR2_X1 U5174 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_77), .ZN(n4793) );
  OAI21_X1 U5175 ( .B1(n4795), .B2(n4794), .A(n4793), .ZN(n4799) );
  XNOR2_X1 U5176 ( .A(n4796), .B(keyinput_79), .ZN(n4798) );
  XNOR2_X1 U5177 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_78), .ZN(n4797) );
  NAND3_X1 U5178 ( .A1(n4799), .A2(n4798), .A3(n4797), .ZN(n4803) );
  XNOR2_X1 U5179 ( .A(n4996), .B(keyinput_80), .ZN(n4802) );
  XOR2_X1 U5180 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_81), .Z(n4801) );
  XNOR2_X1 U5181 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_82), .ZN(n4800) );
  AOI211_X1 U5182 ( .C1(n4803), .C2(n4802), .A(n4801), .B(n4800), .ZN(n4810)
         );
  XNOR2_X1 U5183 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_83), .ZN(n4809) );
  XNOR2_X1 U5184 ( .A(n4804), .B(keyinput_85), .ZN(n4807) );
  XNOR2_X1 U5185 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_84), .ZN(n4806) );
  XNOR2_X1 U5186 ( .A(n2899), .B(keyinput_86), .ZN(n4805) );
  NOR3_X1 U5187 ( .A1(n4807), .A2(n4806), .A3(n4805), .ZN(n4808) );
  OAI21_X1 U5188 ( .B1(n4810), .B2(n4809), .A(n4808), .ZN(n4814) );
  INV_X1 U5189 ( .A(D_REG_2__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U5190 ( .A(n5076), .B(keyinput_89), .ZN(n4813) );
  XOR2_X1 U5191 ( .A(D_REG_0__SCAN_IN), .B(keyinput_87), .Z(n4812) );
  XNOR2_X1 U5192 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .ZN(n4811) );
  NAND4_X1 U5193 ( .A1(n4814), .A2(n4813), .A3(n4812), .A4(n4811), .ZN(n4828)
         );
  OAI22_X1 U5194 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_91), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput_92), .ZN(n4825) );
  INV_X1 U5195 ( .A(keyinput_90), .ZN(n4820) );
  INV_X1 U5196 ( .A(D_REG_3__SCAN_IN), .ZN(n5077) );
  AOI22_X1 U5197 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput_93), .B1(n5077), .B2(
        keyinput_90), .ZN(n4818) );
  AOI22_X1 U5198 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput_95), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput_92), .ZN(n4817) );
  AOI22_X1 U5199 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput_97), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput_94), .ZN(n4816) );
  AOI22_X1 U5200 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_91), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput_96), .ZN(n4815) );
  NAND4_X1 U5201 ( .A1(n4818), .A2(n4817), .A3(n4816), .A4(n4815), .ZN(n4819)
         );
  AOI21_X1 U5202 ( .B1(n4820), .B2(D_REG_3__SCAN_IN), .A(n4819), .ZN(n4821) );
  OAI21_X1 U5203 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput_97), .A(n4821), .ZN(
        n4824) );
  OAI22_X1 U5204 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput_93), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput_95), .ZN(n4823) );
  OAI22_X1 U5205 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput_96), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput_94), .ZN(n4822) );
  NOR4_X1 U5206 ( .A1(n4825), .A2(n4824), .A3(n4823), .A4(n4822), .ZN(n4827)
         );
  XNOR2_X1 U5207 ( .A(D_REG_11__SCAN_IN), .B(keyinput_98), .ZN(n4826) );
  AOI21_X1 U5208 ( .B1(n4828), .B2(n4827), .A(n4826), .ZN(n4831) );
  XNOR2_X1 U5209 ( .A(D_REG_12__SCAN_IN), .B(keyinput_99), .ZN(n4830) );
  XNOR2_X1 U5210 ( .A(D_REG_13__SCAN_IN), .B(keyinput_100), .ZN(n4829) );
  OAI21_X1 U5211 ( .B1(n4831), .B2(n4830), .A(n4829), .ZN(n4835) );
  INV_X1 U5212 ( .A(D_REG_14__SCAN_IN), .ZN(n5083) );
  XNOR2_X1 U5213 ( .A(n5083), .B(keyinput_101), .ZN(n4834) );
  INV_X1 U5214 ( .A(D_REG_15__SCAN_IN), .ZN(n5084) );
  XNOR2_X1 U5215 ( .A(n5084), .B(keyinput_102), .ZN(n4833) );
  XNOR2_X1 U5216 ( .A(D_REG_16__SCAN_IN), .B(keyinput_103), .ZN(n4832) );
  AOI211_X1 U5217 ( .C1(n4835), .C2(n4834), .A(n4833), .B(n4832), .ZN(n4838)
         );
  INV_X1 U5218 ( .A(D_REG_18__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U5219 ( .A(n5087), .B(keyinput_105), .ZN(n4837) );
  XNOR2_X1 U5220 ( .A(D_REG_17__SCAN_IN), .B(keyinput_104), .ZN(n4836) );
  NOR3_X1 U5221 ( .A1(n4838), .A2(n4837), .A3(n4836), .ZN(n4846) );
  XNOR2_X1 U5222 ( .A(D_REG_21__SCAN_IN), .B(keyinput_108), .ZN(n4845) );
  XNOR2_X1 U5223 ( .A(D_REG_22__SCAN_IN), .B(keyinput_109), .ZN(n4844) );
  INV_X1 U5224 ( .A(D_REG_20__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U5225 ( .A(n5089), .B(keyinput_107), .ZN(n4842) );
  XNOR2_X1 U5226 ( .A(D_REG_19__SCAN_IN), .B(keyinput_106), .ZN(n4841) );
  XNOR2_X1 U5227 ( .A(D_REG_24__SCAN_IN), .B(keyinput_111), .ZN(n4840) );
  XNOR2_X1 U5228 ( .A(D_REG_23__SCAN_IN), .B(keyinput_110), .ZN(n4839) );
  NAND4_X1 U5229 ( .A1(n4842), .A2(n4841), .A3(n4840), .A4(n4839), .ZN(n4843)
         );
  NOR4_X1 U5230 ( .A1(n4846), .A2(n4845), .A3(n4844), .A4(n4843), .ZN(n4852)
         );
  INV_X1 U5231 ( .A(D_REG_25__SCAN_IN), .ZN(n5094) );
  XNOR2_X1 U5232 ( .A(n5094), .B(keyinput_112), .ZN(n4851) );
  INV_X1 U5233 ( .A(D_REG_27__SCAN_IN), .ZN(n5096) );
  XNOR2_X1 U5234 ( .A(n5096), .B(keyinput_114), .ZN(n4849) );
  INV_X1 U5235 ( .A(D_REG_26__SCAN_IN), .ZN(n5095) );
  XNOR2_X1 U5236 ( .A(n5095), .B(keyinput_113), .ZN(n4848) );
  INV_X1 U5237 ( .A(D_REG_28__SCAN_IN), .ZN(n5097) );
  XNOR2_X1 U5238 ( .A(n5097), .B(keyinput_115), .ZN(n4847) );
  NOR3_X1 U5239 ( .A1(n4849), .A2(n4848), .A3(n4847), .ZN(n4850) );
  OAI21_X1 U5240 ( .B1(n4852), .B2(n4851), .A(n4850), .ZN(n4855) );
  XNOR2_X1 U5241 ( .A(D_REG_29__SCAN_IN), .B(keyinput_116), .ZN(n4854) );
  XNOR2_X1 U5242 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n4853) );
  AOI21_X1 U5243 ( .B1(n4855), .B2(n4854), .A(n4853), .ZN(n4859) );
  INV_X1 U5244 ( .A(D_REG_31__SCAN_IN), .ZN(n5100) );
  XNOR2_X1 U5245 ( .A(n5100), .B(keyinput_118), .ZN(n4858) );
  XOR2_X1 U5246 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .Z(n4857) );
  XNOR2_X1 U5247 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .ZN(n4856) );
  OAI211_X1 U5248 ( .C1(n4859), .C2(n4858), .A(n4857), .B(n4856), .ZN(n4863)
         );
  XNOR2_X1 U5249 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n4862) );
  XNOR2_X1 U5250 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_123), .ZN(n4861) );
  XNOR2_X1 U5251 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4860) );
  AOI211_X1 U5252 ( .C1(n4863), .C2(n4862), .A(n4861), .B(n4860), .ZN(n4866)
         );
  XOR2_X1 U5253 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .Z(n4865) );
  XNOR2_X1 U5254 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .ZN(n4864) );
  OAI21_X1 U5255 ( .B1(n4866), .B2(n4865), .A(n4864), .ZN(n5071) );
  XNOR2_X1 U5256 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .ZN(n5070) );
  XOR2_X1 U5257 ( .A(DATAI_30_), .B(keyinput_129), .Z(n4869) );
  XOR2_X1 U5258 ( .A(DATAI_29_), .B(keyinput_130), .Z(n4868) );
  XOR2_X1 U5259 ( .A(DATAI_31_), .B(keyinput_128), .Z(n4867) );
  NAND3_X1 U5260 ( .A1(n4869), .A2(n4868), .A3(n4867), .ZN(n4873) );
  XOR2_X1 U5261 ( .A(DATAI_28_), .B(keyinput_131), .Z(n4872) );
  XOR2_X1 U5262 ( .A(DATAI_27_), .B(keyinput_132), .Z(n4871) );
  XNOR2_X1 U5263 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n4870) );
  NAND4_X1 U5264 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), .ZN(n4876)
         );
  XOR2_X1 U5265 ( .A(DATAI_24_), .B(keyinput_135), .Z(n4875) );
  XNOR2_X1 U5266 ( .A(DATAI_25_), .B(keyinput_134), .ZN(n4874) );
  NAND3_X1 U5267 ( .A1(n4876), .A2(n4875), .A3(n4874), .ZN(n4879) );
  XOR2_X1 U5268 ( .A(DATAI_23_), .B(keyinput_136), .Z(n4878) );
  XOR2_X1 U5269 ( .A(DATAI_22_), .B(keyinput_137), .Z(n4877) );
  NAND3_X1 U5270 ( .A1(n4879), .A2(n4878), .A3(n4877), .ZN(n4882) );
  XNOR2_X1 U5271 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4881) );
  XNOR2_X1 U5272 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n4880) );
  NAND3_X1 U5273 ( .A1(n4882), .A2(n4881), .A3(n4880), .ZN(n4886) );
  XOR2_X1 U5274 ( .A(DATAI_19_), .B(keyinput_140), .Z(n4885) );
  XOR2_X1 U5275 ( .A(DATAI_17_), .B(keyinput_142), .Z(n4884) );
  XNOR2_X1 U5276 ( .A(DATAI_18_), .B(keyinput_141), .ZN(n4883) );
  AOI211_X1 U5277 ( .C1(n4886), .C2(n4885), .A(n4884), .B(n4883), .ZN(n4889)
         );
  XOR2_X1 U5278 ( .A(DATAI_16_), .B(keyinput_143), .Z(n4888) );
  XOR2_X1 U5279 ( .A(DATAI_15_), .B(keyinput_144), .Z(n4887) );
  NOR3_X1 U5280 ( .A1(n4889), .A2(n4888), .A3(n4887), .ZN(n4892) );
  XOR2_X1 U5281 ( .A(DATAI_14_), .B(keyinput_145), .Z(n4891) );
  XNOR2_X1 U5282 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n4890) );
  NOR3_X1 U5283 ( .A1(n4892), .A2(n4891), .A3(n4890), .ZN(n4895) );
  XOR2_X1 U5284 ( .A(DATAI_12_), .B(keyinput_147), .Z(n4894) );
  XOR2_X1 U5285 ( .A(DATAI_11_), .B(keyinput_148), .Z(n4893) );
  NOR3_X1 U5286 ( .A1(n4895), .A2(n4894), .A3(n4893), .ZN(n4898) );
  XNOR2_X1 U5287 ( .A(DATAI_10_), .B(keyinput_149), .ZN(n4897) );
  XOR2_X1 U5288 ( .A(DATAI_9_), .B(keyinput_150), .Z(n4896) );
  OAI21_X1 U5289 ( .B1(n4898), .B2(n4897), .A(n4896), .ZN(n4906) );
  XOR2_X1 U5290 ( .A(DATAI_8_), .B(keyinput_151), .Z(n4905) );
  XOR2_X1 U5291 ( .A(DATAI_7_), .B(keyinput_152), .Z(n4904) );
  XOR2_X1 U5292 ( .A(DATAI_6_), .B(keyinput_153), .Z(n4902) );
  XOR2_X1 U5293 ( .A(DATAI_5_), .B(keyinput_154), .Z(n4901) );
  XNOR2_X1 U5294 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n4900) );
  XNOR2_X1 U5295 ( .A(DATAI_3_), .B(keyinput_156), .ZN(n4899) );
  NOR4_X1 U5296 ( .A1(n4902), .A2(n4901), .A3(n4900), .A4(n4899), .ZN(n4903)
         );
  NAND4_X1 U5297 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4910)
         );
  XNOR2_X1 U5298 ( .A(DATAI_2_), .B(keyinput_157), .ZN(n4909) );
  XNOR2_X1 U5299 ( .A(DATAI_1_), .B(keyinput_158), .ZN(n4908) );
  XNOR2_X1 U5300 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n4907) );
  AOI211_X1 U5301 ( .C1(n4910), .C2(n4909), .A(n4908), .B(n4907), .ZN(n4913)
         );
  XNOR2_X1 U5302 ( .A(STATE_REG_SCAN_IN), .B(keyinput_160), .ZN(n4912) );
  XOR2_X1 U5303 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .Z(n4911) );
  OAI21_X1 U5304 ( .B1(n4913), .B2(n4912), .A(n4911), .ZN(n4917) );
  XNOR2_X1 U5305 ( .A(n4914), .B(keyinput_162), .ZN(n4916) );
  XNOR2_X1 U5306 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_163), .ZN(n4915) );
  NAND3_X1 U5307 ( .A1(n4917), .A2(n4916), .A3(n4915), .ZN(n4920) );
  XOR2_X1 U5308 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .Z(n4919) );
  XNOR2_X1 U5309 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_164), .ZN(n4918) );
  NAND3_X1 U5310 ( .A1(n4920), .A2(n4919), .A3(n4918), .ZN(n4927) );
  XNOR2_X1 U5311 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_166), .ZN(n4926) );
  XNOR2_X1 U5312 ( .A(n4921), .B(keyinput_169), .ZN(n4924) );
  XNOR2_X1 U5313 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_167), .ZN(n4923) );
  XNOR2_X1 U5314 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_168), .ZN(n4922) );
  NAND3_X1 U5315 ( .A1(n4924), .A2(n4923), .A3(n4922), .ZN(n4925) );
  AOI21_X1 U5316 ( .B1(n4927), .B2(n4926), .A(n4925), .ZN(n4931) );
  XOR2_X1 U5317 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .Z(n4930) );
  XNOR2_X1 U5318 ( .A(n4928), .B(keyinput_171), .ZN(n4929) );
  OAI21_X1 U5319 ( .B1(n4931), .B2(n4930), .A(n4929), .ZN(n4934) );
  XNOR2_X1 U5320 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_173), .ZN(n4933) );
  XNOR2_X1 U5321 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_172), .ZN(n4932) );
  NAND3_X1 U5322 ( .A1(n4934), .A2(n4933), .A3(n4932), .ZN(n4938) );
  XNOR2_X1 U5323 ( .A(n4935), .B(keyinput_174), .ZN(n4937) );
  XOR2_X1 U5324 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_175), .Z(n4936) );
  NAND3_X1 U5325 ( .A1(n4938), .A2(n4937), .A3(n4936), .ZN(n4942) );
  XOR2_X1 U5326 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_176), .Z(n4941) );
  XNOR2_X1 U5327 ( .A(n4939), .B(keyinput_177), .ZN(n4940) );
  NAND3_X1 U5328 ( .A1(n4942), .A2(n4941), .A3(n4940), .ZN(n4947) );
  XNOR2_X1 U5329 ( .A(n4943), .B(keyinput_179), .ZN(n4946) );
  XNOR2_X1 U5330 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n4945) );
  XNOR2_X1 U5331 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .ZN(n4944) );
  NAND4_X1 U5332 ( .A1(n4947), .A2(n4946), .A3(n4945), .A4(n4944), .ZN(n4951)
         );
  XOR2_X1 U5333 ( .A(n5167), .B(keyinput_183), .Z(n4950) );
  XNOR2_X1 U5334 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .ZN(n4949) );
  XNOR2_X1 U5335 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_182), .ZN(n4948) );
  NAND4_X1 U5336 ( .A1(n4951), .A2(n4950), .A3(n4949), .A4(n4948), .ZN(n4955)
         );
  XNOR2_X1 U5337 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .ZN(n4954) );
  XNOR2_X1 U5338 ( .A(n4952), .B(keyinput_185), .ZN(n4953) );
  AOI21_X1 U5339 ( .B1(n4955), .B2(n4954), .A(n4953), .ZN(n4958) );
  XNOR2_X1 U5340 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_186), .ZN(n4957) );
  XNOR2_X1 U5341 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_187), .ZN(n4956) );
  OAI21_X1 U5342 ( .B1(n4958), .B2(n4957), .A(n4956), .ZN(n4962) );
  XNOR2_X1 U5343 ( .A(n4959), .B(keyinput_188), .ZN(n4961) );
  XNOR2_X1 U5344 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n4960) );
  AOI21_X1 U5345 ( .B1(n4962), .B2(n4961), .A(n4960), .ZN(n4966) );
  XNOR2_X1 U5346 ( .A(n4963), .B(keyinput_191), .ZN(n4965) );
  XNOR2_X1 U5347 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_190), .ZN(n4964) );
  NOR3_X1 U5348 ( .A1(n4966), .A2(n4965), .A3(n4964), .ZN(n4973) );
  XNOR2_X1 U5349 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_192), .ZN(n4972) );
  XNOR2_X1 U5350 ( .A(n4967), .B(keyinput_194), .ZN(n4970) );
  XNOR2_X1 U5351 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_195), .ZN(n4969) );
  XNOR2_X1 U5352 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_193), .ZN(n4968) );
  NOR3_X1 U5353 ( .A1(n4970), .A2(n4969), .A3(n4968), .ZN(n4971) );
  OAI21_X1 U5354 ( .B1(n4973), .B2(n4972), .A(n4971), .ZN(n4976) );
  XOR2_X1 U5355 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_197), .Z(n4975) );
  XOR2_X1 U5356 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_196), .Z(n4974) );
  NAND3_X1 U5357 ( .A1(n4976), .A2(n4975), .A3(n4974), .ZN(n4979) );
  XNOR2_X1 U5358 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n4978) );
  XNOR2_X1 U5359 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_199), .ZN(n4977) );
  NAND3_X1 U5360 ( .A1(n4979), .A2(n4978), .A3(n4977), .ZN(n4984) );
  XNOR2_X1 U5361 ( .A(n4980), .B(keyinput_200), .ZN(n4983) );
  XNOR2_X1 U5362 ( .A(n4981), .B(keyinput_201), .ZN(n4982) );
  NAND3_X1 U5363 ( .A1(n4984), .A2(n4983), .A3(n4982), .ZN(n4988) );
  XNOR2_X1 U5364 ( .A(n4985), .B(keyinput_203), .ZN(n4987) );
  XNOR2_X1 U5365 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_202), .ZN(n4986) );
  NAND3_X1 U5366 ( .A1(n4988), .A2(n4987), .A3(n4986), .ZN(n4992) );
  XNOR2_X1 U5367 ( .A(n4989), .B(keyinput_204), .ZN(n4991) );
  XNOR2_X1 U5368 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_205), .ZN(n4990) );
  AOI21_X1 U5369 ( .B1(n4992), .B2(n4991), .A(n4990), .ZN(n4995) );
  XNOR2_X1 U5370 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_207), .ZN(n4994) );
  XNOR2_X1 U5371 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_206), .ZN(n4993) );
  NOR3_X1 U5372 ( .A1(n4995), .A2(n4994), .A3(n4993), .ZN(n5000) );
  XNOR2_X1 U5373 ( .A(n4996), .B(keyinput_208), .ZN(n4999) );
  XOR2_X1 U5374 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_209), .Z(n4998) );
  XNOR2_X1 U5375 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_210), .ZN(n4997) );
  OAI211_X1 U5376 ( .C1(n5000), .C2(n4999), .A(n4998), .B(n4997), .ZN(n5007)
         );
  XNOR2_X1 U5377 ( .A(n5001), .B(keyinput_211), .ZN(n5006) );
  XNOR2_X1 U5378 ( .A(n2899), .B(keyinput_214), .ZN(n5005) );
  XNOR2_X1 U5379 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_212), .ZN(n5003) );
  XNOR2_X1 U5380 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n5002) );
  NAND2_X1 U5381 ( .A1(n5003), .A2(n5002), .ZN(n5004) );
  AOI211_X1 U5382 ( .C1(n5007), .C2(n5006), .A(n5005), .B(n5004), .ZN(n5011)
         );
  XNOR2_X1 U5383 ( .A(n5076), .B(keyinput_217), .ZN(n5010) );
  XOR2_X1 U5384 ( .A(D_REG_0__SCAN_IN), .B(keyinput_215), .Z(n5009) );
  XNOR2_X1 U5385 ( .A(D_REG_1__SCAN_IN), .B(keyinput_216), .ZN(n5008) );
  INV_X1 U5386 ( .A(D_REG_10__SCAN_IN), .ZN(n5080) );
  INV_X1 U5387 ( .A(D_REG_7__SCAN_IN), .ZN(n5018) );
  INV_X1 U5388 ( .A(keyinput_222), .ZN(n5017) );
  INV_X1 U5389 ( .A(D_REG_8__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U5390 ( .A1(n5079), .A2(keyinput_223), .B1(n5077), .B2(keyinput_218), .ZN(n5015) );
  INV_X1 U5391 ( .A(D_REG_5__SCAN_IN), .ZN(n5078) );
  AOI22_X1 U5392 ( .A1(n5080), .A2(keyinput_225), .B1(n5078), .B2(keyinput_220), .ZN(n5014) );
  AOI22_X1 U5393 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput_224), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput_222), .ZN(n5013) );
  AOI22_X1 U5394 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_219), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput_221), .ZN(n5012) );
  NAND4_X1 U5395 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(n5016)
         );
  AOI21_X1 U5396 ( .B1(n5018), .B2(n5017), .A(n5016), .ZN(n5019) );
  OAI21_X1 U5397 ( .B1(keyinput_225), .B2(n5080), .A(n5019), .ZN(n5023) );
  OAI22_X1 U5398 ( .A1(keyinput_218), .A2(n5077), .B1(n5078), .B2(keyinput_220), .ZN(n5022) );
  OAI22_X1 U5399 ( .A1(n5079), .A2(keyinput_223), .B1(D_REG_6__SCAN_IN), .B2(
        keyinput_221), .ZN(n5021) );
  OAI22_X1 U5400 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_219), .B1(
        D_REG_9__SCAN_IN), .B2(keyinput_224), .ZN(n5020) );
  NOR4_X1 U5401 ( .A1(n5023), .A2(n5022), .A3(n5021), .A4(n5020), .ZN(n5025)
         );
  XNOR2_X1 U5402 ( .A(D_REG_11__SCAN_IN), .B(keyinput_226), .ZN(n5024) );
  AOI21_X1 U5403 ( .B1(n5026), .B2(n5025), .A(n5024), .ZN(n5029) );
  XNOR2_X1 U5404 ( .A(D_REG_12__SCAN_IN), .B(keyinput_227), .ZN(n5028) );
  INV_X1 U5405 ( .A(D_REG_13__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U5406 ( .A(n5082), .B(keyinput_228), .ZN(n5027) );
  OAI21_X1 U5407 ( .B1(n5029), .B2(n5028), .A(n5027), .ZN(n5033) );
  XNOR2_X1 U5408 ( .A(n5083), .B(keyinput_229), .ZN(n5032) );
  INV_X1 U5409 ( .A(D_REG_16__SCAN_IN), .ZN(n5085) );
  XNOR2_X1 U5410 ( .A(n5085), .B(keyinput_231), .ZN(n5031) );
  XNOR2_X1 U5411 ( .A(D_REG_15__SCAN_IN), .B(keyinput_230), .ZN(n5030) );
  AOI211_X1 U5412 ( .C1(n5033), .C2(n5032), .A(n5031), .B(n5030), .ZN(n5036)
         );
  INV_X1 U5413 ( .A(D_REG_17__SCAN_IN), .ZN(n5086) );
  XNOR2_X1 U5414 ( .A(n5086), .B(keyinput_232), .ZN(n5035) );
  XNOR2_X1 U5415 ( .A(D_REG_18__SCAN_IN), .B(keyinput_233), .ZN(n5034) );
  NOR3_X1 U5416 ( .A1(n5036), .A2(n5035), .A3(n5034), .ZN(n5044) );
  XNOR2_X1 U5417 ( .A(D_REG_19__SCAN_IN), .B(keyinput_234), .ZN(n5043) );
  XNOR2_X1 U5418 ( .A(D_REG_22__SCAN_IN), .B(keyinput_237), .ZN(n5042) );
  INV_X1 U5419 ( .A(D_REG_23__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U5420 ( .A(n5092), .B(keyinput_238), .ZN(n5040) );
  XNOR2_X1 U5421 ( .A(D_REG_20__SCAN_IN), .B(keyinput_235), .ZN(n5039) );
  XNOR2_X1 U5422 ( .A(D_REG_24__SCAN_IN), .B(keyinput_239), .ZN(n5038) );
  XNOR2_X1 U5423 ( .A(D_REG_21__SCAN_IN), .B(keyinput_236), .ZN(n5037) );
  NAND4_X1 U5424 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), .ZN(n5041)
         );
  NOR4_X1 U5425 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n5050)
         );
  XNOR2_X1 U5426 ( .A(n5094), .B(keyinput_240), .ZN(n5049) );
  XNOR2_X1 U5427 ( .A(n5096), .B(keyinput_242), .ZN(n5047) );
  XNOR2_X1 U5428 ( .A(D_REG_26__SCAN_IN), .B(keyinput_241), .ZN(n5046) );
  XNOR2_X1 U5429 ( .A(D_REG_28__SCAN_IN), .B(keyinput_243), .ZN(n5045) );
  NOR3_X1 U5430 ( .A1(n5047), .A2(n5046), .A3(n5045), .ZN(n5048) );
  OAI21_X1 U5431 ( .B1(n5050), .B2(n5049), .A(n5048), .ZN(n5053) );
  XNOR2_X1 U5432 ( .A(D_REG_29__SCAN_IN), .B(keyinput_244), .ZN(n5052) );
  INV_X1 U5433 ( .A(D_REG_30__SCAN_IN), .ZN(n5099) );
  XNOR2_X1 U5434 ( .A(n5099), .B(keyinput_245), .ZN(n5051) );
  AOI21_X1 U5435 ( .B1(n5053), .B2(n5052), .A(n5051), .ZN(n5057) );
  XNOR2_X1 U5436 ( .A(n5100), .B(keyinput_246), .ZN(n5056) );
  XOR2_X1 U5437 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .Z(n5055) );
  XNOR2_X1 U5438 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .ZN(n5054) );
  OAI211_X1 U5439 ( .C1(n5057), .C2(n5056), .A(n5055), .B(n5054), .ZN(n5061)
         );
  XOR2_X1 U5440 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .Z(n5060) );
  XOR2_X1 U5441 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .Z(n5059) );
  XNOR2_X1 U5442 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_250), .ZN(n5058) );
  AOI211_X1 U5443 ( .C1(n5061), .C2(n5060), .A(n5059), .B(n5058), .ZN(n5064)
         );
  XOR2_X1 U5444 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .Z(n5063) );
  XNOR2_X1 U5445 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .ZN(n5062) );
  OAI21_X1 U5446 ( .B1(n5064), .B2(n5063), .A(n5062), .ZN(n5067) );
  XNOR2_X1 U5447 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .ZN(n5066) );
  XNOR2_X1 U5448 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_255), .ZN(n5065) );
  AOI21_X1 U5449 ( .B1(n5067), .B2(n5066), .A(n5065), .ZN(n5069) );
  XNOR2_X1 U5450 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .ZN(n5068) );
  AOI211_X1 U5451 ( .C1(n5071), .C2(n5070), .A(n5069), .B(n5068), .ZN(n5072)
         );
  XOR2_X1 U5452 ( .A(n5073), .B(n5072), .Z(U3344) );
  MUX2_X1 U5453 ( .A(n5137), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5454 ( .A(n5074), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5455 ( .A(n5126), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5456 ( .A(n5206), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U5457 ( .A(n5075), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5458 ( .A(n2800), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  NOR2_X1 U5459 ( .A1(n5101), .A2(n5076), .ZN(U3320) );
  NOR2_X1 U5460 ( .A1(n5101), .A2(n5077), .ZN(U3319) );
  AND2_X1 U5461 ( .A1(n5091), .A2(D_REG_4__SCAN_IN), .ZN(U3318) );
  NOR2_X1 U5462 ( .A1(n5101), .A2(n5078), .ZN(U3317) );
  AND2_X1 U5463 ( .A1(n5091), .A2(D_REG_6__SCAN_IN), .ZN(U3316) );
  AND2_X1 U5464 ( .A1(n5091), .A2(D_REG_7__SCAN_IN), .ZN(U3315) );
  NOR2_X1 U5465 ( .A1(n5101), .A2(n5079), .ZN(U3314) );
  AND2_X1 U5466 ( .A1(n5091), .A2(D_REG_9__SCAN_IN), .ZN(U3313) );
  NOR2_X1 U5467 ( .A1(n5101), .A2(n5080), .ZN(U3312) );
  AND2_X1 U5468 ( .A1(n5091), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  INV_X1 U5469 ( .A(D_REG_12__SCAN_IN), .ZN(n5081) );
  NOR2_X1 U5470 ( .A1(n5101), .A2(n5081), .ZN(U3310) );
  NOR2_X1 U5471 ( .A1(n5101), .A2(n5082), .ZN(U3309) );
  NOR2_X1 U5472 ( .A1(n5101), .A2(n5083), .ZN(U3308) );
  NOR2_X1 U5473 ( .A1(n5101), .A2(n5084), .ZN(U3307) );
  NOR2_X1 U5474 ( .A1(n5101), .A2(n5085), .ZN(U3306) );
  NOR2_X1 U5475 ( .A1(n5101), .A2(n5086), .ZN(U3305) );
  NOR2_X1 U5476 ( .A1(n5101), .A2(n5087), .ZN(U3304) );
  INV_X1 U5477 ( .A(D_REG_19__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U5478 ( .A1(n5101), .A2(n5088), .ZN(U3303) );
  NOR2_X1 U5479 ( .A1(n5101), .A2(n5089), .ZN(U3302) );
  INV_X1 U5480 ( .A(D_REG_21__SCAN_IN), .ZN(n5090) );
  NOR2_X1 U5481 ( .A1(n5101), .A2(n5090), .ZN(U3301) );
  AND2_X1 U5482 ( .A1(n5091), .A2(D_REG_22__SCAN_IN), .ZN(U3300) );
  NOR2_X1 U5483 ( .A1(n5101), .A2(n5092), .ZN(U3299) );
  INV_X1 U5484 ( .A(D_REG_24__SCAN_IN), .ZN(n5093) );
  NOR2_X1 U5485 ( .A1(n5101), .A2(n5093), .ZN(U3298) );
  NOR2_X1 U5486 ( .A1(n5101), .A2(n5094), .ZN(U3297) );
  NOR2_X1 U5487 ( .A1(n5101), .A2(n5095), .ZN(U3296) );
  NOR2_X1 U5488 ( .A1(n5101), .A2(n5096), .ZN(U3295) );
  NOR2_X1 U5489 ( .A1(n5101), .A2(n5097), .ZN(U3294) );
  INV_X1 U5490 ( .A(D_REG_29__SCAN_IN), .ZN(n5098) );
  NOR2_X1 U5491 ( .A1(n5101), .A2(n5098), .ZN(U3293) );
  NOR2_X1 U5492 ( .A1(n5101), .A2(n5099), .ZN(U3292) );
  NOR2_X1 U5493 ( .A1(n5101), .A2(n5100), .ZN(U3291) );
  OAI21_X1 U5494 ( .B1(REG2_REG_0__SCAN_IN), .B2(n5183), .A(n5184), .ZN(n5189)
         );
  AOI21_X1 U5495 ( .B1(n5183), .B2(n5102), .A(n5189), .ZN(n5103) );
  XNOR2_X1 U5496 ( .A(n5103), .B(n5167), .ZN(n5105) );
  AOI22_X1 U5497 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n5196), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n5104) );
  OAI21_X1 U5498 ( .B1(n5106), .B2(n5105), .A(n5104), .ZN(U3240) );
  AOI22_X1 U5499 ( .A1(ADDR_REG_1__SCAN_IN), .A2(n5196), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n5118) );
  AOI21_X1 U5500 ( .B1(n5108), .B2(n5186), .A(n5107), .ZN(n5109) );
  NAND2_X1 U5501 ( .A1(n2795), .A2(n5109), .ZN(n5115) );
  AOI21_X1 U5502 ( .B1(n5112), .B2(n5111), .A(n5110), .ZN(n5113) );
  NAND2_X1 U5503 ( .A1(n5177), .A2(n5113), .ZN(n5114) );
  OAI211_X1 U5504 ( .C1(n5181), .C2(n2675), .A(n5115), .B(n5114), .ZN(n5116)
         );
  INV_X1 U5505 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U5506 ( .A1(n5118), .A2(n5117), .ZN(U3241) );
  AOI211_X1 U5507 ( .C1(n2524), .C2(n5120), .A(n5119), .B(n5200), .ZN(n5122)
         );
  AOI211_X1 U5508 ( .C1(n5196), .C2(ADDR_REG_5__SCAN_IN), .A(n5122), .B(n5121), 
        .ZN(n5128) );
  AOI211_X1 U5509 ( .C1(n2525), .C2(n5124), .A(n5123), .B(n5197), .ZN(n5125)
         );
  AOI21_X1 U5510 ( .B1(n5207), .B2(n5126), .A(n5125), .ZN(n5127) );
  NAND2_X1 U5511 ( .A1(n5128), .A2(n5127), .ZN(U3245) );
  INV_X1 U5512 ( .A(n5129), .ZN(n5130) );
  AOI211_X1 U5513 ( .C1(n5132), .C2(n5131), .A(n5130), .B(n5200), .ZN(n5134)
         );
  AOI211_X1 U5514 ( .C1(n5196), .C2(ADDR_REG_7__SCAN_IN), .A(n5134), .B(n5133), 
        .ZN(n5141) );
  AOI21_X1 U5515 ( .B1(n5136), .B2(n5135), .A(n5197), .ZN(n5139) );
  AOI22_X1 U5516 ( .A1(n5139), .A2(n5138), .B1(n5137), .B2(n5207), .ZN(n5140)
         );
  NAND2_X1 U5517 ( .A1(n5141), .A2(n5140), .ZN(U3247) );
  AOI211_X1 U5518 ( .C1(n2509), .C2(n5143), .A(n5142), .B(n5197), .ZN(n5145)
         );
  AOI211_X1 U5519 ( .C1(n5196), .C2(ADDR_REG_15__SCAN_IN), .A(n5145), .B(n5144), .ZN(n5152) );
  AOI211_X1 U5520 ( .C1(n5148), .C2(n5147), .A(n5146), .B(n5200), .ZN(n5149)
         );
  AOI21_X1 U5521 ( .B1(n5207), .B2(n5150), .A(n5149), .ZN(n5151) );
  NAND2_X1 U5522 ( .A1(n5152), .A2(n5151), .ZN(U3255) );
  OAI21_X1 U5523 ( .B1(n5155), .B2(n5154), .A(n5153), .ZN(n5157) );
  AOI22_X1 U5524 ( .A1(n5157), .A2(n5177), .B1(n5156), .B2(n5207), .ZN(n5166)
         );
  NAND2_X1 U5525 ( .A1(n5159), .A2(n5158), .ZN(n5161) );
  AOI211_X1 U5526 ( .C1(n5162), .C2(n5161), .A(n5160), .B(n5200), .ZN(n5164)
         );
  AOI211_X1 U5527 ( .C1(n5196), .C2(ADDR_REG_17__SCAN_IN), .A(n5164), .B(n5163), .ZN(n5165) );
  NAND2_X1 U5528 ( .A1(n5166), .A2(n5165), .ZN(U3257) );
  INV_X1 U5529 ( .A(n5167), .ZN(n5190) );
  INV_X1 U5530 ( .A(DATAI_0_), .ZN(n5168) );
  AOI22_X1 U5531 ( .A1(STATE_REG_SCAN_IN), .A2(n5190), .B1(n5168), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5532 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n5196), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n5194) );
  AOI21_X1 U5533 ( .B1(n5171), .B2(n5170), .A(n5169), .ZN(n5172) );
  NAND2_X1 U5534 ( .A1(n2795), .A2(n5172), .ZN(n5179) );
  AOI21_X1 U5535 ( .B1(n5175), .B2(n5173), .A(n5174), .ZN(n5176) );
  NAND2_X1 U5536 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  OAI211_X1 U5537 ( .C1(n5181), .C2(n5180), .A(n5179), .B(n5178), .ZN(n5182)
         );
  INV_X1 U5538 ( .A(n5182), .ZN(n5193) );
  NAND3_X1 U5539 ( .A1(n5185), .A2(n5184), .A3(n5183), .ZN(n5192) );
  INV_X1 U5540 ( .A(n5186), .ZN(n5187) );
  AOI22_X1 U5541 ( .A1(n5190), .A2(n5189), .B1(n5188), .B2(n5187), .ZN(n5191)
         );
  NAND3_X1 U5542 ( .A1(n5192), .A2(U4043), .A3(n5191), .ZN(n5208) );
  NAND3_X1 U5543 ( .A1(n5194), .A2(n5193), .A3(n5208), .ZN(U3242) );
  AOI21_X1 U5544 ( .B1(n5196), .B2(ADDR_REG_4__SCAN_IN), .A(n5195), .ZN(n5210)
         );
  AOI211_X1 U5545 ( .C1(n5236), .C2(n5199), .A(n5198), .B(n5197), .ZN(n5205)
         );
  AOI211_X1 U5546 ( .C1(n5203), .C2(n5202), .A(n5201), .B(n5200), .ZN(n5204)
         );
  AOI211_X1 U5547 ( .C1(n5207), .C2(n5206), .A(n5205), .B(n5204), .ZN(n5209)
         );
  NAND3_X1 U5548 ( .A1(n5210), .A2(n5209), .A3(n5208), .ZN(U3244) );
  INV_X1 U5549 ( .A(REG3_REG_0__SCAN_IN), .ZN(n5218) );
  NOR3_X1 U5550 ( .A1(n5213), .A2(n5212), .A3(n5211), .ZN(n5214) );
  NOR2_X1 U5551 ( .A1(n5215), .A2(n5214), .ZN(n5216) );
  AOI22_X1 U5552 ( .A1(n5356), .A2(REG2_REG_0__SCAN_IN), .B1(n5216), .B2(n4545), .ZN(n5217) );
  OAI21_X1 U5553 ( .B1(n5218), .B2(n5307), .A(n5217), .ZN(U3290) );
  OAI22_X1 U5554 ( .A1(U3149), .A2(n5219), .B1(DATAI_1_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5220) );
  INV_X1 U5555 ( .A(n5220), .ZN(U3351) );
  AOI22_X1 U5556 ( .A1(n5352), .A2(n5221), .B1(REG3_REG_1__SCAN_IN), .B2(n5302), .ZN(n5222) );
  OAI221_X1 U5557 ( .B1(n5356), .B2(n5224), .C1(n4545), .C2(n5223), .A(n5222), 
        .ZN(U3289) );
  AOI22_X1 U5558 ( .A1(n5352), .A2(n5225), .B1(REG3_REG_2__SCAN_IN), .B2(n5302), .ZN(n5226) );
  OAI221_X1 U5559 ( .B1(n5356), .B2(n5228), .C1(n4545), .C2(n5227), .A(n5226), 
        .ZN(U3288) );
  AOI22_X1 U5560 ( .A1(n5352), .A2(n5230), .B1(n5302), .B2(n5229), .ZN(n5231)
         );
  OAI221_X1 U5561 ( .B1(n5356), .B2(n5232), .C1(n4545), .C2(n2618), .A(n5231), 
        .ZN(U3287) );
  INV_X1 U5562 ( .A(n5233), .ZN(n5234) );
  NOR2_X1 U5563 ( .A1(n5235), .A2(n5234), .ZN(n5238) );
  AOI22_X1 U5564 ( .A1(n5344), .A2(n5238), .B1(n5236), .B2(n5342), .ZN(U3522)
         );
  INV_X1 U5565 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5237) );
  AOI22_X1 U5566 ( .A1(n5348), .A2(n5238), .B1(n5237), .B2(n5345), .ZN(U3475)
         );
  OAI21_X1 U5567 ( .B1(n5338), .B2(n5240), .A(n5239), .ZN(n5241) );
  AOI21_X1 U5568 ( .B1(n5340), .B2(n5242), .A(n5241), .ZN(n5245) );
  INV_X1 U5569 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5243) );
  AOI22_X1 U5570 ( .A1(n5344), .A2(n5245), .B1(n5243), .B2(n5342), .ZN(U3523)
         );
  INV_X1 U5571 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5244) );
  AOI22_X1 U5572 ( .A1(n5348), .A2(n5245), .B1(n5244), .B2(n5345), .ZN(U3477)
         );
  AOI211_X1 U5573 ( .C1(n5248), .C2(n5340), .A(n5247), .B(n5246), .ZN(n5250)
         );
  AOI22_X1 U5574 ( .A1(n5344), .A2(n5250), .B1(n2810), .B2(n5342), .ZN(U3525)
         );
  INV_X1 U5575 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U5576 ( .A1(n5348), .A2(n5250), .B1(n5249), .B2(n5345), .ZN(U3481)
         );
  INV_X1 U5577 ( .A(n5251), .ZN(n5252) );
  OAI22_X1 U5578 ( .A1(n5253), .A2(n5309), .B1(n5252), .B2(n5307), .ZN(n5254)
         );
  INV_X1 U5579 ( .A(n5254), .ZN(n5255) );
  OAI221_X1 U5580 ( .B1(n5356), .B2(n5256), .C1(n4545), .C2(n2719), .A(n5255), 
        .ZN(U3281) );
  AND3_X1 U5581 ( .A1(n5258), .A2(n5340), .A3(n5257), .ZN(n5259) );
  AOI211_X1 U5582 ( .C1(n5277), .C2(n5261), .A(n5260), .B(n5259), .ZN(n5264)
         );
  AOI22_X1 U5583 ( .A1(n5344), .A2(n5264), .B1(n5262), .B2(n5342), .ZN(U3528)
         );
  INV_X1 U5584 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5263) );
  AOI22_X1 U5585 ( .A1(n5348), .A2(n5264), .B1(n5263), .B2(n5345), .ZN(U3487)
         );
  OAI21_X1 U5586 ( .B1(n5338), .B2(n5266), .A(n5265), .ZN(n5267) );
  AOI21_X1 U5587 ( .B1(n5268), .B2(n5340), .A(n5267), .ZN(n5271) );
  AOI22_X1 U5588 ( .A1(n5344), .A2(n5271), .B1(n5269), .B2(n5342), .ZN(U3529)
         );
  INV_X1 U5589 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5270) );
  AOI22_X1 U5590 ( .A1(n5348), .A2(n5271), .B1(n5270), .B2(n5345), .ZN(U3489)
         );
  NOR2_X1 U5591 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  AOI211_X1 U5592 ( .C1(n5277), .C2(n5276), .A(n5275), .B(n5274), .ZN(n5280)
         );
  AOI22_X1 U5593 ( .A1(n5344), .A2(n5280), .B1(n5278), .B2(n5342), .ZN(U3530)
         );
  INV_X1 U5594 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U5595 ( .A1(n5348), .A2(n5280), .B1(n5279), .B2(n5345), .ZN(U3491)
         );
  AOI22_X1 U5596 ( .A1(n5284), .A2(n5283), .B1(n5282), .B2(n5281), .ZN(n5298)
         );
  NAND2_X1 U5597 ( .A1(n5286), .A2(n5285), .ZN(n5288) );
  NAND2_X1 U5598 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  XOR2_X1 U5599 ( .A(n5290), .B(n5289), .Z(n5292) );
  NOR2_X1 U5600 ( .A1(n5292), .A2(n5291), .ZN(n5293) );
  AOI211_X1 U5601 ( .C1(n5296), .C2(n5295), .A(n5294), .B(n5293), .ZN(n5297)
         );
  OAI211_X1 U5602 ( .C1(n5300), .C2(n5299), .A(n5298), .B(n5297), .ZN(U3231)
         );
  INV_X1 U5603 ( .A(n5301), .ZN(n5304) );
  AOI22_X1 U5604 ( .A1(n5304), .A2(n5352), .B1(n5303), .B2(n5302), .ZN(n5305)
         );
  OAI221_X1 U5605 ( .B1(n5356), .B2(n5306), .C1(n4545), .C2(n2732), .A(n5305), 
        .ZN(U3277) );
  OAI22_X1 U5606 ( .A1(n5310), .A2(n5309), .B1(n5308), .B2(n5307), .ZN(n5311)
         );
  INV_X1 U5607 ( .A(n5311), .ZN(n5312) );
  OAI221_X1 U5608 ( .B1(n5356), .B2(n5314), .C1(n4545), .C2(n5313), .A(n5312), 
        .ZN(U3276) );
  AOI21_X1 U5609 ( .B1(n5340), .B2(n5316), .A(n5315), .ZN(n5319) );
  INV_X1 U5610 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5317) );
  AOI22_X1 U5611 ( .A1(n5344), .A2(n5319), .B1(n5317), .B2(n5342), .ZN(U3533)
         );
  INV_X1 U5612 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5318) );
  AOI22_X1 U5613 ( .A1(n5348), .A2(n5319), .B1(n5318), .B2(n5345), .ZN(U3497)
         );
  OAI21_X1 U5614 ( .B1(n5338), .B2(n5321), .A(n5320), .ZN(n5322) );
  AOI21_X1 U5615 ( .B1(n5340), .B2(n5323), .A(n5322), .ZN(n5326) );
  INV_X1 U5616 ( .A(REG1_REG_17__SCAN_IN), .ZN(n5324) );
  AOI22_X1 U5617 ( .A1(n5344), .A2(n5326), .B1(n5324), .B2(n5342), .ZN(U3535)
         );
  INV_X1 U5618 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5325) );
  AOI22_X1 U5619 ( .A1(n5348), .A2(n5326), .B1(n5325), .B2(n5345), .ZN(U3501)
         );
  OAI22_X1 U5620 ( .A1(U3149), .A2(n5327), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5328) );
  INV_X1 U5621 ( .A(n5328), .ZN(U3334) );
  INV_X1 U5622 ( .A(n5329), .ZN(n5331) );
  AOI211_X1 U5623 ( .C1(n5332), .C2(n5340), .A(n5331), .B(n5330), .ZN(n5335)
         );
  INV_X1 U5624 ( .A(REG1_REG_18__SCAN_IN), .ZN(n5333) );
  AOI22_X1 U5625 ( .A1(n5344), .A2(n5335), .B1(n5333), .B2(n5342), .ZN(U3536)
         );
  INV_X1 U5626 ( .A(REG0_REG_18__SCAN_IN), .ZN(n5334) );
  AOI22_X1 U5627 ( .A1(n5348), .A2(n5335), .B1(n5334), .B2(n5345), .ZN(U3503)
         );
  OAI21_X1 U5628 ( .B1(n5338), .B2(n5337), .A(n5336), .ZN(n5339) );
  AOI21_X1 U5629 ( .B1(n5341), .B2(n5340), .A(n5339), .ZN(n5347) );
  AOI22_X1 U5630 ( .A1(n5344), .A2(n5347), .B1(n5343), .B2(n5342), .ZN(U3537)
         );
  INV_X1 U5631 ( .A(REG0_REG_19__SCAN_IN), .ZN(n5346) );
  AOI22_X1 U5632 ( .A1(n5348), .A2(n5347), .B1(n5346), .B2(n5345), .ZN(U3505)
         );
  AOI22_X1 U5633 ( .A1(n5349), .A2(n5352), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5356), .ZN(n5350) );
  OAI21_X1 U5634 ( .B1(n5356), .B2(n5351), .A(n5350), .ZN(U3261) );
  AOI22_X1 U5635 ( .A1(n5353), .A2(n5352), .B1(n5356), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5354) );
  OAI21_X1 U5636 ( .B1(n5356), .B2(n5355), .A(n5354), .ZN(U3260) );
  NOR2_X1 U3202 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2738)
         );
  NAND2_X1 U2609 ( .A1(n4312), .A2(n4210), .ZN(n4578) );
  INV_X2 U2524 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AND2_X2 U2552 ( .A1(n4328), .A2(n4314), .ZN(n4312) );
  CLKBUF_X1 U2554 ( .A(n4403), .Z(n4423) );
endmodule

