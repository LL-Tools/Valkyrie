

module b21_C_gen_AntiSAT_k_256_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4481, n4482, n4483, n4484, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509;

  OAI21_X1 U4986 ( .B1(n4586), .B2(n5690), .A(n4585), .ZN(n4584) );
  NOR2_X2 U4987 ( .A1(n9593), .A2(n9637), .ZN(n9592) );
  XNOR2_X1 U4990 ( .A(n4803), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U4991 ( .A1(n5557), .A2(n4976), .ZN(n5224) );
  INV_X1 U4992 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6221) );
  NAND2_X2 U4993 ( .A1(n8058), .A2(n7863), .ZN(n8804) );
  OR2_X1 U4994 ( .A1(n8481), .A2(n4900), .ZN(n6164) );
  NAND2_X1 U4996 ( .A1(n4747), .A2(n4523), .ZN(n8748) );
  OR2_X1 U4997 ( .A1(n7635), .A2(n7721), .ZN(n7771) );
  NOR2_X1 U4998 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4909) );
  NAND2_X1 U4999 ( .A1(n7238), .A2(n9876), .ZN(n8286) );
  MUX2_X1 U5000 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5222), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5223) );
  INV_X1 U5001 ( .A(n5928), .ZN(n6024) );
  NAND2_X1 U5003 ( .A1(n7786), .A2(n7505), .ZN(n6252) );
  NAND2_X1 U5004 ( .A1(n4520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5794) );
  INV_X2 U5005 ( .A(n7030), .ZN(n7804) );
  INV_X1 U5006 ( .A(n5281), .ZN(n5316) );
  OR2_X1 U5007 ( .A1(n9183), .A2(n4704), .ZN(n9137) );
  INV_X1 U5008 ( .A(n9847), .ZN(n7300) );
  NAND2_X1 U5009 ( .A1(n5115), .A2(n5114), .ZN(n5403) );
  NAND2_X1 U5010 ( .A1(n6117), .A2(n6116), .ZN(n8888) );
  AND4_X1 U5011 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n9848)
         );
  XNOR2_X1 U5012 ( .A(n5432), .B(n5431), .ZN(n6595) );
  INV_X2 U5013 ( .A(n8696), .ZN(n8788) );
  OR3_X4 U5014 ( .A1(n8199), .A2(n8324), .A3(n8325), .ZN(n4586) );
  NAND4_X1 U5015 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n5292)
         );
  OAI21_X2 U5016 ( .B1(n5374), .B2(n5373), .A(n5110), .ZN(n5389) );
  NAND2_X2 U5017 ( .A1(n4651), .A2(n5105), .ZN(n5374) );
  OR2_X2 U5018 ( .A1(n9719), .A2(n9718), .ZN(n9722) );
  XNOR2_X2 U5019 ( .A(n5794), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6255) );
  AOI21_X2 U5020 ( .B1(n8412), .B2(n8804), .A(n8411), .ZN(n8844) );
  XNOR2_X2 U5021 ( .A(n5685), .B(n5725), .ZN(n8386) );
  OR2_X1 U5023 ( .A1(n7199), .A2(n7198), .ZN(n7295) );
  OAI211_X2 U5024 ( .C1(n5316), .C2(n6526), .A(n5306), .B(n5305), .ZN(n7198)
         );
  NOR2_X1 U5025 ( .A1(n8936), .A2(n8938), .ZN(n5835) );
  AOI21_X2 U5026 ( .B1(n5046), .B2(n5044), .A(n4542), .ZN(n5043) );
  OAI21_X1 U5027 ( .B1(n4811), .B2(n9909), .A(n4783), .ZN(n5760) );
  NAND2_X1 U5028 ( .A1(n4812), .A2(n4784), .ZN(n4811) );
  XNOR2_X1 U5029 ( .A(n4780), .B(n8238), .ZN(n9148) );
  NOR2_X1 U5030 ( .A1(n9154), .A2(n9149), .ZN(n4784) );
  OAI21_X1 U5031 ( .B1(n5723), .B2(n9882), .A(n5722), .ZN(n9154) );
  AOI21_X1 U5032 ( .B1(n6165), .B2(n4951), .A(n4546), .ZN(n4949) );
  NOR2_X1 U5033 ( .A1(n9144), .A2(n9615), .ZN(n9373) );
  NAND2_X1 U5034 ( .A1(n6166), .A2(n4951), .ZN(n4950) );
  NAND2_X1 U5035 ( .A1(n8648), .A2(n8656), .ZN(n8647) );
  AOI21_X1 U5036 ( .B1(n4624), .B2(n4626), .A(n4539), .ZN(n4623) );
  NAND2_X1 U5037 ( .A1(n4496), .A2(n4705), .ZN(n4704) );
  OR2_X1 U5038 ( .A1(n6169), .A2(n4952), .ZN(n4951) );
  NAND2_X1 U5039 ( .A1(n6190), .A2(n6189), .ZN(n8852) );
  NAND2_X1 U5040 ( .A1(n6168), .A2(n6167), .ZN(n8864) );
  NAND2_X2 U5041 ( .A1(n5804), .A2(n5803), .ZN(n8867) );
  NAND2_X1 U5042 ( .A1(n6156), .A2(n6155), .ZN(n8872) );
  AOI21_X1 U5043 ( .B1(n7708), .B2(n7707), .A(n6048), .ZN(n7740) );
  XNOR2_X1 U5044 ( .A(n5626), .B(n5625), .ZN(n7613) );
  NAND2_X1 U5045 ( .A1(n5601), .A2(n5600), .ZN(n9267) );
  NAND2_X1 U5046 ( .A1(n5588), .A2(n5587), .ZN(n9284) );
  NAND2_X1 U5047 ( .A1(n6129), .A2(n6128), .ZN(n8882) );
  INV_X1 U5048 ( .A(n8400), .ZN(n4482) );
  OAI21_X1 U5049 ( .B1(n5586), .B2(n5169), .A(n5171), .ZN(n5599) );
  AND2_X1 U5050 ( .A1(n8129), .A2(n8258), .ZN(n8227) );
  NAND2_X1 U5051 ( .A1(n6021), .A2(n6020), .ZN(n7628) );
  NAND2_X1 U5052 ( .A1(n5439), .A2(n5438), .ZN(n7618) );
  NAND2_X1 U5053 ( .A1(n5456), .A2(n5455), .ZN(n9637) );
  NAND2_X1 U5054 ( .A1(n5423), .A2(n5422), .ZN(n9634) );
  AND2_X1 U5055 ( .A1(n7146), .A2(n7948), .ZN(n7111) );
  NAND2_X1 U5056 ( .A1(n5452), .A2(n4502), .ZN(n5132) );
  NAND2_X1 U5057 ( .A1(n5409), .A2(n5408), .ZN(n7501) );
  NAND2_X2 U5058 ( .A1(n9781), .A2(n7300), .ZN(n8287) );
  NAND2_X1 U5059 ( .A1(n8548), .A2(n7070), .ZN(n7918) );
  AND2_X1 U5060 ( .A1(n5880), .A2(n5879), .ZN(n8822) );
  INV_X1 U5061 ( .A(n9782), .ZN(n9876) );
  NAND2_X1 U5062 ( .A1(n5864), .A2(n5863), .ZN(n9973) );
  OAI211_X1 U5063 ( .C1(n5323), .C2(n6529), .A(n5322), .B(n5321), .ZN(n9847)
         );
  INV_X1 U5064 ( .A(n8442), .ZN(n9967) );
  INV_X2 U5065 ( .A(n6482), .ZN(n7808) );
  INV_X1 U5066 ( .A(n6689), .ZN(n9832) );
  INV_X1 U5067 ( .A(n6917), .ZN(n6818) );
  INV_X2 U5068 ( .A(n5350), .ZN(n5512) );
  INV_X1 U5069 ( .A(n6892), .ZN(n4483) );
  NAND3_X1 U5070 ( .A1(n5832), .A2(n5831), .A3(n5830), .ZN(n6917) );
  BUF_X2 U5071 ( .A(n5844), .Z(n6157) );
  NAND2_X1 U5072 ( .A1(n5094), .A2(n5093), .ZN(n5318) );
  INV_X2 U5073 ( .A(n5860), .ZN(n6070) );
  NAND2_X1 U5074 ( .A1(n5248), .A2(n5247), .ZN(n7799) );
  AND2_X1 U5075 ( .A1(n5688), .A2(n5687), .ZN(n8332) );
  CLKBUF_X1 U5076 ( .A(n5717), .Z(n8382) );
  NAND2_X4 U5077 ( .A1(n4484), .A2(n6668), .ZN(n5860) );
  NAND2_X2 U5078 ( .A1(n6521), .A2(P1_U3084), .ZN(n9548) );
  OR2_X1 U5079 ( .A1(n4643), .A2(n4645), .ZN(n4488) );
  NOR2_X1 U5080 ( .A1(n4958), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4702) );
  AND4_X1 U5081 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n5763)
         );
  AND3_X1 U5082 ( .A1(n5826), .A2(n4904), .A3(n5039), .ZN(n4647) );
  AND2_X1 U5083 ( .A1(n5207), .A2(n5275), .ZN(n4703) );
  INV_X1 U5084 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6219) );
  INV_X1 U5085 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5795) );
  INV_X1 U5086 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6086) );
  NOR2_X1 U5087 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4908) );
  NOR2_X1 U5088 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4907) );
  INV_X1 U5089 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5725) );
  NOR2_X2 U5090 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5826) );
  NOR2_X1 U5091 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5275) );
  INV_X1 U5092 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10434) );
  INV_X1 U5093 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10234) );
  INV_X1 U5094 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5556) );
  INV_X1 U5095 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5486) );
  INV_X2 U5096 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10430) );
  INV_X1 U5097 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5730) );
  BUF_X2 U5098 ( .A(n8406), .Z(n4484) );
  INV_X1 U5099 ( .A(n6100), .ZN(n4486) );
  INV_X1 U5100 ( .A(n6100), .ZN(n4487) );
  NAND2_X1 U5101 ( .A1(n6963), .A2(n7872), .ZN(n4621) );
  NAND2_X1 U5102 ( .A1(n4776), .A2(n4777), .ZN(n5452) );
  AOI21_X1 U5103 ( .B1(n4489), .B2(n4842), .A(n4778), .ZN(n4777) );
  INV_X1 U5104 ( .A(n5127), .ZN(n4778) );
  NAND2_X1 U5105 ( .A1(n4753), .A2(n4495), .ZN(n7833) );
  INV_X1 U5106 ( .A(n5835), .ZN(n7843) );
  OR2_X1 U5107 ( .A1(n9167), .A2(n9182), .ZN(n8308) );
  INV_X1 U5108 ( .A(n4836), .ZN(n4835) );
  INV_X1 U5109 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5769) );
  OAI21_X1 U5110 ( .B1(n4772), .B2(n4771), .A(n5193), .ZN(n4770) );
  INV_X1 U5111 ( .A(n5652), .ZN(n4771) );
  OAI211_X1 U5112 ( .C1(n5035), .C2(n4663), .A(n4661), .B(n4660), .ZN(n5099)
         );
  NAND2_X1 U5113 ( .A1(n4662), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4661) );
  INV_X1 U5114 ( .A(n5034), .ZN(n4662) );
  NOR2_X1 U5115 ( .A1(n7752), .A2(n4925), .ZN(n4924) );
  INV_X1 U5116 ( .A(n6065), .ZN(n4925) );
  NOR2_X1 U5117 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4906) );
  NOR2_X1 U5118 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4904) );
  INV_X1 U5119 ( .A(n8643), .ZN(n5031) );
  AOI21_X1 U5120 ( .B1(n5043), .B2(n5045), .A(n8688), .ZN(n5041) );
  NOR2_X1 U5121 ( .A1(n8705), .A2(n5047), .ZN(n5046) );
  INV_X1 U5122 ( .A(n5048), .ZN(n5047) );
  NOR2_X1 U5123 ( .A1(n8398), .A2(n5067), .ZN(n5066) );
  INV_X1 U5124 ( .A(n8396), .ZN(n5067) );
  OR2_X1 U5125 ( .A1(n8907), .A2(n7781), .ZN(n7901) );
  OR2_X1 U5126 ( .A1(n7721), .A2(n7743), .ZN(n7983) );
  OR2_X1 U5127 ( .A1(n7628), .A2(n7709), .ZN(n7977) );
  NAND2_X1 U5128 ( .A1(n5914), .A2(n5014), .ZN(n7950) );
  AND2_X1 U5129 ( .A1(n5015), .A2(n5913), .ZN(n5014) );
  NAND2_X1 U5130 ( .A1(n5769), .A2(n5798), .ZN(n5063) );
  INV_X1 U5131 ( .A(n4575), .ZN(n5770) );
  NAND2_X1 U5132 ( .A1(n4490), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6217) );
  INV_X1 U5133 ( .A(n4683), .ZN(n4682) );
  OAI21_X1 U5134 ( .B1(n4853), .B2(n4684), .A(n9039), .ZN(n4683) );
  INV_X1 U5135 ( .A(n6450), .ZN(n4857) );
  AND2_X1 U5136 ( .A1(n8981), .A2(n4856), .ZN(n4855) );
  OR2_X1 U5137 ( .A1(n9029), .A2(n4857), .ZN(n4856) );
  AND2_X1 U5138 ( .A1(n4853), .A2(n4684), .ZN(n4685) );
  OAI21_X1 U5139 ( .B1(n4508), .B2(n4884), .A(n6407), .ZN(n4883) );
  NOR2_X1 U5140 ( .A1(n4884), .A2(n4881), .ZN(n4880) );
  INV_X1 U5141 ( .A(n7621), .ZN(n4881) );
  AND2_X1 U5142 ( .A1(n5217), .A2(n5218), .ZN(n4976) );
  INV_X1 U5143 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5218) );
  OAI21_X1 U5144 ( .B1(n9192), .B2(n5665), .A(n5666), .ZN(n9176) );
  OR2_X1 U5145 ( .A1(n5643), .A2(n8991), .ZN(n5657) );
  NOR2_X1 U5146 ( .A1(n5624), .A2(n4985), .ZN(n4984) );
  INV_X1 U5147 ( .A(n5608), .ZN(n4985) );
  INV_X1 U5148 ( .A(n7799), .ZN(n5250) );
  INV_X1 U5149 ( .A(n5691), .ZN(n9168) );
  XNOR2_X1 U5150 ( .A(n7854), .B(n7853), .ZN(n7852) );
  INV_X1 U5151 ( .A(n5519), .ZN(n4847) );
  AND2_X1 U5152 ( .A1(n5434), .A2(n5433), .ZN(n5436) );
  AOI21_X1 U5153 ( .B1(n4841), .B2(n4843), .A(n4540), .ZN(n4840) );
  INV_X1 U5154 ( .A(n5074), .ZN(n4841) );
  INV_X1 U5155 ( .A(SI_11_), .ZN(n5120) );
  NAND2_X1 U5156 ( .A1(n6258), .A2(n6197), .ZN(n4916) );
  OR2_X1 U5157 ( .A1(n6266), .A2(n6242), .ZN(n6251) );
  AND2_X1 U5158 ( .A1(n4720), .A2(n4719), .ZN(n6768) );
  NAND2_X1 U5159 ( .A1(n6724), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4719) );
  AND4_X1 U5160 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n8630)
         );
  AOI21_X1 U5161 ( .B1(n4634), .B2(n4629), .A(n4538), .ZN(n4628) );
  INV_X1 U5162 ( .A(n4751), .ZN(n4750) );
  OAI21_X1 U5163 ( .B1(n4752), .B2(n7828), .A(n8003), .ZN(n4751) );
  NAND2_X1 U5164 ( .A1(n4749), .A2(n4748), .ZN(n4747) );
  INV_X1 U5165 ( .A(n4752), .ZN(n4748) );
  OR2_X1 U5166 ( .A1(n8897), .A2(n8811), .ZN(n4642) );
  OR2_X1 U5167 ( .A1(n8775), .A2(n8399), .ZN(n4640) );
  AND3_X1 U5168 ( .A1(n6108), .A2(n6107), .A3(n6106), .ZN(n8765) );
  OR2_X1 U5169 ( .A1(n10004), .A2(n7794), .ZN(n7908) );
  AND3_X1 U5170 ( .A1(n7070), .A2(n9967), .A3(n8822), .ZN(n4666) );
  AND2_X1 U5171 ( .A1(n8547), .A2(n6965), .ZN(n4620) );
  NAND2_X1 U5172 ( .A1(n5860), .A2(n6521), .ZN(n6100) );
  NAND2_X1 U5173 ( .A1(n5860), .A2(n7856), .ZN(n5847) );
  INV_X1 U5174 ( .A(n8416), .ZN(n8841) );
  NAND2_X1 U5175 ( .A1(n8410), .A2(n8409), .ZN(n8411) );
  NAND2_X1 U5176 ( .A1(n8404), .A2(n4506), .ZN(n4614) );
  AND2_X1 U5177 ( .A1(n4927), .A2(n6253), .ZN(n10013) );
  INV_X1 U5178 ( .A(n6267), .ZN(n6253) );
  NOR2_X1 U5179 ( .A1(n5800), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U5180 ( .A1(n5800), .A2(n5802), .ZN(n6668) );
  MUX2_X1 U5181 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5801), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5802) );
  NAND2_X1 U5182 ( .A1(n4895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5801) );
  OR2_X1 U5183 ( .A1(n4646), .A2(n4644), .ZN(n4895) );
  XNOR2_X1 U5184 ( .A(n5799), .B(n5798), .ZN(n8406) );
  NAND2_X1 U5185 ( .A1(n6225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5799) );
  OR2_X1 U5186 ( .A1(n5792), .A2(n5771), .ZN(n5796) );
  NAND2_X1 U5187 ( .A1(n6590), .A2(n6589), .ZN(n6588) );
  NAND2_X1 U5188 ( .A1(n8989), .A2(n8990), .ZN(n4693) );
  OR2_X1 U5189 ( .A1(n7141), .A2(n7140), .ZN(n7458) );
  AND2_X1 U5190 ( .A1(n7460), .A2(n7685), .ZN(n7679) );
  AND2_X1 U5191 ( .A1(n5261), .A2(n5260), .ZN(n9170) );
  INV_X1 U5192 ( .A(n5683), .ZN(n4979) );
  AND2_X1 U5193 ( .A1(n8308), .A2(n8318), .ZN(n9161) );
  AND2_X1 U5194 ( .A1(n4988), .A2(n4517), .ZN(n4986) );
  NAND2_X1 U5195 ( .A1(n5672), .A2(n5671), .ZN(n9385) );
  AOI21_X1 U5196 ( .B1(n8052), .B2(n4505), .A(n4738), .ZN(n4737) );
  OAI21_X1 U5197 ( .B1(n8055), .B2(n8784), .A(n8066), .ZN(n4738) );
  MUX2_X1 U5198 ( .A(n7916), .B(n7915), .S(n8053), .Z(n7931) );
  NAND2_X1 U5199 ( .A1(n4572), .A2(n4571), .ZN(n7947) );
  NAND2_X1 U5200 ( .A1(n4600), .A2(n8200), .ZN(n4599) );
  NOR2_X1 U5201 ( .A1(n8128), .A2(n9625), .ZN(n4598) );
  NAND2_X1 U5202 ( .A1(n4602), .A2(n8198), .ZN(n4601) );
  AND2_X1 U5203 ( .A1(n8264), .A2(n8261), .ZN(n4597) );
  NOR2_X1 U5204 ( .A1(n4592), .A2(n4589), .ZN(n4588) );
  AOI211_X1 U5205 ( .C1(n8154), .C2(n4596), .A(n4595), .B(n4593), .ZN(n4592)
         );
  NAND2_X1 U5206 ( .A1(n8163), .A2(n4590), .ZN(n4589) );
  NOR2_X1 U5207 ( .A1(n8096), .A2(n5710), .ZN(n4596) );
  MUX2_X1 U5208 ( .A(n8030), .B(n8029), .S(n8053), .Z(n8031) );
  NAND2_X1 U5209 ( .A1(n4838), .A2(n4833), .ZN(n4832) );
  INV_X1 U5210 ( .A(n7836), .ZN(n4833) );
  NAND2_X1 U5211 ( .A1(n6892), .A2(n6917), .ZN(n7937) );
  INV_X1 U5212 ( .A(n4886), .ZN(n4884) );
  NOR2_X1 U5213 ( .A1(n4770), .A2(n4768), .ZN(n4767) );
  INV_X1 U5214 ( .A(n5181), .ZN(n4768) );
  INV_X1 U5215 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5133) );
  INV_X1 U5216 ( .A(SI_13_), .ZN(n10456) );
  NOR2_X1 U5217 ( .A1(n7507), .A2(n4935), .ZN(n4934) );
  INV_X1 U5218 ( .A(n6004), .ZN(n4935) );
  INV_X1 U5219 ( .A(n4934), .ZN(n4930) );
  INV_X1 U5220 ( .A(n8057), .ZN(n4577) );
  NOR2_X1 U5221 ( .A1(n8867), .A2(n8872), .ZN(n4898) );
  OR2_X1 U5222 ( .A1(n8867), .A2(n8472), .ZN(n8020) );
  OR2_X1 U5223 ( .A1(n4672), .A2(n8882), .ZN(n4671) );
  NAND2_X1 U5224 ( .A1(n8732), .A2(n4673), .ZN(n4672) );
  NAND2_X1 U5225 ( .A1(n8796), .A2(n8803), .ZN(n8776) );
  NAND2_X1 U5226 ( .A1(n4548), .A2(n7968), .ZN(n4745) );
  NOR2_X1 U5227 ( .A1(n7961), .A2(n7960), .ZN(n5002) );
  NAND2_X1 U5228 ( .A1(n4604), .A2(n7271), .ZN(n7379) );
  INV_X1 U5229 ( .A(n7273), .ZN(n4604) );
  AND2_X1 U5230 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5881) );
  NAND2_X1 U5231 ( .A1(n4483), .A2(n6818), .ZN(n7935) );
  AND2_X1 U5232 ( .A1(n7940), .A2(n7938), .ZN(n7869) );
  OR2_X1 U5233 ( .A1(n8901), .A2(n7826), .ZN(n8779) );
  AOI21_X1 U5234 ( .B1(n9947), .B2(n9941), .A(n9949), .ZN(n6976) );
  INV_X1 U5235 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U5236 ( .A1(n4956), .A2(n6086), .ZN(n4955) );
  INV_X1 U5237 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4956) );
  INV_X1 U5238 ( .A(n4647), .ZN(n4643) );
  INV_X1 U5239 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U5240 ( .A1(n7236), .A2(n4527), .ZN(n6347) );
  INV_X1 U5241 ( .A(n6530), .ZN(n4699) );
  OR2_X1 U5242 ( .A1(n9385), .A2(n9199), .ZN(n8362) );
  INV_X1 U5243 ( .A(n8161), .ZN(n4826) );
  NOR2_X1 U5244 ( .A1(n4826), .A2(n4827), .ZN(n4825) );
  INV_X1 U5245 ( .A(n9289), .ZN(n4827) );
  OR2_X1 U5246 ( .A1(n9409), .A2(n9263), .ZN(n8091) );
  OR2_X1 U5247 ( .A1(n9284), .A2(n9293), .ZN(n8298) );
  NAND2_X1 U5248 ( .A1(n8251), .A2(n8099), .ZN(n4817) );
  NOR2_X1 U5249 ( .A1(n9083), .A2(n8962), .ZN(n4707) );
  NAND2_X1 U5250 ( .A1(n5232), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5493) );
  INV_X1 U5251 ( .A(n5477), .ZN(n5232) );
  NOR2_X1 U5252 ( .A1(n8256), .A2(n4814), .ZN(n4813) );
  INV_X1 U5253 ( .A(n5324), .ZN(n4962) );
  AND2_X1 U5254 ( .A1(n4700), .A2(n5556), .ZN(n4695) );
  INV_X1 U5255 ( .A(n8386), .ZN(n5716) );
  INV_X1 U5256 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5240) );
  INV_X1 U5257 ( .A(n5224), .ZN(n5243) );
  INV_X1 U5258 ( .A(n5256), .ZN(n4838) );
  AOI21_X1 U5259 ( .B1(n5256), .B2(n4837), .A(n4561), .ZN(n4836) );
  INV_X1 U5260 ( .A(n5201), .ZN(n4837) );
  NAND2_X1 U5261 ( .A1(n5200), .A2(n5199), .ZN(n5669) );
  AND2_X1 U5262 ( .A1(n5193), .A2(n5192), .ZN(n5652) );
  NAND3_X1 U5263 ( .A1(n4696), .A2(n4888), .A3(n4695), .ZN(n4891) );
  AND2_X1 U5264 ( .A1(n5076), .A2(n4889), .ZN(n4888) );
  NAND2_X1 U5265 ( .A1(n5612), .A2(n5181), .ZN(n5626) );
  NAND2_X1 U5266 ( .A1(n5684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5686) );
  OAI21_X1 U5267 ( .B1(n5553), .B2(n5552), .A(n5161), .ZN(n5572) );
  AND2_X1 U5268 ( .A1(n5166), .A2(n5165), .ZN(n5571) );
  AOI21_X1 U5269 ( .B1(n4758), .B2(n4503), .A(n4756), .ZN(n4755) );
  AND2_X1 U5270 ( .A1(n5147), .A2(n5146), .ZN(n5501) );
  INV_X1 U5271 ( .A(n4759), .ZN(n4758) );
  OAI21_X1 U5272 ( .B1(n4762), .B2(n4503), .A(n5142), .ZN(n4759) );
  INV_X1 U5273 ( .A(n5119), .ZN(n4844) );
  OR2_X1 U5274 ( .A1(n5469), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U5275 ( .A1(n5359), .A2(n5103), .ZN(n4651) );
  AOI21_X1 U5276 ( .B1(n5098), .B2(n5000), .A(n4534), .ZN(n4999) );
  INV_X1 U5277 ( .A(n6016), .ZN(n4932) );
  NAND2_X1 U5278 ( .A1(n8507), .A2(n6154), .ZN(n6159) );
  NAND2_X1 U5279 ( .A1(n4920), .A2(n4918), .ZN(n4657) );
  AND2_X1 U5280 ( .A1(n4919), .A2(n7780), .ZN(n4918) );
  NAND2_X1 U5281 ( .A1(n4921), .A2(n4923), .ZN(n4919) );
  OR2_X1 U5282 ( .A1(n6250), .A2(n6249), .ZN(n6258) );
  NAND2_X1 U5283 ( .A1(n7186), .A2(n5956), .ZN(n4947) );
  INV_X1 U5284 ( .A(n5956), .ZN(n4948) );
  AND2_X1 U5285 ( .A1(n8061), .A2(n7892), .ZN(n6267) );
  NOR2_X1 U5286 ( .A1(n8483), .A2(n4653), .ZN(n6166) );
  NAND2_X1 U5287 ( .A1(n4655), .A2(n4654), .ZN(n4653) );
  INV_X1 U5288 ( .A(n8482), .ZN(n4654) );
  NAND2_X1 U5289 ( .A1(n8485), .A2(n8472), .ZN(n4655) );
  AND4_X1 U5290 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n8534)
         );
  OR2_X1 U5291 ( .A1(n6748), .A2(n6747), .ZN(n4720) );
  OR2_X1 U5292 ( .A1(n6768), .A2(n6767), .ZN(n4718) );
  NOR2_X1 U5293 ( .A1(n8591), .A2(n4563), .ZN(n8593) );
  NAND2_X1 U5294 ( .A1(n8593), .A2(n8594), .ZN(n8606) );
  NOR2_X1 U5295 ( .A1(n8635), .A2(n8841), .ZN(n8624) );
  NAND2_X1 U5296 ( .A1(n8650), .A2(n8640), .ZN(n8635) );
  NOR2_X1 U5297 ( .A1(n5030), .A2(n8024), .ZN(n4754) );
  NOR2_X1 U5298 ( .A1(n8655), .A2(n8656), .ZN(n8654) );
  AND2_X1 U5299 ( .A1(n8025), .A2(n8028), .ZN(n8675) );
  INV_X1 U5300 ( .A(n8401), .ZN(n4626) );
  INV_X1 U5301 ( .A(n5046), .ZN(n5045) );
  NAND2_X1 U5302 ( .A1(n5042), .A2(n5041), .ZN(n8682) );
  INV_X1 U5303 ( .A(n8720), .ZN(n5044) );
  OAI21_X1 U5304 ( .B1(n5011), .B2(n7896), .A(n5007), .ZN(n8706) );
  NAND2_X1 U5305 ( .A1(n8872), .A2(n5012), .ZN(n5048) );
  AND3_X1 U5306 ( .A1(n8016), .A2(n8008), .A3(n7829), .ZN(n5011) );
  NAND2_X1 U5307 ( .A1(n5008), .A2(n8748), .ZN(n5013) );
  NAND2_X1 U5308 ( .A1(n8016), .A2(n7829), .ZN(n8720) );
  AOI22_X1 U5309 ( .A1(n4510), .A2(n8734), .B1(n8534), .B2(n8732), .ZN(n8714)
         );
  NAND2_X1 U5310 ( .A1(n8714), .A2(n8720), .ZN(n8713) );
  NAND2_X1 U5311 ( .A1(n4509), .A2(n4637), .ZN(n4636) );
  INV_X1 U5312 ( .A(n8399), .ZN(n4637) );
  NAND2_X1 U5313 ( .A1(n4635), .A2(n4509), .ZN(n4634) );
  INV_X1 U5314 ( .A(n4638), .ZN(n4635) );
  NAND2_X1 U5315 ( .A1(n4482), .A2(n8757), .ZN(n4752) );
  AND2_X1 U5316 ( .A1(n8805), .A2(n7828), .ZN(n8781) );
  AOI21_X1 U5317 ( .B1(n7990), .B2(n5066), .A(n4518), .ZN(n5064) );
  AOI21_X1 U5318 ( .B1(n5026), .B2(n7902), .A(n5027), .ZN(n5025) );
  NAND2_X1 U5319 ( .A1(n7728), .A2(n5026), .ZN(n5024) );
  INV_X1 U5320 ( .A(n7901), .ZN(n5027) );
  AND2_X1 U5321 ( .A1(n8779), .A2(n7999), .ZN(n8806) );
  OR2_X1 U5322 ( .A1(n7767), .A2(n7990), .ZN(n8397) );
  OR2_X1 U5323 ( .A1(n7728), .A2(n7902), .ZN(n7761) );
  NAND2_X1 U5324 ( .A1(n7588), .A2(n4526), .ZN(n7630) );
  NAND2_X1 U5325 ( .A1(n7560), .A2(n5072), .ZN(n7588) );
  NOR2_X1 U5326 ( .A1(n7970), .A2(n5073), .ZN(n5072) );
  INV_X1 U5327 ( .A(n7559), .ZN(n5073) );
  AND2_X1 U5328 ( .A1(n7973), .A2(n7972), .ZN(n7970) );
  NAND2_X1 U5329 ( .A1(n5052), .A2(n5050), .ZN(n5078) );
  NAND2_X1 U5330 ( .A1(n5051), .A2(n7518), .ZN(n5050) );
  NAND2_X1 U5331 ( .A1(n5053), .A2(n4531), .ZN(n5052) );
  INV_X1 U5332 ( .A(n7879), .ZN(n5051) );
  NAND2_X1 U5333 ( .A1(n5078), .A2(n7520), .ZN(n7560) );
  AND4_X1 U5334 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n7794)
         );
  NAND2_X1 U5335 ( .A1(n5006), .A2(n7485), .ZN(n5005) );
  INV_X1 U5336 ( .A(n7477), .ZN(n5006) );
  AND4_X1 U5337 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n7793)
         );
  NAND2_X1 U5338 ( .A1(n7379), .A2(n5049), .ZN(n5053) );
  NOR2_X1 U5339 ( .A1(n7485), .A2(n5054), .ZN(n5049) );
  INV_X1 U5340 ( .A(n7378), .ZN(n5054) );
  NAND2_X1 U5341 ( .A1(n7107), .A2(n4619), .ZN(n5056) );
  AND2_X1 U5342 ( .A1(n4551), .A2(n7106), .ZN(n4619) );
  AND2_X1 U5343 ( .A1(n5059), .A2(n4550), .ZN(n5057) );
  NAND2_X1 U5344 ( .A1(n7266), .A2(n5060), .ZN(n5059) );
  INV_X1 U5345 ( .A(n7108), .ZN(n5060) );
  AND4_X1 U5346 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(n7381)
         );
  AND2_X1 U5347 ( .A1(n6555), .A2(n8942), .ZN(n8809) );
  NAND2_X1 U5348 ( .A1(n6926), .A2(n7873), .ZN(n6929) );
  NAND2_X1 U5349 ( .A1(n5846), .A2(n4649), .ZN(n8442) );
  OAI21_X1 U5350 ( .B1(n5847), .B2(n6526), .A(n4650), .ZN(n4648) );
  AND4_X1 U5351 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n6915)
         );
  NAND2_X1 U5352 ( .A1(n6668), .A2(n6555), .ZN(n8762) );
  INV_X1 U5353 ( .A(n8809), .ZN(n8764) );
  OR2_X1 U5354 ( .A1(n10024), .A2(n7892), .ZN(n6973) );
  INV_X1 U5355 ( .A(n8762), .ZN(n8810) );
  NAND2_X1 U5356 ( .A1(n8042), .A2(n8036), .ZN(n8643) );
  NAND2_X1 U5357 ( .A1(n8647), .A2(n8403), .ZN(n8644) );
  NOR2_X1 U5358 ( .A1(n8404), .A2(n4506), .ZN(n4616) );
  NAND2_X1 U5359 ( .A1(n5021), .A2(n5020), .ZN(n5019) );
  INV_X1 U5360 ( .A(n7349), .ZN(n5021) );
  INV_X1 U5361 ( .A(n10024), .ZN(n10014) );
  INV_X1 U5362 ( .A(n6941), .ZN(n6821) );
  NOR2_X1 U5363 ( .A1(n5063), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U5364 ( .A1(n6218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6241) );
  AND2_X1 U5365 ( .A1(n5892), .A2(n5878), .ZN(n6724) );
  OR2_X1 U5366 ( .A1(n5826), .A2(n5771), .ZN(n5834) );
  AND2_X1 U5367 ( .A1(n6493), .A2(n6487), .ZN(n4876) );
  OR2_X1 U5368 ( .A1(n7668), .A2(n7667), .ZN(n4886) );
  INV_X1 U5369 ( .A(n6384), .ZN(n4885) );
  AND2_X1 U5370 ( .A1(n7544), .A2(n6376), .ZN(n7620) );
  NAND2_X1 U5371 ( .A1(n5236), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5631) );
  OR2_X1 U5372 ( .A1(n6468), .A2(n4867), .ZN(n4866) );
  INV_X1 U5373 ( .A(n8965), .ZN(n4867) );
  OR2_X1 U5374 ( .A1(n5562), .A2(n5561), .ZN(n5576) );
  AOI21_X1 U5375 ( .B1(n4855), .B2(n4857), .A(n4535), .ZN(n4853) );
  NAND2_X1 U5376 ( .A1(n4852), .A2(n4685), .ZN(n9037) );
  NAND2_X1 U5377 ( .A1(n6588), .A2(n6287), .ZN(n6599) );
  AND3_X1 U5378 ( .A1(n5549), .A2(n5548), .A3(n5547), .ZN(n6433) );
  AND4_X1 U5380 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n9836)
         );
  XNOR2_X1 U5381 ( .A(n6868), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6864) );
  OR2_X1 U5382 ( .A1(n9556), .A2(n9555), .ZN(n4794) );
  OR2_X1 U5383 ( .A1(n5390), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5469) );
  OR2_X1 U5384 ( .A1(n7000), .A2(n6999), .ZN(n4796) );
  AND2_X1 U5385 ( .A1(n4796), .A2(n4795), .ZN(n7141) );
  NAND2_X1 U5386 ( .A1(n7139), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4795) );
  NOR2_X1 U5387 ( .A1(n9129), .A2(n4789), .ZN(n9732) );
  AND2_X1 U5388 ( .A1(n9121), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4789) );
  OR2_X1 U5389 ( .A1(n6275), .A2(n7555), .ZN(n6620) );
  OR2_X1 U5390 ( .A1(n9732), .A2(n9733), .ZN(n4788) );
  NAND2_X1 U5391 ( .A1(n5557), .A2(n5217), .ZN(n5221) );
  NAND2_X1 U5392 ( .A1(n5238), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U5393 ( .A1(n4957), .A2(n5651), .ZN(n9192) );
  AOI21_X1 U5394 ( .B1(n4984), .B2(n4492), .A(n4532), .ZN(n4983) );
  AND2_X1 U5395 ( .A1(n8091), .A2(n8166), .ZN(n9240) );
  OR2_X1 U5396 ( .A1(n9295), .A2(n9309), .ZN(n9270) );
  NOR2_X1 U5397 ( .A1(n9317), .A2(n4815), .ZN(n4820) );
  INV_X1 U5398 ( .A(n8099), .ZN(n4815) );
  INV_X1 U5399 ( .A(n4989), .ZN(n4988) );
  OAI21_X1 U5400 ( .B1(n5483), .B2(n4990), .A(n4996), .ZN(n4989) );
  NAND2_X1 U5401 ( .A1(n4516), .A2(n4994), .ZN(n4990) );
  NOR2_X1 U5402 ( .A1(n5483), .A2(n4993), .ZN(n4992) );
  INV_X1 U5403 ( .A(n4994), .ZN(n4993) );
  OR2_X1 U5404 ( .A1(n8254), .A2(n8278), .ZN(n8230) );
  NAND2_X1 U5405 ( .A1(n9637), .A2(n9089), .ZN(n4994) );
  AND2_X1 U5406 ( .A1(n4973), .A2(n8127), .ZN(n4972) );
  NAND2_X1 U5407 ( .A1(n4974), .A2(n8126), .ZN(n4973) );
  NAND2_X1 U5408 ( .A1(n7118), .A2(n8255), .ZN(n9760) );
  NAND2_X1 U5409 ( .A1(n7799), .A2(n5249), .ZN(n5511) );
  AND2_X1 U5410 ( .A1(n9538), .A2(n7799), .ZN(n5350) );
  AND2_X1 U5411 ( .A1(n5249), .A2(n5250), .ZN(n5284) );
  INV_X1 U5412 ( .A(n8333), .ZN(n9798) );
  OR2_X1 U5413 ( .A1(n6503), .A2(P1_U3084), .ZN(n7239) );
  NAND2_X1 U5414 ( .A1(n6275), .A2(n6496), .ZN(n7009) );
  XNOR2_X1 U5415 ( .A(n4828), .B(n7858), .ZN(n8194) );
  OAI21_X1 U5416 ( .B1(n7852), .B2(n4829), .A(n7855), .ZN(n4828) );
  XNOR2_X1 U5417 ( .A(n5244), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U5418 ( .A1(n5247), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5244) );
  XNOR2_X1 U5419 ( .A(n7852), .B(SI_30_), .ZN(n8935) );
  NAND2_X1 U5420 ( .A1(n5686), .A2(n10434), .ZN(n5688) );
  XNOR2_X1 U5421 ( .A(n5572), .B(n5571), .ZN(n7444) );
  NAND2_X1 U5422 ( .A1(n4761), .A2(n5136), .ZN(n5485) );
  NAND2_X1 U5423 ( .A1(n5132), .A2(n4762), .ZN(n4761) );
  NAND2_X1 U5424 ( .A1(n4845), .A2(n5119), .ZN(n5419) );
  NAND2_X1 U5425 ( .A1(n5403), .A2(n5074), .ZN(n4845) );
  NAND2_X1 U5426 ( .A1(n6572), .A2(n5891), .ZN(n4658) );
  NAND2_X1 U5427 ( .A1(n8443), .A2(n8445), .ZN(n8444) );
  NAND2_X1 U5428 ( .A1(n6103), .A2(n6102), .ZN(n8897) );
  NOR2_X1 U5429 ( .A1(n4915), .A2(n4917), .ZN(n4911) );
  NOR2_X1 U5430 ( .A1(n6246), .A2(n6197), .ZN(n4917) );
  INV_X1 U5431 ( .A(n6258), .ZN(n4914) );
  NAND2_X1 U5432 ( .A1(n4940), .A2(n4937), .ZN(n7057) );
  AOI21_X1 U5433 ( .B1(n4939), .B2(n4938), .A(n4530), .ZN(n4937) );
  NAND2_X1 U5434 ( .A1(n7077), .A2(n4936), .ZN(n4940) );
  OR2_X1 U5435 ( .A1(n7187), .A2(n7186), .ZN(n7184) );
  NAND2_X1 U5436 ( .A1(n7468), .A2(n7469), .ZN(n7467) );
  INV_X1 U5437 ( .A(n7483), .ZN(n10012) );
  INV_X1 U5438 ( .A(n8526), .ZN(n8498) );
  OAI21_X1 U5439 ( .B1(n6251), .B2(n6244), .A(n8821), .ZN(n8503) );
  NAND2_X1 U5440 ( .A1(n4942), .A2(n5906), .ZN(n7075) );
  NAND2_X1 U5441 ( .A1(n6259), .A2(n6256), .ZN(n8505) );
  AND2_X1 U5442 ( .A1(n4736), .A2(n7553), .ZN(n4734) );
  INV_X1 U5443 ( .A(n4505), .ZN(n4736) );
  NAND2_X1 U5444 ( .A1(n4498), .A2(n7553), .ZN(n4735) );
  AND2_X1 U5445 ( .A1(n7832), .A2(n7831), .ZN(n8416) );
  NAND2_X1 U5446 ( .A1(n6007), .A2(n6006), .ZN(n7586) );
  NAND2_X1 U5447 ( .A1(n5058), .A2(n7108), .ZN(n7267) );
  INV_X1 U5448 ( .A(n8821), .ZN(n8800) );
  NAND2_X1 U5449 ( .A1(n4618), .A2(n8404), .ZN(n4612) );
  NAND2_X1 U5450 ( .A1(n8642), .A2(n4606), .ZN(n4605) );
  NOR2_X1 U5451 ( .A1(n5069), .A2(n4607), .ZN(n4606) );
  INV_X1 U5452 ( .A(n4616), .ZN(n4607) );
  INV_X1 U5453 ( .A(n4609), .ZN(n4608) );
  OAI21_X1 U5454 ( .B1(n5069), .B2(n4536), .A(n10052), .ZN(n4609) );
  INV_X1 U5455 ( .A(n4614), .ZN(n4613) );
  NAND2_X1 U5456 ( .A1(n7236), .A2(n7234), .ZN(n6338) );
  NOR2_X1 U5457 ( .A1(n6493), .A2(n4874), .ZN(n4871) );
  AND2_X1 U5458 ( .A1(n4873), .A2(n4877), .ZN(n4872) );
  INV_X1 U5459 ( .A(n4878), .ZN(n4877) );
  NAND2_X1 U5460 ( .A1(n4876), .A2(n4874), .ZN(n4873) );
  OAI21_X1 U5461 ( .B1(n6493), .B2(n6487), .A(n9056), .ZN(n4878) );
  INV_X1 U5462 ( .A(n4876), .ZN(n4875) );
  NAND2_X1 U5463 ( .A1(n4687), .A2(n4686), .ZN(n7823) );
  AOI21_X1 U5464 ( .B1(n4688), .B2(n4691), .A(n4537), .ZN(n4686) );
  NAND2_X1 U5465 ( .A1(n8941), .A2(n8193), .ZN(n5258) );
  XNOR2_X1 U5466 ( .A(n6290), .B(n7804), .ZN(n6601) );
  NAND2_X1 U5467 ( .A1(n6803), .A2(n6307), .ZN(n7022) );
  AND2_X1 U5468 ( .A1(n4693), .A2(n4524), .ZN(n9059) );
  AND2_X1 U5469 ( .A1(n9789), .A2(n4481), .ZN(n4565) );
  INV_X1 U5470 ( .A(n9398), .ZN(n9196) );
  INV_X1 U5471 ( .A(n9762), .ZN(n9091) );
  OR2_X1 U5472 ( .A1(n7679), .A2(n7461), .ZN(n7462) );
  INV_X1 U5473 ( .A(n9136), .ZN(n9143) );
  AND2_X1 U5474 ( .A1(n4980), .A2(n4978), .ZN(n9159) );
  INV_X1 U5475 ( .A(n9385), .ZN(n9189) );
  NAND2_X1 U5476 ( .A1(n5560), .A2(n5559), .ZN(n9434) );
  OR2_X1 U5477 ( .A1(n7032), .A2(n9789), .ZN(n9361) );
  NAND2_X1 U5478 ( .A1(n8386), .A2(n8243), .ZN(n7011) );
  NAND2_X1 U5479 ( .A1(n9148), .A2(n9885), .ZN(n4812) );
  OR2_X1 U5480 ( .A1(n7945), .A2(n8053), .ZN(n4571) );
  AND2_X1 U5481 ( .A1(n4570), .A2(n7958), .ZN(n7965) );
  OAI21_X1 U5482 ( .B1(n8125), .B2(n8124), .A(n4603), .ZN(n4602) );
  AND2_X1 U5483 ( .A1(n8129), .A2(n8123), .ZN(n4603) );
  OAI21_X1 U5484 ( .B1(n8120), .B2(n8256), .A(n8119), .ZN(n4600) );
  NAND2_X1 U5485 ( .A1(n8137), .A2(n4597), .ZN(n8142) );
  AOI21_X1 U5486 ( .B1(n8000), .B2(n7999), .A(n7998), .ZN(n8005) );
  NOR2_X1 U5487 ( .A1(n4529), .A2(n4591), .ZN(n4590) );
  NOR2_X1 U5488 ( .A1(n8303), .A2(n8198), .ZN(n4591) );
  NAND2_X1 U5489 ( .A1(n8298), .A2(n4594), .ZN(n4593) );
  AND2_X1 U5490 ( .A1(n9270), .A2(n8198), .ZN(n4594) );
  MUX2_X1 U5491 ( .A(n8012), .B(n8011), .S(n8034), .Z(n8013) );
  NAND2_X1 U5492 ( .A1(n8162), .A2(n4588), .ZN(n8164) );
  OR2_X1 U5493 ( .A1(n9228), .A2(n8992), .ZN(n8092) );
  INV_X1 U5494 ( .A(n4574), .ZN(n4573) );
  OAI21_X1 U5495 ( .B1(n8035), .B2(n8034), .A(n8042), .ZN(n4574) );
  NOR2_X1 U5496 ( .A1(n8882), .A2(n8535), .ZN(n5055) );
  AOI21_X1 U5497 ( .B1(n5669), .B2(n4834), .A(n4831), .ZN(n4830) );
  NOR2_X1 U5498 ( .A1(n4835), .A2(n7836), .ZN(n4834) );
  OAI21_X1 U5499 ( .B1(n4835), .B2(n4832), .A(n7835), .ZN(n4831) );
  INV_X1 U5500 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5149) );
  INV_X1 U5501 ( .A(n5501), .ZN(n4756) );
  INV_X1 U5502 ( .A(n5431), .ZN(n4846) );
  INV_X1 U5503 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5123) );
  NOR2_X1 U5504 ( .A1(n5333), .A2(n5317), .ZN(n4998) );
  INV_X1 U5505 ( .A(n5097), .ZN(n5000) );
  INV_X1 U5506 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U5507 ( .A1(n10486), .A2(n5080), .ZN(n5037) );
  INV_X1 U5508 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5509 ( .A1(n5081), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5033) );
  INV_X1 U5510 ( .A(SI_12_), .ZN(n10212) );
  INV_X1 U5511 ( .A(SI_9_), .ZN(n10145) );
  INV_X1 U5512 ( .A(n5907), .ZN(n4941) );
  AND2_X1 U5513 ( .A1(n8485), .A2(n6161), .ZN(n4900) );
  NAND2_X1 U5514 ( .A1(n7648), .A2(n4715), .ZN(n8552) );
  OR2_X1 U5515 ( .A1(n7649), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4715) );
  NOR2_X1 U5516 ( .A1(n8734), .A2(n5010), .ZN(n5008) );
  INV_X1 U5517 ( .A(n8006), .ZN(n5010) );
  NAND2_X1 U5518 ( .A1(n5009), .A2(n5012), .ZN(n8016) );
  AND2_X1 U5519 ( .A1(n4634), .A2(n4633), .ZN(n4632) );
  INV_X1 U5520 ( .A(n5055), .ZN(n4633) );
  NOR2_X1 U5521 ( .A1(n5055), .A2(n4630), .ZN(n4629) );
  INV_X1 U5522 ( .A(n4636), .ZN(n4630) );
  NOR2_X1 U5523 ( .A1(n7824), .A2(n5028), .ZN(n5026) );
  INV_X1 U5524 ( .A(n7986), .ZN(n5028) );
  OR2_X1 U5525 ( .A1(n5945), .A2(n5944), .ZN(n5962) );
  NAND2_X1 U5526 ( .A1(n7270), .A2(n7269), .ZN(n7273) );
  AND2_X1 U5527 ( .A1(n7909), .A2(n7956), .ZN(n7278) );
  NAND2_X1 U5528 ( .A1(n5860), .A2(n4512), .ZN(n4650) );
  INV_X1 U5529 ( .A(n7873), .ZN(n7930) );
  NAND2_X1 U5530 ( .A1(n9967), .A2(n8549), .ZN(n7917) );
  NAND2_X1 U5531 ( .A1(n7935), .A2(n7937), .ZN(n5038) );
  NOR2_X1 U5532 ( .A1(n7771), .A2(n8912), .ZN(n7772) );
  INV_X1 U5533 ( .A(n5063), .ZN(n5061) );
  NAND2_X1 U5534 ( .A1(n5770), .A2(n5769), .ZN(n6225) );
  INV_X1 U5535 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5039) );
  NOR2_X1 U5536 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  OR2_X1 U5537 ( .A1(n5911), .A2(n5910), .ZN(n5924) );
  INV_X1 U5538 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5909) );
  NOR2_X1 U5539 ( .A1(n4682), .A2(n4685), .ZN(n4680) );
  AOI21_X1 U5540 ( .B1(n4682), .B2(n4684), .A(n4499), .ZN(n4679) );
  NAND2_X1 U5541 ( .A1(n7020), .A2(n6312), .ZN(n7229) );
  NOR2_X1 U5542 ( .A1(n9267), .A2(n9409), .ZN(n4713) );
  NOR2_X1 U5543 ( .A1(n9228), .A2(n4712), .ZN(n4711) );
  INV_X1 U5544 ( .A(n4713), .ZN(n4712) );
  INV_X1 U5545 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5457) );
  OR2_X1 U5546 ( .A1(n5458), .A2(n5457), .ZN(n5477) );
  INV_X1 U5547 ( .A(n5417), .ZN(n4974) );
  NOR2_X1 U5548 ( .A1(n4975), .A2(n4971), .ZN(n4970) );
  INV_X1 U5549 ( .A(n8126), .ZN(n4975) );
  INV_X1 U5550 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5394) );
  OR2_X1 U5551 ( .A1(n5395), .A2(n5394), .ZN(n5410) );
  NAND2_X1 U5552 ( .A1(n5716), .A2(n9814), .ZN(n6498) );
  NAND2_X1 U5553 ( .A1(n9280), .A2(n9504), .ZN(n9264) );
  AND2_X1 U5554 ( .A1(n9508), .A2(n9294), .ZN(n9280) );
  OR2_X1 U5555 ( .A1(n9434), .A2(n9325), .ZN(n9311) );
  INV_X1 U5556 ( .A(n9807), .ZN(n9803) );
  OAI21_X1 U5557 ( .B1(n6547), .B2(P1_D_REG_1__SCAN_IN), .A(n6550), .ZN(n7006)
         );
  INV_X1 U5558 ( .A(SI_30_), .ZN(n4829) );
  NAND2_X1 U5559 ( .A1(n4766), .A2(n4765), .ZN(n5668) );
  OR2_X1 U5560 ( .A1(n4770), .A2(n4559), .ZN(n4765) );
  AOI21_X1 U5561 ( .B1(n4774), .B2(n5184), .A(n4773), .ZN(n4772) );
  INV_X1 U5562 ( .A(n5188), .ZN(n4773) );
  NOR2_X1 U5563 ( .A1(n5639), .A2(n4775), .ZN(n4774) );
  INV_X1 U5564 ( .A(n5183), .ZN(n4775) );
  AND2_X1 U5565 ( .A1(n5181), .A2(n5180), .ZN(n5609) );
  NAND2_X1 U5566 ( .A1(n5724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5689) );
  INV_X1 U5567 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5521) );
  OR2_X1 U5568 ( .A1(n5503), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5504) );
  INV_X1 U5569 ( .A(n5136), .ZN(n4760) );
  NOR2_X1 U5570 ( .A1(n5137), .A2(n4763), .ZN(n4762) );
  INV_X1 U5571 ( .A(n5131), .ZN(n4763) );
  INV_X1 U5572 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U5573 ( .A1(n4652), .A2(n5102), .ZN(n5359) );
  NAND2_X1 U5574 ( .A1(n5208), .A2(n4959), .ZN(n4958) );
  INV_X1 U5575 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4959) );
  NOR2_X1 U5576 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5207) );
  NAND2_X1 U5577 ( .A1(n4703), .A2(n5208), .ZN(n5335) );
  NAND2_X1 U5578 ( .A1(n7467), .A2(n4934), .ZN(n4933) );
  NOR2_X1 U5579 ( .A1(n5906), .A2(n4941), .ZN(n4938) );
  NAND2_X1 U5580 ( .A1(n7740), .A2(n7741), .ZN(n7739) );
  NAND2_X1 U5581 ( .A1(n4901), .A2(n6160), .ZN(n8481) );
  INV_X1 U5582 ( .A(n6159), .ZN(n4901) );
  AND2_X1 U5583 ( .A1(n6114), .A2(n6099), .ZN(n4656) );
  AND2_X1 U5584 ( .A1(n5976), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5993) );
  AND2_X1 U5585 ( .A1(n6075), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6091) );
  AND2_X1 U5586 ( .A1(n6091), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6104) );
  INV_X1 U5587 ( .A(n4924), .ZN(n4923) );
  AOI21_X1 U5588 ( .B1(n4924), .B2(n4922), .A(n4544), .ZN(n4921) );
  INV_X1 U5589 ( .A(n7741), .ZN(n4922) );
  INV_X1 U5590 ( .A(n8469), .ZN(n4952) );
  AOI21_X1 U5591 ( .B1(n4931), .B2(n4930), .A(n4929), .ZN(n4928) );
  INV_X1 U5592 ( .A(n6034), .ZN(n4929) );
  AND2_X1 U5593 ( .A1(n8416), .A2(n8634), .ZN(n8044) );
  NAND2_X1 U5594 ( .A1(n8048), .A2(n7865), .ZN(n4578) );
  NAND2_X1 U5595 ( .A1(n7890), .A2(n7892), .ZN(n4739) );
  AND3_X1 U5596 ( .A1(n7848), .A2(n7847), .A3(n7846), .ZN(n8530) );
  AND4_X1 U5597 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n8472)
         );
  AND4_X1 U5598 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(n7581)
         );
  AND4_X1 U5599 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n7268)
         );
  AND4_X1 U5600 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n7110)
         );
  AND4_X1 U5601 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n6914)
         );
  NOR2_X1 U5602 ( .A1(n6694), .A2(n4511), .ZN(n6665) );
  OR2_X1 U5603 ( .A1(n6665), .A2(n6664), .ZN(n4724) );
  NAND2_X1 U5604 ( .A1(n4724), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U5605 ( .A1(n6729), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U5606 ( .A1(n6711), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4717) );
  NOR2_X1 U5607 ( .A1(n6777), .A2(n4728), .ZN(n6789) );
  AND2_X1 U5608 ( .A1(n6721), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4728) );
  NOR2_X1 U5609 ( .A1(n6789), .A2(n6788), .ZN(n6787) );
  NOR2_X1 U5610 ( .A1(n7091), .A2(n4730), .ZN(n7093) );
  AND2_X1 U5611 ( .A1(n7092), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4730) );
  NOR2_X1 U5612 ( .A1(n7094), .A2(n7093), .ZN(n7166) );
  NOR2_X1 U5613 ( .A1(n7166), .A2(n4729), .ZN(n7169) );
  AND2_X1 U5614 ( .A1(n7174), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5615 ( .A1(n7169), .A2(n7168), .ZN(n7322) );
  NAND2_X1 U5616 ( .A1(n7324), .A2(n7325), .ZN(n7425) );
  NAND2_X1 U5617 ( .A1(n7425), .A2(n4716), .ZN(n7427) );
  OR2_X1 U5618 ( .A1(n7426), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U5619 ( .A1(n7427), .A2(n7428), .ZN(n7648) );
  AND2_X1 U5620 ( .A1(n5761), .A2(n4905), .ZN(n5762) );
  NOR2_X1 U5621 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5761) );
  NOR2_X1 U5622 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4905) );
  XNOR2_X1 U5623 ( .A(n4726), .B(n4725), .ZN(n8612) );
  INV_X1 U5624 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n4725) );
  NAND2_X1 U5625 ( .A1(n8606), .A2(n4564), .ZN(n4726) );
  AND4_X1 U5626 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n8657)
         );
  NOR2_X1 U5627 ( .A1(n8668), .A2(n8852), .ZN(n8650) );
  INV_X1 U5628 ( .A(n4671), .ZN(n4670) );
  NAND2_X1 U5629 ( .A1(n4896), .A2(n8672), .ZN(n8668) );
  OR2_X1 U5630 ( .A1(n6171), .A2(n6170), .ZN(n6179) );
  NAND2_X1 U5631 ( .A1(n8728), .A2(n4898), .ZN(n8699) );
  NAND2_X1 U5632 ( .A1(n8728), .A2(n5009), .ZN(n8715) );
  NOR2_X1 U5633 ( .A1(n8777), .A2(n4671), .ZN(n8728) );
  NOR3_X1 U5634 ( .A1(n8777), .A2(n8882), .A3(n8888), .ZN(n8743) );
  OR2_X1 U5635 ( .A1(n8776), .A2(n8897), .ZN(n8777) );
  NOR2_X1 U5636 ( .A1(n8777), .A2(n8888), .ZN(n8768) );
  NOR2_X1 U5637 ( .A1(n4482), .A2(n4639), .ZN(n4638) );
  INV_X1 U5638 ( .A(n4642), .ZN(n4639) );
  AND2_X1 U5639 ( .A1(n7772), .A2(n7773), .ZN(n8796) );
  AND2_X1 U5640 ( .A1(n7983), .A2(n7982), .ZN(n7980) );
  INV_X1 U5641 ( .A(n7980), .ZN(n7884) );
  OR2_X1 U5642 ( .A1(n6008), .A2(n7327), .ZN(n6022) );
  INV_X1 U5643 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U5644 ( .A1(n7571), .A2(n9578), .ZN(n7590) );
  OR2_X1 U5645 ( .A1(n7590), .A2(n7628), .ZN(n7635) );
  OAI211_X1 U5646 ( .C1(n4745), .C2(n4743), .A(n4742), .B(n7579), .ZN(n7631)
         );
  NAND2_X1 U5647 ( .A1(n7477), .A2(n4514), .ZN(n4744) );
  NOR2_X1 U5648 ( .A1(n7521), .A2(n10012), .ZN(n7523) );
  AND2_X1 U5649 ( .A1(n7968), .A2(n7967), .ZN(n7881) );
  NAND2_X1 U5650 ( .A1(n7878), .A2(n4491), .ZN(n5003) );
  OR2_X1 U5651 ( .A1(n7386), .A2(n10004), .ZN(n7521) );
  NAND2_X1 U5652 ( .A1(n7379), .A2(n7378), .ZN(n7486) );
  NAND2_X1 U5653 ( .A1(n7351), .A2(n9998), .ZN(n7386) );
  INV_X1 U5654 ( .A(n7278), .ZN(n7271) );
  NAND2_X1 U5655 ( .A1(n7274), .A2(n7950), .ZN(n7356) );
  NOR2_X1 U5656 ( .A1(n7150), .A2(n5023), .ZN(n7349) );
  AND2_X1 U5657 ( .A1(n7349), .A2(n9992), .ZN(n7351) );
  OR2_X1 U5658 ( .A1(n7149), .A2(n7155), .ZN(n7150) );
  NAND2_X1 U5659 ( .A1(n4667), .A2(n9967), .ZN(n6969) );
  AND4_X1 U5660 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n6964)
         );
  NAND2_X1 U5661 ( .A1(n6823), .A2(n6822), .ZN(n6926) );
  AND4_X1 U5662 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(n6892)
         );
  INV_X1 U5663 ( .A(n7869), .ZN(n6902) );
  INV_X1 U5664 ( .A(n5038), .ZN(n7870) );
  NAND2_X1 U5665 ( .A1(n7839), .A2(n7838), .ZN(n8837) );
  NAND2_X1 U5666 ( .A1(n6199), .A2(n6198), .ZN(n8847) );
  NAND2_X1 U5667 ( .A1(n6178), .A2(n6177), .ZN(n8858) );
  NAND2_X1 U5668 ( .A1(n6142), .A2(n6141), .ZN(n8877) );
  OR2_X1 U5669 ( .A1(n6252), .A2(n7868), .ZN(n10024) );
  NOR2_X1 U5670 ( .A1(n6896), .A2(n4668), .ZN(n6970) );
  NAND2_X1 U5671 ( .A1(n9967), .A2(n7070), .ZN(n4668) );
  INV_X1 U5672 ( .A(n6978), .ZN(n6981) );
  NOR2_X1 U5673 ( .A1(n6977), .A2(n6976), .ZN(n6982) );
  INV_X1 U5674 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U5675 ( .A1(n4954), .A2(n5793), .ZN(n4953) );
  INV_X1 U5676 ( .A(n4955), .ZN(n4954) );
  OR3_X1 U5677 ( .A1(n5989), .A2(P2_IR_REG_11__SCAN_IN), .A3(n5988), .ZN(n6005) );
  INV_X1 U5678 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U5679 ( .A1(n7856), .A2(n5082), .ZN(n5817) );
  INV_X1 U5680 ( .A(n9058), .ZN(n4874) );
  NAND2_X1 U5681 ( .A1(n6463), .A2(n9037), .ZN(n4869) );
  OAI21_X1 U5682 ( .B1(n4852), .B2(n4684), .A(n4682), .ZN(n6463) );
  NAND2_X1 U5683 ( .A1(n4869), .A2(n6468), .ZN(n8966) );
  AOI21_X1 U5684 ( .B1(n4547), .B2(n9046), .A(n4861), .ZN(n4860) );
  AND2_X1 U5685 ( .A1(n4862), .A2(n9047), .ZN(n4861) );
  NOR2_X1 U5686 ( .A1(n9047), .A2(n9046), .ZN(n4863) );
  AOI21_X1 U5687 ( .B1(n4692), .B2(n4690), .A(n4689), .ZN(n4688) );
  INV_X1 U5688 ( .A(n6487), .ZN(n4689) );
  INV_X1 U5689 ( .A(n8990), .ZN(n4690) );
  INV_X1 U5690 ( .A(n4692), .ZN(n4691) );
  NAND2_X1 U5691 ( .A1(n5281), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5692 ( .A1(n5315), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4697) );
  INV_X1 U5693 ( .A(n9001), .ZN(n6416) );
  INV_X1 U5694 ( .A(n5508), .ZN(n5233) );
  NAND2_X1 U5695 ( .A1(n9004), .A2(n8999), .ZN(n9013) );
  AND2_X1 U5696 ( .A1(n6349), .A2(n7409), .ZN(n7436) );
  AND2_X1 U5697 ( .A1(n6282), .A2(n4677), .ZN(n6590) );
  NAND2_X1 U5698 ( .A1(n5235), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U5699 ( .A1(n9012), .A2(n4860), .ZN(n4675) );
  AOI21_X1 U5700 ( .B1(n4860), .B2(n4863), .A(n4859), .ZN(n4858) );
  INV_X1 U5701 ( .A(n8974), .ZN(n4859) );
  NAND2_X1 U5702 ( .A1(n7620), .A2(n7621), .ZN(n7619) );
  OR2_X1 U5703 ( .A1(n5410), .A2(n7495), .ZN(n5425) );
  OR2_X1 U5704 ( .A1(n6298), .A2(n6297), .ZN(n6302) );
  NAND2_X1 U5705 ( .A1(n9013), .A2(n9014), .ZN(n9012) );
  AND2_X1 U5706 ( .A1(n9058), .A2(n4524), .ZN(n4692) );
  INV_X1 U5707 ( .A(n4883), .ZN(n4882) );
  OAI21_X1 U5708 ( .B1(n8954), .B2(n6405), .A(n6409), .ZN(n9069) );
  OR4_X1 U5709 ( .A1(n8242), .A2(n8374), .A3(n8241), .A4(n8240), .ZN(n8244) );
  INV_X1 U5710 ( .A(n5511), .ZN(n5285) );
  NOR2_X1 U5711 ( .A1(n6864), .A2(n6865), .ZN(n6863) );
  NAND2_X1 U5712 ( .A1(n9661), .A2(n4790), .ZN(n9675) );
  NAND2_X1 U5713 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  NOR2_X1 U5714 ( .A1(n9693), .A2(n4800), .ZN(n9116) );
  AND2_X1 U5715 ( .A1(n6637), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4800) );
  NAND2_X1 U5716 ( .A1(n9116), .A2(n9115), .ZN(n9114) );
  NOR2_X1 U5717 ( .A1(n9702), .A2(n4802), .ZN(n9717) );
  AND2_X1 U5718 ( .A1(n9707), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4802) );
  NOR2_X1 U5719 ( .A1(n9717), .A2(n9716), .ZN(n9714) );
  NOR2_X1 U5720 ( .A1(n9714), .A2(n4801), .ZN(n6843) );
  AND2_X1 U5721 ( .A1(n6850), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4801) );
  NAND2_X1 U5722 ( .A1(n6843), .A2(n6842), .ZN(n6996) );
  NAND2_X1 U5723 ( .A1(n5691), .A2(n5690), .ZN(n9136) );
  AND2_X1 U5724 ( .A1(n5266), .A2(n5265), .ZN(n9182) );
  OAI21_X1 U5725 ( .B1(n9214), .B2(n9215), .A(n8311), .ZN(n9195) );
  AND2_X1 U5726 ( .A1(n8310), .A2(n8316), .ZN(n9194) );
  NAND2_X1 U5727 ( .A1(n9195), .A2(n9194), .ZN(n9193) );
  AND2_X1 U5728 ( .A1(n5680), .A2(n5679), .ZN(n9199) );
  NAND2_X1 U5729 ( .A1(n9280), .A2(n4709), .ZN(n9209) );
  NOR2_X1 U5730 ( .A1(n9394), .A2(n4710), .ZN(n4709) );
  INV_X1 U5731 ( .A(n4711), .ZN(n4710) );
  NAND2_X1 U5732 ( .A1(n9280), .A2(n4713), .ZN(n9245) );
  NAND2_X1 U5733 ( .A1(n4824), .A2(n4822), .ZN(n9241) );
  INV_X1 U5734 ( .A(n4823), .ZN(n4822) );
  AND2_X1 U5735 ( .A1(n8303), .A2(n8210), .ZN(n9257) );
  NAND2_X1 U5736 ( .A1(n9288), .A2(n5712), .ZN(n9271) );
  AND2_X1 U5737 ( .A1(n5595), .A2(n5594), .ZN(n9293) );
  AND2_X1 U5738 ( .A1(n9270), .A2(n8153), .ZN(n9289) );
  NAND2_X1 U5739 ( .A1(n9290), .A2(n9289), .ZN(n9288) );
  NAND2_X1 U5740 ( .A1(n4819), .A2(n4818), .ZN(n9303) );
  INV_X1 U5741 ( .A(n4816), .ZN(n4818) );
  OAI21_X1 U5742 ( .B1(n9317), .B2(n4817), .A(n8253), .ZN(n4816) );
  AND2_X1 U5743 ( .A1(n9592), .A2(n4556), .ZN(n9333) );
  NAND2_X1 U5744 ( .A1(n9592), .A2(n4707), .ZN(n9357) );
  NAND2_X1 U5745 ( .A1(n9592), .A2(n9533), .ZN(n7661) );
  OR2_X1 U5746 ( .A1(n9617), .A2(n7618), .ZN(n9593) );
  INV_X1 U5747 ( .A(n8227), .ZN(n5449) );
  NAND2_X1 U5748 ( .A1(n5230), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5441) );
  INV_X1 U5749 ( .A(n5425), .ZN(n5230) );
  OR2_X1 U5750 ( .A1(n9616), .A2(n9634), .ZN(n9617) );
  NOR2_X1 U5751 ( .A1(n5387), .A2(n5701), .ZN(n5702) );
  AND2_X1 U5752 ( .A1(n5349), .A2(n5348), .ZN(n7209) );
  NOR2_X1 U5753 ( .A1(n9779), .A2(n4962), .ZN(n4961) );
  NAND2_X1 U5754 ( .A1(n8110), .A2(n8287), .ZN(n9778) );
  NOR2_X1 U5755 ( .A1(n7295), .A2(n9847), .ZN(n9776) );
  AND2_X1 U5756 ( .A1(n9776), .A2(n9860), .ZN(n9774) );
  INV_X1 U5757 ( .A(n8213), .ZN(n4967) );
  NOR2_X1 U5758 ( .A1(n8333), .A2(n7012), .ZN(n9793) );
  NAND2_X1 U5759 ( .A1(n9806), .A2(n9807), .ZN(n9805) );
  NOR2_X1 U5760 ( .A1(n9804), .A2(n9796), .ZN(n9806) );
  INV_X1 U5761 ( .A(n9882), .ZN(n9808) );
  OR2_X1 U5762 ( .A1(n7010), .A2(n7009), .ZN(n9800) );
  NAND2_X1 U5763 ( .A1(n5655), .A2(n5654), .ZN(n9201) );
  AND4_X1 U5764 ( .A1(n5370), .A2(n5369), .A3(n5368), .A4(n5367), .ZN(n9887)
         );
  NAND2_X2 U5765 ( .A1(n5378), .A2(n5377), .ZN(n9893) );
  OR2_X1 U5766 ( .A1(n8245), .A2(n6872), .ZN(n9888) );
  NOR2_X1 U5767 ( .A1(n5757), .A2(n7239), .ZN(n7008) );
  XNOR2_X1 U5768 ( .A(n7837), .B(n5206), .ZN(n7830) );
  OAI21_X1 U5769 ( .B1(n5669), .B2(n4838), .A(n4836), .ZN(n7837) );
  XNOR2_X1 U5770 ( .A(n4764), .B(n5256), .ZN(n8941) );
  NAND2_X1 U5771 ( .A1(n5669), .A2(n5201), .ZN(n4764) );
  XNOR2_X1 U5772 ( .A(n5736), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5773 ( .A1(n5735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5736) );
  XNOR2_X1 U5774 ( .A(n5653), .B(n5652), .ZN(n7749) );
  NAND2_X1 U5775 ( .A1(n4769), .A2(n4772), .ZN(n5653) );
  NAND2_X1 U5776 ( .A1(n5626), .A2(n4774), .ZN(n4769) );
  NAND2_X1 U5777 ( .A1(n5729), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U5778 ( .A1(n5731), .A2(n5730), .ZN(n5735) );
  OAI21_X1 U5779 ( .B1(n5626), .B2(n5184), .A(n5183), .ZN(n5640) );
  XNOR2_X1 U5780 ( .A(n4890), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U5781 ( .A1(n4891), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4890) );
  XNOR2_X1 U5782 ( .A(n5755), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U5783 ( .A1(n5727), .A2(n5076), .ZN(n5754) );
  INV_X1 U5784 ( .A(n5724), .ZN(n5727) );
  XNOR2_X1 U5785 ( .A(n5689), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8376) );
  NAND2_X1 U5786 ( .A1(n5132), .A2(n5131), .ZN(n5465) );
  AND2_X1 U5787 ( .A1(n5437), .A2(n5453), .ZN(n7139) );
  NAND2_X1 U5788 ( .A1(n4839), .A2(n4840), .ZN(n5432) );
  NAND2_X1 U5789 ( .A1(n4779), .A2(n4843), .ZN(n4839) );
  INV_X1 U5790 ( .A(n5403), .ZN(n4779) );
  XNOR2_X1 U5791 ( .A(n5403), .B(n5074), .ZN(n6572) );
  NAND2_X1 U5792 ( .A1(n5001), .A2(n5097), .ZN(n5334) );
  NAND2_X1 U5793 ( .A1(n5318), .A2(n5095), .ZN(n5001) );
  AND3_X1 U5794 ( .A1(n5035), .A2(n5034), .A3(SI_0_), .ZN(n5291) );
  XNOR2_X1 U5795 ( .A(n6241), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6554) );
  AND2_X1 U5796 ( .A1(n8511), .A2(n8545), .ZN(n5022) );
  NAND2_X1 U5797 ( .A1(n7075), .A2(n5907), .ZN(n7251) );
  NAND2_X1 U5798 ( .A1(n4933), .A2(n6016), .ZN(n7604) );
  XNOR2_X1 U5799 ( .A(n6159), .B(n6158), .ZN(n8483) );
  NAND2_X1 U5800 ( .A1(n4657), .A2(n6099), .ZN(n8453) );
  OR2_X1 U5801 ( .A1(n5847), .A2(n6530), .ZN(n5830) );
  OR2_X1 U5802 ( .A1(n6100), .A2(n5829), .ZN(n5831) );
  NAND2_X1 U5803 ( .A1(n7308), .A2(n5820), .ZN(n6912) );
  AND2_X1 U5804 ( .A1(n6052), .A2(n6051), .ZN(n7748) );
  AND3_X1 U5805 ( .A1(n6080), .A2(n6079), .A3(n6078), .ZN(n7781) );
  AND4_X1 U5806 ( .A1(n6044), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(n7743)
         );
  INV_X1 U5807 ( .A(n8510), .ZN(n8500) );
  NAND2_X1 U5808 ( .A1(n7739), .A2(n6065), .ZN(n7753) );
  NAND2_X1 U5809 ( .A1(n8444), .A2(n5859), .ZN(n7065) );
  NAND2_X1 U5810 ( .A1(n4945), .A2(n4943), .ZN(n7791) );
  INV_X1 U5811 ( .A(n4944), .ZN(n4943) );
  NAND2_X1 U5812 ( .A1(n7187), .A2(n4946), .ZN(n4945) );
  NAND2_X1 U5813 ( .A1(n6090), .A2(n6089), .ZN(n8901) );
  NOR2_X1 U5814 ( .A1(n8524), .A2(n8764), .ZN(n8510) );
  NAND2_X1 U5815 ( .A1(n5890), .A2(n5889), .ZN(n7077) );
  INV_X1 U5816 ( .A(n8505), .ZN(n8517) );
  XNOR2_X1 U5817 ( .A(n6047), .B(n6045), .ZN(n7708) );
  AND2_X1 U5818 ( .A1(n6270), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8526) );
  NAND2_X1 U5819 ( .A1(n6040), .A2(n6039), .ZN(n7721) );
  INV_X1 U5820 ( .A(n8529), .ZN(n8492) );
  INV_X1 U5821 ( .A(n6964), .ZN(n8548) );
  INV_X1 U5822 ( .A(n4720), .ZN(n6746) );
  INV_X1 U5823 ( .A(n4718), .ZN(n6766) );
  NOR2_X1 U5824 ( .A1(n6787), .A2(n4727), .ZN(n6716) );
  AND2_X1 U5825 ( .A1(n6718), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4727) );
  NOR2_X1 U5826 ( .A1(n6716), .A2(n6715), .ZN(n6946) );
  AND2_X1 U5827 ( .A1(n6669), .A2(n6668), .ZN(n8611) );
  INV_X1 U5828 ( .A(n9935), .ZN(n9930) );
  NAND2_X1 U5829 ( .A1(n7860), .A2(n7859), .ZN(n8834) );
  INV_X1 U5830 ( .A(n8837), .ZN(n8625) );
  INV_X1 U5831 ( .A(n8847), .ZN(n8640) );
  AOI211_X1 U5832 ( .C1(n8810), .C2(n8634), .A(n8633), .B(n8632), .ZN(n8850)
         );
  NAND2_X1 U5833 ( .A1(n4753), .A2(n5029), .ZN(n8631) );
  NAND2_X1 U5834 ( .A1(n8682), .A2(n8401), .ZN(n8666) );
  OAI21_X1 U5835 ( .B1(n5042), .B2(n4626), .A(n4624), .ZN(n8664) );
  NAND2_X1 U5836 ( .A1(n5040), .A2(n5043), .ZN(n8684) );
  OR2_X1 U5837 ( .A1(n8714), .A2(n5045), .ZN(n5040) );
  AND2_X1 U5838 ( .A1(n8709), .A2(n8708), .ZN(n8870) );
  NAND2_X1 U5839 ( .A1(n8713), .A2(n5048), .ZN(n8698) );
  NAND2_X1 U5840 ( .A1(n8748), .A2(n8006), .ZN(n8735) );
  INV_X1 U5841 ( .A(n8877), .ZN(n8732) );
  AND2_X1 U5842 ( .A1(n4747), .A2(n4750), .ZN(n8750) );
  NAND2_X1 U5843 ( .A1(n4627), .A2(n4634), .ZN(n8742) );
  OR2_X1 U5844 ( .A1(n8775), .A2(n4636), .ZN(n4627) );
  NAND2_X1 U5845 ( .A1(n4640), .A2(n4642), .ZN(n8772) );
  NOR2_X1 U5846 ( .A1(n8781), .A2(n4752), .ZN(n8761) );
  NAND2_X1 U5847 ( .A1(n8397), .A2(n8396), .ZN(n8795) );
  NAND2_X1 U5848 ( .A1(n6072), .A2(n6071), .ZN(n8907) );
  NAND2_X1 U5849 ( .A1(n7761), .A2(n7986), .ZN(n7825) );
  INV_X1 U5850 ( .A(n7748), .ZN(n8912) );
  AND2_X1 U5851 ( .A1(n7588), .A2(n7587), .ZN(n7589) );
  NAND2_X1 U5852 ( .A1(n7560), .A2(n7559), .ZN(n7561) );
  AND2_X1 U5853 ( .A1(n5974), .A2(n5973), .ZN(n7483) );
  NAND2_X1 U5854 ( .A1(n5005), .A2(n7908), .ZN(n7514) );
  NAND2_X1 U5855 ( .A1(n7487), .A2(n7879), .ZN(n7519) );
  NAND2_X1 U5856 ( .A1(n5053), .A2(n7484), .ZN(n7487) );
  AND2_X1 U5857 ( .A1(n5056), .A2(n5057), .ZN(n7348) );
  NOR2_X1 U5858 ( .A1(n8422), .A2(n5019), .ZN(n5018) );
  NAND2_X1 U5859 ( .A1(n7107), .A2(n7106), .ZN(n7156) );
  OAI211_X1 U5860 ( .C1(n6525), .C2(n5847), .A(n4665), .B(n4664), .ZN(n6941)
         );
  NAND2_X1 U5861 ( .A1(n5860), .A2(n4493), .ZN(n4665) );
  OR2_X1 U5862 ( .A1(n5860), .A2(n4741), .ZN(n4664) );
  INV_X1 U5863 ( .A(n8818), .ZN(n8826) );
  NAND2_X1 U5864 ( .A1(n8696), .A2(n6816), .ZN(n8823) );
  NAND2_X1 U5865 ( .A1(n9943), .A2(n6243), .ZN(n8821) );
  INV_X1 U5866 ( .A(n8823), .ZN(n8620) );
  AND2_X2 U5867 ( .A1(n6982), .A2(n6978), .ZN(n10052) );
  NAND2_X1 U5868 ( .A1(n8843), .A2(n8844), .ZN(n5069) );
  NAND2_X1 U5869 ( .A1(n8642), .A2(n4616), .ZN(n4615) );
  AND2_X1 U5870 ( .A1(n4611), .A2(n4614), .ZN(n4610) );
  OR2_X1 U5871 ( .A1(n8642), .A2(n4617), .ZN(n4611) );
  NOR2_X1 U5872 ( .A1(n9987), .A2(n5016), .ZN(n9988) );
  NAND2_X1 U5873 ( .A1(n5019), .A2(n5017), .ZN(n5016) );
  NOR2_X1 U5874 ( .A1(n6554), .A2(P2_U3152), .ZN(n9948) );
  OR2_X1 U5875 ( .A1(n5773), .A2(n5771), .ZN(n5772) );
  AND2_X1 U5876 ( .A1(n8932), .A2(n5775), .ZN(n8938) );
  XNOR2_X1 U5877 ( .A(n6222), .B(n6221), .ZN(n7615) );
  NAND2_X1 U5878 ( .A1(n6220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6222) );
  INV_X1 U5879 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7788) );
  INV_X1 U5880 ( .A(n6255), .ZN(n7505) );
  INV_X1 U5881 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7448) );
  XNOR2_X1 U5882 ( .A(n5791), .B(n5790), .ZN(n8061) );
  INV_X1 U5883 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5790) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7316) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7130) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7045) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6839) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6802) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6574) );
  INV_X1 U5890 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6561) );
  INV_X1 U5891 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6546) );
  INV_X1 U5892 ( .A(n5826), .ZN(n5827) );
  AND4_X1 U5893 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n9875)
         );
  NAND2_X1 U5894 ( .A1(n4694), .A2(n4886), .ZN(n8954) );
  NAND2_X1 U5895 ( .A1(n7619), .A2(n4508), .ZN(n4694) );
  NAND2_X1 U5896 ( .A1(n4865), .A2(n4868), .ZN(n8968) );
  INV_X1 U5897 ( .A(n4869), .ZN(n4865) );
  OAI21_X1 U5898 ( .B1(n9012), .B2(n4863), .A(n4860), .ZN(n8975) );
  NAND2_X1 U5899 ( .A1(n4854), .A2(n6450), .ZN(n8982) );
  NAND2_X1 U5900 ( .A1(n9030), .A2(n9029), .ZN(n4854) );
  OAI21_X1 U5901 ( .B1(n6471), .B2(n6470), .A(n9021), .ZN(n8989) );
  INV_X1 U5902 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9016) );
  AND4_X1 U5903 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n9762)
         );
  NAND2_X1 U5904 ( .A1(n5574), .A2(n5573), .ZN(n9295) );
  NAND2_X1 U5905 ( .A1(n7619), .A2(n6384), .ZN(n7670) );
  INV_X1 U5906 ( .A(n4681), .ZN(n9036) );
  AOI21_X1 U5907 ( .B1(n4852), .B2(n4853), .A(n4684), .ZN(n4681) );
  NAND2_X1 U5908 ( .A1(n4887), .A2(n7491), .ZN(n7543) );
  NAND2_X1 U5909 ( .A1(n6293), .A2(n6292), .ZN(n6294) );
  NAND2_X1 U5910 ( .A1(n9012), .A2(n6429), .ZN(n9049) );
  NAND2_X1 U5911 ( .A1(n6326), .A2(n6325), .ZN(n7236) );
  NAND2_X1 U5912 ( .A1(n7020), .A2(n4533), .ZN(n6326) );
  NAND2_X1 U5913 ( .A1(n6507), .A2(n7237), .ZN(n9076) );
  NAND2_X1 U5914 ( .A1(n4693), .A2(n4692), .ZN(n9057) );
  AND2_X1 U5915 ( .A1(n6512), .A2(n6502), .ZN(n9056) );
  AND4_X1 U5916 ( .A1(n5516), .A2(n5515), .A3(n5514), .A4(n5513), .ZN(n9080)
         );
  NAND2_X1 U5917 ( .A1(n5491), .A2(n5490), .ZN(n9083) );
  INV_X1 U5918 ( .A(n9067), .ZN(n9082) );
  INV_X1 U5919 ( .A(n9056), .ZN(n9085) );
  NAND2_X1 U5920 ( .A1(n4587), .A2(n4507), .ZN(n8246) );
  OR2_X1 U5921 ( .A1(n8204), .A2(n8203), .ZN(n4587) );
  OR2_X1 U5922 ( .A1(n8202), .A2(n8201), .ZN(n8373) );
  INV_X1 U5923 ( .A(n9199), .ZN(n9164) );
  NAND2_X1 U5924 ( .A1(n5664), .A2(n5663), .ZN(n9216) );
  NAND2_X1 U5925 ( .A1(n5637), .A2(n5636), .ZN(n9242) );
  OR2_X1 U5926 ( .A1(n9229), .A2(n5659), .ZN(n5637) );
  NAND2_X1 U5927 ( .A1(n5623), .A2(n5622), .ZN(n9413) );
  INV_X1 U5928 ( .A(n9293), .ZN(n9412) );
  INV_X1 U5929 ( .A(n9887), .ZN(n9864) );
  INV_X1 U5930 ( .A(n9848), .ZN(n9865) );
  INV_X1 U5931 ( .A(n8334), .ZN(n9096) );
  INV_X1 U5932 ( .A(n4794), .ZN(n9554) );
  NAND2_X1 U5933 ( .A1(n9663), .A2(n9662), .ZN(n9661) );
  AND2_X1 U5934 ( .A1(n4794), .A2(n4793), .ZN(n9663) );
  NAND2_X1 U5935 ( .A1(n6634), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U5936 ( .A1(n6617), .A2(n6618), .ZN(n6840) );
  NAND2_X1 U5937 ( .A1(n9114), .A2(n4797), .ZN(n6617) );
  NAND2_X1 U5938 ( .A1(n4799), .A2(n4798), .ZN(n4797) );
  INV_X1 U5939 ( .A(n4796), .ZN(n7138) );
  INV_X1 U5940 ( .A(n7458), .ZN(n7457) );
  INV_X1 U5941 ( .A(n9735), .ZN(n9715) );
  INV_X1 U5942 ( .A(n4788), .ZN(n9731) );
  INV_X2 U5943 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n10486) );
  XNOR2_X1 U5944 ( .A(n4786), .B(n4785), .ZN(n8084) );
  INV_X1 U5945 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4785) );
  NAND2_X1 U5946 ( .A1(n4788), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U5947 ( .A1(n8077), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4787) );
  AND2_X1 U5948 ( .A1(n6624), .A2(n6623), .ZN(n9744) );
  NAND2_X1 U5949 ( .A1(n4782), .A2(n4781), .ZN(n4780) );
  AOI21_X1 U5950 ( .B1(n4978), .B2(n9178), .A(n4981), .ZN(n4781) );
  NAND2_X1 U5951 ( .A1(n4977), .A2(n4978), .ZN(n4782) );
  AND2_X1 U5952 ( .A1(n5650), .A2(n5649), .ZN(n9398) );
  OAI21_X1 U5953 ( .B1(n9258), .B2(n4492), .A(n5608), .ZN(n9238) );
  NAND2_X1 U5954 ( .A1(n4821), .A2(n8099), .ZN(n9316) );
  OR2_X1 U5955 ( .A1(n9340), .A2(n8251), .ZN(n4821) );
  NAND2_X1 U5956 ( .A1(n5543), .A2(n5542), .ZN(n9329) );
  NAND2_X1 U5957 ( .A1(n4991), .A2(n4988), .ZN(n7659) );
  INV_X1 U5958 ( .A(n9089), .ZN(n9474) );
  NAND2_X1 U5959 ( .A1(n4987), .A2(n4994), .ZN(n7598) );
  OR2_X1 U5960 ( .A1(n4995), .A2(n4516), .ZN(n4987) );
  NAND2_X1 U5961 ( .A1(n7336), .A2(n5417), .ZN(n9614) );
  INV_X1 U5962 ( .A(n9361), .ZN(n9755) );
  AND2_X1 U5963 ( .A1(n5558), .A2(n5724), .ZN(n9789) );
  INV_X1 U5964 ( .A(n5557), .ZN(n5554) );
  NAND2_X1 U5965 ( .A1(n4964), .A2(n5324), .ZN(n9773) );
  NAND2_X1 U5966 ( .A1(n5350), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U5967 ( .A1(n9816), .A2(n9785), .ZN(n9337) );
  AND2_X1 U5968 ( .A1(n8196), .A2(n8195), .ZN(n9482) );
  AND2_X1 U5969 ( .A1(n8192), .A2(n8191), .ZN(n9486) );
  OR2_X1 U5970 ( .A1(n9378), .A2(n9377), .ZN(n9379) );
  INV_X1 U5971 ( .A(n9201), .ZN(n9494) );
  INV_X1 U5972 ( .A(n9284), .ZN(n9508) );
  INV_X1 U5973 ( .A(n9083), .ZN(n9528) );
  INV_X1 U5974 ( .A(n5249), .ZN(n9538) );
  MUX2_X1 U5975 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5246), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5248) );
  NAND2_X1 U5976 ( .A1(n5735), .A2(n5732), .ZN(n7719) );
  OR2_X1 U5977 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  INV_X1 U5978 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U5979 ( .A1(n5688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5685) );
  INV_X1 U5980 ( .A(n8332), .ZN(n8243) );
  INV_X1 U5981 ( .A(n8376), .ZN(n7446) );
  INV_X1 U5982 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10432) );
  INV_X1 U5983 ( .A(n9789), .ZN(n9814) );
  INV_X1 U5984 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10360) );
  AND2_X1 U5985 ( .A1(n5473), .A2(n5503), .ZN(n7685) );
  INV_X1 U5986 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10387) );
  INV_X1 U5987 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10419) );
  INV_X1 U5988 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6559) );
  INV_X1 U5989 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U5990 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4803) );
  NOR2_X1 U5991 ( .A1(n10083), .A2(n10491), .ZN(n10109) );
  AOI21_X1 U5992 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10107), .ZN(n10106) );
  NOR2_X1 U5993 ( .A1(n10106), .A2(n10105), .ZN(n10104) );
  AOI21_X1 U5994 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10104), .ZN(n10103) );
  OAI21_X1 U5995 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10101), .ZN(n10099) );
  NAND2_X1 U5996 ( .A1(n7184), .A2(n5956), .ZN(n7160) );
  NAND2_X1 U5997 ( .A1(n4913), .A2(n4914), .ZN(n4912) );
  NAND2_X1 U5998 ( .A1(n7467), .A2(n6004), .ZN(n7508) );
  AND2_X1 U5999 ( .A1(n4732), .A2(n4733), .ZN(n4568) );
  OR2_X1 U6000 ( .A1(n4740), .A2(n8070), .ZN(n4569) );
  NAND2_X1 U6001 ( .A1(n4894), .A2(n4892), .ZN(P2_U3549) );
  OR2_X1 U6002 ( .A1(n10052), .A2(n4893), .ZN(n4892) );
  INV_X1 U6003 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4893) );
  OAI211_X1 U6004 ( .C1(n8845), .C2(n5070), .A(n5071), .B(n5068), .ZN(P2_U3517) );
  NAND2_X1 U6005 ( .A1(n10032), .A2(n10029), .ZN(n5070) );
  NAND2_X1 U6006 ( .A1(n10030), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6007 ( .A1(n5069), .A2(n10032), .ZN(n5068) );
  OAI21_X1 U6008 ( .B1(n9189), .B2(n9067), .A(n6515), .ZN(n6516) );
  INV_X1 U6009 ( .A(n4809), .ZN(n4808) );
  NAND2_X1 U6010 ( .A1(n4811), .A2(n9928), .ZN(n4810) );
  OAI22_X1 U6011 ( .A1(n5690), .A2(n9478), .B1(n9928), .B2(n9376), .ZN(n4809)
         );
  NAND2_X1 U6012 ( .A1(n9909), .A2(n5758), .ZN(n4783) );
  XNOR2_X1 U6013 ( .A(n6217), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6254) );
  AND2_X1 U6014 ( .A1(n4840), .A2(n4846), .ZN(n4489) );
  OR3_X1 U6015 ( .A1(n4488), .A2(n4515), .A3(n4953), .ZN(n4490) );
  AND2_X1 U6016 ( .A1(n4545), .A2(n7908), .ZN(n4491) );
  AND2_X1 U6017 ( .A1(n9267), .A2(n9421), .ZN(n4492) );
  NOR2_X1 U6018 ( .A1(n5122), .A2(n4844), .ZN(n4843) );
  XNOR2_X1 U6019 ( .A(n5099), .B(SI_5_), .ZN(n5333) );
  AND2_X1 U6020 ( .A1(n6521), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4493) );
  INV_X1 U6021 ( .A(n7824), .ZN(n7990) );
  INV_X1 U6022 ( .A(n8404), .ZN(n4617) );
  AOI21_X1 U6023 ( .B1(n9140), .B2(n8371), .A(n9482), .ZN(n8325) );
  INV_X1 U6024 ( .A(n8325), .ZN(n4582) );
  AND2_X1 U6025 ( .A1(n4963), .A2(n8216), .ZN(n4494) );
  AND2_X1 U6026 ( .A1(n5029), .A2(n8042), .ZN(n4495) );
  AND2_X1 U6027 ( .A1(n5690), .A2(n9486), .ZN(n4496) );
  AND2_X1 U6028 ( .A1(n4707), .A2(n4706), .ZN(n4497) );
  AND2_X1 U6029 ( .A1(n4739), .A2(n4737), .ZN(n4498) );
  NOR2_X1 U6030 ( .A1(n4868), .A2(n8965), .ZN(n4499) );
  AND2_X1 U6031 ( .A1(n7275), .A2(n7950), .ZN(n4500) );
  AND2_X1 U6032 ( .A1(n4898), .A2(n4897), .ZN(n4501) );
  INV_X1 U6033 ( .A(n6308), .ZN(n7806) );
  INV_X1 U6034 ( .A(n8872), .ZN(n5009) );
  AND2_X1 U6035 ( .A1(n5131), .A2(n5130), .ZN(n4502) );
  OR2_X1 U6036 ( .A1(n5484), .A2(n4760), .ZN(n4503) );
  NAND2_X1 U6037 ( .A1(n5341), .A2(n5340), .ZN(n9784) );
  INV_X1 U6038 ( .A(n7878), .ZN(n7485) );
  XNOR2_X1 U6039 ( .A(n8852), .B(n8630), .ZN(n8656) );
  INV_X1 U6040 ( .A(n8656), .ZN(n5032) );
  AND2_X1 U6041 ( .A1(n4722), .A2(n4721), .ZN(n4504) );
  AND2_X1 U6042 ( .A1(n8055), .A2(n8784), .ZN(n4505) );
  NOR2_X1 U6043 ( .A1(n8847), .A2(n8532), .ZN(n4506) );
  AND3_X1 U6044 ( .A1(n4583), .A2(n4580), .A3(n8373), .ZN(n4507) );
  NOR2_X1 U6045 ( .A1(n6389), .A2(n4885), .ZN(n4508) );
  NAND2_X1 U6046 ( .A1(n8888), .A2(n8751), .ZN(n4509) );
  AND2_X1 U6047 ( .A1(n4631), .A2(n4628), .ZN(n4510) );
  AND2_X1 U6048 ( .A1(n6660), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4511) );
  AND2_X1 U6049 ( .A1(n6521), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U6050 ( .A1(n7155), .A2(n8546), .ZN(n4513) );
  AND2_X1 U6051 ( .A1(n7968), .A2(n4491), .ZN(n4514) );
  OR2_X1 U6052 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4515) );
  NOR2_X1 U6053 ( .A1(n9637), .A2(n9089), .ZN(n4516) );
  OR2_X1 U6054 ( .A1(n9083), .A2(n9458), .ZN(n4517) );
  INV_X1 U6055 ( .A(n7337), .ZN(n4971) );
  AND2_X1 U6056 ( .A1(n8901), .A2(n8536), .ZN(n4518) );
  AND2_X1 U6057 ( .A1(n8966), .A2(n8965), .ZN(n4519) );
  OR3_X1 U6058 ( .A1(n4488), .A2(n4955), .A3(n4515), .ZN(n4520) );
  OR3_X1 U6059 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_1__SCAN_IN), .ZN(n4521) );
  OR3_X1 U6060 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4522) );
  AND2_X1 U6061 ( .A1(n4750), .A2(n8749), .ZN(n4523) );
  NAND2_X1 U6062 ( .A1(n6478), .A2(n6477), .ZN(n4524) );
  AND2_X1 U6063 ( .A1(n4718), .A2(n4717), .ZN(n4525) );
  NAND2_X1 U6064 ( .A1(n8858), .A2(n8657), .ZN(n8028) );
  AND2_X1 U6065 ( .A1(n7883), .A2(n7587), .ZN(n4526) );
  AND2_X1 U6066 ( .A1(n7234), .A2(n6333), .ZN(n4527) );
  NOR2_X1 U6067 ( .A1(n8654), .A2(n8038), .ZN(n4528) );
  NOR2_X1 U6068 ( .A1(n8155), .A2(n8161), .ZN(n4529) );
  INV_X1 U6069 ( .A(n9267), .ZN(n9504) );
  AND2_X1 U6070 ( .A1(n5923), .A2(n5922), .ZN(n4530) );
  AND2_X1 U6071 ( .A1(n8362), .A2(n8317), .ZN(n9178) );
  INV_X1 U6072 ( .A(n6429), .ZN(n4862) );
  AND2_X1 U6073 ( .A1(n7518), .A2(n7484), .ZN(n4531) );
  AND2_X1 U6074 ( .A1(n9409), .A2(n9413), .ZN(n4532) );
  AND2_X1 U6075 ( .A1(n6312), .A2(n6317), .ZN(n4533) );
  INV_X1 U6076 ( .A(n8962), .ZN(n9533) );
  NAND2_X1 U6077 ( .A1(n5475), .A2(n5474), .ZN(n8962) );
  NOR2_X1 U6078 ( .A1(n9161), .A2(n4979), .ZN(n4978) );
  NAND2_X1 U6079 ( .A1(n9280), .A2(n4711), .ZN(n4714) );
  OR2_X1 U6080 ( .A1(n9267), .A2(n5713), .ZN(n8303) );
  INV_X1 U6081 ( .A(n8303), .ZN(n4595) );
  AND2_X1 U6082 ( .A1(n5099), .A2(SI_5_), .ZN(n4534) );
  AND2_X1 U6083 ( .A1(n4703), .A2(n4702), .ZN(n5346) );
  INV_X1 U6084 ( .A(n4843), .ZN(n4842) );
  OR2_X1 U6085 ( .A1(n8847), .A2(n8658), .ZN(n8042) );
  NAND2_X1 U6086 ( .A1(n5527), .A2(n5526), .ZN(n9453) );
  INV_X1 U6087 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5771) );
  INV_X1 U6088 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5798) );
  AND2_X1 U6089 ( .A1(n6457), .A2(n6456), .ZN(n4535) );
  NOR2_X1 U6090 ( .A1(n4613), .A2(n10019), .ZN(n4536) );
  NOR2_X1 U6091 ( .A1(n7813), .A2(n7812), .ZN(n4537) );
  AND2_X1 U6092 ( .A1(n8882), .A2(n8535), .ZN(n4538) );
  INV_X1 U6093 ( .A(n4915), .ZN(n4913) );
  NAND2_X1 U6094 ( .A1(n4916), .A2(n6257), .ZN(n4915) );
  NOR2_X1 U6095 ( .A1(n8858), .A2(n8533), .ZN(n4539) );
  AND2_X1 U6096 ( .A1(n5121), .A2(SI_11_), .ZN(n4540) );
  NAND2_X1 U6097 ( .A1(n5013), .A2(n5011), .ZN(n4541) );
  NOR2_X1 U6098 ( .A1(n8867), .A2(n8723), .ZN(n4542) );
  OR2_X1 U6099 ( .A1(n8888), .A2(n8464), .ZN(n8003) );
  OR2_X1 U6100 ( .A1(n6912), .A2(n6936), .ZN(n4543) );
  AND2_X1 U6101 ( .A1(n6084), .A2(n6083), .ZN(n4544) );
  NAND2_X1 U6102 ( .A1(n7483), .A2(n8542), .ZN(n4545) );
  NOR2_X1 U6103 ( .A1(n8470), .A2(n8469), .ZN(n4546) );
  OR2_X1 U6104 ( .A1(n9047), .A2(n4862), .ZN(n4547) );
  INV_X1 U6105 ( .A(n4703), .ZN(n5319) );
  INV_X1 U6106 ( .A(n5069), .ZN(n4618) );
  NAND2_X1 U6107 ( .A1(n4746), .A2(n5002), .ZN(n4548) );
  NOR2_X1 U6108 ( .A1(n6166), .A2(n6165), .ZN(n4549) );
  NAND4_X1 U6109 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n8547)
         );
  OR2_X1 U6110 ( .A1(n5023), .A2(n5015), .ZN(n4550) );
  AND4_X1 U6111 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n7358)
         );
  INV_X1 U6112 ( .A(n7358), .ZN(n5015) );
  AND2_X1 U6113 ( .A1(n7266), .A2(n4513), .ZN(n4551) );
  AND2_X1 U6114 ( .A1(n5387), .A2(n5371), .ZN(n4552) );
  AND2_X1 U6115 ( .A1(n9161), .A2(n8186), .ZN(n4553) );
  AND2_X1 U6116 ( .A1(n6371), .A2(n7491), .ZN(n4554) );
  AND2_X1 U6117 ( .A1(n7976), .A2(n7974), .ZN(n4555) );
  INV_X1 U6118 ( .A(n4625), .ZN(n4624) );
  OAI21_X1 U6119 ( .B1(n5041), .B2(n4626), .A(n8665), .ZN(n4625) );
  AND2_X1 U6120 ( .A1(n4497), .A2(n9338), .ZN(n4556) );
  OR2_X1 U6121 ( .A1(n8877), .A2(n8534), .ZN(n8008) );
  NOR2_X1 U6122 ( .A1(n7605), .A2(n4932), .ZN(n4931) );
  AND2_X1 U6123 ( .A1(n4501), .A2(n4670), .ZN(n4557) );
  INV_X1 U6124 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6125 ( .A1(n5258), .A2(n5257), .ZN(n9167) );
  INV_X1 U6126 ( .A(n9167), .ZN(n4705) );
  NOR2_X1 U6127 ( .A1(n4488), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n6068) );
  INV_X1 U6128 ( .A(n6462), .ZN(n4684) );
  OAI22_X1 U6129 ( .A1(n8496), .A2(n8495), .B1(n6127), .B2(n6126), .ZN(n8461)
         );
  INV_X1 U6130 ( .A(n8864), .ZN(n4897) );
  OR2_X1 U6131 ( .A1(n9893), .A2(n9875), .ZN(n8255) );
  INV_X1 U6132 ( .A(n8255), .ZN(n4814) );
  NAND2_X1 U6133 ( .A1(n9592), .A2(n4497), .ZN(n4708) );
  AND2_X1 U6134 ( .A1(n4821), .A2(n4820), .ZN(n4558) );
  NAND2_X1 U6135 ( .A1(n4640), .A2(n4638), .ZN(n4641) );
  AND2_X1 U6136 ( .A1(n4774), .A2(n5652), .ZN(n4559) );
  NAND2_X1 U6137 ( .A1(n5226), .A2(n5225), .ZN(n8307) );
  INV_X1 U6138 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n4791) );
  INV_X1 U6139 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n4798) );
  INV_X1 U6140 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U6141 ( .A1(n5506), .A2(n5505), .ZN(n9364) );
  INV_X1 U6142 ( .A(n9364), .ZN(n4706) );
  AND4_X1 U6143 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n8736)
         );
  INV_X1 U6144 ( .A(n8736), .ZN(n5012) );
  INV_X1 U6145 ( .A(n8888), .ZN(n4673) );
  AND2_X1 U6146 ( .A1(n4933), .A2(n4931), .ZN(n4560) );
  AND2_X1 U6147 ( .A1(n5204), .A2(n5203), .ZN(n4561) );
  AND2_X1 U6148 ( .A1(n8289), .A2(n8108), .ZN(n9779) );
  AND2_X1 U6149 ( .A1(n5372), .A2(n5371), .ZN(n4562) );
  INV_X1 U6150 ( .A(n6252), .ZN(n4927) );
  AND2_X2 U6151 ( .A1(n6982), .A2(n6981), .ZN(n10032) );
  AND2_X2 U6152 ( .A1(n7008), .A2(n6585), .ZN(n9911) );
  NAND2_X1 U6153 ( .A1(n8386), .A2(n9789), .ZN(n8200) );
  AND2_X1 U6154 ( .A1(n7568), .A2(n9576), .ZN(n10019) );
  INV_X1 U6155 ( .A(n5294), .ZN(n6602) );
  AND2_X1 U6156 ( .A1(n8592), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4563) );
  INV_X1 U6157 ( .A(n4926), .ZN(n6936) );
  NAND2_X1 U6158 ( .A1(n4483), .A2(n7864), .ZN(n4926) );
  OR2_X1 U6159 ( .A1(n8607), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4564) );
  INV_X1 U6160 ( .A(n9671), .ZN(n4792) );
  INV_X1 U6161 ( .A(n6660), .ZN(n4741) );
  XNOR2_X1 U6162 ( .A(n5360), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9113) );
  INV_X1 U6163 ( .A(n9113), .ZN(n4799) );
  INV_X1 U6164 ( .A(n7892), .ZN(n8784) );
  XNOR2_X1 U6165 ( .A(n5796), .B(n5795), .ZN(n7892) );
  INV_X1 U6166 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4663) );
  OAI21_X1 U6167 ( .B1(n5520), .B2(n4847), .A(n5152), .ZN(n5538) );
  NAND2_X1 U6168 ( .A1(n5389), .A2(n5079), .ZN(n5115) );
  NAND2_X1 U6169 ( .A1(n5610), .A2(n5609), .ZN(n5612) );
  NAND2_X1 U6170 ( .A1(n8033), .A2(n4573), .ZN(n8043) );
  NAND2_X1 U6171 ( .A1(n4576), .A2(n8056), .ZN(n8062) );
  NAND2_X2 U6172 ( .A1(n9030), .A2(n4855), .ZN(n4852) );
  NAND2_X1 U6173 ( .A1(n7410), .A2(n7412), .ZN(n6349) );
  NAND3_X1 U6174 ( .A1(n6344), .A2(n6339), .A3(n6345), .ZN(n7410) );
  NAND2_X1 U6175 ( .A1(n6417), .A2(n6416), .ZN(n9004) );
  NAND2_X1 U6176 ( .A1(n4675), .A2(n4858), .ZN(n4674) );
  NAND2_X1 U6177 ( .A1(n7494), .A2(n7492), .ZN(n4887) );
  NAND2_X1 U6178 ( .A1(n6295), .A2(n6294), .ZN(n6686) );
  NAND3_X1 U6179 ( .A1(n8247), .A2(n8387), .A3(n4565), .ZN(n8393) );
  NAND2_X1 U6180 ( .A1(n4566), .A2(n8188), .ZN(n8199) );
  NAND2_X1 U6181 ( .A1(n8187), .A2(n4553), .ZN(n4566) );
  NAND2_X1 U6182 ( .A1(n5148), .A2(n5147), .ZN(n5520) );
  NAND2_X1 U6183 ( .A1(n5167), .A2(n5166), .ZN(n5586) );
  OAI21_X1 U6184 ( .B1(n5599), .B2(n5598), .A(n5175), .ZN(n5610) );
  NAND2_X1 U6185 ( .A1(n5344), .A2(n5100), .ZN(n4652) );
  NAND2_X1 U6186 ( .A1(n5083), .A2(n5817), .ZN(n5085) );
  XNOR2_X1 U6187 ( .A(n5085), .B(n5084), .ZN(n5280) );
  AOI21_X2 U6189 ( .B1(n8094), .B2(n8302), .A(n8093), .ZN(n8361) );
  NAND2_X1 U6190 ( .A1(n4567), .A2(n7979), .ZN(n7981) );
  NAND2_X1 U6191 ( .A1(n7975), .A2(n4555), .ZN(n4567) );
  NAND3_X1 U6192 ( .A1(n8007), .A2(n8010), .A3(n8006), .ZN(n8009) );
  NAND2_X1 U6193 ( .A1(n4569), .A2(n4568), .ZN(P2_U3244) );
  NAND3_X1 U6194 ( .A1(n7957), .A2(n7955), .A3(n7956), .ZN(n4570) );
  NAND3_X1 U6195 ( .A1(n7944), .A2(n7942), .A3(n7943), .ZN(n4572) );
  NAND4_X1 U6196 ( .A1(n4647), .A2(n5768), .A3(n5763), .A4(n5762), .ZN(n4575)
         );
  OAI21_X1 U6197 ( .B1(n8050), .B2(n4578), .A(n4577), .ZN(n4576) );
  NAND2_X1 U6198 ( .A1(n4997), .A2(n4999), .ZN(n5344) );
  NAND2_X1 U6199 ( .A1(n5572), .A2(n5571), .ZN(n5167) );
  NAND2_X1 U6200 ( .A1(n5156), .A2(n5155), .ZN(n5553) );
  NAND2_X1 U6201 ( .A1(n4757), .A2(n4755), .ZN(n5148) );
  NAND2_X1 U6202 ( .A1(n5597), .A2(n5596), .ZN(n9258) );
  NAND2_X1 U6203 ( .A1(n7397), .A2(n8218), .ZN(n5372) );
  AOI21_X2 U6204 ( .B1(n9750), .B2(n5402), .A(n5401), .ZN(n7338) );
  NAND2_X1 U6205 ( .A1(n4995), .A2(n4992), .ZN(n4991) );
  OAI21_X2 U6206 ( .B1(n9305), .B2(n5570), .A(n5569), .ZN(n9287) );
  NAND2_X1 U6207 ( .A1(n5518), .A2(n5517), .ZN(n9332) );
  NAND2_X1 U6208 ( .A1(n7532), .A2(n5451), .ZN(n9591) );
  NAND2_X1 U6209 ( .A1(n4810), .A2(n4808), .ZN(P1_U3552) );
  NAND2_X1 U6210 ( .A1(n9208), .A2(n9215), .ZN(n4957) );
  NAND2_X1 U6211 ( .A1(n4579), .A2(n5086), .ZN(n5274) );
  NAND2_X1 U6212 ( .A1(n5279), .A2(n5280), .ZN(n4579) );
  INV_X1 U6213 ( .A(n9591), .ZN(n4995) );
  NAND2_X1 U6214 ( .A1(n4991), .A2(n4986), .ZN(n5500) );
  OAI22_X1 U6215 ( .A1(n9225), .A2(n5638), .B1(n9228), .B2(n9242), .ZN(n9208)
         );
  NAND2_X1 U6216 ( .A1(n5450), .A2(n5449), .ZN(n7532) );
  NOR2_X2 U6217 ( .A1(n9159), .A2(n9158), .ZN(n9380) );
  NAND2_X1 U6218 ( .A1(n4980), .A2(n5683), .ZN(n9157) );
  NAND2_X1 U6219 ( .A1(n4581), .A2(n8198), .ZN(n4580) );
  OAI21_X1 U6220 ( .B1(n4586), .B2(n8306), .A(n4582), .ZN(n4581) );
  NAND2_X1 U6221 ( .A1(n4584), .A2(n8200), .ZN(n4583) );
  NAND2_X1 U6222 ( .A1(n8324), .A2(n8207), .ZN(n4585) );
  NAND3_X1 U6223 ( .A1(n4601), .A2(n4599), .A3(n4598), .ZN(n8137) );
  AND2_X2 U6224 ( .A1(n4700), .A2(n4696), .ZN(n5557) );
  AND2_X2 U6225 ( .A1(n4702), .A2(n4703), .ZN(n4696) );
  XNOR2_X1 U6226 ( .A(n5292), .B(n8333), .ZN(n9807) );
  OAI211_X1 U6227 ( .C1(n4612), .C2(n8642), .A(n4608), .B(n4605), .ZN(n4894)
         );
  NAND2_X1 U6228 ( .A1(n4615), .A2(n4610), .ZN(n8845) );
  NAND2_X1 U6229 ( .A1(n4621), .A2(n6965), .ZN(n7105) );
  NAND2_X1 U6230 ( .A1(n4621), .A2(n4620), .ZN(n7106) );
  INV_X1 U6231 ( .A(n5042), .ZN(n4622) );
  OAI21_X1 U6232 ( .B1(n4622), .B2(n4625), .A(n4623), .ZN(n8648) );
  NAND2_X1 U6233 ( .A1(n8775), .A2(n4632), .ZN(n4631) );
  INV_X1 U6234 ( .A(n4641), .ZN(n8893) );
  NAND2_X1 U6235 ( .A1(n7917), .A2(n7923), .ZN(n7873) );
  NAND3_X1 U6236 ( .A1(n5763), .A2(n5762), .A3(n5061), .ZN(n4644) );
  NAND2_X1 U6237 ( .A1(n5762), .A2(n5763), .ZN(n4645) );
  NAND2_X1 U6238 ( .A1(n5768), .A2(n4647), .ZN(n4646) );
  AND2_X1 U6239 ( .A1(n5826), .A2(n4904), .ZN(n5876) );
  INV_X1 U6240 ( .A(n4648), .ZN(n4649) );
  NAND2_X1 U6241 ( .A1(n4657), .A2(n4656), .ZN(n8450) );
  NAND2_X2 U6242 ( .A1(n4658), .A2(n5961), .ZN(n10004) );
  NAND2_X1 U6243 ( .A1(n4928), .A2(n4659), .ZN(n6047) );
  NAND3_X1 U6244 ( .A1(n4931), .A2(n7469), .A3(n7468), .ZN(n4659) );
  INV_X2 U6245 ( .A(n7856), .ZN(n6521) );
  NAND3_X1 U6246 ( .A1(n5035), .A2(n5034), .A3(P2_DATAO_REG_5__SCAN_IN), .ZN(
        n4660) );
  NAND2_X2 U6247 ( .A1(n5033), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5034) );
  NAND2_X2 U6248 ( .A1(n5037), .A2(n5036), .ZN(n5035) );
  INV_X1 U6249 ( .A(n6896), .ZN(n4667) );
  NAND2_X1 U6250 ( .A1(n4667), .A2(n4666), .ZN(n7149) );
  INV_X1 U6251 ( .A(n8777), .ZN(n4669) );
  NAND2_X1 U6252 ( .A1(n4557), .A2(n4669), .ZN(n4899) );
  NAND2_X2 U6253 ( .A1(n4674), .A2(n6442), .ZN(n9030) );
  INV_X1 U6254 ( .A(n7801), .ZN(n6318) );
  NAND3_X1 U6255 ( .A1(n6284), .A2(n6285), .A3(n4676), .ZN(n6589) );
  NAND2_X1 U6256 ( .A1(n7801), .A2(n7012), .ZN(n4676) );
  NAND2_X1 U6257 ( .A1(n6482), .A2(n9804), .ZN(n4677) );
  AND2_X4 U6258 ( .A1(n7801), .A2(n6277), .ZN(n6482) );
  OR2_X2 U6259 ( .A1(n7022), .A2(n7023), .ZN(n7020) );
  INV_X1 U6260 ( .A(n4852), .ZN(n4678) );
  OAI21_X1 U6261 ( .B1(n4678), .B2(n4680), .A(n4679), .ZN(n4864) );
  NAND2_X1 U6262 ( .A1(n8989), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U6263 ( .A1(n4695), .A2(n4696), .ZN(n5724) );
  NAND3_X1 U6264 ( .A1(n4698), .A2(n5283), .A3(n4697), .ZN(n8333) );
  AND2_X2 U6265 ( .A1(n5488), .A2(n7856), .ZN(n5315) );
  NOR2_X2 U6266 ( .A1(n5213), .A2(n4701), .ZN(n4700) );
  NAND4_X1 U6267 ( .A1(n5521), .A2(n5486), .A3(n10234), .A4(n10430), .ZN(n4701) );
  NOR2_X1 U6268 ( .A1(n9183), .A2(n9167), .ZN(n5691) );
  INV_X1 U6269 ( .A(n4708), .ZN(n9359) );
  INV_X1 U6270 ( .A(n4714), .ZN(n9227) );
  INV_X1 U6271 ( .A(n4724), .ZN(n6707) );
  INV_X1 U6272 ( .A(n4722), .ZN(n6758) );
  INV_X1 U6273 ( .A(n6757), .ZN(n4721) );
  INV_X1 U6274 ( .A(n4731), .ZN(n4732) );
  OAI21_X1 U6275 ( .B1(n7862), .B2(n4735), .A(n8069), .ZN(n4731) );
  NAND3_X1 U6276 ( .A1(n7862), .A2(n4737), .A3(n4734), .ZN(n4733) );
  NAND2_X1 U6277 ( .A1(n8065), .A2(n8064), .ZN(n4740) );
  NAND3_X1 U6278 ( .A1(n7477), .A2(n4514), .A3(n7970), .ZN(n4742) );
  INV_X1 U6279 ( .A(n7970), .ZN(n4743) );
  NAND2_X1 U6280 ( .A1(n7564), .A2(n7970), .ZN(n7580) );
  NAND2_X1 U6281 ( .A1(n4744), .A2(n4745), .ZN(n7564) );
  NAND2_X1 U6282 ( .A1(n7878), .A2(n4491), .ZN(n4746) );
  INV_X1 U6283 ( .A(n8805), .ZN(n4749) );
  NAND2_X1 U6284 ( .A1(n7274), .A2(n4500), .ZN(n7277) );
  NAND2_X1 U6285 ( .A1(n7277), .A2(n7954), .ZN(n7276) );
  NAND2_X1 U6286 ( .A1(n8674), .A2(n8028), .ZN(n8655) );
  NAND2_X1 U6287 ( .A1(n8674), .A2(n4754), .ZN(n4753) );
  INV_X1 U6288 ( .A(n7833), .ZN(n8405) );
  NAND2_X1 U6289 ( .A1(n5132), .A2(n4758), .ZN(n4757) );
  OAI21_X1 U6290 ( .B1(n5132), .B2(n4503), .A(n4758), .ZN(n5502) );
  NAND2_X1 U6291 ( .A1(n5612), .A2(n4767), .ZN(n4766) );
  NAND2_X1 U6292 ( .A1(n5403), .A2(n4489), .ZN(n4776) );
  NOR2_X1 U6293 ( .A1(n7036), .A2(n4807), .ZN(n4804) );
  OAI21_X1 U6294 ( .B1(n8213), .B2(n4807), .A(n8285), .ZN(n4806) );
  OAI21_X2 U6295 ( .B1(n4804), .B2(n4806), .A(n8338), .ZN(n8110) );
  NAND2_X1 U6296 ( .A1(n4805), .A2(n8336), .ZN(n8292) );
  NAND2_X1 U6297 ( .A1(n7036), .A2(n8213), .ZN(n4805) );
  INV_X1 U6298 ( .A(n8336), .ZN(n4807) );
  NAND2_X1 U6299 ( .A1(n4813), .A2(n7118), .ZN(n9624) );
  NAND2_X1 U6300 ( .A1(n5702), .A2(n7394), .ZN(n7118) );
  NAND2_X1 U6301 ( .A1(n8257), .A2(n9624), .ZN(n5703) );
  NAND2_X1 U6302 ( .A1(n9340), .A2(n4820), .ZN(n4819) );
  NAND2_X1 U6303 ( .A1(n9290), .A2(n4825), .ZN(n4824) );
  OAI21_X1 U6304 ( .B1(n4826), .B2(n5712), .A(n8303), .ZN(n4823) );
  NAND2_X2 U6305 ( .A1(n9221), .A2(n8165), .ZN(n9214) );
  AOI21_X2 U6306 ( .B1(n7655), .B2(n8265), .A(n8254), .ZN(n9347) );
  OAI21_X2 U6307 ( .B1(n7596), .B2(n8229), .A(n8139), .ZN(n7655) );
  NAND2_X1 U6308 ( .A1(n9603), .A2(n8260), .ZN(n7596) );
  NAND2_X1 U6309 ( .A1(n5707), .A2(n8261), .ZN(n9601) );
  NAND2_X1 U6310 ( .A1(n9239), .A2(n8091), .ZN(n9223) );
  NAND2_X1 U6311 ( .A1(n5700), .A2(n5699), .ZN(n7396) );
  NAND2_X1 U6312 ( .A1(n5708), .A2(n8249), .ZN(n9340) );
  INV_X1 U6313 ( .A(n5333), .ZN(n5098) );
  AOI21_X2 U6314 ( .B1(n9303), .B2(n9304), .A(n5710), .ZN(n9290) );
  XNOR2_X1 U6315 ( .A(n5280), .B(n5279), .ZN(n6530) );
  NOR2_X2 U6316 ( .A1(n7398), .A2(n9893), .ZN(n9751) );
  NOR2_X2 U6317 ( .A1(n9201), .A2(n9209), .ZN(n9200) );
  OR2_X2 U6318 ( .A1(n9223), .A2(n9224), .ZN(n9221) );
  OR2_X2 U6319 ( .A1(n9601), .A2(n9600), .ZN(n9603) );
  OR2_X1 U6320 ( .A1(n7396), .A2(n8218), .ZN(n7394) );
  INV_X1 U6321 ( .A(n4830), .ZN(n7854) );
  NAND3_X1 U6322 ( .A1(n4850), .A2(n4849), .A3(n4848), .ZN(n5088) );
  NAND3_X1 U6323 ( .A1(n5033), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_DATAO_REG_2__SCAN_IN), .ZN(n4848) );
  NAND3_X1 U6324 ( .A1(n5037), .A2(n5036), .A3(P1_DATAO_REG_2__SCAN_IN), .ZN(
        n4849) );
  NAND3_X1 U6325 ( .A1(n5035), .A2(P2_DATAO_REG_2__SCAN_IN), .A3(n5034), .ZN(
        n4850) );
  NAND2_X1 U6326 ( .A1(n4864), .A2(n4866), .ZN(n9022) );
  INV_X1 U6327 ( .A(n6468), .ZN(n4868) );
  OAI211_X1 U6328 ( .C1(n9059), .C2(n4875), .A(n4872), .B(n4870), .ZN(n6518)
         );
  NAND2_X1 U6329 ( .A1(n9059), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U6330 ( .A1(n7620), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U6331 ( .A1(n4879), .A2(n4882), .ZN(n6401) );
  NAND2_X1 U6332 ( .A1(n4887), .A2(n4554), .ZN(n7544) );
  INV_X1 U6333 ( .A(n4891), .ZN(n5733) );
  NAND2_X1 U6334 ( .A1(n6347), .A2(n6343), .ZN(n6339) );
  INV_X1 U6335 ( .A(n4899), .ZN(n4896) );
  NAND2_X1 U6336 ( .A1(n4902), .A2(n6935), .ZN(n8443) );
  NAND3_X1 U6337 ( .A1(n4543), .A2(n6934), .A3(n4903), .ZN(n4902) );
  NAND2_X1 U6338 ( .A1(n5833), .A2(n6938), .ZN(n4903) );
  NAND2_X1 U6339 ( .A1(n8430), .A2(n4911), .ZN(n4910) );
  OAI211_X1 U6340 ( .C1(n8430), .C2(n4912), .A(n4910), .B(n6273), .ZN(P2_U3222) );
  OAI21_X1 U6341 ( .B1(n7740), .B2(n4923), .A(n4921), .ZN(n7779) );
  NAND2_X1 U6342 ( .A1(n7740), .A2(n4921), .ZN(n4920) );
  INV_X2 U6343 ( .A(n7864), .ZN(n7306) );
  NAND2_X4 U6344 ( .A1(n6267), .A2(n4927), .ZN(n7864) );
  NOR2_X1 U6345 ( .A1(n7250), .A2(n4941), .ZN(n4936) );
  INV_X1 U6346 ( .A(n7077), .ZN(n4942) );
  INV_X1 U6347 ( .A(n7250), .ZN(n4939) );
  OAI21_X1 U6348 ( .B1(n4947), .B2(n7159), .A(n5970), .ZN(n4944) );
  NOR2_X1 U6349 ( .A1(n7159), .A2(n4948), .ZN(n4946) );
  NAND2_X1 U6350 ( .A1(n4950), .A2(n4949), .ZN(n8520) );
  NOR2_X1 U6351 ( .A1(n4488), .A2(n4955), .ZN(n5792) );
  NOR2_X1 U6352 ( .A1(n5319), .A2(n4958), .ZN(n5337) );
  NAND2_X1 U6353 ( .A1(n7291), .A2(n8216), .ZN(n4964) );
  OAI21_X1 U6354 ( .B1(n4961), .B2(n5075), .A(n4960), .ZN(n7208) );
  NAND2_X1 U6355 ( .A1(n7291), .A2(n4494), .ZN(n4960) );
  INV_X1 U6356 ( .A(n5075), .ZN(n4963) );
  NAND2_X1 U6357 ( .A1(n5372), .A2(n4552), .ZN(n7121) );
  NAND2_X1 U6358 ( .A1(n7121), .A2(n5388), .ZN(n9750) );
  NAND2_X1 U6359 ( .A1(n7029), .A2(n5295), .ZN(n7196) );
  NAND2_X1 U6360 ( .A1(n4968), .A2(n4967), .ZN(n7029) );
  OAI211_X1 U6361 ( .C1(n4968), .C2(n4966), .A(n4965), .B(n7195), .ZN(n5308)
         );
  NAND2_X1 U6362 ( .A1(n8213), .A2(n5295), .ZN(n4965) );
  INV_X1 U6363 ( .A(n5295), .ZN(n4966) );
  INV_X1 U6364 ( .A(n7027), .ZN(n4968) );
  NAND2_X1 U6365 ( .A1(n7338), .A2(n7337), .ZN(n7336) );
  NAND2_X1 U6366 ( .A1(n4969), .A2(n4972), .ZN(n7530) );
  NAND2_X1 U6367 ( .A1(n7338), .A2(n4970), .ZN(n4969) );
  NAND2_X1 U6368 ( .A1(n5682), .A2(n5681), .ZN(n4980) );
  INV_X1 U6369 ( .A(n5682), .ZN(n4977) );
  AND2_X1 U6370 ( .A1(n9167), .A2(n9088), .ZN(n4981) );
  NAND2_X1 U6371 ( .A1(n9258), .A2(n4984), .ZN(n4982) );
  NAND2_X1 U6372 ( .A1(n4982), .A2(n4983), .ZN(n9225) );
  OR2_X1 U6373 ( .A1(n8962), .A2(n9605), .ZN(n4996) );
  NAND2_X1 U6374 ( .A1(n5318), .A2(n4998), .ZN(n4997) );
  NAND2_X1 U6375 ( .A1(n7477), .A2(n4491), .ZN(n5004) );
  NAND3_X1 U6376 ( .A1(n5004), .A2(n5003), .A3(n7959), .ZN(n7563) );
  NAND3_X1 U6377 ( .A1(n8748), .A2(n7829), .A3(n5008), .ZN(n5007) );
  INV_X1 U6378 ( .A(n5013), .ZN(n8733) );
  NAND2_X1 U6379 ( .A1(n5914), .A2(n5913), .ZN(n5023) );
  NAND2_X1 U6380 ( .A1(n5023), .A2(n7358), .ZN(n7949) );
  XNOR2_X1 U6381 ( .A(n5023), .B(n6157), .ZN(n5923) );
  NAND2_X1 U6382 ( .A1(n5023), .A2(n10013), .ZN(n5017) );
  AOI21_X1 U6383 ( .B1(n8620), .B2(n5023), .A(n5018), .ZN(n7116) );
  AOI21_X1 U6384 ( .B1(n7150), .B2(n5023), .A(n10024), .ZN(n5020) );
  AOI21_X1 U6385 ( .B1(n8492), .B2(n5023), .A(n5022), .ZN(n7254) );
  NAND2_X1 U6386 ( .A1(n5025), .A2(n5024), .ZN(n8807) );
  NAND2_X1 U6387 ( .A1(n5031), .A2(n8038), .ZN(n5029) );
  NAND2_X1 U6388 ( .A1(n5031), .A2(n5032), .ZN(n5030) );
  INV_X1 U6389 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5036) );
  INV_X2 U6390 ( .A(n7856), .ZN(n5194) );
  NAND2_X1 U6391 ( .A1(n5038), .A2(n8420), .ZN(n6820) );
  XNOR2_X1 U6392 ( .A(n7870), .B(n7221), .ZN(n8426) );
  XNOR2_X1 U6393 ( .A(n7870), .B(n5819), .ZN(n9959) );
  NAND3_X1 U6394 ( .A1(n5763), .A2(n5876), .A3(n5762), .ZN(n6049) );
  NAND2_X1 U6395 ( .A1(n8714), .A2(n5043), .ZN(n5042) );
  NAND3_X1 U6396 ( .A1(n5056), .A2(n7355), .A3(n5057), .ZN(n7270) );
  NAND3_X1 U6397 ( .A1(n7106), .A2(n7107), .A3(n4513), .ZN(n5058) );
  NAND2_X1 U6398 ( .A1(n5770), .A2(n5062), .ZN(n5800) );
  NAND2_X1 U6399 ( .A1(n7767), .A2(n5066), .ZN(n5065) );
  NAND2_X1 U6400 ( .A1(n5065), .A2(n5064), .ZN(n8775) );
  NAND2_X1 U6401 ( .A1(n6252), .A2(n7892), .ZN(n6831) );
  INV_X1 U6402 ( .A(n6599), .ZN(n6293) );
  NAND2_X1 U6403 ( .A1(n5243), .A2(n5242), .ZN(n5247) );
  AND2_X1 U6404 ( .A1(n7532), .A2(n7531), .ZN(n9647) );
  INV_X1 U6405 ( .A(n5668), .ZN(n5200) );
  NAND2_X4 U6406 ( .A1(n6498), .A2(n6497), .ZN(n7030) );
  NAND2_X1 U6407 ( .A1(n5737), .A2(n5753), .ZN(n6547) );
  INV_X1 U6408 ( .A(n6562), .ZN(n5721) );
  OAI21_X1 U6409 ( .B1(n6966), .B2(n7872), .A(n7918), .ZN(n7109) );
  INV_X1 U6410 ( .A(n6601), .ZN(n6292) );
  INV_X1 U6411 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5987) );
  INV_X1 U6412 ( .A(n5851), .ZN(n6095) );
  INV_X1 U6413 ( .A(n8223), .ZN(n5387) );
  CLKBUF_X3 U6414 ( .A(n5284), .Z(n5674) );
  AND2_X1 U6415 ( .A1(n5119), .A2(n5118), .ZN(n5074) );
  AND2_X1 U6416 ( .A1(n9865), .A2(n9784), .ZN(n5075) );
  INV_X1 U6417 ( .A(n9779), .ZN(n5342) );
  AND3_X1 U6418 ( .A1(n10434), .A2(n5726), .A3(n5725), .ZN(n5076) );
  OR2_X1 U6419 ( .A1(n5690), .A2(n9532), .ZN(n5077) );
  AND2_X1 U6420 ( .A1(n5114), .A2(n5113), .ZN(n5079) );
  INV_X1 U6421 ( .A(n9818), .ZN(n9350) );
  NAND2_X2 U6422 ( .A1(n7032), .A2(n9800), .ZN(n9816) );
  INV_X1 U6423 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5214) );
  INV_X1 U6424 ( .A(n7355), .ZN(n7275) );
  INV_X1 U6425 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5765) );
  NOR2_X1 U6426 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  INV_X1 U6427 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5944) );
  INV_X1 U6428 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U6429 ( .A1(n6162), .A2(n8484), .ZN(n6163) );
  INV_X1 U6430 ( .A(n8938), .ZN(n5784) );
  NOR2_X1 U6431 ( .A1(n5962), .A2(n10462), .ZN(n5976) );
  AND2_X1 U6432 ( .A1(n6237), .A2(n9941), .ZN(n6972) );
  INV_X1 U6433 ( .A(n5616), .ZN(n5236) );
  INV_X1 U6434 ( .A(n5545), .ZN(n5234) );
  INV_X1 U6435 ( .A(n5576), .ZN(n5235) );
  INV_X1 U6436 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5492) );
  INV_X1 U6437 ( .A(n8307), .ZN(n5690) );
  NOR2_X1 U6438 ( .A1(n7719), .A2(n7617), .ZN(n5752) );
  INV_X1 U6439 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5241) );
  INV_X1 U6440 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5728) );
  INV_X1 U6441 ( .A(SI_22_), .ZN(n10375) );
  INV_X1 U6442 ( .A(SI_19_), .ZN(n5157) );
  INV_X1 U6443 ( .A(SI_15_), .ZN(n5138) );
  INV_X1 U6444 ( .A(SI_10_), .ZN(n10198) );
  NOR2_X1 U6445 ( .A1(n6053), .A2(n5777), .ZN(n6075) );
  INV_X1 U6446 ( .A(n8452), .ZN(n6114) );
  INV_X1 U6447 ( .A(n7078), .ZN(n5906) );
  OR2_X1 U6448 ( .A1(n8852), .A2(n8402), .ZN(n8403) );
  OR2_X1 U6449 ( .A1(n8864), .A2(n8707), .ZN(n8401) );
  INV_X1 U6450 ( .A(n7902), .ZN(n7727) );
  NAND2_X1 U6451 ( .A1(n8531), .A2(n8618), .ZN(n8409) );
  INV_X1 U6452 ( .A(n6308), .ZN(n6489) );
  INV_X1 U6453 ( .A(n6485), .ZN(n6486) );
  NAND2_X1 U6454 ( .A1(n5234), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5562) );
  OR2_X1 U6455 ( .A1(n5673), .A2(n5239), .ZN(n5260) );
  OR2_X1 U6456 ( .A1(n5589), .A2(n8983), .ZN(n5602) );
  OR2_X1 U6457 ( .A1(n5493), .A2(n5492), .ZN(n5508) );
  AND2_X1 U6458 ( .A1(n5657), .A2(n5644), .ZN(n9211) );
  OR2_X1 U6459 ( .A1(n5488), .A2(n5282), .ZN(n5283) );
  NOR2_X2 U6460 ( .A1(n9295), .A2(n9311), .ZN(n9294) );
  AND2_X1 U6461 ( .A1(n5716), .A2(n8332), .ZN(n6608) );
  AND2_X1 U6462 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  AND2_X1 U6463 ( .A1(n6260), .A2(n6206), .ZN(n8638) );
  OR2_X1 U6464 ( .A1(n6179), .A2(n10182), .ZN(n6205) );
  INV_X1 U6465 ( .A(n8511), .ZN(n8499) );
  INV_X1 U6466 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10462) );
  INV_X1 U6467 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7327) );
  INV_X1 U6468 ( .A(n9929), .ZN(n9934) );
  INV_X1 U6469 ( .A(n8675), .ZN(n8665) );
  OR2_X1 U6470 ( .A1(n6022), .A2(n10277), .ZN(n6053) );
  INV_X1 U6471 ( .A(n6830), .ZN(n6555) );
  INV_X1 U6472 ( .A(n8061), .ZN(n7868) );
  AND2_X1 U6473 ( .A1(n7943), .A2(n7948), .ZN(n7876) );
  AND2_X1 U6474 ( .A1(n6227), .A2(n7750), .ZN(n9941) );
  NAND2_X1 U6475 ( .A1(n5233), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U6476 ( .A1(n7436), .A2(n7437), .ZN(n7435) );
  OR2_X1 U6477 ( .A1(n7006), .A2(n6583), .ZN(n6591) );
  OR2_X1 U6478 ( .A1(n5602), .A2(n9040), .ZN(n5616) );
  OR2_X1 U6479 ( .A1(n5528), .A2(n9016), .ZN(n5545) );
  INV_X1 U6480 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7495) );
  INV_X1 U6481 ( .A(n9436), .ZN(n9309) );
  AND2_X1 U6482 ( .A1(n8127), .A2(n8126), .ZN(n9625) );
  OR2_X1 U6483 ( .A1(n7011), .A2(n4481), .ZN(n9615) );
  AND2_X1 U6484 ( .A1(n6608), .A2(n6872), .ZN(n9866) );
  OR2_X1 U6485 ( .A1(n7011), .A2(n9814), .ZN(n5759) );
  INV_X1 U6486 ( .A(n9892), .ZN(n9902) );
  OR2_X1 U6487 ( .A1(n9896), .A2(n8332), .ZN(n7010) );
  INV_X1 U6488 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9534) );
  OR3_X1 U6489 ( .A1(n7615), .A2(n7717), .A3(n6240), .ZN(n6519) );
  NOR2_X1 U6490 ( .A1(n8524), .A2(n8762), .ZN(n8511) );
  AND2_X1 U6491 ( .A1(n6205), .A2(n6180), .ZN(n8670) );
  INV_X1 U6492 ( .A(n6251), .ZN(n6259) );
  AND4_X1 U6493 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n8658)
         );
  AND4_X1 U6494 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n8464)
         );
  AND4_X1 U6495 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n7709)
         );
  AND2_X1 U6496 ( .A1(n6663), .A2(n6662), .ZN(n9929) );
  NOR2_X1 U6497 ( .A1(n8041), .A2(n8044), .ZN(n8404) );
  AND2_X1 U6498 ( .A1(n7765), .A2(n7725), .ZN(n8911) );
  AND2_X1 U6499 ( .A1(n8696), .A2(n6817), .ZN(n8792) );
  NAND2_X1 U6500 ( .A1(n6824), .A2(n8821), .ZN(n8696) );
  NOR2_X1 U6501 ( .A1(n9945), .A2(n6238), .ZN(n6978) );
  AND2_X1 U6502 ( .A1(n8813), .A2(n8812), .ZN(n8904) );
  INV_X1 U6503 ( .A(n10019), .ZN(n10029) );
  AND2_X1 U6504 ( .A1(n6519), .A2(n9948), .ZN(n9943) );
  AND2_X1 U6505 ( .A1(n5971), .A2(n5960), .ZN(n7092) );
  INV_X1 U6506 ( .A(n9062), .ZN(n9074) );
  INV_X1 U6507 ( .A(n9079), .ZN(n9064) );
  OR2_X1 U6508 ( .A1(n9060), .A2(n5659), .ZN(n5664) );
  INV_X1 U6509 ( .A(n5674), .ZN(n5659) );
  AND4_X1 U6510 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n9627)
         );
  NOR2_X1 U6511 ( .A1(n8081), .A2(n8382), .ZN(n9735) );
  NAND2_X1 U6512 ( .A1(n6619), .A2(n8382), .ZN(n9739) );
  INV_X1 U6513 ( .A(n9748), .ZN(n9134) );
  INV_X1 U6514 ( .A(n9615), .ZN(n9794) );
  AND2_X1 U6515 ( .A1(n8156), .A2(n8281), .ZN(n9304) );
  AND2_X1 U6516 ( .A1(n8100), .A2(n8099), .ZN(n9339) );
  INV_X1 U6517 ( .A(n9888), .ZN(n9863) );
  AND2_X1 U6518 ( .A1(n5715), .A2(n8205), .ZN(n9882) );
  AND2_X1 U6519 ( .A1(n7031), .A2(n7030), .ZN(n9791) );
  INV_X1 U6520 ( .A(n9800), .ZN(n9787) );
  NAND2_X1 U6521 ( .A1(n9797), .A2(n5759), .ZN(n9892) );
  NAND2_X1 U6522 ( .A1(n9812), .A2(n9896), .ZN(n9885) );
  AND2_X1 U6523 ( .A1(n7006), .A2(n7010), .ZN(n6585) );
  AND2_X1 U6524 ( .A1(n5539), .A2(n5525), .ZN(n9121) );
  AND2_X1 U6525 ( .A1(n5407), .A2(n5420), .ZN(n6850) );
  XNOR2_X1 U6526 ( .A(n5318), .B(n5317), .ZN(n6528) );
  NOR2_X1 U6527 ( .A1(n10498), .A2(n10072), .ZN(n10073) );
  NOR2_X1 U6528 ( .A1(n6519), .A2(P2_U3152), .ZN(n6652) );
  INV_X1 U6529 ( .A(n8617), .ZN(n9932) );
  AND2_X1 U6530 ( .A1(n6272), .A2(n6271), .ZN(n6273) );
  INV_X1 U6531 ( .A(n8503), .ZN(n8529) );
  INV_X1 U6532 ( .A(n8658), .ZN(n8532) );
  INV_X1 U6533 ( .A(n8765), .ZN(n8811) );
  INV_X1 U6534 ( .A(n7268), .ZN(n8545) );
  NAND2_X1 U6535 ( .A1(n6669), .A2(n6657), .ZN(n9935) );
  INV_X1 U6536 ( .A(n8611), .ZN(n9933) );
  INV_X1 U6537 ( .A(n8816), .ZN(n8629) );
  NAND2_X1 U6538 ( .A1(n8696), .A2(n6901), .ZN(n8818) );
  INV_X1 U6539 ( .A(n10052), .ZN(n10050) );
  INV_X1 U6540 ( .A(n10032), .ZN(n10030) );
  NAND2_X1 U6541 ( .A1(n9943), .A2(n9942), .ZN(n9946) );
  INV_X1 U6542 ( .A(n6254), .ZN(n7786) );
  INV_X1 U6543 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6988) );
  CLKBUF_X1 U6544 ( .A(n8944), .Z(n8949) );
  NAND2_X1 U6545 ( .A1(n7237), .A2(n6501), .ZN(n9067) );
  INV_X1 U6546 ( .A(n9182), .ZN(n9088) );
  OAI21_X1 U6547 ( .B1(n9259), .B2(n5659), .A(n5607), .ZN(n9421) );
  INV_X1 U6548 ( .A(n9627), .ZN(n9606) );
  INV_X1 U6549 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U6550 ( .A1(n6621), .A2(n6620), .ZN(n9748) );
  NAND2_X1 U6551 ( .A1(n9816), .A2(n9791), .ZN(n9818) );
  INV_X1 U6552 ( .A(n9928), .ZN(n9925) );
  AND2_X2 U6553 ( .A1(n6585), .A2(n6584), .ZN(n9928) );
  INV_X1 U6554 ( .A(n9228), .ZN(n9499) );
  INV_X1 U6555 ( .A(n9329), .ZN(n9520) );
  INV_X1 U6556 ( .A(n9911), .ZN(n9909) );
  INV_X1 U6557 ( .A(n7009), .ZN(n6552) );
  NAND2_X1 U6558 ( .A1(n6552), .A2(n6547), .ZN(n9823) );
  INV_X1 U6559 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10171) );
  INV_X1 U6560 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7445) );
  INV_X1 U6561 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10393) );
  INV_X1 U6562 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6573) );
  NOR2_X1 U6563 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  OAI21_X1 U6564 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10098), .ZN(n10096) );
  AND2_X2 U6565 ( .A1(n6652), .A2(n6520), .ZN(P2_U3966) );
  INV_X1 U6566 ( .A(n9095), .ZN(P1_U4006) );
  INV_X4 U6567 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U6568 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5758) );
  INV_X2 U6569 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6570 ( .A1(n5291), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5083) );
  AND2_X1 U6571 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5082) );
  INV_X1 U6572 ( .A(SI_1_), .ZN(n5084) );
  MUX2_X1 U6573 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5194), .Z(n5279) );
  NAND2_X1 U6574 ( .A1(n5085), .A2(SI_1_), .ZN(n5086) );
  INV_X1 U6575 ( .A(SI_2_), .ZN(n5087) );
  XNOR2_X1 U6576 ( .A(n5088), .B(n5087), .ZN(n5273) );
  NAND2_X1 U6577 ( .A1(n5274), .A2(n5273), .ZN(n5090) );
  NAND2_X1 U6578 ( .A1(n5088), .A2(SI_2_), .ZN(n5089) );
  NAND2_X1 U6579 ( .A1(n5090), .A2(n5089), .ZN(n5303) );
  MUX2_X1 U6580 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5194), .Z(n5092) );
  INV_X1 U6581 ( .A(SI_3_), .ZN(n5091) );
  XNOR2_X1 U6582 ( .A(n5092), .B(n5091), .ZN(n5302) );
  NAND2_X1 U6583 ( .A1(n5303), .A2(n5302), .ZN(n5094) );
  NAND2_X1 U6584 ( .A1(n5092), .A2(SI_3_), .ZN(n5093) );
  MUX2_X1 U6585 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5194), .Z(n5096) );
  XNOR2_X1 U6586 ( .A(n5096), .B(SI_4_), .ZN(n5317) );
  INV_X1 U6587 ( .A(n5317), .ZN(n5095) );
  NAND2_X1 U6588 ( .A1(n5096), .A2(SI_4_), .ZN(n5097) );
  MUX2_X1 U6589 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6521), .Z(n5101) );
  XNOR2_X1 U6590 ( .A(n5101), .B(SI_6_), .ZN(n5343) );
  INV_X1 U6591 ( .A(n5343), .ZN(n5100) );
  NAND2_X1 U6592 ( .A1(n5101), .A2(SI_6_), .ZN(n5102) );
  MUX2_X1 U6593 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6521), .Z(n5104) );
  XNOR2_X1 U6594 ( .A(n5104), .B(SI_7_), .ZN(n5358) );
  INV_X1 U6595 ( .A(n5358), .ZN(n5103) );
  NAND2_X1 U6596 ( .A1(n5104), .A2(SI_7_), .ZN(n5105) );
  MUX2_X1 U6597 ( .A(n6546), .B(n6544), .S(n6521), .Z(n5107) );
  INV_X1 U6598 ( .A(SI_8_), .ZN(n5106) );
  NAND2_X1 U6599 ( .A1(n5107), .A2(n5106), .ZN(n5110) );
  INV_X1 U6600 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6601 ( .A1(n5108), .A2(SI_8_), .ZN(n5109) );
  NAND2_X1 U6602 ( .A1(n5110), .A2(n5109), .ZN(n5373) );
  MUX2_X1 U6603 ( .A(n6561), .B(n6559), .S(n6521), .Z(n5111) );
  NAND2_X1 U6604 ( .A1(n5111), .A2(n10145), .ZN(n5114) );
  INV_X1 U6605 ( .A(n5111), .ZN(n5112) );
  NAND2_X1 U6606 ( .A1(n5112), .A2(SI_9_), .ZN(n5113) );
  MUX2_X1 U6607 ( .A(n6574), .B(n6573), .S(n6521), .Z(n5116) );
  NAND2_X1 U6608 ( .A1(n5116), .A2(n10198), .ZN(n5119) );
  INV_X1 U6609 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U6610 ( .A1(n5117), .A2(SI_10_), .ZN(n5118) );
  MUX2_X1 U6611 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6521), .Z(n5121) );
  XNOR2_X1 U6612 ( .A(n5121), .B(n5120), .ZN(n5418) );
  INV_X1 U6613 ( .A(n5418), .ZN(n5122) );
  MUX2_X1 U6614 ( .A(n5123), .B(n10419), .S(n6521), .Z(n5124) );
  NAND2_X1 U6615 ( .A1(n5124), .A2(n10212), .ZN(n5127) );
  INV_X1 U6616 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6617 ( .A1(n5125), .A2(SI_12_), .ZN(n5126) );
  NAND2_X1 U6618 ( .A1(n5127), .A2(n5126), .ZN(n5431) );
  MUX2_X1 U6619 ( .A(n6802), .B(n10387), .S(n6521), .Z(n5128) );
  NAND2_X1 U6620 ( .A1(n5128), .A2(n10456), .ZN(n5131) );
  INV_X1 U6621 ( .A(n5128), .ZN(n5129) );
  NAND2_X1 U6622 ( .A1(n5129), .A2(SI_13_), .ZN(n5130) );
  MUX2_X1 U6623 ( .A(n6839), .B(n5133), .S(n5194), .Z(n5134) );
  XNOR2_X1 U6624 ( .A(n5134), .B(SI_14_), .ZN(n5464) );
  INV_X1 U6625 ( .A(n5464), .ZN(n5137) );
  INV_X1 U6626 ( .A(n5134), .ZN(n5135) );
  NAND2_X1 U6627 ( .A1(n5135), .A2(SI_14_), .ZN(n5136) );
  MUX2_X1 U6628 ( .A(n6988), .B(n10393), .S(n6521), .Z(n5139) );
  NAND2_X1 U6629 ( .A1(n5139), .A2(n5138), .ZN(n5142) );
  INV_X1 U6630 ( .A(n5139), .ZN(n5140) );
  NAND2_X1 U6631 ( .A1(n5140), .A2(SI_15_), .ZN(n5141) );
  NAND2_X1 U6632 ( .A1(n5142), .A2(n5141), .ZN(n5484) );
  MUX2_X1 U6633 ( .A(n7045), .B(n10360), .S(n6521), .Z(n5144) );
  INV_X1 U6634 ( .A(SI_16_), .ZN(n5143) );
  NAND2_X1 U6635 ( .A1(n5144), .A2(n5143), .ZN(n5147) );
  INV_X1 U6636 ( .A(n5144), .ZN(n5145) );
  NAND2_X1 U6637 ( .A1(n5145), .A2(SI_16_), .ZN(n5146) );
  MUX2_X1 U6638 ( .A(n7130), .B(n5149), .S(n6521), .Z(n5150) );
  XNOR2_X1 U6639 ( .A(n5150), .B(SI_17_), .ZN(n5519) );
  INV_X1 U6640 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6641 ( .A1(n5151), .A2(SI_17_), .ZN(n5152) );
  MUX2_X1 U6642 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6521), .Z(n5154) );
  XNOR2_X1 U6643 ( .A(n5154), .B(SI_18_), .ZN(n5537) );
  INV_X1 U6644 ( .A(n5537), .ZN(n5153) );
  NAND2_X1 U6645 ( .A1(n5538), .A2(n5153), .ZN(n5156) );
  NAND2_X1 U6646 ( .A1(n5154), .A2(SI_18_), .ZN(n5155) );
  MUX2_X1 U6647 ( .A(n7316), .B(n10432), .S(n6521), .Z(n5158) );
  NAND2_X1 U6648 ( .A1(n5158), .A2(n5157), .ZN(n5161) );
  INV_X1 U6649 ( .A(n5158), .ZN(n5159) );
  NAND2_X1 U6650 ( .A1(n5159), .A2(SI_19_), .ZN(n5160) );
  NAND2_X1 U6651 ( .A1(n5161), .A2(n5160), .ZN(n5552) );
  MUX2_X1 U6652 ( .A(n7448), .B(n7445), .S(n6521), .Z(n5163) );
  INV_X1 U6653 ( .A(SI_20_), .ZN(n5162) );
  NAND2_X1 U6654 ( .A1(n5163), .A2(n5162), .ZN(n5166) );
  INV_X1 U6655 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6656 ( .A1(n5164), .A2(SI_20_), .ZN(n5165) );
  MUX2_X1 U6657 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5194), .Z(n5170) );
  INV_X1 U6658 ( .A(SI_21_), .ZN(n5168) );
  XNOR2_X1 U6659 ( .A(n5170), .B(n5168), .ZN(n5585) );
  INV_X1 U6660 ( .A(n5585), .ZN(n5169) );
  NAND2_X1 U6661 ( .A1(n5170), .A2(SI_21_), .ZN(n5171) );
  MUX2_X1 U6662 ( .A(n7788), .B(n10392), .S(n6521), .Z(n5172) );
  NAND2_X1 U6663 ( .A1(n5172), .A2(n10375), .ZN(n5175) );
  INV_X1 U6664 ( .A(n5172), .ZN(n5173) );
  NAND2_X1 U6665 ( .A1(n5173), .A2(SI_22_), .ZN(n5174) );
  NAND2_X1 U6666 ( .A1(n5175), .A2(n5174), .ZN(n5598) );
  INV_X1 U6667 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5177) );
  INV_X1 U6668 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5176) );
  MUX2_X1 U6669 ( .A(n5177), .B(n5176), .S(n6521), .Z(n5178) );
  INV_X1 U6670 ( .A(SI_23_), .ZN(n10220) );
  NAND2_X1 U6671 ( .A1(n5178), .A2(n10220), .ZN(n5181) );
  INV_X1 U6672 ( .A(n5178), .ZN(n5179) );
  NAND2_X1 U6673 ( .A1(n5179), .A2(SI_23_), .ZN(n5180) );
  MUX2_X1 U6674 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6521), .Z(n5182) );
  INV_X1 U6675 ( .A(SI_24_), .ZN(n10446) );
  XNOR2_X1 U6676 ( .A(n5182), .B(n10446), .ZN(n5625) );
  INV_X1 U6677 ( .A(n5625), .ZN(n5184) );
  NAND2_X1 U6678 ( .A1(n5182), .A2(SI_24_), .ZN(n5183) );
  INV_X1 U6679 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7718) );
  INV_X1 U6680 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10184) );
  MUX2_X1 U6681 ( .A(n7718), .B(n10184), .S(n6521), .Z(n5185) );
  INV_X1 U6682 ( .A(SI_25_), .ZN(n10461) );
  NAND2_X1 U6683 ( .A1(n5185), .A2(n10461), .ZN(n5188) );
  INV_X1 U6684 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6685 ( .A1(n5186), .A2(SI_25_), .ZN(n5187) );
  NAND2_X1 U6686 ( .A1(n5188), .A2(n5187), .ZN(n5639) );
  INV_X1 U6687 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U6688 ( .A(n5189), .B(n10171), .S(n6521), .Z(n5190) );
  NAND2_X1 U6689 ( .A1(n5190), .A2(n10373), .ZN(n5193) );
  INV_X1 U6690 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U6691 ( .A1(n5191), .A2(SI_26_), .ZN(n5192) );
  INV_X1 U6692 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5195) );
  MUX2_X1 U6693 ( .A(n5195), .B(n10181), .S(n5194), .Z(n5196) );
  INV_X1 U6694 ( .A(SI_27_), .ZN(n10148) );
  NAND2_X1 U6695 ( .A1(n5196), .A2(n10148), .ZN(n5201) );
  INV_X1 U6696 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6697 ( .A1(n5197), .A2(SI_27_), .ZN(n5198) );
  NAND2_X1 U6698 ( .A1(n5201), .A2(n5198), .ZN(n5667) );
  INV_X1 U6699 ( .A(n5667), .ZN(n5199) );
  INV_X1 U6700 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5202) );
  INV_X1 U6701 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10150) );
  MUX2_X1 U6702 ( .A(n5202), .B(n10150), .S(n6521), .Z(n5204) );
  XNOR2_X1 U6703 ( .A(n5204), .B(SI_28_), .ZN(n5256) );
  INV_X1 U6704 ( .A(SI_28_), .ZN(n5203) );
  MUX2_X1 U6705 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6521), .Z(n7834) );
  INV_X1 U6706 ( .A(SI_29_), .ZN(n5205) );
  XNOR2_X1 U6707 ( .A(n7834), .B(n5205), .ZN(n5206) );
  NOR2_X1 U6708 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5212) );
  NOR2_X1 U6709 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5211) );
  NOR2_X1 U6710 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5210) );
  NOR2_X1 U6711 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5209) );
  NAND4_X1 U6712 ( .A1(n5212), .A2(n5211), .A3(n5210), .A4(n5209), .ZN(n5213)
         );
  NAND4_X1 U6713 ( .A1(n10434), .A2(n5726), .A3(n5556), .A4(n5725), .ZN(n5216)
         );
  NAND4_X1 U6714 ( .A1(n4889), .A2(n5214), .A3(n5730), .A4(n5728), .ZN(n5215)
         );
  NAND2_X1 U6715 ( .A1(n5224), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5219) );
  MUX2_X1 U6716 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5219), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5220) );
  NAND2_X1 U6717 ( .A1(n5243), .A2(n5240), .ZN(n5245) );
  NAND2_X1 U6718 ( .A1(n5220), .A2(n5245), .ZN(n5717) );
  NAND2_X1 U6719 ( .A1(n5221), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5222) );
  NAND2_X2 U6720 ( .A1(n5224), .A2(n5223), .ZN(n8381) );
  NAND2_X2 U6721 ( .A1(n5717), .A2(n8381), .ZN(n5488) );
  AND2_X2 U6722 ( .A1(n5488), .A2(n6521), .ZN(n5281) );
  INV_X4 U6723 ( .A(n5316), .ZN(n8193) );
  NAND2_X1 U6724 ( .A1(n7830), .A2(n8193), .ZN(n5226) );
  CLKBUF_X3 U6725 ( .A(n5315), .Z(n5627) );
  NAND2_X1 U6726 ( .A1(n5627), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5225) );
  NAND3_X1 U6727 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5351) );
  INV_X1 U6728 ( .A(n5351), .ZN(n5227) );
  NAND2_X1 U6729 ( .A1(n5227), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5364) );
  INV_X1 U6730 ( .A(n5364), .ZN(n5228) );
  NAND2_X1 U6731 ( .A1(n5228), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5380) );
  INV_X1 U6732 ( .A(n5380), .ZN(n5229) );
  NAND2_X1 U6733 ( .A1(n5229), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5395) );
  INV_X1 U6734 ( .A(n5441), .ZN(n5231) );
  NAND2_X1 U6735 ( .A1(n5231), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5458) );
  INV_X1 U6736 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5561) );
  INV_X1 U6737 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8983) );
  INV_X1 U6738 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9040) );
  INV_X1 U6739 ( .A(n5631), .ZN(n5237) );
  NAND2_X1 U6740 ( .A1(n5237), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5643) );
  INV_X1 U6741 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8991) );
  INV_X1 U6742 ( .A(n5657), .ZN(n5238) );
  NAND2_X1 U6743 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5239) );
  INV_X1 U6744 ( .A(n5260), .ZN(n9150) );
  NAND2_X1 U6745 ( .A1(n5245), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6746 ( .A1(n9150), .A2(n5284), .ZN(n5255) );
  INV_X1 U6747 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9376) );
  AND2_X4 U6748 ( .A1(n5250), .A2(n9538), .ZN(n6562) );
  NAND2_X1 U6749 ( .A1(n6563), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6750 ( .A1(n6564), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5251) );
  OAI211_X1 U6751 ( .C1(n9376), .C2(n5721), .A(n5252), .B(n5251), .ZN(n5253)
         );
  INV_X1 U6752 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6753 ( .A1(n5255), .A2(n5254), .ZN(n9163) );
  XNOR2_X1 U6754 ( .A(n8307), .B(n9163), .ZN(n8238) );
  NAND2_X1 U6755 ( .A1(n5627), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5257) );
  INV_X1 U6756 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6510) );
  INV_X1 U6757 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5259) );
  OAI21_X1 U6758 ( .B1(n5673), .B2(n6510), .A(n5259), .ZN(n5261) );
  NAND2_X1 U6759 ( .A1(n9170), .A2(n5674), .ZN(n5266) );
  INV_X1 U6760 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U6761 ( .A1(n6563), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6762 ( .A1(n6564), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5262) );
  OAI211_X1 U6763 ( .C1(n9381), .C2(n5721), .A(n5263), .B(n5262), .ZN(n5264)
         );
  INV_X1 U6764 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6765 ( .A1(n6562), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6766 ( .A1(n5284), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5271) );
  INV_X1 U6767 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5267) );
  OR2_X1 U6768 ( .A1(n5511), .A2(n5267), .ZN(n5270) );
  INV_X1 U6769 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5268) );
  AND4_X2 U6770 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n5294)
         );
  XNOR2_X1 U6771 ( .A(n5274), .B(n5273), .ZN(n6525) );
  NAND2_X1 U6772 ( .A1(n5315), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5278) );
  INV_X2 U6773 ( .A(n5488), .ZN(n6610) );
  OR2_X1 U6774 ( .A1(n5275), .A2(n9534), .ZN(n5276) );
  XNOR2_X1 U6775 ( .A(n5276), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U6776 ( .A1(n6610), .A2(n6886), .ZN(n5277) );
  OAI211_X1 U6777 ( .C1(n5316), .C2(n6525), .A(n5278), .B(n5277), .ZN(n6689)
         );
  NAND2_X1 U6778 ( .A1(n6602), .A2(n9832), .ZN(n8340) );
  NAND2_X1 U6779 ( .A1(n5294), .A2(n6689), .ZN(n8336) );
  AND2_X2 U6780 ( .A1(n8340), .A2(n8336), .ZN(n8213) );
  NAND2_X1 U6781 ( .A1(n5285), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U6782 ( .A1(n5350), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U6783 ( .A1(n6562), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6784 ( .A1(n5284), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5693) );
  INV_X1 U6785 ( .A(n6868), .ZN(n5282) );
  NAND2_X1 U6786 ( .A1(n5284), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6787 ( .A1(n5285), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6788 ( .A1(n6562), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6789 ( .A1(n5350), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5286) );
  NAND4_X2 U6790 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n9804)
         );
  INV_X1 U6791 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U6792 ( .A(n5291), .B(n5290), .ZN(n9550) );
  MUX2_X1 U6793 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9550), .S(n5488), .Z(n7012) );
  AND2_X1 U6794 ( .A1(n9804), .A2(n7012), .ZN(n9802) );
  NAND2_X1 U6795 ( .A1(n9803), .A2(n9802), .ZN(n9801) );
  NAND2_X1 U6796 ( .A1(n9096), .A2(n8333), .ZN(n5293) );
  NAND2_X1 U6797 ( .A1(n9801), .A2(n5293), .ZN(n7027) );
  NAND2_X1 U6798 ( .A1(n5294), .A2(n9832), .ZN(n5295) );
  NAND2_X1 U6799 ( .A1(n6562), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5301) );
  INV_X1 U6800 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U6801 ( .A1(n5674), .A2(n6806), .ZN(n5300) );
  INV_X1 U6802 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5296) );
  OR2_X1 U6803 ( .A1(n5511), .A2(n5296), .ZN(n5299) );
  INV_X1 U6804 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5297) );
  OR2_X1 U6805 ( .A1(n5512), .A2(n5297), .ZN(n5298) );
  AND4_X2 U6806 ( .A1(n5301), .A2(n5300), .A3(n5299), .A4(n5298), .ZN(n9849)
         );
  XNOR2_X1 U6807 ( .A(n5303), .B(n5302), .ZN(n6526) );
  NAND2_X1 U6808 ( .A1(n5627), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6809 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4521), .ZN(n5304) );
  XNOR2_X1 U6810 ( .A(n5304), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U6811 ( .A1(n6610), .A2(n6634), .ZN(n5305) );
  NAND2_X1 U6812 ( .A1(n9849), .A2(n7198), .ZN(n8338) );
  INV_X1 U6813 ( .A(n9849), .ZN(n9094) );
  INV_X1 U6814 ( .A(n7198), .ZN(n9840) );
  NAND2_X1 U6815 ( .A1(n9094), .A2(n9840), .ZN(n8285) );
  NAND2_X1 U6816 ( .A1(n8338), .A2(n8285), .ZN(n7195) );
  NAND2_X1 U6817 ( .A1(n9849), .A2(n9840), .ZN(n5307) );
  NAND2_X1 U6818 ( .A1(n5308), .A2(n5307), .ZN(n7291) );
  INV_X1 U6819 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6820 ( .A(n5309), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U6821 ( .A1(n5674), .A2(n7294), .ZN(n5314) );
  NAND2_X1 U6822 ( .A1(n6562), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5313) );
  OR2_X1 U6823 ( .A1(n5511), .A2(n4791), .ZN(n5312) );
  INV_X1 U6824 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5310) );
  OR2_X1 U6825 ( .A1(n5512), .A2(n5310), .ZN(n5311) );
  INV_X1 U6826 ( .A(n5315), .ZN(n5323) );
  INV_X1 U6827 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U6828 ( .A1(n8193), .A2(n6528), .ZN(n5322) );
  NAND2_X1 U6829 ( .A1(n5319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5320) );
  XNOR2_X1 U6830 ( .A(n5320), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9671) );
  NAND2_X1 U6831 ( .A1(n6610), .A2(n9671), .ZN(n5321) );
  NAND2_X1 U6832 ( .A1(n9836), .A2(n9847), .ZN(n9777) );
  INV_X2 U6833 ( .A(n9836), .ZN(n9781) );
  NAND2_X1 U6834 ( .A1(n9836), .A2(n7300), .ZN(n5324) );
  NAND2_X1 U6835 ( .A1(n6562), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5332) );
  INV_X1 U6836 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6837 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5325) );
  NAND2_X1 U6838 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  AND2_X1 U6839 ( .A1(n5351), .A2(n5327), .ZN(n9786) );
  NAND2_X1 U6840 ( .A1(n5674), .A2(n9786), .ZN(n5331) );
  INV_X1 U6841 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6615) );
  OR2_X1 U6842 ( .A1(n5511), .A2(n6615), .ZN(n5330) );
  INV_X1 U6843 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6844 ( .A1(n5512), .A2(n5328), .ZN(n5329) );
  XNOR2_X1 U6845 ( .A(n5334), .B(n5333), .ZN(n6533) );
  NAND2_X1 U6846 ( .A1(n6533), .A2(n8193), .ZN(n5341) );
  NAND2_X1 U6847 ( .A1(n5335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5336) );
  MUX2_X1 U6848 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5336), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5339) );
  INV_X1 U6849 ( .A(n5337), .ZN(n5338) );
  AND2_X1 U6850 ( .A1(n5339), .A2(n5338), .ZN(n6635) );
  AOI22_X1 U6851 ( .A1(n5315), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6610), .B2(
        n6635), .ZN(n5340) );
  NAND2_X1 U6852 ( .A1(n9848), .A2(n9784), .ZN(n8289) );
  INV_X1 U6853 ( .A(n9784), .ZN(n9860) );
  NAND2_X1 U6854 ( .A1(n9865), .A2(n9860), .ZN(n8108) );
  XNOR2_X1 U6855 ( .A(n5344), .B(n5343), .ZN(n6536) );
  NAND2_X1 U6856 ( .A1(n6536), .A2(n8193), .ZN(n5349) );
  NOR2_X1 U6857 ( .A1(n5337), .A2(n9534), .ZN(n5345) );
  MUX2_X1 U6858 ( .A(n9534), .B(n5345), .S(P1_IR_REG_6__SCAN_IN), .Z(n5347) );
  OR2_X1 U6859 ( .A1(n5347), .A2(n5346), .ZN(n9697) );
  INV_X1 U6860 ( .A(n9697), .ZN(n6637) );
  AOI22_X1 U6861 ( .A1(n5627), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6610), .B2(
        n6637), .ZN(n5348) );
  NAND2_X1 U6862 ( .A1(n5350), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6863 ( .A1(n6563), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5355) );
  INV_X1 U6864 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U6865 ( .A1(n5351), .A2(n7241), .ZN(n5352) );
  AND2_X1 U6866 ( .A1(n5364), .A2(n5352), .ZN(n7246) );
  NAND2_X1 U6867 ( .A1(n5674), .A2(n7246), .ZN(n5354) );
  NAND2_X1 U6868 ( .A1(n6562), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5353) );
  NAND4_X1 U6869 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n9782)
         );
  NAND2_X1 U6870 ( .A1(n7209), .A2(n9782), .ZN(n8283) );
  INV_X1 U6871 ( .A(n7209), .ZN(n7238) );
  NAND2_X1 U6872 ( .A1(n8283), .A2(n8286), .ZN(n8219) );
  NAND2_X1 U6873 ( .A1(n7208), .A2(n8219), .ZN(n7207) );
  OR2_X1 U6874 ( .A1(n9782), .A2(n7238), .ZN(n5357) );
  NAND2_X1 U6875 ( .A1(n7207), .A2(n5357), .ZN(n7397) );
  XNOR2_X1 U6876 ( .A(n5359), .B(n5358), .ZN(n6540) );
  NAND2_X1 U6877 ( .A1(n6540), .A2(n8193), .ZN(n5362) );
  OR2_X1 U6878 ( .A1(n5346), .A2(n9534), .ZN(n5360) );
  AOI22_X1 U6879 ( .A1(n5627), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6610), .B2(
        n9113), .ZN(n5361) );
  NAND2_X1 U6880 ( .A1(n5362), .A2(n5361), .ZN(n9879) );
  NAND2_X1 U6881 ( .A1(n6562), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5370) );
  INV_X1 U6882 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6883 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  AND2_X1 U6884 ( .A1(n5380), .A2(n5365), .ZN(n7401) );
  NAND2_X1 U6885 ( .A1(n5674), .A2(n7401), .ZN(n5369) );
  OR2_X1 U6886 ( .A1(n5511), .A2(n4798), .ZN(n5368) );
  INV_X1 U6887 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5366) );
  OR2_X1 U6888 ( .A1(n5512), .A2(n5366), .ZN(n5367) );
  OR2_X1 U6889 ( .A1(n9879), .A2(n9887), .ZN(n8284) );
  NAND2_X1 U6890 ( .A1(n9879), .A2(n9887), .ZN(n8273) );
  NAND2_X1 U6891 ( .A1(n8284), .A2(n8273), .ZN(n8218) );
  OR2_X1 U6892 ( .A1(n9879), .A2(n9864), .ZN(n5371) );
  XNOR2_X1 U6893 ( .A(n5374), .B(n5373), .ZN(n6543) );
  NAND2_X1 U6894 ( .A1(n6543), .A2(n8193), .ZN(n5378) );
  NAND2_X1 U6895 ( .A1(n5346), .A2(n5375), .ZN(n5390) );
  NAND2_X1 U6896 ( .A1(n5390), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5376) );
  XNOR2_X1 U6897 ( .A(n5376), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U6898 ( .A1(n5627), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6610), .B2(
        n6847), .ZN(n5377) );
  NAND2_X1 U6899 ( .A1(n6562), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5386) );
  INV_X1 U6900 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6901 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  AND2_X1 U6902 ( .A1(n5395), .A2(n5381), .ZN(n7418) );
  NAND2_X1 U6903 ( .A1(n5674), .A2(n7418), .ZN(n5385) );
  INV_X1 U6904 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7123) );
  OR2_X1 U6905 ( .A1(n5511), .A2(n7123), .ZN(n5384) );
  INV_X1 U6906 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5382) );
  OR2_X1 U6907 ( .A1(n5512), .A2(n5382), .ZN(n5383) );
  NAND2_X1 U6908 ( .A1(n9893), .A2(n9875), .ZN(n8274) );
  AND2_X1 U6909 ( .A1(n8255), .A2(n8274), .ZN(n8223) );
  INV_X1 U6910 ( .A(n9875), .ZN(n9093) );
  NAND2_X1 U6911 ( .A1(n9893), .A2(n9093), .ZN(n5388) );
  XNOR2_X1 U6912 ( .A(n5389), .B(n5079), .ZN(n6558) );
  NAND2_X1 U6913 ( .A1(n6558), .A2(n8193), .ZN(n5393) );
  NAND2_X1 U6914 ( .A1(n5469), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5391) );
  XNOR2_X1 U6915 ( .A(n5391), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U6916 ( .A1(n5627), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6610), .B2(
        n9707), .ZN(n5392) );
  NAND2_X1 U6917 ( .A1(n5393), .A2(n5392), .ZN(n9769) );
  NAND2_X1 U6918 ( .A1(n6563), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6919 ( .A1(n6562), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6920 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  AND2_X1 U6921 ( .A1(n5410), .A2(n5396), .ZN(n9756) );
  NAND2_X1 U6922 ( .A1(n5674), .A2(n9756), .ZN(n5398) );
  NAND2_X1 U6923 ( .A1(n5350), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5397) );
  NAND4_X1 U6924 ( .A1(n5400), .A2(n5399), .A3(n5398), .A4(n5397), .ZN(n9092)
         );
  OR2_X1 U6925 ( .A1(n9769), .A2(n9092), .ZN(n5402) );
  AND2_X1 U6926 ( .A1(n9769), .A2(n9092), .ZN(n5401) );
  NAND2_X1 U6927 ( .A1(n6572), .A2(n8193), .ZN(n5409) );
  NAND2_X1 U6928 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5434) );
  INV_X1 U6929 ( .A(n5434), .ZN(n5405) );
  NAND2_X1 U6930 ( .A1(n5405), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5407) );
  INV_X1 U6931 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6932 ( .A1(n5434), .A2(n5406), .ZN(n5420) );
  AOI22_X1 U6933 ( .A1(n5627), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6610), .B2(
        n6850), .ZN(n5408) );
  NAND2_X1 U6934 ( .A1(n6562), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6935 ( .A1(n5410), .A2(n7495), .ZN(n5411) );
  AND2_X1 U6936 ( .A1(n5425), .A2(n5411), .ZN(n7496) );
  NAND2_X1 U6937 ( .A1(n5674), .A2(n7496), .ZN(n5415) );
  INV_X1 U6938 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7340) );
  OR2_X1 U6939 ( .A1(n5511), .A2(n7340), .ZN(n5414) );
  INV_X1 U6940 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5412) );
  OR2_X1 U6941 ( .A1(n5512), .A2(n5412), .ZN(n5413) );
  OR2_X1 U6942 ( .A1(n7501), .A2(n9762), .ZN(n8123) );
  NAND2_X1 U6943 ( .A1(n7501), .A2(n9762), .ZN(n8119) );
  NAND2_X1 U6944 ( .A1(n8123), .A2(n8119), .ZN(n7337) );
  OR2_X1 U6945 ( .A1(n7501), .A2(n9091), .ZN(n5417) );
  XNOR2_X1 U6946 ( .A(n5419), .B(n5418), .ZN(n6570) );
  NAND2_X1 U6947 ( .A1(n6570), .A2(n8193), .ZN(n5423) );
  NAND2_X1 U6948 ( .A1(n5420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5421) );
  XNOR2_X1 U6949 ( .A(n5421), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U6950 ( .A1(n5627), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6610), .B2(
        n6997), .ZN(n5422) );
  NAND2_X1 U6951 ( .A1(n6564), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5430) );
  INV_X1 U6952 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9622) );
  OR2_X1 U6953 ( .A1(n5511), .A2(n9622), .ZN(n5429) );
  INV_X1 U6954 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6955 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  AND2_X1 U6956 ( .A1(n5441), .A2(n5426), .ZN(n9620) );
  NAND2_X1 U6957 ( .A1(n5674), .A2(n9620), .ZN(n5428) );
  NAND2_X1 U6958 ( .A1(n6562), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5427) );
  NAND4_X1 U6959 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n9090)
         );
  NAND2_X1 U6960 ( .A1(n9634), .A2(n9090), .ZN(n8126) );
  OR2_X1 U6961 ( .A1(n9634), .A2(n9090), .ZN(n8127) );
  INV_X1 U6962 ( .A(n7530), .ZN(n5450) );
  NAND2_X1 U6963 ( .A1(n6595), .A2(n5281), .ZN(n5439) );
  NOR2_X1 U6964 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5467) );
  OR2_X1 U6965 ( .A1(n5467), .A2(n9534), .ZN(n5433) );
  INV_X1 U6966 ( .A(n5436), .ZN(n5435) );
  NAND2_X1 U6967 ( .A1(n5435), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6968 ( .A1(n5436), .A2(n10234), .ZN(n5453) );
  AOI22_X1 U6969 ( .A1(n5627), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6610), .B2(
        n7139), .ZN(n5438) );
  INV_X1 U6970 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6971 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  AND2_X1 U6972 ( .A1(n5458), .A2(n5442), .ZN(n7625) );
  NAND2_X1 U6973 ( .A1(n5674), .A2(n7625), .ZN(n5448) );
  NAND2_X1 U6974 ( .A1(n6562), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5447) );
  INV_X1 U6975 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5443) );
  OR2_X1 U6976 ( .A1(n5511), .A2(n5443), .ZN(n5446) );
  INV_X1 U6977 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5444) );
  OR2_X1 U6978 ( .A1(n5512), .A2(n5444), .ZN(n5445) );
  OR2_X1 U6979 ( .A1(n7618), .A2(n9627), .ZN(n8129) );
  NAND2_X1 U6980 ( .A1(n7618), .A2(n9627), .ZN(n8258) );
  NAND2_X1 U6981 ( .A1(n7618), .A2(n9606), .ZN(n5451) );
  XNOR2_X1 U6982 ( .A(n5452), .B(n4502), .ZN(n6800) );
  NAND2_X1 U6983 ( .A1(n6800), .A2(n5281), .ZN(n5456) );
  NAND2_X1 U6984 ( .A1(n5453), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5454) );
  XNOR2_X1 U6985 ( .A(n5454), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7451) );
  AOI22_X1 U6986 ( .A1(n6610), .A2(n7451), .B1(n5627), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6987 ( .A1(n6564), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6988 ( .A1(n6563), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6989 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  AND2_X1 U6990 ( .A1(n5477), .A2(n5459), .ZN(n9597) );
  NAND2_X1 U6991 ( .A1(n5674), .A2(n9597), .ZN(n5461) );
  NAND2_X1 U6992 ( .A1(n6562), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5460) );
  NAND4_X1 U6993 ( .A1(n5463), .A2(n5462), .A3(n5461), .A4(n5460), .ZN(n9089)
         );
  XNOR2_X1 U6994 ( .A(n5465), .B(n5464), .ZN(n6798) );
  NAND2_X1 U6995 ( .A1(n6798), .A2(n8193), .ZN(n5475) );
  INV_X1 U6996 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5466) );
  INV_X1 U6997 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U6998 ( .A1(n5467), .A2(n10234), .A3(n5466), .A4(n10437), .ZN(n5468) );
  NOR2_X1 U6999 ( .A1(n5469), .A2(n5468), .ZN(n5472) );
  OR2_X1 U7000 ( .A1(n5472), .A2(n9534), .ZN(n5470) );
  INV_X1 U7001 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5471) );
  MUX2_X1 U7002 ( .A(n5470), .B(P1_IR_REG_31__SCAN_IN), .S(n5471), .Z(n5473)
         );
  NAND2_X1 U7003 ( .A1(n5472), .A2(n5471), .ZN(n5503) );
  AOI22_X1 U7004 ( .A1(n5627), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6610), .B2(
        n7685), .ZN(n5474) );
  NAND2_X1 U7005 ( .A1(n6564), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U7006 ( .A1(n6563), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5481) );
  INV_X1 U7007 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7008 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  AND2_X1 U7009 ( .A1(n5493), .A2(n5478), .ZN(n8957) );
  NAND2_X1 U7010 ( .A1(n5674), .A2(n8957), .ZN(n5480) );
  NAND2_X1 U7011 ( .A1(n6562), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5479) );
  NAND4_X1 U7012 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n9605)
         );
  AND2_X1 U7013 ( .A1(n8962), .A2(n9605), .ZN(n5483) );
  XNOR2_X1 U7014 ( .A(n5485), .B(n5484), .ZN(n6986) );
  NAND2_X1 U7015 ( .A1(n6986), .A2(n8193), .ZN(n5491) );
  NAND2_X1 U7016 ( .A1(n5503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5487) );
  XNOR2_X1 U7017 ( .A(n5487), .B(n5486), .ZN(n7697) );
  OAI22_X1 U7018 ( .A1(n5323), .A2(n10393), .B1(n7697), .B2(n5488), .ZN(n5489)
         );
  INV_X1 U7019 ( .A(n5489), .ZN(n5490) );
  NAND2_X1 U7020 ( .A1(n6563), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7021 ( .A1(n6562), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7022 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  AND2_X1 U7023 ( .A1(n5508), .A2(n5494), .ZN(n9075) );
  NAND2_X1 U7024 ( .A1(n5674), .A2(n9075), .ZN(n5496) );
  NAND2_X1 U7025 ( .A1(n6564), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5495) );
  NAND4_X1 U7026 ( .A1(n5498), .A2(n5497), .A3(n5496), .A4(n5495), .ZN(n9458)
         );
  NAND2_X1 U7027 ( .A1(n9083), .A2(n9458), .ZN(n5499) );
  NAND2_X1 U7028 ( .A1(n5500), .A2(n5499), .ZN(n9349) );
  XNOR2_X1 U7029 ( .A(n5502), .B(n5501), .ZN(n7043) );
  NAND2_X1 U7030 ( .A1(n7043), .A2(n8193), .ZN(n5506) );
  NAND2_X1 U7031 ( .A1(n5504), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5522) );
  XNOR2_X1 U7032 ( .A(n5522), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8076) );
  AOI22_X1 U7033 ( .A1(n5627), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8076), .B2(
        n6610), .ZN(n5505) );
  INV_X1 U7034 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7035 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  AND2_X1 U7036 ( .A1(n5528), .A2(n5509), .ZN(n9351) );
  NAND2_X1 U7037 ( .A1(n9351), .A2(n5674), .ZN(n5516) );
  NAND2_X1 U7038 ( .A1(n6562), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5515) );
  INV_X1 U7039 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5510) );
  OR2_X1 U7040 ( .A1(n5511), .A2(n5510), .ZN(n5514) );
  INV_X1 U7041 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9523) );
  OR2_X1 U7042 ( .A1(n5512), .A2(n9523), .ZN(n5513) );
  OR2_X1 U7043 ( .A1(n9364), .A2(n9080), .ZN(n8270) );
  NAND2_X1 U7044 ( .A1(n9364), .A2(n9080), .ZN(n8249) );
  NAND2_X1 U7045 ( .A1(n8270), .A2(n8249), .ZN(n9346) );
  NAND2_X1 U7046 ( .A1(n9349), .A2(n9346), .ZN(n5518) );
  INV_X1 U7047 ( .A(n9080), .ZN(n9341) );
  NAND2_X1 U7048 ( .A1(n9364), .A2(n9341), .ZN(n5517) );
  XNOR2_X1 U7049 ( .A(n5520), .B(n5519), .ZN(n7046) );
  NAND2_X1 U7050 ( .A1(n7046), .A2(n8193), .ZN(n5527) );
  NAND2_X1 U7051 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  NAND2_X1 U7052 ( .A1(n5523), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7053 ( .A1(n5524), .A2(n10430), .ZN(n5539) );
  OR2_X1 U7054 ( .A1(n5524), .A2(n10430), .ZN(n5525) );
  AOI22_X1 U7055 ( .A1(n9121), .A2(n6610), .B1(n5627), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7056 ( .A1(n5528), .A2(n9016), .ZN(n5529) );
  NAND2_X1 U7057 ( .A1(n5545), .A2(n5529), .ZN(n9334) );
  NAND2_X1 U7058 ( .A1(n6563), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7059 ( .A1(n6564), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5530) );
  AND2_X1 U7060 ( .A1(n5531), .A2(n5530), .ZN(n5533) );
  NAND2_X1 U7061 ( .A1(n6562), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5532) );
  OAI211_X1 U7062 ( .C1(n9334), .C2(n5659), .A(n5533), .B(n5532), .ZN(n9459)
         );
  OR2_X1 U7063 ( .A1(n9453), .A2(n9459), .ZN(n5534) );
  NAND2_X1 U7064 ( .A1(n9332), .A2(n5534), .ZN(n5536) );
  NAND2_X1 U7065 ( .A1(n9453), .A2(n9459), .ZN(n5535) );
  NAND2_X1 U7066 ( .A1(n5536), .A2(n5535), .ZN(n9318) );
  XNOR2_X1 U7067 ( .A(n5538), .B(n5537), .ZN(n7226) );
  NAND2_X1 U7068 ( .A1(n7226), .A2(n8193), .ZN(n5543) );
  NAND2_X1 U7069 ( .A1(n5539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5540) );
  XNOR2_X1 U7070 ( .A(n5540), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8077) );
  INV_X1 U7071 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10389) );
  NOR2_X1 U7072 ( .A1(n5323), .A2(n10389), .ZN(n5541) );
  AOI21_X1 U7073 ( .B1(n8077), .B2(n6610), .A(n5541), .ZN(n5542) );
  INV_X1 U7074 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7075 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  NAND2_X1 U7076 ( .A1(n5562), .A2(n5546), .ZN(n9319) );
  OR2_X1 U7077 ( .A1(n9319), .A2(n5659), .ZN(n5549) );
  AOI22_X1 U7078 ( .A1(n6562), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6563), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7079 ( .A1(n6564), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5547) );
  OR2_X1 U7080 ( .A1(n9329), .A2(n6433), .ZN(n8152) );
  NAND2_X1 U7081 ( .A1(n9329), .A2(n6433), .ZN(n8253) );
  NAND2_X1 U7082 ( .A1(n8152), .A2(n8253), .ZN(n9317) );
  NAND2_X1 U7083 ( .A1(n9318), .A2(n9317), .ZN(n5551) );
  INV_X1 U7084 ( .A(n6433), .ZN(n9435) );
  NAND2_X1 U7085 ( .A1(n9329), .A2(n9435), .ZN(n5550) );
  NAND2_X1 U7086 ( .A1(n5551), .A2(n5550), .ZN(n9305) );
  XNOR2_X1 U7087 ( .A(n5553), .B(n5552), .ZN(n7314) );
  NAND2_X1 U7088 ( .A1(n7314), .A2(n8193), .ZN(n5560) );
  NAND2_X1 U7089 ( .A1(n5554), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5555) );
  MUX2_X1 U7090 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5555), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5558) );
  AOI22_X1 U7091 ( .A1(n5627), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6610), .B2(
        n9789), .ZN(n5559) );
  NAND2_X1 U7092 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  AND2_X1 U7093 ( .A1(n5576), .A2(n5563), .ZN(n9306) );
  NAND2_X1 U7094 ( .A1(n9306), .A2(n5674), .ZN(n5568) );
  INV_X1 U7095 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U7096 ( .A1(n6564), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7097 ( .A1(n6563), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5564) );
  OAI211_X1 U7098 ( .C1(n9442), .C2(n5721), .A(n5565), .B(n5564), .ZN(n5566)
         );
  INV_X1 U7099 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7100 ( .A1(n5568), .A2(n5567), .ZN(n9444) );
  AND2_X1 U7101 ( .A1(n9434), .A2(n9444), .ZN(n5570) );
  OR2_X1 U7102 ( .A1(n9434), .A2(n9444), .ZN(n5569) );
  NAND2_X1 U7103 ( .A1(n7444), .A2(n8193), .ZN(n5574) );
  NAND2_X1 U7104 ( .A1(n5627), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5573) );
  INV_X1 U7105 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7106 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  NAND2_X1 U7107 ( .A1(n5589), .A2(n5577), .ZN(n9296) );
  OR2_X1 U7108 ( .A1(n9296), .A2(n5659), .ZN(n5582) );
  INV_X1 U7109 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U7110 ( .A1(n6564), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7111 ( .A1(n6563), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5578) );
  OAI211_X1 U7112 ( .C1(n9432), .C2(n5721), .A(n5579), .B(n5578), .ZN(n5580)
         );
  INV_X1 U7113 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7114 ( .A1(n5582), .A2(n5581), .ZN(n9436) );
  NOR2_X1 U7115 ( .A1(n9295), .A2(n9436), .ZN(n5584) );
  NAND2_X1 U7116 ( .A1(n9295), .A2(n9436), .ZN(n5583) );
  OAI21_X1 U7117 ( .B1(n9287), .B2(n5584), .A(n5583), .ZN(n9275) );
  XNOR2_X1 U7118 ( .A(n5586), .B(n5585), .ZN(n7475) );
  NAND2_X1 U7119 ( .A1(n7475), .A2(n8193), .ZN(n5588) );
  NAND2_X1 U7120 ( .A1(n5627), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7121 ( .A1(n5589), .A2(n8983), .ZN(n5590) );
  NAND2_X1 U7122 ( .A1(n5602), .A2(n5590), .ZN(n9276) );
  OR2_X1 U7123 ( .A1(n9276), .A2(n5659), .ZN(n5595) );
  INV_X1 U7124 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U7125 ( .A1(n6563), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7126 ( .A1(n6564), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7127 ( .C1(n5721), .C2(n9427), .A(n5592), .B(n5591), .ZN(n5593)
         );
  INV_X1 U7128 ( .A(n5593), .ZN(n5594) );
  NAND2_X1 U7129 ( .A1(n9284), .A2(n9293), .ZN(n9254) );
  NAND2_X1 U7130 ( .A1(n8298), .A2(n9254), .ZN(n9274) );
  NAND2_X1 U7131 ( .A1(n9275), .A2(n9274), .ZN(n5597) );
  NAND2_X1 U7132 ( .A1(n9284), .A2(n9412), .ZN(n5596) );
  XNOR2_X1 U7133 ( .A(n5599), .B(n5598), .ZN(n7551) );
  NAND2_X1 U7134 ( .A1(n7551), .A2(n8193), .ZN(n5601) );
  NAND2_X1 U7135 ( .A1(n5627), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7136 ( .A1(n5602), .A2(n9040), .ZN(n5603) );
  NAND2_X1 U7137 ( .A1(n5616), .A2(n5603), .ZN(n9259) );
  INV_X1 U7138 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U7139 ( .A1(n6564), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7140 ( .A1(n6563), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5604) );
  OAI211_X1 U7141 ( .C1(n9419), .C2(n5721), .A(n5605), .B(n5604), .ZN(n5606)
         );
  INV_X1 U7142 ( .A(n5606), .ZN(n5607) );
  OR2_X1 U7143 ( .A1(n9267), .A2(n9421), .ZN(n5608) );
  OR2_X1 U7144 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  NAND2_X1 U7145 ( .A1(n5612), .A2(n5611), .ZN(n7552) );
  NAND2_X1 U7146 ( .A1(n7552), .A2(n8193), .ZN(n5614) );
  NAND2_X1 U7147 ( .A1(n5627), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5613) );
  NAND2_X2 U7148 ( .A1(n5614), .A2(n5613), .ZN(n9409) );
  INV_X1 U7149 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7150 ( .A1(n5616), .A2(n5615), .ZN(n5617) );
  NAND2_X1 U7151 ( .A1(n5631), .A2(n5617), .ZN(n9247) );
  OR2_X1 U7152 ( .A1(n9247), .A2(n5659), .ZN(n5623) );
  INV_X1 U7153 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7154 ( .A1(n6563), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7155 ( .A1(n6564), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5618) );
  OAI211_X1 U7156 ( .C1(n5620), .C2(n5721), .A(n5619), .B(n5618), .ZN(n5621)
         );
  INV_X1 U7157 ( .A(n5621), .ZN(n5622) );
  NOR2_X1 U7158 ( .A1(n9409), .A2(n9413), .ZN(n5624) );
  NAND2_X1 U7159 ( .A1(n7613), .A2(n8193), .ZN(n5629) );
  NAND2_X1 U7160 ( .A1(n5627), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5628) );
  NAND2_X2 U7161 ( .A1(n5629), .A2(n5628), .ZN(n9228) );
  INV_X1 U7162 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7163 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  NAND2_X1 U7164 ( .A1(n5643), .A2(n5632), .ZN(n9229) );
  INV_X1 U7165 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U7166 ( .A1(n6563), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7167 ( .A1(n6564), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5633) );
  OAI211_X1 U7168 ( .C1(n5721), .C2(n9405), .A(n5634), .B(n5633), .ZN(n5635)
         );
  INV_X1 U7169 ( .A(n5635), .ZN(n5636) );
  AND2_X1 U7170 ( .A1(n9228), .A2(n9242), .ZN(n5638) );
  XNOR2_X1 U7171 ( .A(n5640), .B(n5639), .ZN(n7716) );
  NAND2_X1 U7172 ( .A1(n7716), .A2(n8193), .ZN(n5642) );
  NAND2_X1 U7173 ( .A1(n5627), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5641) );
  NAND2_X2 U7174 ( .A1(n5642), .A2(n5641), .ZN(n9394) );
  NAND2_X1 U7175 ( .A1(n5643), .A2(n8991), .ZN(n5644) );
  NAND2_X1 U7176 ( .A1(n9211), .A2(n5284), .ZN(n5650) );
  INV_X1 U7177 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7178 ( .A1(n6564), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7179 ( .A1(n6563), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5645) );
  OAI211_X1 U7180 ( .C1(n5647), .C2(n5721), .A(n5646), .B(n5645), .ZN(n5648)
         );
  INV_X1 U7181 ( .A(n5648), .ZN(n5649) );
  OR2_X2 U7182 ( .A1(n9394), .A2(n9398), .ZN(n8311) );
  NAND2_X1 U7183 ( .A1(n9394), .A2(n9398), .ZN(n8178) );
  NAND2_X1 U7184 ( .A1(n8311), .A2(n8178), .ZN(n9215) );
  OR2_X1 U7185 ( .A1(n9394), .A2(n9196), .ZN(n5651) );
  NAND2_X1 U7186 ( .A1(n7749), .A2(n8193), .ZN(n5655) );
  NAND2_X1 U7187 ( .A1(n5627), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5654) );
  INV_X1 U7188 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7189 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U7190 ( .A1(n5673), .A2(n5658), .ZN(n9060) );
  INV_X1 U7191 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U7192 ( .A1(n6564), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7193 ( .A1(n6563), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5660) );
  OAI211_X1 U7194 ( .C1(n9391), .C2(n5721), .A(n5661), .B(n5660), .ZN(n5662)
         );
  INV_X1 U7195 ( .A(n5662), .ZN(n5663) );
  NOR2_X1 U7196 ( .A1(n9201), .A2(n9216), .ZN(n5665) );
  NAND2_X1 U7197 ( .A1(n9201), .A2(n9216), .ZN(n5666) );
  INV_X1 U7198 ( .A(n9176), .ZN(n5682) );
  NAND2_X1 U7199 ( .A1(n5668), .A2(n5667), .ZN(n5670) );
  NAND2_X1 U7200 ( .A1(n5670), .A2(n5669), .ZN(n8945) );
  NAND2_X1 U7201 ( .A1(n8945), .A2(n8193), .ZN(n5672) );
  NAND2_X1 U7202 ( .A1(n5627), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5671) );
  XNOR2_X1 U7203 ( .A(n5673), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U7204 ( .A1(n9186), .A2(n5674), .ZN(n5680) );
  INV_X1 U7205 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7206 ( .A1(n6563), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7207 ( .A1(n6564), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5675) );
  OAI211_X1 U7208 ( .C1(n5721), .C2(n5677), .A(n5676), .B(n5675), .ZN(n5678)
         );
  INV_X1 U7209 ( .A(n5678), .ZN(n5679) );
  NAND2_X1 U7210 ( .A1(n9385), .A2(n9199), .ZN(n8317) );
  INV_X1 U7211 ( .A(n9178), .ZN(n5681) );
  OR2_X1 U7212 ( .A1(n9385), .A2(n9164), .ZN(n5683) );
  NAND2_X1 U7213 ( .A1(n9167), .A2(n9182), .ZN(n8318) );
  NAND2_X1 U7214 ( .A1(n5689), .A2(n5726), .ZN(n5684) );
  NAND2_X1 U7215 ( .A1(n8386), .A2(n9814), .ZN(n6276) );
  OR2_X1 U7216 ( .A1(n5686), .A2(n10434), .ZN(n5687) );
  NAND2_X2 U7217 ( .A1(n8332), .A2(n7446), .ZN(n6497) );
  MUX2_X1 U7218 ( .A(n6276), .B(n6498), .S(n6497), .Z(n9812) );
  OR2_X1 U7219 ( .A1(n8200), .A2(n4481), .ZN(n9896) );
  INV_X1 U7220 ( .A(n9394), .ZN(n9213) );
  NAND2_X1 U7221 ( .A1(n9793), .A2(n9832), .ZN(n7199) );
  NAND2_X1 U7222 ( .A1(n9774), .A2(n7209), .ZN(n7400) );
  OR2_X1 U7223 ( .A1(n7400), .A2(n9879), .ZN(n7398) );
  INV_X1 U7224 ( .A(n9769), .ZN(n9903) );
  AND2_X1 U7225 ( .A1(n9751), .A2(n9903), .ZN(n9752) );
  INV_X1 U7226 ( .A(n7501), .ZN(n7371) );
  NAND2_X1 U7227 ( .A1(n9752), .A2(n7371), .ZN(n9616) );
  INV_X1 U7228 ( .A(n9453), .ZN(n9338) );
  NAND2_X1 U7229 ( .A1(n9333), .A2(n9520), .ZN(n9325) );
  NAND2_X1 U7230 ( .A1(n9200), .A2(n9189), .ZN(n9183) );
  AOI21_X1 U7231 ( .B1(n8307), .B2(n9168), .A(n9615), .ZN(n5692) );
  AND2_X1 U7232 ( .A1(n5692), .A2(n9136), .ZN(n9149) );
  INV_X1 U7233 ( .A(n7012), .ZN(n9796) );
  AND4_X1 U7234 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n8334)
         );
  NAND2_X1 U7235 ( .A1(n8334), .A2(n8333), .ZN(n5697) );
  NAND2_X1 U7236 ( .A1(n9805), .A2(n5697), .ZN(n7036) );
  AND2_X1 U7237 ( .A1(n8289), .A2(n9777), .ZN(n7213) );
  AND2_X1 U7238 ( .A1(n7213), .A2(n8286), .ZN(n8344) );
  NAND2_X1 U7239 ( .A1(n9778), .A2(n8344), .ZN(n5700) );
  INV_X1 U7240 ( .A(n8108), .ZN(n5698) );
  NAND2_X1 U7241 ( .A1(n8286), .A2(n5698), .ZN(n8345) );
  AND2_X1 U7242 ( .A1(n8345), .A2(n8283), .ZN(n5699) );
  INV_X1 U7243 ( .A(n8273), .ZN(n5701) );
  INV_X1 U7244 ( .A(n9092), .ZN(n9889) );
  OR2_X1 U7245 ( .A1(n9769), .A2(n9889), .ZN(n8212) );
  NAND2_X1 U7246 ( .A1(n8123), .A2(n8212), .ZN(n8256) );
  NAND2_X1 U7247 ( .A1(n9769), .A2(n9889), .ZN(n8211) );
  NAND2_X1 U7248 ( .A1(n8119), .A2(n8211), .ZN(n8124) );
  NAND2_X1 U7249 ( .A1(n8124), .A2(n8123), .ZN(n9623) );
  INV_X1 U7250 ( .A(n9090), .ZN(n7499) );
  NAND2_X1 U7251 ( .A1(n9634), .A2(n7499), .ZN(n8130) );
  AND2_X1 U7252 ( .A1(n9623), .A2(n8130), .ZN(n8257) );
  OR2_X1 U7253 ( .A1(n9634), .A2(n7499), .ZN(n5704) );
  NAND2_X1 U7254 ( .A1(n5703), .A2(n5704), .ZN(n7533) );
  NAND2_X1 U7255 ( .A1(n7533), .A2(n8227), .ZN(n5707) );
  INV_X1 U7256 ( .A(n5704), .ZN(n5705) );
  NAND2_X1 U7257 ( .A1(n8258), .A2(n5705), .ZN(n5706) );
  AND2_X1 U7258 ( .A1(n5706), .A2(n8129), .ZN(n8261) );
  OR2_X1 U7259 ( .A1(n9637), .A2(n9474), .ZN(n8134) );
  NAND2_X1 U7260 ( .A1(n9637), .A2(n9474), .ZN(n8260) );
  NAND2_X1 U7261 ( .A1(n8134), .A2(n8260), .ZN(n9600) );
  INV_X1 U7262 ( .A(n9605), .ZN(n8135) );
  XNOR2_X1 U7263 ( .A(n8962), .B(n8135), .ZN(n8229) );
  OR2_X1 U7264 ( .A1(n8962), .A2(n8135), .ZN(n8139) );
  INV_X1 U7265 ( .A(n9458), .ZN(n8960) );
  NAND2_X1 U7266 ( .A1(n9083), .A2(n8960), .ZN(n8265) );
  AND2_X1 U7267 ( .A1(n9528), .A2(n9458), .ZN(n8254) );
  NAND2_X1 U7268 ( .A1(n9347), .A2(n8270), .ZN(n5708) );
  INV_X1 U7269 ( .A(n9459), .ZN(n9356) );
  AND2_X1 U7270 ( .A1(n9453), .A2(n9356), .ZN(n8251) );
  OR2_X1 U7271 ( .A1(n9453), .A2(n9356), .ZN(n8099) );
  INV_X1 U7272 ( .A(n9444), .ZN(n5709) );
  OR2_X1 U7273 ( .A1(n9434), .A2(n5709), .ZN(n8156) );
  NAND2_X1 U7274 ( .A1(n9434), .A2(n5709), .ZN(n8281) );
  INV_X1 U7275 ( .A(n8281), .ZN(n5710) );
  NAND2_X1 U7276 ( .A1(n9295), .A2(n9309), .ZN(n8153) );
  INV_X1 U7277 ( .A(n9270), .ZN(n5711) );
  NOR2_X1 U7278 ( .A1(n9274), .A2(n5711), .ZN(n5712) );
  INV_X1 U7279 ( .A(n9421), .ZN(n5713) );
  NAND2_X1 U7280 ( .A1(n9267), .A2(n5713), .ZN(n8210) );
  AND2_X1 U7281 ( .A1(n8210), .A2(n9254), .ZN(n8161) );
  INV_X1 U7282 ( .A(n9413), .ZN(n9263) );
  NAND2_X1 U7283 ( .A1(n9409), .A2(n9263), .ZN(n8166) );
  NAND2_X1 U7284 ( .A1(n9241), .A2(n9240), .ZN(n9239) );
  INV_X1 U7285 ( .A(n9242), .ZN(n8992) );
  XNOR2_X1 U7286 ( .A(n9228), .B(n8992), .ZN(n9224) );
  NAND2_X1 U7287 ( .A1(n9228), .A2(n8992), .ZN(n8165) );
  INV_X1 U7288 ( .A(n9216), .ZN(n8995) );
  OR2_X1 U7289 ( .A1(n9201), .A2(n8995), .ZN(n8310) );
  NAND2_X1 U7290 ( .A1(n9201), .A2(n8995), .ZN(n8316) );
  NAND2_X1 U7291 ( .A1(n9193), .A2(n8310), .ZN(n9179) );
  NAND2_X1 U7292 ( .A1(n9179), .A2(n9178), .ZN(n9177) );
  NAND2_X1 U7293 ( .A1(n9177), .A2(n8362), .ZN(n9162) );
  NAND2_X1 U7294 ( .A1(n9162), .A2(n9161), .ZN(n9160) );
  NAND2_X1 U7295 ( .A1(n9160), .A2(n8308), .ZN(n5714) );
  XNOR2_X1 U7296 ( .A(n5714), .B(n8238), .ZN(n5723) );
  NAND2_X1 U7297 ( .A1(n5716), .A2(n9789), .ZN(n5715) );
  NAND2_X1 U7298 ( .A1(n8332), .A2(n4481), .ZN(n8205) );
  INV_X1 U7299 ( .A(n8382), .ZN(n6872) );
  INV_X1 U7300 ( .A(n6608), .ZN(n8245) );
  INV_X1 U7301 ( .A(P1_B_REG_SCAN_IN), .ZN(n8385) );
  NOR2_X1 U7302 ( .A1(n8381), .A2(n8385), .ZN(n5718) );
  NOR2_X1 U7303 ( .A1(n9888), .A2(n5718), .ZN(n9139) );
  INV_X1 U7304 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U7305 ( .A1(n6563), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7306 ( .A1(n6564), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5719) );
  OAI211_X1 U7307 ( .C1(n5721), .C2(n9374), .A(n5720), .B(n5719), .ZN(n9087)
         );
  AOI22_X1 U7308 ( .A1(n9088), .A2(n9866), .B1(n9139), .B2(n9087), .ZN(n5722)
         );
  NAND2_X1 U7309 ( .A1(n5733), .A2(n5728), .ZN(n5729) );
  NAND2_X1 U7310 ( .A1(n7719), .A2(P1_B_REG_SCAN_IN), .ZN(n5734) );
  MUX2_X1 U7311 ( .A(n5734), .B(P1_B_REG_SCAN_IN), .S(n5738), .Z(n5737) );
  INV_X1 U7312 ( .A(n5753), .ZN(n7760) );
  INV_X1 U7313 ( .A(n5738), .ZN(n7617) );
  NAND2_X1 U7314 ( .A1(n7760), .A2(n7617), .ZN(n6548) );
  OAI21_X1 U7315 ( .B1(n6547), .B2(P1_D_REG_0__SCAN_IN), .A(n6548), .ZN(n5751)
         );
  INV_X1 U7316 ( .A(n6547), .ZN(n5749) );
  NOR4_X1 U7317 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5742) );
  NOR4_X1 U7318 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5741) );
  NOR4_X1 U7319 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5740) );
  NOR4_X1 U7320 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5739) );
  AND4_X1 U7321 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n5748)
         );
  NOR2_X1 U7322 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n5746) );
  NOR4_X1 U7323 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5745) );
  NOR4_X1 U7324 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5744) );
  NOR4_X1 U7325 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5743) );
  AND4_X1 U7326 ( .A1(n5746), .A2(n5745), .A3(n5744), .A4(n5743), .ZN(n5747)
         );
  NAND2_X1 U7327 ( .A1(n5748), .A2(n5747), .ZN(n6494) );
  NAND2_X1 U7328 ( .A1(n5749), .A2(n6494), .ZN(n5750) );
  NAND2_X1 U7329 ( .A1(n5751), .A2(n5750), .ZN(n5757) );
  NAND2_X2 U7330 ( .A1(n5753), .A2(n5752), .ZN(n6275) );
  NAND2_X1 U7331 ( .A1(n7446), .A2(n9814), .ZN(n8378) );
  NAND2_X1 U7332 ( .A1(n5754), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5755) );
  AOI21_X1 U7333 ( .B1(n6608), .B2(n8378), .A(n7555), .ZN(n5756) );
  NAND2_X1 U7334 ( .A1(n6275), .A2(n5756), .ZN(n6503) );
  NAND2_X1 U7335 ( .A1(n7760), .A2(n7719), .ZN(n6550) );
  OR2_X1 U7336 ( .A1(n7011), .A2(n7446), .ZN(n9797) );
  NAND2_X1 U7337 ( .A1(n9911), .A2(n9892), .ZN(n9532) );
  NAND2_X1 U7338 ( .A1(n5760), .A2(n5077), .ZN(P1_U3520) );
  NOR2_X1 U7339 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5764) );
  NAND4_X1 U7340 ( .A1(n5764), .A2(n5795), .A3(n6086), .A4(n5793), .ZN(n5767)
         );
  NAND4_X1 U7341 ( .A1(n6216), .A2(n6221), .A3(n6219), .A4(n5765), .ZN(n5766)
         );
  XNOR2_X2 U7342 ( .A(n5772), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8936) );
  INV_X1 U7343 ( .A(n5773), .ZN(n8932) );
  NAND2_X1 U7344 ( .A1(n5800), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5774) );
  MUX2_X1 U7345 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5774), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5775) );
  NOR2_X2 U7346 ( .A1(n8936), .A2(n5784), .ZN(n5849) );
  INV_X1 U7347 ( .A(n5849), .ZN(n5928) );
  NAND2_X1 U7348 ( .A1(n5975), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5788) );
  INV_X2 U7349 ( .A(n7843), .ZN(n7845) );
  NAND2_X1 U7350 ( .A1(n7845), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5787) );
  AND2_X2 U7351 ( .A1(n8936), .A2(n8938), .ZN(n5851) );
  NAND2_X1 U7352 ( .A1(n5881), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7353 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5776) );
  NOR2_X1 U7354 ( .A1(n5915), .A2(n5776), .ZN(n5929) );
  NAND2_X1 U7355 ( .A1(n5929), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7356 ( .A1(n5993), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7357 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5777) );
  NAND2_X1 U7358 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(n6104), .ZN(n6118) );
  INV_X1 U7359 ( .A(n6118), .ZN(n5778) );
  NAND2_X1 U7360 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n5778), .ZN(n6130) );
  INV_X1 U7361 ( .A(n6130), .ZN(n5779) );
  NAND2_X1 U7362 ( .A1(n5779), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6144) );
  INV_X1 U7363 ( .A(n6144), .ZN(n5780) );
  NAND2_X1 U7364 ( .A1(n5780), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6146) );
  INV_X1 U7365 ( .A(n6146), .ZN(n5781) );
  NAND2_X1 U7366 ( .A1(n5781), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5806) );
  INV_X1 U7367 ( .A(n5806), .ZN(n5782) );
  NAND2_X1 U7368 ( .A1(n5782), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6171) );
  INV_X1 U7369 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10400) );
  NAND2_X1 U7370 ( .A1(n5806), .A2(n10400), .ZN(n5783) );
  AND2_X1 U7371 ( .A1(n6171), .A2(n5783), .ZN(n8701) );
  NAND2_X1 U7372 ( .A1(n6261), .A2(n8701), .ZN(n5786) );
  AND2_X2 U7373 ( .A1(n8936), .A2(n5784), .ZN(n5848) );
  CLKBUF_X3 U7374 ( .A(n5848), .Z(n7844) );
  NAND2_X1 U7375 ( .A1(n7844), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7376 ( .A1(n5796), .A2(n5795), .ZN(n5789) );
  NAND2_X1 U7377 ( .A1(n5789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  MUX2_X1 U7378 ( .A(n7868), .B(n6831), .S(n7505), .Z(n5797) );
  INV_X2 U7379 ( .A(n5797), .ZN(n5844) );
  INV_X2 U7380 ( .A(n5847), .ZN(n5891) );
  NAND2_X1 U7381 ( .A1(n7613), .A2(n5891), .ZN(n5804) );
  NAND2_X1 U7382 ( .A1(n4487), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5803) );
  XOR2_X1 U7383 ( .A(n6157), .B(n8867), .Z(n8485) );
  NAND2_X1 U7384 ( .A1(n7845), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7385 ( .A1(n6024), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5809) );
  INV_X1 U7386 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U7387 ( .A1(n6146), .A2(n10211), .ZN(n5805) );
  AND2_X1 U7388 ( .A1(n5806), .A2(n5805), .ZN(n8718) );
  NAND2_X1 U7389 ( .A1(n6261), .A2(n8718), .ZN(n5808) );
  NAND2_X1 U7390 ( .A1(n7844), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5807) );
  OR2_X1 U7391 ( .A1(n8736), .A2(n7306), .ZN(n8482) );
  NAND2_X1 U7392 ( .A1(n5851), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7393 ( .A1(n5849), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7394 ( .A1(n5848), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7395 ( .A1(n5835), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5811) );
  INV_X1 U7396 ( .A(n6914), .ZN(n8551) );
  NAND2_X1 U7397 ( .A1(n7856), .A2(SI_0_), .ZN(n5816) );
  INV_X1 U7398 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7399 ( .A1(n5816), .A2(n5815), .ZN(n5818) );
  AND2_X1 U7400 ( .A1(n5818), .A2(n5817), .ZN(n8950) );
  MUX2_X1 U7401 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8950), .S(n5860), .Z(n9950) );
  NAND2_X1 U7402 ( .A1(n8551), .A2(n9950), .ZN(n8420) );
  INV_X1 U7403 ( .A(n8420), .ZN(n5819) );
  NAND2_X1 U7404 ( .A1(n5819), .A2(n7864), .ZN(n7308) );
  INV_X1 U7405 ( .A(n9950), .ZN(n7305) );
  NAND2_X1 U7406 ( .A1(n5797), .A2(n7305), .ZN(n5820) );
  NAND2_X1 U7407 ( .A1(n5851), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7408 ( .A1(n5849), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7409 ( .A1(n5835), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7410 ( .A1(n5848), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7411 ( .A1(n6912), .A2(n6936), .ZN(n5833) );
  NAND2_X1 U7412 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5825) );
  MUX2_X1 U7413 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5825), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5828) );
  NAND2_X1 U7414 ( .A1(n5828), .A2(n5827), .ZN(n6658) );
  INV_X1 U7415 ( .A(n6658), .ZN(n6679) );
  NAND2_X1 U7416 ( .A1(n6070), .A2(n6679), .ZN(n5832) );
  INV_X1 U7417 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5829) );
  XNOR2_X1 U7418 ( .A(n5844), .B(n6818), .ZN(n6938) );
  XNOR2_X1 U7419 ( .A(n5834), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6660) );
  XNOR2_X1 U7420 ( .A(n5844), .B(n6821), .ZN(n5841) );
  NAND2_X1 U7421 ( .A1(n5851), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7422 ( .A1(n5849), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7423 ( .A1(n5848), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7424 ( .A1(n5835), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5836) );
  OR2_X1 U7425 ( .A1(n6915), .A2(n7306), .ZN(n5840) );
  NAND2_X1 U7426 ( .A1(n5841), .A2(n5840), .ZN(n6934) );
  INV_X1 U7427 ( .A(n5840), .ZN(n5843) );
  INV_X1 U7428 ( .A(n5841), .ZN(n5842) );
  NAND2_X1 U7429 ( .A1(n5843), .A2(n5842), .ZN(n6935) );
  NAND2_X1 U7430 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4522), .ZN(n5845) );
  XNOR2_X1 U7431 ( .A(n5845), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U7432 ( .A1(n6070), .A2(n6729), .ZN(n5846) );
  XNOR2_X1 U7433 ( .A(n5844), .B(n8442), .ZN(n5857) );
  INV_X2 U7434 ( .A(n7843), .ZN(n6200) );
  NAND2_X1 U7435 ( .A1(n5848), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7436 ( .A1(n5849), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5853) );
  INV_X1 U7437 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7438 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  NAND3_X1 U7439 ( .A1(n5854), .A2(n5853), .A3(n5852), .ZN(n5855) );
  AOI21_X2 U7440 ( .B1(n6200), .B2(P2_REG0_REG_3__SCAN_IN), .A(n5855), .ZN(
        n6927) );
  OR2_X1 U7441 ( .A1(n6927), .A2(n7306), .ZN(n5856) );
  XNOR2_X1 U7442 ( .A(n5857), .B(n5856), .ZN(n8445) );
  INV_X1 U7443 ( .A(n5856), .ZN(n5858) );
  NAND2_X1 U7444 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  INV_X1 U7445 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6532) );
  OR2_X1 U7446 ( .A1(n5876), .A2(n5771), .ZN(n5861) );
  XNOR2_X1 U7447 ( .A(n5861), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6727) );
  INV_X1 U7448 ( .A(n6727), .ZN(n6765) );
  OAI22_X1 U7449 ( .A1(n6100), .A2(n6532), .B1(n5860), .B2(n6765), .ZN(n5862)
         );
  INV_X1 U7450 ( .A(n5862), .ZN(n5864) );
  NAND2_X1 U7451 ( .A1(n6528), .A2(n5891), .ZN(n5863) );
  INV_X2 U7452 ( .A(n9973), .ZN(n7070) );
  XNOR2_X1 U7453 ( .A(n6157), .B(n7070), .ZN(n5871) );
  NAND2_X1 U7454 ( .A1(n6024), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7455 ( .A1(n7844), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5868) );
  NOR2_X1 U7456 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5865) );
  NOR2_X1 U7457 ( .A1(n5881), .A2(n5865), .ZN(n6930) );
  NAND2_X1 U7458 ( .A1(n5851), .A2(n6930), .ZN(n5867) );
  NAND2_X1 U7459 ( .A1(n6200), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5866) );
  OR2_X1 U7460 ( .A1(n6964), .A2(n7306), .ZN(n5870) );
  NAND2_X1 U7461 ( .A1(n5871), .A2(n5870), .ZN(n7063) );
  NAND2_X1 U7462 ( .A1(n7065), .A2(n7063), .ZN(n5874) );
  INV_X1 U7463 ( .A(n5870), .ZN(n5873) );
  INV_X1 U7464 ( .A(n5871), .ZN(n5872) );
  NAND2_X1 U7465 ( .A1(n5873), .A2(n5872), .ZN(n7064) );
  NAND2_X1 U7466 ( .A1(n5874), .A2(n7064), .ZN(n6907) );
  NAND2_X1 U7467 ( .A1(n6533), .A2(n5891), .ZN(n5880) );
  INV_X1 U7468 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7469 ( .A1(n5876), .A2(n5875), .ZN(n5911) );
  NAND2_X1 U7470 ( .A1(n5911), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7471 ( .A1(n5877), .A2(n5909), .ZN(n5892) );
  OR2_X1 U7472 ( .A1(n5877), .A2(n5909), .ZN(n5878) );
  AOI22_X1 U7473 ( .A1(n4486), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6070), .B2(
        n6724), .ZN(n5879) );
  XNOR2_X1 U7474 ( .A(n8822), .B(n6157), .ZN(n5888) );
  NAND2_X1 U7475 ( .A1(n7845), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7476 ( .A1(n5975), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5884) );
  OAI21_X1 U7477 ( .B1(n5881), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5915), .ZN(
        n8820) );
  INV_X1 U7478 ( .A(n8820), .ZN(n6908) );
  NAND2_X1 U7479 ( .A1(n5851), .A2(n6908), .ZN(n5883) );
  NAND2_X1 U7480 ( .A1(n7844), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5882) );
  AND2_X1 U7481 ( .A1(n8547), .A2(n7864), .ZN(n5886) );
  XNOR2_X1 U7482 ( .A(n5888), .B(n5886), .ZN(n6906) );
  NAND2_X1 U7483 ( .A1(n6907), .A2(n6906), .ZN(n5890) );
  INV_X1 U7484 ( .A(n5886), .ZN(n5887) );
  OR2_X1 U7485 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  NAND2_X1 U7486 ( .A1(n6536), .A2(n5891), .ZN(n5896) );
  INV_X1 U7487 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U7488 ( .A1(n5892), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5893) );
  XNOR2_X1 U7489 ( .A(n5893), .B(n5908), .ZN(n6776) );
  OAI22_X1 U7490 ( .A1(n6100), .A2(n6539), .B1(n5860), .B2(n6776), .ZN(n5894)
         );
  INV_X1 U7491 ( .A(n5894), .ZN(n5895) );
  NAND2_X1 U7492 ( .A1(n5896), .A2(n5895), .ZN(n7155) );
  XNOR2_X1 U7493 ( .A(n7155), .B(n6211), .ZN(n5901) );
  NAND2_X1 U7494 ( .A1(n5975), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7495 ( .A1(n7844), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5899) );
  XNOR2_X1 U7496 ( .A(n5915), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n7152) );
  NAND2_X1 U7497 ( .A1(n5851), .A2(n7152), .ZN(n5898) );
  NAND2_X1 U7498 ( .A1(n7845), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5897) );
  OR2_X1 U7499 ( .A1(n7110), .A2(n7306), .ZN(n5902) );
  NAND2_X1 U7500 ( .A1(n5901), .A2(n5902), .ZN(n5907) );
  INV_X1 U7501 ( .A(n5901), .ZN(n5904) );
  INV_X1 U7502 ( .A(n5902), .ZN(n5903) );
  NAND2_X1 U7503 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  NAND2_X1 U7504 ( .A1(n5907), .A2(n5905), .ZN(n7078) );
  NAND2_X1 U7505 ( .A1(n6540), .A2(n5891), .ZN(n5914) );
  NAND2_X1 U7506 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  NAND2_X1 U7507 ( .A1(n5924), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5912) );
  XNOR2_X1 U7508 ( .A(n5912), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7509 ( .A1(n4487), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6070), .B2(
        n6721), .ZN(n5913) );
  NAND2_X1 U7510 ( .A1(n6024), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7511 ( .A1(n7845), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5920) );
  INV_X1 U7512 ( .A(n5915), .ZN(n5916) );
  AOI21_X1 U7513 ( .B1(n5916), .B2(P2_REG3_REG_6__SCAN_IN), .A(
        P2_REG3_REG_7__SCAN_IN), .ZN(n5917) );
  OR2_X1 U7514 ( .A1(n5917), .A2(n5929), .ZN(n7252) );
  INV_X1 U7515 ( .A(n7252), .ZN(n7114) );
  NAND2_X1 U7516 ( .A1(n6261), .A2(n7114), .ZN(n5919) );
  NAND2_X1 U7517 ( .A1(n7844), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5918) );
  NOR2_X1 U7518 ( .A1(n7358), .A2(n7306), .ZN(n5922) );
  XNOR2_X1 U7519 ( .A(n5923), .B(n5922), .ZN(n7250) );
  NAND2_X1 U7520 ( .A1(n6543), .A2(n5891), .ZN(n5927) );
  NOR2_X1 U7521 ( .A1(n5924), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5941) );
  OR2_X1 U7522 ( .A1(n5941), .A2(n5771), .ZN(n5925) );
  XNOR2_X1 U7523 ( .A(n5925), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6718) );
  AOI22_X1 U7524 ( .A1(n4487), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6070), .B2(
        n6718), .ZN(n5926) );
  NAND2_X1 U7525 ( .A1(n5927), .A2(n5926), .ZN(n7353) );
  XNOR2_X1 U7526 ( .A(n7353), .B(n6211), .ZN(n5935) );
  INV_X2 U7527 ( .A(n5928), .ZN(n5975) );
  NAND2_X1 U7528 ( .A1(n5975), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7529 ( .A1(n7844), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5933) );
  OR2_X1 U7530 ( .A1(n5929), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5930) );
  AND2_X1 U7531 ( .A1(n5945), .A2(n5930), .ZN(n7352) );
  NAND2_X1 U7532 ( .A1(n6261), .A2(n7352), .ZN(n5932) );
  NAND2_X1 U7533 ( .A1(n7845), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5931) );
  NOR2_X1 U7534 ( .A1(n7268), .A2(n7306), .ZN(n5936) );
  XNOR2_X1 U7535 ( .A(n5935), .B(n5936), .ZN(n7056) );
  NAND2_X1 U7536 ( .A1(n7057), .A2(n7056), .ZN(n5939) );
  INV_X1 U7537 ( .A(n5935), .ZN(n5937) );
  NAND2_X1 U7538 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  NAND2_X1 U7539 ( .A1(n5939), .A2(n5938), .ZN(n7187) );
  NAND2_X1 U7540 ( .A1(n6558), .A2(n5891), .ZN(n5943) );
  INV_X1 U7541 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7542 ( .A1(n5941), .A2(n5940), .ZN(n5989) );
  NAND2_X1 U7543 ( .A1(n5989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5957) );
  XNOR2_X1 U7544 ( .A(n5957), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6952) );
  AOI22_X1 U7545 ( .A1(n4487), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6070), .B2(
        n6952), .ZN(n5942) );
  NAND2_X1 U7546 ( .A1(n5943), .A2(n5942), .ZN(n7377) );
  XNOR2_X1 U7547 ( .A(n7377), .B(n6211), .ZN(n5951) );
  NAND2_X1 U7548 ( .A1(n5975), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7549 ( .A1(n7844), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7550 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  AND2_X1 U7551 ( .A1(n5962), .A2(n5946), .ZN(n7285) );
  NAND2_X1 U7552 ( .A1(n6261), .A2(n7285), .ZN(n5948) );
  NAND2_X1 U7553 ( .A1(n7845), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7554 ( .A1(n7381), .A2(n7306), .ZN(n5952) );
  NAND2_X1 U7555 ( .A1(n5951), .A2(n5952), .ZN(n5956) );
  INV_X1 U7556 ( .A(n5951), .ZN(n5954) );
  INV_X1 U7557 ( .A(n5952), .ZN(n5953) );
  NAND2_X1 U7558 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7559 ( .A1(n5956), .A2(n5955), .ZN(n7186) );
  NAND2_X1 U7560 ( .A1(n5957), .A2(n5986), .ZN(n5958) );
  NAND2_X1 U7561 ( .A1(n5958), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7562 ( .A1(n5959), .A2(n5987), .ZN(n5971) );
  OR2_X1 U7563 ( .A1(n5959), .A2(n5987), .ZN(n5960) );
  AOI22_X1 U7564 ( .A1(n4487), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6070), .B2(
        n7092), .ZN(n5961) );
  XNOR2_X1 U7565 ( .A(n10004), .B(n6157), .ZN(n5969) );
  NAND2_X1 U7566 ( .A1(n5975), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7567 ( .A1(n7844), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5966) );
  AND2_X1 U7568 ( .A1(n5962), .A2(n10462), .ZN(n5963) );
  NOR2_X1 U7569 ( .A1(n5976), .A2(n5963), .ZN(n7388) );
  NAND2_X1 U7570 ( .A1(n6261), .A2(n7388), .ZN(n5965) );
  NAND2_X1 U7571 ( .A1(n7845), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5964) );
  NOR2_X1 U7572 ( .A1(n7794), .A2(n7306), .ZN(n5968) );
  XNOR2_X1 U7573 ( .A(n5969), .B(n5968), .ZN(n7159) );
  NAND2_X1 U7574 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  NAND2_X1 U7575 ( .A1(n6570), .A2(n5891), .ZN(n5974) );
  NAND2_X1 U7576 ( .A1(n5971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U7577 ( .A(n5972), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7174) );
  AOI22_X1 U7578 ( .A1(n4487), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6070), .B2(
        n7174), .ZN(n5973) );
  XNOR2_X1 U7579 ( .A(n7483), .B(n6211), .ZN(n5984) );
  NAND2_X1 U7580 ( .A1(n5975), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7581 ( .A1(n7844), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5980) );
  NOR2_X1 U7582 ( .A1(n5976), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5977) );
  OR2_X1 U7583 ( .A1(n5993), .A2(n5977), .ZN(n7792) );
  INV_X1 U7584 ( .A(n7792), .ZN(n7481) );
  NAND2_X1 U7585 ( .A1(n6261), .A2(n7481), .ZN(n5979) );
  NAND2_X1 U7586 ( .A1(n7845), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5978) );
  NAND4_X1 U7587 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n8542)
         );
  NAND2_X1 U7588 ( .A1(n8542), .A2(n7864), .ZN(n5982) );
  XNOR2_X1 U7589 ( .A(n5984), .B(n5982), .ZN(n7790) );
  INV_X1 U7590 ( .A(n5982), .ZN(n5983) );
  AND2_X1 U7591 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  AOI21_X2 U7592 ( .B1(n7791), .B2(n7790), .A(n5985), .ZN(n7468) );
  NAND2_X1 U7593 ( .A1(n6595), .A2(n5891), .ZN(n5992) );
  NAND2_X1 U7594 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7595 ( .A1(n6005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5990) );
  XNOR2_X1 U7596 ( .A(n5990), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7323) );
  AOI22_X1 U7597 ( .A1(n4487), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6070), .B2(
        n7323), .ZN(n5991) );
  NAND2_X1 U7598 ( .A1(n5992), .A2(n5991), .ZN(n7558) );
  XNOR2_X1 U7599 ( .A(n7558), .B(n6211), .ZN(n5999) );
  NAND2_X1 U7600 ( .A1(n6024), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7601 ( .A1(n7844), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5997) );
  OR2_X1 U7602 ( .A1(n5993), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5994) );
  AND2_X1 U7603 ( .A1(n6008), .A2(n5994), .ZN(n7524) );
  NAND2_X1 U7604 ( .A1(n6261), .A2(n7524), .ZN(n5996) );
  NAND2_X1 U7605 ( .A1(n7845), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5995) );
  OR2_X1 U7606 ( .A1(n7793), .A2(n7306), .ZN(n6000) );
  NAND2_X1 U7607 ( .A1(n5999), .A2(n6000), .ZN(n6004) );
  INV_X1 U7608 ( .A(n5999), .ZN(n6002) );
  INV_X1 U7609 ( .A(n6000), .ZN(n6001) );
  NAND2_X1 U7610 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  AND2_X1 U7611 ( .A1(n6004), .A2(n6003), .ZN(n7469) );
  NAND2_X1 U7612 ( .A1(n6800), .A2(n5891), .ZN(n6007) );
  OAI21_X1 U7613 ( .B1(n6005), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U7614 ( .A(n6018), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7426) );
  AOI22_X1 U7615 ( .A1(n4487), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6070), .B2(
        n7426), .ZN(n6006) );
  XNOR2_X1 U7616 ( .A(n7586), .B(n6157), .ZN(n6015) );
  NAND2_X1 U7617 ( .A1(n6024), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7618 ( .A1(n7844), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7619 ( .A1(n6008), .A2(n7327), .ZN(n6009) );
  AND2_X1 U7620 ( .A1(n6022), .A2(n6009), .ZN(n7509) );
  NAND2_X1 U7621 ( .A1(n6261), .A2(n7509), .ZN(n6011) );
  NAND2_X1 U7622 ( .A1(n6200), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6010) );
  NOR2_X1 U7623 ( .A1(n7581), .A2(n7306), .ZN(n6014) );
  XNOR2_X1 U7624 ( .A(n6015), .B(n6014), .ZN(n7507) );
  NAND2_X1 U7625 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  NAND2_X1 U7626 ( .A1(n6798), .A2(n5891), .ZN(n6021) );
  INV_X1 U7627 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7628 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  NAND2_X1 U7629 ( .A1(n6019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6036) );
  XNOR2_X1 U7630 ( .A(n6036), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7649) );
  AOI22_X1 U7631 ( .A1(n4487), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7649), .B2(
        n6070), .ZN(n6020) );
  XNOR2_X1 U7632 ( .A(n7628), .B(n6211), .ZN(n6029) );
  NAND2_X1 U7633 ( .A1(n6022), .A2(n10277), .ZN(n6023) );
  AND2_X1 U7634 ( .A1(n6053), .A2(n6023), .ZN(n7606) );
  NAND2_X1 U7635 ( .A1(n6261), .A2(n7606), .ZN(n6028) );
  NAND2_X1 U7636 ( .A1(n6024), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7637 ( .A1(n7844), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7638 ( .A1(n6200), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6025) );
  OR2_X1 U7639 ( .A1(n7709), .A2(n7306), .ZN(n6030) );
  NAND2_X1 U7640 ( .A1(n6029), .A2(n6030), .ZN(n6034) );
  INV_X1 U7641 ( .A(n6029), .ZN(n6032) );
  INV_X1 U7642 ( .A(n6030), .ZN(n6031) );
  NAND2_X1 U7643 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  NAND2_X1 U7644 ( .A1(n6034), .A2(n6033), .ZN(n7605) );
  NAND2_X1 U7645 ( .A1(n6986), .A2(n5891), .ZN(n6040) );
  INV_X1 U7646 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7647 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U7648 ( .A1(n6037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7649 ( .A(n6038), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8561) );
  AOI22_X1 U7650 ( .A1(n8561), .A2(n6070), .B1(n4487), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6039) );
  XNOR2_X1 U7651 ( .A(n7721), .B(n6157), .ZN(n6045) );
  NAND2_X1 U7652 ( .A1(n6024), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7653 ( .A1(n7844), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6043) );
  XNOR2_X1 U7654 ( .A(n6053), .B(P2_REG3_REG_15__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U7655 ( .A1(n6261), .A2(n7712), .ZN(n6042) );
  NAND2_X1 U7656 ( .A1(n6200), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6041) );
  NOR2_X1 U7657 ( .A1(n7743), .A2(n7306), .ZN(n7707) );
  INV_X1 U7658 ( .A(n6045), .ZN(n6046) );
  NOR2_X1 U7659 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  NAND2_X1 U7660 ( .A1(n7043), .A2(n5891), .ZN(n6052) );
  NAND2_X1 U7661 ( .A1(n6049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6050) );
  XNOR2_X1 U7662 ( .A(n6050), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8578) );
  AOI22_X1 U7663 ( .A1(n4487), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6070), .B2(
        n8578), .ZN(n6051) );
  XNOR2_X1 U7664 ( .A(n7748), .B(n6157), .ZN(n6060) );
  NAND2_X1 U7665 ( .A1(n6024), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6059) );
  INV_X1 U7666 ( .A(n6053), .ZN(n6054) );
  AOI21_X1 U7667 ( .B1(n6054), .B2(P2_REG3_REG_15__SCAN_IN), .A(
        P2_REG3_REG_16__SCAN_IN), .ZN(n6055) );
  OR2_X1 U7668 ( .A1(n6055), .A2(n6075), .ZN(n7732) );
  INV_X1 U7669 ( .A(n7732), .ZN(n7745) );
  NAND2_X1 U7670 ( .A1(n7745), .A2(n6261), .ZN(n6058) );
  NAND2_X1 U7671 ( .A1(n7844), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7672 ( .A1(n7845), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6056) );
  NAND4_X1 U7673 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n8537)
         );
  NAND2_X1 U7674 ( .A1(n8537), .A2(n7864), .ZN(n6061) );
  NAND2_X1 U7675 ( .A1(n6060), .A2(n6061), .ZN(n6065) );
  INV_X1 U7676 ( .A(n6060), .ZN(n6063) );
  INV_X1 U7677 ( .A(n6061), .ZN(n6062) );
  NAND2_X1 U7678 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  AND2_X1 U7679 ( .A1(n6065), .A2(n6064), .ZN(n7741) );
  NAND2_X1 U7680 ( .A1(n7046), .A2(n5891), .ZN(n6072) );
  NAND2_X1 U7681 ( .A1(n4488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6066) );
  MUX2_X1 U7682 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6066), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n6067) );
  INV_X1 U7683 ( .A(n6067), .ZN(n6069) );
  NOR2_X1 U7684 ( .A1(n6069), .A2(n6068), .ZN(n8592) );
  AOI22_X1 U7685 ( .A1(n4487), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6070), .B2(
        n8592), .ZN(n6071) );
  XNOR2_X1 U7686 ( .A(n8907), .B(n6211), .ZN(n6081) );
  NAND2_X1 U7687 ( .A1(n5975), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7688 ( .A1(n6200), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6073) );
  AND2_X1 U7689 ( .A1(n6074), .A2(n6073), .ZN(n6080) );
  NOR2_X1 U7690 ( .A1(n6075), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6076) );
  OR2_X1 U7691 ( .A1(n6091), .A2(n6076), .ZN(n7768) );
  INV_X1 U7692 ( .A(n7768), .ZN(n6077) );
  NAND2_X1 U7693 ( .A1(n6077), .A2(n6261), .ZN(n6079) );
  NAND2_X1 U7694 ( .A1(n7844), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6078) );
  INV_X1 U7695 ( .A(n7781), .ZN(n8808) );
  NAND2_X1 U7696 ( .A1(n8808), .A2(n7864), .ZN(n6082) );
  XNOR2_X1 U7697 ( .A(n6081), .B(n6082), .ZN(n7752) );
  INV_X1 U7698 ( .A(n6081), .ZN(n6084) );
  INV_X1 U7699 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7700 ( .A1(n7226), .A2(n5891), .ZN(n6090) );
  INV_X1 U7701 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7227) );
  INV_X1 U7702 ( .A(n6068), .ZN(n6085) );
  NAND2_X1 U7703 ( .A1(n6085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6087) );
  XNOR2_X1 U7704 ( .A(n6087), .B(n6086), .ZN(n8590) );
  OAI22_X1 U7705 ( .A1(n6100), .A2(n7227), .B1(n5860), .B2(n8590), .ZN(n6088)
         );
  INV_X1 U7706 ( .A(n6088), .ZN(n6089) );
  XNOR2_X1 U7707 ( .A(n8901), .B(n6157), .ZN(n6098) );
  NOR2_X1 U7708 ( .A1(n6091), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7709 ( .A1(n6104), .A2(n6092), .ZN(n8799) );
  AOI22_X1 U7710 ( .A1(n6200), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n6024), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7711 ( .A1(n7844), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6093) );
  OAI211_X1 U7712 ( .C1(n8799), .C2(n6095), .A(n6094), .B(n6093), .ZN(n8536)
         );
  NAND2_X1 U7713 ( .A1(n8536), .A2(n7864), .ZN(n6096) );
  XNOR2_X1 U7714 ( .A(n6098), .B(n6096), .ZN(n7780) );
  INV_X1 U7715 ( .A(n6096), .ZN(n6097) );
  NAND2_X1 U7716 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  NAND2_X1 U7717 ( .A1(n7314), .A2(n5891), .ZN(n6103) );
  OAI22_X1 U7718 ( .A1(n6100), .A2(n7316), .B1(n7892), .B2(n5860), .ZN(n6101)
         );
  INV_X1 U7719 ( .A(n6101), .ZN(n6102) );
  XNOR2_X1 U7720 ( .A(n8897), .B(n6211), .ZN(n6109) );
  OR2_X1 U7721 ( .A1(n6104), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6105) );
  AND2_X1 U7722 ( .A1(n6105), .A2(n6118), .ZN(n8787) );
  NAND2_X1 U7723 ( .A1(n8787), .A2(n6261), .ZN(n6108) );
  AOI22_X1 U7724 ( .A1(n6200), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n6024), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7725 ( .A1(n7844), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7726 ( .A1(n8811), .A2(n7864), .ZN(n6110) );
  NAND2_X1 U7727 ( .A1(n6109), .A2(n6110), .ZN(n6115) );
  INV_X1 U7728 ( .A(n6109), .ZN(n6112) );
  INV_X1 U7729 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7730 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  NAND2_X1 U7731 ( .A1(n6115), .A2(n6113), .ZN(n8452) );
  NAND2_X1 U7732 ( .A1(n8450), .A2(n6115), .ZN(n8496) );
  NAND2_X1 U7733 ( .A1(n7444), .A2(n5891), .ZN(n6117) );
  NAND2_X1 U7734 ( .A1(n4487), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6116) );
  XNOR2_X1 U7735 ( .A(n8888), .B(n6157), .ZN(n6124) );
  NAND2_X1 U7736 ( .A1(n6024), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7737 ( .A1(n7845), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6122) );
  INV_X1 U7738 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10429) );
  NAND2_X1 U7739 ( .A1(n10429), .A2(n6118), .ZN(n6119) );
  AND2_X1 U7740 ( .A1(n6119), .A2(n6130), .ZN(n8769) );
  NAND2_X1 U7741 ( .A1(n6261), .A2(n8769), .ZN(n6121) );
  NAND2_X1 U7742 ( .A1(n7844), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6120) );
  NOR2_X1 U7743 ( .A1(n8464), .A2(n7306), .ZN(n6125) );
  XNOR2_X1 U7744 ( .A(n6124), .B(n6125), .ZN(n8495) );
  INV_X1 U7745 ( .A(n6124), .ZN(n6127) );
  INV_X1 U7746 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7747 ( .A1(n7475), .A2(n5891), .ZN(n6129) );
  NAND2_X1 U7748 ( .A1(n4487), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7749 ( .A(n8882), .B(n6157), .ZN(n6138) );
  NAND2_X1 U7750 ( .A1(n6024), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7751 ( .A1(n6200), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6134) );
  INV_X1 U7752 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U7753 ( .A1(n10483), .A2(n6130), .ZN(n6131) );
  AND2_X1 U7754 ( .A1(n6144), .A2(n6131), .ZN(n8745) );
  NAND2_X1 U7755 ( .A1(n6261), .A2(n8745), .ZN(n6133) );
  NAND2_X1 U7756 ( .A1(n7844), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6132) );
  NAND4_X1 U7757 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n8535)
         );
  NAND2_X1 U7758 ( .A1(n8535), .A2(n7864), .ZN(n6136) );
  XNOR2_X1 U7759 ( .A(n6138), .B(n6136), .ZN(n8462) );
  NAND2_X1 U7760 ( .A1(n8461), .A2(n8462), .ZN(n6140) );
  INV_X1 U7761 ( .A(n6136), .ZN(n6137) );
  NAND2_X1 U7762 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  NAND2_X1 U7763 ( .A1(n6140), .A2(n6139), .ZN(n6153) );
  NAND2_X1 U7764 ( .A1(n7551), .A2(n5891), .ZN(n6142) );
  NAND2_X1 U7765 ( .A1(n4487), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7766 ( .A(n8877), .B(n6211), .ZN(n6151) );
  XNOR2_X1 U7767 ( .A(n6153), .B(n6151), .ZN(n8509) );
  NAND2_X1 U7768 ( .A1(n6200), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7769 ( .A1(n5975), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6149) );
  INV_X1 U7770 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7771 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  AND2_X1 U7772 ( .A1(n6146), .A2(n6145), .ZN(n8730) );
  NAND2_X1 U7773 ( .A1(n6261), .A2(n8730), .ZN(n6148) );
  NAND2_X1 U7774 ( .A1(n7844), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6147) );
  OR2_X1 U7775 ( .A1(n8534), .A2(n7306), .ZN(n8508) );
  NAND2_X1 U7776 ( .A1(n8509), .A2(n8508), .ZN(n8507) );
  INV_X1 U7777 ( .A(n6151), .ZN(n6152) );
  OR2_X1 U7778 ( .A1(n6153), .A2(n6152), .ZN(n6154) );
  NAND2_X1 U7779 ( .A1(n7552), .A2(n5891), .ZN(n6156) );
  NAND2_X1 U7780 ( .A1(n4487), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6155) );
  XNOR2_X1 U7781 ( .A(n8872), .B(n6157), .ZN(n6160) );
  INV_X1 U7782 ( .A(n6160), .ZN(n6158) );
  INV_X1 U7783 ( .A(n8472), .ZN(n8723) );
  NAND2_X1 U7784 ( .A1(n8723), .A2(n7864), .ZN(n6161) );
  INV_X1 U7785 ( .A(n8485), .ZN(n6162) );
  INV_X1 U7786 ( .A(n6161), .ZN(n8484) );
  NAND2_X1 U7787 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7788 ( .A1(n7716), .A2(n5891), .ZN(n6168) );
  NAND2_X1 U7789 ( .A1(n4487), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6167) );
  XNOR2_X1 U7790 ( .A(n8864), .B(n6157), .ZN(n6169) );
  INV_X1 U7791 ( .A(n6169), .ZN(n8470) );
  NAND2_X1 U7792 ( .A1(n7845), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7793 ( .A1(n6024), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6175) );
  INV_X1 U7794 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7795 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  AND2_X1 U7796 ( .A1(n6179), .A2(n6172), .ZN(n8692) );
  NAND2_X1 U7797 ( .A1(n6261), .A2(n8692), .ZN(n6174) );
  NAND2_X1 U7798 ( .A1(n7844), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6173) );
  NAND4_X1 U7799 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n8707)
         );
  NAND2_X1 U7800 ( .A1(n8707), .A2(n7864), .ZN(n8469) );
  NAND2_X1 U7801 ( .A1(n7749), .A2(n5891), .ZN(n6178) );
  NAND2_X1 U7802 ( .A1(n4487), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6177) );
  XNOR2_X1 U7803 ( .A(n8858), .B(n6211), .ZN(n6186) );
  NAND2_X1 U7804 ( .A1(n7845), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7805 ( .A1(n5975), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6183) );
  INV_X1 U7806 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U7807 ( .A1(n6179), .A2(n10182), .ZN(n6180) );
  NAND2_X1 U7808 ( .A1(n6261), .A2(n8670), .ZN(n6182) );
  NAND2_X1 U7809 ( .A1(n7844), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6181) );
  OR2_X1 U7810 ( .A1(n8657), .A2(n7306), .ZN(n6185) );
  NOR2_X1 U7811 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  AOI21_X1 U7812 ( .B1(n6186), .B2(n6185), .A(n6187), .ZN(n8519) );
  NAND2_X1 U7813 ( .A1(n8520), .A2(n8519), .ZN(n8518) );
  INV_X1 U7814 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7815 ( .A1(n8518), .A2(n6188), .ZN(n8432) );
  NAND2_X1 U7816 ( .A1(n8945), .A2(n5891), .ZN(n6190) );
  NAND2_X1 U7817 ( .A1(n4487), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6189) );
  XNOR2_X1 U7818 ( .A(n8852), .B(n6211), .ZN(n6196) );
  NAND2_X1 U7819 ( .A1(n6200), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7820 ( .A1(n5975), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7821 ( .A(n6205), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7822 ( .A1(n6261), .A2(n8651), .ZN(n6192) );
  NAND2_X1 U7823 ( .A1(n7844), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6191) );
  OR2_X1 U7824 ( .A1(n8630), .A2(n7306), .ZN(n6195) );
  NOR2_X1 U7825 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  AOI21_X1 U7826 ( .B1(n6196), .B2(n6195), .A(n6197), .ZN(n8431) );
  NAND2_X1 U7827 ( .A1(n8432), .A2(n8431), .ZN(n8430) );
  NAND2_X1 U7828 ( .A1(n8941), .A2(n5891), .ZN(n6199) );
  NAND2_X1 U7829 ( .A1(n4487), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7830 ( .A1(n6200), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7831 ( .A1(n5975), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6209) );
  INV_X1 U7832 ( .A(n6205), .ZN(n6202) );
  AND2_X1 U7833 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6201) );
  NAND2_X1 U7834 ( .A1(n6202), .A2(n6201), .ZN(n6260) );
  INV_X1 U7835 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6204) );
  INV_X1 U7836 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6203) );
  OAI21_X1 U7837 ( .B1(n6205), .B2(n6204), .A(n6203), .ZN(n6206) );
  NAND2_X1 U7838 ( .A1(n6261), .A2(n8638), .ZN(n6208) );
  NAND2_X1 U7839 ( .A1(n7844), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6207) );
  OR2_X1 U7840 ( .A1(n8658), .A2(n7306), .ZN(n6212) );
  XNOR2_X1 U7841 ( .A(n6212), .B(n6211), .ZN(n6247) );
  INV_X1 U7842 ( .A(n6247), .ZN(n6248) );
  INV_X1 U7843 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9947) );
  NAND3_X1 U7844 ( .A1(n6216), .A2(n6219), .A3(n6221), .ZN(n6213) );
  OAI21_X1 U7845 ( .B1(n4490), .B2(n6213), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6214) );
  MUX2_X1 U7846 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6214), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6215) );
  NAND2_X1 U7847 ( .A1(n6215), .A2(n4575), .ZN(n7717) );
  NAND2_X1 U7848 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  NAND2_X1 U7849 ( .A1(n6241), .A2(n6219), .ZN(n6220) );
  INV_X1 U7850 ( .A(P2_B_REG_SCAN_IN), .ZN(n10172) );
  XOR2_X1 U7851 ( .A(n7615), .B(n10172), .Z(n6223) );
  NAND2_X1 U7852 ( .A1(n7717), .A2(n6223), .ZN(n6227) );
  NAND2_X1 U7853 ( .A1(n4575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6224) );
  MUX2_X1 U7854 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6224), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6226) );
  NAND2_X1 U7855 ( .A1(n6226), .A2(n6225), .ZN(n6240) );
  INV_X1 U7856 ( .A(n6240), .ZN(n7750) );
  AND2_X1 U7857 ( .A1(n7717), .A2(n6240), .ZN(n9949) );
  NOR4_X1 U7858 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6236) );
  OR4_X1 U7859 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6233) );
  NOR4_X1 U7860 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6231) );
  NOR4_X1 U7861 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6230) );
  NOR4_X1 U7862 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6229) );
  NOR4_X1 U7863 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6228) );
  NAND4_X1 U7864 ( .A1(n6231), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(n6232)
         );
  NOR4_X1 U7865 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6233), .A4(n6232), .ZN(n6235) );
  NOR4_X1 U7866 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6234) );
  NAND3_X1 U7867 ( .A1(n6236), .A2(n6235), .A3(n6234), .ZN(n6237) );
  AND2_X1 U7868 ( .A1(n7615), .A2(n6240), .ZN(n9945) );
  INV_X1 U7869 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9944) );
  AND2_X1 U7870 ( .A1(n9941), .A2(n9944), .ZN(n6238) );
  NOR2_X1 U7871 ( .A1(n6972), .A2(n6981), .ZN(n6239) );
  NAND2_X1 U7872 ( .A1(n6976), .A2(n6239), .ZN(n6266) );
  INV_X2 U7873 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U7874 ( .A(n9943), .ZN(n6242) );
  NOR2_X1 U7875 ( .A1(n6252), .A2(n8061), .ZN(n6816) );
  INV_X1 U7876 ( .A(n6816), .ZN(n6244) );
  INV_X1 U7877 ( .A(n6973), .ZN(n6243) );
  NOR3_X1 U7878 ( .A1(n8640), .A2(n6248), .A3(n8492), .ZN(n6245) );
  AOI21_X1 U7879 ( .B1(n8640), .B2(n6248), .A(n6245), .ZN(n6246) );
  NOR3_X1 U7880 ( .A1(n8640), .A2(n6247), .A3(n8492), .ZN(n6250) );
  NOR2_X1 U7881 ( .A1(n8847), .A2(n6248), .ZN(n6249) );
  NAND2_X1 U7882 ( .A1(n6254), .A2(n6255), .ZN(n6830) );
  NOR2_X1 U7883 ( .A1(n10013), .A2(n6555), .ZN(n6256) );
  OAI21_X1 U7884 ( .B1(n8640), .B2(n8529), .A(n8505), .ZN(n6257) );
  NAND2_X1 U7885 ( .A1(n6259), .A2(n6267), .ZN(n8524) );
  NAND2_X1 U7886 ( .A1(n5975), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7887 ( .A1(n7845), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6264) );
  INV_X1 U7888 ( .A(n6260), .ZN(n8414) );
  NAND2_X1 U7889 ( .A1(n6261), .A2(n8414), .ZN(n6263) );
  NAND2_X1 U7890 ( .A1(n7844), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6262) );
  NAND4_X1 U7891 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n8634)
         );
  INV_X1 U7892 ( .A(n6668), .ZN(n8942) );
  INV_X1 U7893 ( .A(n8630), .ZN(n8402) );
  AOI22_X1 U7894 ( .A1(n8511), .A2(n8634), .B1(n8510), .B2(n8402), .ZN(n6272)
         );
  NAND2_X1 U7895 ( .A1(n6266), .A2(n6973), .ZN(n6916) );
  NOR2_X1 U7896 ( .A1(n6830), .A2(n6267), .ZN(n6268) );
  NOR2_X1 U7897 ( .A1(n6268), .A2(n6554), .ZN(n6269) );
  NAND2_X1 U7898 ( .A1(n6519), .A2(n6269), .ZN(n6813) );
  INV_X1 U7899 ( .A(n6813), .ZN(n8067) );
  NAND2_X1 U7900 ( .A1(n6916), .A2(n8067), .ZN(n6270) );
  AOI22_X1 U7901 ( .A1(n8526), .A2(n8638), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6271) );
  INV_X1 U7902 ( .A(n6497), .ZN(n6274) );
  NAND2_X2 U7903 ( .A1(n6275), .A2(n6274), .ZN(n6308) );
  INV_X2 U7904 ( .A(n6308), .ZN(n6394) );
  AND2_X4 U7905 ( .A1(n6275), .A2(n6497), .ZN(n7801) );
  OR2_X1 U7906 ( .A1(n6276), .A2(n4481), .ZN(n6277) );
  AOI22_X1 U7907 ( .A1(n9228), .A2(n6489), .B1(n6482), .B2(n9242), .ZN(n6469)
         );
  INV_X1 U7908 ( .A(n6469), .ZN(n6471) );
  NAND2_X1 U7909 ( .A1(n9228), .A2(n7801), .ZN(n6279) );
  NAND2_X1 U7910 ( .A1(n9242), .A2(n7806), .ZN(n6278) );
  NAND2_X1 U7911 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  XNOR2_X1 U7912 ( .A(n6280), .B(n7030), .ZN(n6470) );
  INV_X1 U7913 ( .A(n6275), .ZN(n6281) );
  AOI22_X1 U7914 ( .A1(n6394), .A2(n7012), .B1(n6281), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7915 ( .A1(n6394), .A2(n9804), .ZN(n6285) );
  INV_X1 U7916 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6283) );
  OR2_X1 U7917 ( .A1(n6275), .A2(n6283), .ZN(n6284) );
  INV_X1 U7918 ( .A(n6589), .ZN(n6286) );
  NAND2_X1 U7919 ( .A1(n6286), .A2(n7030), .ZN(n6287) );
  NAND2_X1 U7920 ( .A1(n7801), .A2(n8333), .ZN(n6289) );
  NAND2_X1 U7921 ( .A1(n6394), .A2(n5292), .ZN(n6288) );
  NAND2_X1 U7922 ( .A1(n6289), .A2(n6288), .ZN(n6290) );
  NAND2_X1 U7923 ( .A1(n6599), .A2(n6601), .ZN(n6291) );
  OAI22_X1 U7924 ( .A1(n8334), .A2(n7808), .B1(n9798), .B2(n6308), .ZN(n6598)
         );
  NAND2_X1 U7925 ( .A1(n6291), .A2(n6598), .ZN(n6295) );
  INV_X1 U7926 ( .A(n6686), .ZN(n6301) );
  OAI22_X1 U7927 ( .A1(n5294), .A2(n6308), .B1(n9832), .B2(n6318), .ZN(n6296)
         );
  XNOR2_X1 U7928 ( .A(n6296), .B(n7030), .ZN(n6298) );
  OAI22_X1 U7929 ( .A1(n7808), .A2(n5294), .B1(n9832), .B2(n6308), .ZN(n6297)
         );
  NAND2_X1 U7930 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  NAND2_X1 U7931 ( .A1(n6302), .A2(n6299), .ZN(n6687) );
  INV_X1 U7932 ( .A(n6687), .ZN(n6300) );
  NAND2_X1 U7933 ( .A1(n6301), .A2(n6300), .ZN(n6684) );
  NAND2_X1 U7934 ( .A1(n6684), .A2(n6302), .ZN(n6804) );
  OAI22_X1 U7935 ( .A1(n9849), .A2(n6308), .B1(n9840), .B2(n6318), .ZN(n6303)
         );
  XNOR2_X1 U7936 ( .A(n6303), .B(n7804), .ZN(n6304) );
  OAI22_X1 U7937 ( .A1(n7808), .A2(n9849), .B1(n9840), .B2(n6308), .ZN(n6305)
         );
  XNOR2_X1 U7938 ( .A(n6304), .B(n6305), .ZN(n6805) );
  NAND2_X1 U7939 ( .A1(n6804), .A2(n6805), .ZN(n6803) );
  INV_X1 U7940 ( .A(n6304), .ZN(n6306) );
  OR2_X1 U7941 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  OAI22_X1 U7942 ( .A1(n9836), .A2(n6308), .B1(n7300), .B2(n6318), .ZN(n6309)
         );
  XNOR2_X1 U7943 ( .A(n6309), .B(n7030), .ZN(n6311) );
  OAI22_X1 U7944 ( .A1(n7808), .A2(n9836), .B1(n7300), .B2(n6308), .ZN(n6310)
         );
  XNOR2_X1 U7945 ( .A(n6311), .B(n6310), .ZN(n7023) );
  NAND2_X1 U7946 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  NAND2_X1 U7947 ( .A1(n7801), .A2(n9784), .ZN(n6313) );
  OAI21_X1 U7948 ( .B1(n9848), .B2(n6308), .A(n6313), .ZN(n6314) );
  XNOR2_X1 U7949 ( .A(n6314), .B(n7030), .ZN(n7230) );
  OR2_X1 U7950 ( .A1(n9848), .A2(n7808), .ZN(n6316) );
  NAND2_X1 U7951 ( .A1(n6394), .A2(n9784), .ZN(n6315) );
  NAND2_X1 U7952 ( .A1(n6316), .A2(n6315), .ZN(n6322) );
  NAND2_X1 U7953 ( .A1(n7230), .A2(n6322), .ZN(n6317) );
  OAI22_X1 U7954 ( .A1(n7209), .A2(n6318), .B1(n9876), .B2(n6308), .ZN(n6319)
         );
  XNOR2_X1 U7955 ( .A(n6319), .B(n7804), .ZN(n6327) );
  NAND2_X1 U7956 ( .A1(n6482), .A2(n9782), .ZN(n6321) );
  OR2_X1 U7957 ( .A1(n7209), .A2(n6308), .ZN(n6320) );
  AND2_X1 U7958 ( .A1(n6321), .A2(n6320), .ZN(n6328) );
  NAND2_X1 U7959 ( .A1(n6327), .A2(n6328), .ZN(n7232) );
  INV_X1 U7960 ( .A(n7230), .ZN(n6323) );
  INV_X1 U7961 ( .A(n6322), .ZN(n7259) );
  NAND2_X1 U7962 ( .A1(n6323), .A2(n7259), .ZN(n6324) );
  AND2_X1 U7963 ( .A1(n7232), .A2(n6324), .ZN(n6325) );
  INV_X1 U7964 ( .A(n6327), .ZN(n6330) );
  INV_X1 U7965 ( .A(n6328), .ZN(n6329) );
  NAND2_X1 U7966 ( .A1(n6330), .A2(n6329), .ZN(n7234) );
  NAND2_X1 U7967 ( .A1(n9879), .A2(n7806), .ZN(n6332) );
  NAND2_X1 U7968 ( .A1(n6482), .A2(n9864), .ZN(n6331) );
  NAND2_X1 U7969 ( .A1(n6332), .A2(n6331), .ZN(n7048) );
  INV_X1 U7970 ( .A(n7048), .ZN(n6333) );
  NAND2_X1 U7971 ( .A1(n9879), .A2(n7801), .ZN(n6335) );
  NAND2_X1 U7972 ( .A1(n9864), .A2(n7806), .ZN(n6334) );
  NAND2_X1 U7973 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  XNOR2_X1 U7974 ( .A(n6336), .B(n7030), .ZN(n6343) );
  NOR2_X1 U7975 ( .A1(n7808), .A2(n9875), .ZN(n6337) );
  AOI21_X1 U7976 ( .B1(n9893), .B2(n6489), .A(n6337), .ZN(n6345) );
  NAND2_X1 U7977 ( .A1(n6338), .A2(n7048), .ZN(n6344) );
  NAND2_X1 U7978 ( .A1(n9893), .A2(n7801), .ZN(n6341) );
  NAND2_X1 U7979 ( .A1(n9093), .A2(n6489), .ZN(n6340) );
  NAND2_X1 U7980 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  XNOR2_X1 U7981 ( .A(n6342), .B(n7030), .ZN(n7412) );
  INV_X1 U7982 ( .A(n6343), .ZN(n7049) );
  NAND2_X1 U7983 ( .A1(n6344), .A2(n7049), .ZN(n6348) );
  INV_X1 U7984 ( .A(n6345), .ZN(n6346) );
  NAND3_X1 U7985 ( .A1(n6348), .A2(n6347), .A3(n6346), .ZN(n7409) );
  NAND2_X1 U7986 ( .A1(n9769), .A2(n7801), .ZN(n6351) );
  NAND2_X1 U7987 ( .A1(n6394), .A2(n9092), .ZN(n6350) );
  NAND2_X1 U7988 ( .A1(n6351), .A2(n6350), .ZN(n6352) );
  XNOR2_X1 U7989 ( .A(n6352), .B(n7030), .ZN(n6354) );
  NOR2_X1 U7990 ( .A1(n9889), .A2(n7808), .ZN(n6353) );
  AOI21_X1 U7991 ( .B1(n9769), .B2(n6489), .A(n6353), .ZN(n6355) );
  XNOR2_X1 U7992 ( .A(n6354), .B(n6355), .ZN(n7437) );
  INV_X1 U7993 ( .A(n6354), .ZN(n6356) );
  NAND2_X1 U7994 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  NAND2_X1 U7995 ( .A1(n7435), .A2(n6357), .ZN(n7494) );
  NAND2_X1 U7996 ( .A1(n7501), .A2(n7801), .ZN(n6359) );
  NAND2_X1 U7997 ( .A1(n9091), .A2(n6489), .ZN(n6358) );
  NAND2_X1 U7998 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  XNOR2_X1 U7999 ( .A(n6360), .B(n7030), .ZN(n6363) );
  NAND2_X1 U8000 ( .A1(n7501), .A2(n6489), .ZN(n6362) );
  NAND2_X1 U8001 ( .A1(n6482), .A2(n9091), .ZN(n6361) );
  NAND2_X1 U8002 ( .A1(n6362), .A2(n6361), .ZN(n6364) );
  NAND2_X1 U8003 ( .A1(n6363), .A2(n6364), .ZN(n7492) );
  INV_X1 U8004 ( .A(n6363), .ZN(n6366) );
  INV_X1 U8005 ( .A(n6364), .ZN(n6365) );
  NAND2_X1 U8006 ( .A1(n6366), .A2(n6365), .ZN(n7491) );
  NAND2_X1 U8007 ( .A1(n9634), .A2(n7801), .ZN(n6368) );
  NAND2_X1 U8008 ( .A1(n6394), .A2(n9090), .ZN(n6367) );
  NAND2_X1 U8009 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  XNOR2_X1 U8010 ( .A(n6369), .B(n7804), .ZN(n6372) );
  NOR2_X1 U8011 ( .A1(n7499), .A2(n7808), .ZN(n6370) );
  AOI21_X1 U8012 ( .B1(n9634), .B2(n6489), .A(n6370), .ZN(n6373) );
  XNOR2_X1 U8013 ( .A(n6372), .B(n6373), .ZN(n7542) );
  INV_X1 U8014 ( .A(n7542), .ZN(n6371) );
  INV_X1 U8015 ( .A(n6372), .ZN(n6375) );
  INV_X1 U8016 ( .A(n6373), .ZN(n6374) );
  NAND2_X1 U8017 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  NAND2_X1 U8018 ( .A1(n7618), .A2(n7801), .ZN(n6378) );
  NAND2_X1 U8019 ( .A1(n9606), .A2(n7806), .ZN(n6377) );
  NAND2_X1 U8020 ( .A1(n6378), .A2(n6377), .ZN(n6379) );
  XNOR2_X1 U8021 ( .A(n6379), .B(n7030), .ZN(n6381) );
  NOR2_X1 U8022 ( .A1(n7808), .A2(n9627), .ZN(n6380) );
  AOI21_X1 U8023 ( .B1(n7618), .B2(n6489), .A(n6380), .ZN(n6382) );
  XNOR2_X1 U8024 ( .A(n6381), .B(n6382), .ZN(n7621) );
  INV_X1 U8025 ( .A(n6381), .ZN(n6383) );
  NAND2_X1 U8026 ( .A1(n6383), .A2(n6382), .ZN(n6384) );
  NAND2_X1 U8027 ( .A1(n9637), .A2(n7801), .ZN(n6386) );
  NAND2_X1 U8028 ( .A1(n6394), .A2(n9089), .ZN(n6385) );
  NAND2_X1 U8029 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  XNOR2_X1 U8030 ( .A(n6387), .B(n7804), .ZN(n7668) );
  NOR2_X1 U8031 ( .A1(n9474), .A2(n7808), .ZN(n6388) );
  AOI21_X1 U8032 ( .B1(n9637), .B2(n6489), .A(n6388), .ZN(n7667) );
  AND2_X1 U8033 ( .A1(n7668), .A2(n7667), .ZN(n6389) );
  NAND2_X1 U8034 ( .A1(n8962), .A2(n7801), .ZN(n6391) );
  NAND2_X1 U8035 ( .A1(n6394), .A2(n9605), .ZN(n6390) );
  NAND2_X1 U8036 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  XNOR2_X1 U8037 ( .A(n6392), .B(n7804), .ZN(n8952) );
  NOR2_X1 U8038 ( .A1(n8135), .A2(n7808), .ZN(n6393) );
  AOI21_X1 U8039 ( .B1(n8962), .B2(n6489), .A(n6393), .ZN(n6398) );
  NAND2_X1 U8040 ( .A1(n8952), .A2(n6398), .ZN(n6407) );
  NAND2_X1 U8041 ( .A1(n9083), .A2(n7801), .ZN(n6396) );
  NAND2_X1 U8042 ( .A1(n6394), .A2(n9458), .ZN(n6395) );
  NAND2_X1 U8043 ( .A1(n6396), .A2(n6395), .ZN(n6397) );
  XNOR2_X1 U8044 ( .A(n6397), .B(n7804), .ZN(n6406) );
  INV_X1 U8045 ( .A(n8952), .ZN(n6399) );
  INV_X1 U8046 ( .A(n6398), .ZN(n8951) );
  NAND2_X1 U8047 ( .A1(n6399), .A2(n8951), .ZN(n6404) );
  AND2_X1 U8048 ( .A1(n6406), .A2(n6404), .ZN(n6400) );
  NAND2_X1 U8049 ( .A1(n6401), .A2(n6400), .ZN(n9068) );
  NAND2_X1 U8050 ( .A1(n9083), .A2(n7806), .ZN(n6403) );
  NAND2_X1 U8051 ( .A1(n6482), .A2(n9458), .ZN(n6402) );
  NAND2_X1 U8052 ( .A1(n6403), .A2(n6402), .ZN(n9071) );
  NAND2_X1 U8053 ( .A1(n9068), .A2(n9071), .ZN(n6410) );
  INV_X1 U8054 ( .A(n6404), .ZN(n6405) );
  INV_X1 U8055 ( .A(n6406), .ZN(n6408) );
  AND2_X1 U8056 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  NAND2_X1 U8057 ( .A1(n6410), .A2(n9069), .ZN(n9000) );
  INV_X1 U8058 ( .A(n9000), .ZN(n6417) );
  NAND2_X1 U8059 ( .A1(n9364), .A2(n7801), .ZN(n6412) );
  NAND2_X1 U8060 ( .A1(n9341), .A2(n6489), .ZN(n6411) );
  NAND2_X1 U8061 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  XNOR2_X1 U8062 ( .A(n6413), .B(n7030), .ZN(n6418) );
  NAND2_X1 U8063 ( .A1(n9364), .A2(n6489), .ZN(n6415) );
  OR2_X1 U8064 ( .A1(n9080), .A2(n7808), .ZN(n6414) );
  NAND2_X1 U8065 ( .A1(n6415), .A2(n6414), .ZN(n6419) );
  AND2_X1 U8066 ( .A1(n6418), .A2(n6419), .ZN(n9001) );
  INV_X1 U8067 ( .A(n6418), .ZN(n6421) );
  INV_X1 U8068 ( .A(n6419), .ZN(n6420) );
  NAND2_X1 U8069 ( .A1(n6421), .A2(n6420), .ZN(n8999) );
  NAND2_X1 U8070 ( .A1(n9453), .A2(n7801), .ZN(n6423) );
  NAND2_X1 U8071 ( .A1(n9459), .A2(n6489), .ZN(n6422) );
  NAND2_X1 U8072 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  XNOR2_X1 U8073 ( .A(n6424), .B(n7030), .ZN(n6426) );
  AND2_X1 U8074 ( .A1(n6482), .A2(n9459), .ZN(n6425) );
  AOI21_X1 U8075 ( .B1(n9453), .B2(n7806), .A(n6425), .ZN(n6427) );
  XNOR2_X1 U8076 ( .A(n6426), .B(n6427), .ZN(n9014) );
  INV_X1 U8077 ( .A(n6426), .ZN(n6428) );
  NAND2_X1 U8078 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  NAND2_X1 U8079 ( .A1(n9329), .A2(n7801), .ZN(n6431) );
  OR2_X1 U8080 ( .A1(n6433), .A2(n6308), .ZN(n6430) );
  NAND2_X1 U8081 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  XNOR2_X1 U8082 ( .A(n6432), .B(n7804), .ZN(n9047) );
  NOR2_X1 U8083 ( .A1(n6433), .A2(n7808), .ZN(n6434) );
  AOI21_X1 U8084 ( .B1(n9329), .B2(n7806), .A(n6434), .ZN(n9046) );
  NAND2_X1 U8085 ( .A1(n9434), .A2(n7801), .ZN(n6436) );
  NAND2_X1 U8086 ( .A1(n9444), .A2(n6489), .ZN(n6435) );
  NAND2_X1 U8087 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  XNOR2_X1 U8088 ( .A(n6437), .B(n7030), .ZN(n6439) );
  AND2_X1 U8089 ( .A1(n9444), .A2(n6482), .ZN(n6438) );
  AOI21_X1 U8090 ( .B1(n9434), .B2(n7806), .A(n6438), .ZN(n6440) );
  XNOR2_X1 U8091 ( .A(n6439), .B(n6440), .ZN(n8974) );
  INV_X1 U8092 ( .A(n6439), .ZN(n6441) );
  NAND2_X1 U8093 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  NAND2_X1 U8094 ( .A1(n9295), .A2(n7801), .ZN(n6444) );
  NAND2_X1 U8095 ( .A1(n9436), .A2(n6489), .ZN(n6443) );
  NAND2_X1 U8096 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  XNOR2_X1 U8097 ( .A(n6445), .B(n7030), .ZN(n6447) );
  AND2_X1 U8098 ( .A1(n9436), .A2(n6482), .ZN(n6446) );
  AOI21_X1 U8099 ( .B1(n9295), .B2(n7806), .A(n6446), .ZN(n6448) );
  XNOR2_X1 U8100 ( .A(n6447), .B(n6448), .ZN(n9029) );
  INV_X1 U8101 ( .A(n6447), .ZN(n6449) );
  NAND2_X1 U8102 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  NAND2_X1 U8103 ( .A1(n9284), .A2(n7801), .ZN(n6452) );
  NAND2_X1 U8104 ( .A1(n9412), .A2(n6489), .ZN(n6451) );
  NAND2_X1 U8105 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  XNOR2_X1 U8106 ( .A(n6453), .B(n7030), .ZN(n6455) );
  NOR2_X1 U8107 ( .A1(n9293), .A2(n7808), .ZN(n6454) );
  AOI21_X1 U8108 ( .B1(n9284), .B2(n6489), .A(n6454), .ZN(n6456) );
  XNOR2_X1 U8109 ( .A(n6455), .B(n6456), .ZN(n8981) );
  INV_X1 U8110 ( .A(n6455), .ZN(n6457) );
  AND2_X1 U8111 ( .A1(n9421), .A2(n6482), .ZN(n6458) );
  AOI21_X1 U8112 ( .B1(n9267), .B2(n7806), .A(n6458), .ZN(n6462) );
  NAND2_X1 U8113 ( .A1(n9267), .A2(n7801), .ZN(n6460) );
  NAND2_X1 U8114 ( .A1(n9421), .A2(n6489), .ZN(n6459) );
  NAND2_X1 U8115 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  XNOR2_X1 U8116 ( .A(n6461), .B(n7030), .ZN(n9039) );
  NAND2_X1 U8117 ( .A1(n9409), .A2(n7801), .ZN(n6465) );
  NAND2_X1 U8118 ( .A1(n9413), .A2(n7806), .ZN(n6464) );
  NAND2_X1 U8119 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  XNOR2_X1 U8120 ( .A(n6466), .B(n7030), .ZN(n6468) );
  AND2_X1 U8121 ( .A1(n9413), .A2(n6482), .ZN(n6467) );
  AOI21_X1 U8122 ( .B1(n9409), .B2(n6489), .A(n6467), .ZN(n8965) );
  XNOR2_X1 U8123 ( .A(n6470), .B(n6469), .ZN(n9023) );
  NAND2_X1 U8124 ( .A1(n9022), .A2(n9023), .ZN(n9021) );
  OAI22_X1 U8125 ( .A1(n9213), .A2(n6308), .B1(n9398), .B2(n7808), .ZN(n6476)
         );
  NAND2_X1 U8126 ( .A1(n9394), .A2(n7801), .ZN(n6473) );
  NAND2_X1 U8127 ( .A1(n9196), .A2(n7806), .ZN(n6472) );
  NAND2_X1 U8128 ( .A1(n6473), .A2(n6472), .ZN(n6474) );
  XNOR2_X1 U8129 ( .A(n6474), .B(n7030), .ZN(n6475) );
  XOR2_X1 U8130 ( .A(n6476), .B(n6475), .Z(n8990) );
  INV_X1 U8131 ( .A(n6475), .ZN(n6478) );
  INV_X1 U8132 ( .A(n6476), .ZN(n6477) );
  NAND2_X1 U8133 ( .A1(n9201), .A2(n7801), .ZN(n6480) );
  NAND2_X1 U8134 ( .A1(n9216), .A2(n7806), .ZN(n6479) );
  NAND2_X1 U8135 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  XNOR2_X1 U8136 ( .A(n6481), .B(n7030), .ZN(n6484) );
  AND2_X1 U8137 ( .A1(n9216), .A2(n6482), .ZN(n6483) );
  AOI21_X1 U8138 ( .B1(n9201), .B2(n7806), .A(n6483), .ZN(n6485) );
  XNOR2_X1 U8139 ( .A(n6484), .B(n6485), .ZN(n9058) );
  NAND2_X1 U8140 ( .A1(n6484), .A2(n6486), .ZN(n6487) );
  NOR2_X1 U8141 ( .A1(n9199), .A2(n7808), .ZN(n6488) );
  AOI21_X1 U8142 ( .B1(n9385), .B2(n6489), .A(n6488), .ZN(n7800) );
  NAND2_X1 U8143 ( .A1(n9385), .A2(n7801), .ZN(n6491) );
  OR2_X1 U8144 ( .A1(n9199), .A2(n6308), .ZN(n6490) );
  NAND2_X1 U8145 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  XNOR2_X1 U8146 ( .A(n6492), .B(n7030), .ZN(n7813) );
  XOR2_X1 U8147 ( .A(n7800), .B(n7813), .Z(n6493) );
  INV_X1 U8148 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10361) );
  NOR2_X1 U8149 ( .A1(n6494), .A2(n10361), .ZN(n6495) );
  OAI21_X1 U8150 ( .B1(n6547), .B2(n6495), .A(n6548), .ZN(n6583) );
  NOR2_X1 U8151 ( .A1(n7555), .A2(P1_U3084), .ZN(n6496) );
  NOR2_X1 U8152 ( .A1(n6591), .A2(n7009), .ZN(n6512) );
  NOR2_X1 U8153 ( .A1(n9892), .A2(n6608), .ZN(n6502) );
  OR2_X1 U8154 ( .A1(n6498), .A2(n6497), .ZN(n7031) );
  AND2_X1 U8155 ( .A1(n9797), .A2(n7031), .ZN(n6499) );
  NOR2_X1 U8156 ( .A1(n7009), .A2(n6499), .ZN(n6500) );
  NAND2_X1 U8157 ( .A1(n6591), .A2(n6500), .ZN(n7237) );
  NOR2_X1 U8158 ( .A1(n7239), .A2(n9902), .ZN(n6501) );
  NAND2_X1 U8159 ( .A1(n6591), .A2(n6502), .ZN(n6505) );
  INV_X1 U8160 ( .A(n6503), .ZN(n6504) );
  NAND2_X1 U8161 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  NAND2_X1 U8162 ( .A1(n6506), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6507) );
  INV_X1 U8163 ( .A(n6591), .ZN(n6509) );
  OR2_X1 U8164 ( .A1(n7009), .A2(n7031), .ZN(n8383) );
  NOR2_X1 U8165 ( .A1(n8383), .A2(n8382), .ZN(n6508) );
  NAND2_X1 U8166 ( .A1(n6509), .A2(n6508), .ZN(n9062) );
  OAI22_X1 U8167 ( .A1(n8995), .A2(n9062), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6510), .ZN(n6514) );
  NOR2_X1 U8168 ( .A1(n7031), .A2(n6872), .ZN(n6511) );
  NAND2_X1 U8169 ( .A1(n6512), .A2(n6511), .ZN(n9079) );
  NOR2_X1 U8170 ( .A1(n9182), .A2(n9079), .ZN(n6513) );
  AOI211_X1 U8171 ( .C1(n9186), .C2(n9076), .A(n6514), .B(n6513), .ZN(n6515)
         );
  INV_X1 U8172 ( .A(n6516), .ZN(n6517) );
  NAND2_X1 U8173 ( .A1(n6518), .A2(n6517), .ZN(P1_U3212) );
  OR2_X2 U8174 ( .A1(n6620), .A2(P1_U3084), .ZN(n9095) );
  INV_X1 U8175 ( .A(n6554), .ZN(n6520) );
  NAND2_X1 U8176 ( .A1(n7856), .A2(P1_U3084), .ZN(n9541) );
  INV_X1 U8177 ( .A(n9541), .ZN(n9545) );
  AOI22_X1 U8178 ( .A1(n9545), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n6868), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6522) );
  OAI21_X1 U8179 ( .B1(n6530), .B2(n9548), .A(n6522), .ZN(P1_U3352) );
  AOI22_X1 U8180 ( .A1(n9545), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6886), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6523) );
  OAI21_X1 U8181 ( .B1(n6525), .B2(n9548), .A(n6523), .ZN(P1_U3351) );
  NAND2_X1 U8182 ( .A1(n7856), .A2(P2_U3152), .ZN(n8944) );
  NOR2_X1 U8183 ( .A1(n7856), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8947) );
  AOI22_X1 U8184 ( .A1(n8947), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6729), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6524) );
  OAI21_X1 U8185 ( .B1(n6526), .B2(n8944), .A(n6524), .ZN(P2_U3355) );
  INV_X1 U8186 ( .A(n8947), .ZN(n7789) );
  OAI222_X1 U8187 ( .A1(n7789), .A2(n4851), .B1(n8944), .B2(n6525), .C1(
        P2_U3152), .C2(n4741), .ZN(P2_U3356) );
  INV_X1 U8188 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6527) );
  INV_X1 U8189 ( .A(n6634), .ZN(n9559) );
  OAI222_X1 U8190 ( .A1(n9541), .A2(n6527), .B1(n9548), .B2(n6526), .C1(
        P1_U3084), .C2(n9559), .ZN(P1_U3350) );
  INV_X1 U8191 ( .A(n6528), .ZN(n6531) );
  OAI222_X1 U8192 ( .A1(n9541), .A2(n6529), .B1(n9548), .B2(n6531), .C1(
        P1_U3084), .C2(n4792), .ZN(P1_U3349) );
  OAI222_X1 U8193 ( .A1(n7789), .A2(n5829), .B1(n8949), .B2(n6530), .C1(
        P2_U3152), .C2(n6658), .ZN(P2_U3357) );
  OAI222_X1 U8194 ( .A1(n7789), .A2(n6532), .B1(n8949), .B2(n6531), .C1(
        P2_U3152), .C2(n6765), .ZN(P2_U3354) );
  INV_X1 U8195 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6534) );
  INV_X1 U8196 ( .A(n6533), .ZN(n6535) );
  INV_X1 U8197 ( .A(n6635), .ZN(n9682) );
  OAI222_X1 U8198 ( .A1(n9541), .A2(n6534), .B1(n9548), .B2(n6535), .C1(
        P1_U3084), .C2(n9682), .ZN(P1_U3348) );
  INV_X1 U8199 ( .A(n6724), .ZN(n6756) );
  OAI222_X1 U8200 ( .A1(n7789), .A2(n4663), .B1(n8949), .B2(n6535), .C1(
        P2_U3152), .C2(n6756), .ZN(P2_U3353) );
  INV_X1 U8201 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6537) );
  INV_X1 U8202 ( .A(n6536), .ZN(n6538) );
  OAI222_X1 U8203 ( .A1(n9541), .A2(n6537), .B1(n9548), .B2(n6538), .C1(
        P1_U3084), .C2(n9697), .ZN(P1_U3347) );
  OAI222_X1 U8204 ( .A1(n7789), .A2(n6539), .B1(n8949), .B2(n6538), .C1(
        P2_U3152), .C2(n6776), .ZN(P2_U3352) );
  INV_X1 U8205 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10405) );
  INV_X1 U8206 ( .A(n6540), .ZN(n6541) );
  OAI222_X1 U8207 ( .A1(n9541), .A2(n10405), .B1(n9548), .B2(n6541), .C1(
        P1_U3084), .C2(n4799), .ZN(P1_U3346) );
  INV_X1 U8208 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6542) );
  INV_X1 U8209 ( .A(n6721), .ZN(n6786) );
  OAI222_X1 U8210 ( .A1(n7789), .A2(n6542), .B1(n8949), .B2(n6541), .C1(
        P2_U3152), .C2(n6786), .ZN(P2_U3351) );
  INV_X1 U8211 ( .A(n6543), .ZN(n6545) );
  INV_X1 U8212 ( .A(n6847), .ZN(n6645) );
  OAI222_X1 U8213 ( .A1(n9541), .A2(n6544), .B1(n9548), .B2(n6545), .C1(
        P1_U3084), .C2(n6645), .ZN(P1_U3345) );
  INV_X1 U8214 ( .A(n6718), .ZN(n6797) );
  OAI222_X1 U8215 ( .A1(n7789), .A2(n6546), .B1(n8949), .B2(n6545), .C1(
        P2_U3152), .C2(n6797), .ZN(P2_U3350) );
  INV_X1 U8216 ( .A(n6548), .ZN(n6549) );
  AOI22_X1 U8217 ( .A1(n9823), .A2(n10361), .B1(n6552), .B2(n6549), .ZN(
        P1_U3440) );
  INV_X1 U8218 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6553) );
  INV_X1 U8219 ( .A(n6550), .ZN(n6551) );
  AOI22_X1 U8220 ( .A1(n9823), .A2(n6553), .B1(n6552), .B2(n6551), .ZN(
        P1_U3441) );
  NAND2_X1 U8221 ( .A1(n6554), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8070) );
  INV_X1 U8222 ( .A(n8070), .ZN(n7553) );
  NAND2_X1 U8223 ( .A1(n9943), .A2(n6555), .ZN(n6556) );
  NAND2_X1 U8224 ( .A1(n6556), .A2(n5860), .ZN(n6557) );
  OAI21_X1 U8225 ( .B1(n9943), .B2(n7553), .A(n6557), .ZN(n8617) );
  NOR2_X1 U8226 ( .A1(n9932), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8227 ( .A(n6558), .ZN(n6560) );
  INV_X1 U8228 ( .A(n9707), .ZN(n6848) );
  OAI222_X1 U8229 ( .A1(n9541), .A2(n6559), .B1(n9548), .B2(n6560), .C1(n6848), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8230 ( .A(n6952), .ZN(n6745) );
  OAI222_X1 U8231 ( .A1(n7789), .A2(n6561), .B1(n8949), .B2(n6560), .C1(n6745), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8232 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U8233 ( .A1(n6562), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U8234 ( .A1(n6563), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U8235 ( .A1(n6564), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6565) );
  NAND3_X1 U8236 ( .A1(n6567), .A2(n6566), .A3(n6565), .ZN(n9140) );
  NAND2_X1 U8237 ( .A1(P1_U4006), .A2(n9140), .ZN(n6568) );
  OAI21_X1 U8238 ( .B1(P1_U4006), .B2(n6569), .A(n6568), .ZN(P1_U3586) );
  INV_X1 U8239 ( .A(n6570), .ZN(n6582) );
  AOI22_X1 U8240 ( .A1(n7174), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8947), .ZN(n6571) );
  OAI21_X1 U8241 ( .B1(n6582), .B2(n8944), .A(n6571), .ZN(P2_U3347) );
  INV_X1 U8242 ( .A(n6572), .ZN(n6575) );
  INV_X1 U8243 ( .A(n6850), .ZN(n9726) );
  OAI222_X1 U8244 ( .A1(n9541), .A2(n6573), .B1(n9548), .B2(n6575), .C1(n9726), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8245 ( .A(n7092), .ZN(n6961) );
  OAI222_X1 U8246 ( .A1(P2_U3152), .A2(n6961), .B1(n8949), .B2(n6575), .C1(
        n6574), .C2(n7789), .ZN(P2_U3348) );
  INV_X1 U8247 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6581) );
  AND2_X1 U8248 ( .A1(n9804), .A2(n9796), .ZN(n8330) );
  NOR2_X1 U8249 ( .A1(n9806), .A2(n8330), .ZN(n8215) );
  NAND2_X1 U8250 ( .A1(n7031), .A2(n7011), .ZN(n6576) );
  OR2_X1 U8251 ( .A1(n8215), .A2(n6576), .ZN(n6578) );
  NAND2_X1 U8252 ( .A1(n9096), .A2(n9863), .ZN(n6577) );
  NAND2_X1 U8253 ( .A1(n6578), .A2(n6577), .ZN(n7014) );
  INV_X1 U8254 ( .A(n7014), .ZN(n6579) );
  OAI21_X1 U8255 ( .B1(n9796), .B2(n7011), .A(n6579), .ZN(n6586) );
  NAND2_X1 U8256 ( .A1(n6586), .A2(n9911), .ZN(n6580) );
  OAI21_X1 U8257 ( .B1(n9911), .B2(n6581), .A(n6580), .ZN(P1_U3454) );
  INV_X1 U8258 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10438) );
  INV_X1 U8259 ( .A(n6997), .ZN(n6853) );
  OAI222_X1 U8260 ( .A1(n9541), .A2(n10438), .B1(n9548), .B2(n6582), .C1(n6853), .C2(P1_U3084), .ZN(P1_U3342) );
  NOR2_X1 U8261 ( .A1(n6583), .A2(n7239), .ZN(n6584) );
  NAND2_X1 U8262 ( .A1(n6586), .A2(n9928), .ZN(n6587) );
  OAI21_X1 U8263 ( .B1(n9928), .B2(n6283), .A(n6587), .ZN(P1_U3523) );
  AOI22_X1 U8264 ( .A1(n9064), .A2(n9096), .B1(n9082), .B2(n7012), .ZN(n6594)
         );
  OAI21_X1 U8265 ( .B1(n6590), .B2(n6589), .A(n6588), .ZN(n6873) );
  AOI21_X1 U8266 ( .B1(n6591), .B2(n9902), .A(n7239), .ZN(n6592) );
  NAND2_X1 U8267 ( .A1(n6592), .A2(n7237), .ZN(n6688) );
  AOI22_X1 U8268 ( .A1(n6873), .A2(n9056), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6688), .ZN(n6593) );
  NAND2_X1 U8269 ( .A1(n6594), .A2(n6593), .ZN(P1_U3230) );
  INV_X1 U8270 ( .A(n6595), .ZN(n6649) );
  AOI22_X1 U8271 ( .A1(n7323), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8947), .ZN(n6596) );
  OAI21_X1 U8272 ( .B1(n6649), .B2(n8944), .A(n6596), .ZN(P2_U3346) );
  NAND2_X1 U8273 ( .A1(P2_U3966), .A2(n5012), .ZN(n6597) );
  OAI21_X1 U8274 ( .B1(P2_U3966), .B2(n5176), .A(n6597), .ZN(P2_U3575) );
  XNOR2_X1 U8275 ( .A(n6599), .B(n6598), .ZN(n6600) );
  XOR2_X1 U8276 ( .A(n6601), .B(n6600), .Z(n6606) );
  AOI22_X1 U8277 ( .A1(n9064), .A2(n6602), .B1(n9074), .B2(n9804), .ZN(n6605)
         );
  NAND2_X1 U8278 ( .A1(n8333), .A2(n9892), .ZN(n9826) );
  NOR2_X1 U8279 ( .A1(n6688), .A2(n9826), .ZN(n6603) );
  AOI21_X1 U8280 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6688), .A(n6603), .ZN(
        n6604) );
  OAI211_X1 U8281 ( .C1(n6606), .C2(n9085), .A(n6605), .B(n6604), .ZN(P1_U3220) );
  INV_X1 U8282 ( .A(n7555), .ZN(n6607) );
  NAND2_X1 U8283 ( .A1(n6608), .A2(n6607), .ZN(n6609) );
  NAND2_X1 U8284 ( .A1(n6620), .A2(n6609), .ZN(n6622) );
  OR2_X1 U8285 ( .A1(n6622), .A2(n6610), .ZN(n9097) );
  NAND2_X1 U8286 ( .A1(n9097), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8287 ( .A(n8381), .ZN(n9098) );
  NAND2_X1 U8288 ( .A1(n9098), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9547) );
  NOR2_X1 U8289 ( .A1(n6622), .A2(n9547), .ZN(n6619) );
  INV_X1 U8290 ( .A(n6619), .ZN(n8081) );
  NOR2_X1 U8291 ( .A1(n6847), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6611) );
  AOI21_X1 U8292 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6847), .A(n6611), .ZN(
        n6618) );
  NOR2_X1 U8293 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n9113), .ZN(n6612) );
  AOI21_X1 U8294 ( .B1(n9113), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6612), .ZN(
        n9115) );
  NAND2_X1 U8295 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6865) );
  AOI21_X1 U8296 ( .B1(n6868), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6863), .ZN(
        n6883) );
  XNOR2_X1 U8297 ( .A(n6886), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6882) );
  NOR2_X1 U8298 ( .A1(n6883), .A2(n6882), .ZN(n6881) );
  AOI21_X1 U8299 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6886), .A(n6881), .ZN(
        n9556) );
  NAND2_X1 U8300 ( .A1(n6634), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6613) );
  OAI21_X1 U8301 ( .B1(n6634), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6613), .ZN(
        n9555) );
  NOR2_X1 U8302 ( .A1(n9671), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6614) );
  AOI21_X1 U8303 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9671), .A(n6614), .ZN(
        n9662) );
  XNOR2_X1 U8304 ( .A(n6635), .B(n6615), .ZN(n9674) );
  AOI22_X1 U8305 ( .A1(n9675), .A2(n9674), .B1(n6615), .B2(n9682), .ZN(n9691)
         );
  INV_X1 U8306 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6616) );
  MUX2_X1 U8307 ( .A(n6616), .B(P1_REG2_REG_6__SCAN_IN), .S(n9697), .Z(n9690)
         );
  AND2_X1 U8308 ( .A1(n9691), .A2(n9690), .ZN(n9693) );
  OAI21_X1 U8309 ( .B1(n6618), .B2(n6617), .A(n6840), .ZN(n6647) );
  INV_X1 U8310 ( .A(P1_U3083), .ZN(n6621) );
  NAND2_X1 U8311 ( .A1(n9134), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6644) );
  INV_X1 U8312 ( .A(n6622), .ZN(n6624) );
  NOR2_X1 U8313 ( .A1(n8382), .A2(P1_U3084), .ZN(n9542) );
  AND2_X1 U8314 ( .A1(n9542), .A2(n8381), .ZN(n6623) );
  OR2_X1 U8315 ( .A1(n6847), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U8316 ( .A1(n6847), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U8317 ( .A1(n6626), .A2(n6625), .ZN(n6640) );
  OR2_X1 U8318 ( .A1(n9113), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U8319 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n9113), .ZN(n6627) );
  AOI21_X1 U8320 ( .B1(n9113), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6627), .ZN(
        n9109) );
  NOR2_X1 U8321 ( .A1(n9671), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6628) );
  AOI21_X1 U8322 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9671), .A(n6628), .ZN(
        n9666) );
  INV_X1 U8323 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6629) );
  XNOR2_X1 U8324 ( .A(n6886), .B(n6629), .ZN(n6879) );
  INV_X1 U8325 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6630) );
  XNOR2_X1 U8326 ( .A(n6868), .B(n6630), .ZN(n6861) );
  AND2_X1 U8327 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6860) );
  NAND2_X1 U8328 ( .A1(n6861), .A2(n6860), .ZN(n6859) );
  NAND2_X1 U8329 ( .A1(n6868), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8330 ( .A1(n6859), .A2(n6631), .ZN(n6878) );
  NAND2_X1 U8331 ( .A1(n6879), .A2(n6878), .ZN(n6877) );
  INV_X1 U8332 ( .A(n6877), .ZN(n6632) );
  AOI21_X1 U8333 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n6886), .A(n6632), .ZN(
        n9553) );
  NAND2_X1 U8334 ( .A1(n6634), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6633) );
  OAI21_X1 U8335 ( .B1(n6634), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6633), .ZN(
        n9552) );
  NOR2_X1 U8336 ( .A1(n9553), .A2(n9552), .ZN(n9551) );
  AOI21_X1 U8337 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6634), .A(n9551), .ZN(
        n9665) );
  NAND2_X1 U8338 ( .A1(n9666), .A2(n9665), .ZN(n9664) );
  OAI21_X1 U8339 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9671), .A(n9664), .ZN(
        n9677) );
  XNOR2_X1 U8340 ( .A(n6635), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9678) );
  NOR2_X1 U8341 ( .A1(n9677), .A2(n9678), .ZN(n9676) );
  AOI21_X1 U8342 ( .B1(n6635), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9676), .ZN(
        n9689) );
  INV_X1 U8343 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6636) );
  MUX2_X1 U8344 ( .A(n6636), .B(P1_REG1_REG_6__SCAN_IN), .S(n9697), .Z(n9688)
         );
  NAND2_X1 U8345 ( .A1(n9689), .A2(n9688), .ZN(n9687) );
  OAI21_X1 U8346 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6637), .A(n9687), .ZN(
        n9110) );
  NAND2_X1 U8347 ( .A1(n9109), .A2(n9110), .ZN(n9108) );
  NAND2_X1 U8348 ( .A1(n6638), .A2(n9108), .ZN(n6639) );
  NOR2_X1 U8349 ( .A1(n6640), .A2(n6639), .ZN(n6846) );
  AOI21_X1 U8350 ( .B1(n6640), .B2(n6639), .A(n6846), .ZN(n6642) );
  NAND2_X1 U8351 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7414) );
  INV_X1 U8352 ( .A(n7414), .ZN(n6641) );
  AOI21_X1 U8353 ( .B1(n9744), .B2(n6642), .A(n6641), .ZN(n6643) );
  OAI211_X1 U8354 ( .C1(n9739), .C2(n6645), .A(n6644), .B(n6643), .ZN(n6646)
         );
  AOI21_X1 U8355 ( .B1(n9735), .B2(n6647), .A(n6646), .ZN(n6648) );
  INV_X1 U8356 ( .A(n6648), .ZN(P1_U3249) );
  INV_X1 U8357 ( .A(n7139), .ZN(n6995) );
  OAI222_X1 U8358 ( .A1(n9541), .A2(n10419), .B1(n9548), .B2(n6649), .C1(
        P1_U3084), .C2(n6995), .ZN(P1_U3341) );
  NAND2_X1 U8359 ( .A1(n9413), .A2(P1_U4006), .ZN(n6650) );
  OAI21_X1 U8360 ( .B1(P1_U4006), .B2(n5177), .A(n6650), .ZN(P1_U3578) );
  INV_X1 U8361 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8427) );
  MUX2_X1 U8362 ( .A(n8427), .B(P2_REG2_REG_1__SCAN_IN), .S(n6658), .Z(n6680)
         );
  NAND3_X1 U8363 ( .A1(n6680), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U8364 ( .A1(n6679), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6701) );
  INV_X1 U8365 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6895) );
  MUX2_X1 U8366 ( .A(n6895), .B(P2_REG2_REG_2__SCAN_IN), .S(n6660), .Z(n6700)
         );
  AOI21_X1 U8367 ( .B1(n6702), .B2(n6701), .A(n6700), .ZN(n6699) );
  AOI21_X1 U8368 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6660), .A(n6699), .ZN(
        n6731) );
  INV_X1 U8369 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6651) );
  MUX2_X1 U8370 ( .A(n6651), .B(P2_REG2_REG_3__SCAN_IN), .S(n6729), .Z(n6730)
         );
  XNOR2_X1 U8371 ( .A(n6731), .B(n6730), .ZN(n6672) );
  NAND2_X1 U8372 ( .A1(n9943), .A2(n6830), .ZN(n6654) );
  INV_X1 U8373 ( .A(n6652), .ZN(n6653) );
  NAND3_X1 U8374 ( .A1(n6654), .A2(n8070), .A3(n6653), .ZN(n6663) );
  NAND2_X1 U8375 ( .A1(n6663), .A2(n5860), .ZN(n6656) );
  INV_X1 U8376 ( .A(P2_U3966), .ZN(n6655) );
  NAND2_X1 U8377 ( .A1(n6656), .A2(n6655), .ZN(n6669) );
  NOR2_X1 U8378 ( .A1(n6668), .A2(n4484), .ZN(n6657) );
  NOR2_X1 U8379 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5850), .ZN(n6667) );
  XNOR2_X1 U8380 ( .A(n6658), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6675) );
  AND2_X1 U8381 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6674) );
  NAND2_X1 U8382 ( .A1(n6675), .A2(n6674), .ZN(n6673) );
  INV_X1 U8383 ( .A(n6673), .ZN(n6659) );
  AOI21_X1 U8384 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6679), .A(n6659), .ZN(
        n6696) );
  XNOR2_X1 U8385 ( .A(n6660), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6695) );
  NOR2_X1 U8386 ( .A1(n6696), .A2(n6695), .ZN(n6694) );
  NAND2_X1 U8387 ( .A1(n6729), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6661) );
  OAI21_X1 U8388 ( .B1(n6729), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6661), .ZN(
        n6664) );
  AND2_X1 U8389 ( .A1(n5860), .A2(n4484), .ZN(n6662) );
  AOI211_X1 U8390 ( .C1(n6665), .C2(n6664), .A(n6707), .B(n9934), .ZN(n6666)
         );
  AOI211_X1 U8391 ( .C1(n9932), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6667), .B(
        n6666), .ZN(n6671) );
  NAND2_X1 U8392 ( .A1(n8611), .A2(n6729), .ZN(n6670) );
  OAI211_X1 U8393 ( .C1(n6672), .C2(n9935), .A(n6671), .B(n6670), .ZN(P2_U3248) );
  INV_X1 U8394 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10063) );
  OAI211_X1 U8395 ( .C1(n6675), .C2(n6674), .A(n9929), .B(n6673), .ZN(n6677)
         );
  INV_X1 U8396 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10338) );
  NAND2_X1 U8397 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6676) );
  OAI211_X1 U8398 ( .C1(n10063), .C2(n8617), .A(n6677), .B(n6676), .ZN(n6678)
         );
  AOI21_X1 U8399 ( .B1(n6679), .B2(n8611), .A(n6678), .ZN(n6683) );
  AND2_X1 U8400 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6681) );
  OAI211_X1 U8401 ( .C1(n6681), .C2(n6680), .A(n9930), .B(n6702), .ZN(n6682)
         );
  NAND2_X1 U8402 ( .A1(n6683), .A2(n6682), .ZN(P2_U3246) );
  INV_X1 U8403 ( .A(n6684), .ZN(n6685) );
  AOI21_X1 U8404 ( .B1(n6687), .B2(n6686), .A(n6685), .ZN(n6692) );
  AOI22_X1 U8405 ( .A1(n9064), .A2(n9094), .B1(n9074), .B2(n9096), .ZN(n6691)
         );
  AOI22_X1 U8406 ( .A1(n9082), .A2(n6689), .B1(n6688), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6690) );
  OAI211_X1 U8407 ( .C1(n6692), .C2(n9085), .A(n6691), .B(n6690), .ZN(P1_U3235) );
  INV_X1 U8408 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6693) );
  NOR2_X1 U8409 ( .A1(n8617), .A2(n6693), .ZN(n6698) );
  AOI211_X1 U8410 ( .C1(n6696), .C2(n6695), .A(n6694), .B(n9934), .ZN(n6697)
         );
  AOI211_X1 U8411 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(P2_U3152), .A(n6698), .B(
        n6697), .ZN(n6706) );
  INV_X1 U8412 ( .A(n6699), .ZN(n6704) );
  NAND3_X1 U8413 ( .A1(n6702), .A2(n6701), .A3(n6700), .ZN(n6703) );
  NAND3_X1 U8414 ( .A1(n9930), .A2(n6704), .A3(n6703), .ZN(n6705) );
  OAI211_X1 U8415 ( .C1(n9933), .C2(n4741), .A(n6706), .B(n6705), .ZN(P2_U3247) );
  NOR2_X1 U8416 ( .A1(n5944), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7188) );
  INV_X1 U8417 ( .A(n6776), .ZN(n6711) );
  NAND2_X1 U8418 ( .A1(n6727), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6708) );
  OAI21_X1 U8419 ( .B1(n6727), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6708), .ZN(
        n6757) );
  AOI21_X1 U8420 ( .B1(n6727), .B2(P2_REG1_REG_4__SCAN_IN), .A(n4504), .ZN(
        n6748) );
  NAND2_X1 U8421 ( .A1(n6724), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8422 ( .B1(n6724), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6709), .ZN(
        n6747) );
  INV_X1 U8423 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6710) );
  MUX2_X1 U8424 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6710), .S(n6776), .Z(n6767)
         );
  NAND2_X1 U8425 ( .A1(n6721), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6712) );
  OAI21_X1 U8426 ( .B1(n6721), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6712), .ZN(
        n6778) );
  NOR2_X1 U8427 ( .A1(n4525), .A2(n6778), .ZN(n6777) );
  INV_X1 U8428 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6713) );
  MUX2_X1 U8429 ( .A(n6713), .B(P2_REG1_REG_8__SCAN_IN), .S(n6718), .Z(n6788)
         );
  INV_X1 U8430 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6714) );
  MUX2_X1 U8431 ( .A(n6714), .B(P2_REG1_REG_9__SCAN_IN), .S(n6952), .Z(n6715)
         );
  AOI211_X1 U8432 ( .C1(n6716), .C2(n6715), .A(n6946), .B(n9934), .ZN(n6717)
         );
  AOI211_X1 U8433 ( .C1(n9932), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7188), .B(
        n6717), .ZN(n6744) );
  NAND2_X1 U8434 ( .A1(n6718), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6738) );
  INV_X1 U8435 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6719) );
  MUX2_X1 U8436 ( .A(n6719), .B(P2_REG2_REG_8__SCAN_IN), .S(n6718), .Z(n6720)
         );
  INV_X1 U8437 ( .A(n6720), .ZN(n6793) );
  NAND2_X1 U8438 ( .A1(n6721), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6737) );
  INV_X1 U8439 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6722) );
  MUX2_X1 U8440 ( .A(n6722), .B(P2_REG2_REG_7__SCAN_IN), .S(n6721), .Z(n6723)
         );
  INV_X1 U8441 ( .A(n6723), .ZN(n6783) );
  INV_X1 U8442 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6736) );
  MUX2_X1 U8443 ( .A(n6736), .B(P2_REG2_REG_6__SCAN_IN), .S(n6776), .Z(n6772)
         );
  NAND2_X1 U8444 ( .A1(n6724), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6735) );
  INV_X1 U8445 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6725) );
  MUX2_X1 U8446 ( .A(n6725), .B(P2_REG2_REG_5__SCAN_IN), .S(n6724), .Z(n6726)
         );
  INV_X1 U8447 ( .A(n6726), .ZN(n6752) );
  NAND2_X1 U8448 ( .A1(n6727), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6734) );
  INV_X1 U8449 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6728) );
  MUX2_X1 U8450 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6728), .S(n6727), .Z(n6761)
         );
  NAND2_X1 U8451 ( .A1(n6729), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6733) );
  OR2_X1 U8452 ( .A1(n6731), .A2(n6730), .ZN(n6732) );
  NAND2_X1 U8453 ( .A1(n6733), .A2(n6732), .ZN(n6762) );
  NAND2_X1 U8454 ( .A1(n6761), .A2(n6762), .ZN(n6760) );
  NAND2_X1 U8455 ( .A1(n6734), .A2(n6760), .ZN(n6753) );
  NAND2_X1 U8456 ( .A1(n6752), .A2(n6753), .ZN(n6751) );
  NAND2_X1 U8457 ( .A1(n6735), .A2(n6751), .ZN(n6773) );
  NAND2_X1 U8458 ( .A1(n6772), .A2(n6773), .ZN(n6771) );
  OAI21_X1 U8459 ( .B1(n6776), .B2(n6736), .A(n6771), .ZN(n6782) );
  NAND2_X1 U8460 ( .A1(n6783), .A2(n6782), .ZN(n6781) );
  NAND2_X1 U8461 ( .A1(n6737), .A2(n6781), .ZN(n6794) );
  NAND2_X1 U8462 ( .A1(n6793), .A2(n6794), .ZN(n6792) );
  NAND2_X1 U8463 ( .A1(n6738), .A2(n6792), .ZN(n6742) );
  INV_X1 U8464 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6739) );
  MUX2_X1 U8465 ( .A(n6739), .B(P2_REG2_REG_9__SCAN_IN), .S(n6952), .Z(n6740)
         );
  INV_X1 U8466 ( .A(n6740), .ZN(n6741) );
  NAND2_X1 U8467 ( .A1(n6741), .A2(n6742), .ZN(n6953) );
  OAI211_X1 U8468 ( .C1(n6742), .C2(n6741), .A(n9930), .B(n6953), .ZN(n6743)
         );
  OAI211_X1 U8469 ( .C1(n9933), .C2(n6745), .A(n6744), .B(n6743), .ZN(P2_U3254) );
  INV_X1 U8470 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U8471 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10232), .ZN(n6750) );
  AOI211_X1 U8472 ( .C1(n6748), .C2(n6747), .A(n6746), .B(n9934), .ZN(n6749)
         );
  AOI211_X1 U8473 ( .C1(n9932), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6750), .B(
        n6749), .ZN(n6755) );
  OAI211_X1 U8474 ( .C1(n6753), .C2(n6752), .A(n9930), .B(n6751), .ZN(n6754)
         );
  OAI211_X1 U8475 ( .C1(n9933), .C2(n6756), .A(n6755), .B(n6754), .ZN(P2_U3250) );
  INV_X1 U8476 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U8477 ( .A1(n10403), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7067) );
  AOI211_X1 U8478 ( .C1(n6758), .C2(n6757), .A(n4504), .B(n9934), .ZN(n6759)
         );
  AOI211_X1 U8479 ( .C1(n9932), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7067), .B(
        n6759), .ZN(n6764) );
  OAI211_X1 U8480 ( .C1(n6762), .C2(n6761), .A(n9930), .B(n6760), .ZN(n6763)
         );
  OAI211_X1 U8481 ( .C1(n9933), .C2(n6765), .A(n6764), .B(n6763), .ZN(P2_U3249) );
  NAND2_X1 U8482 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7079) );
  INV_X1 U8483 ( .A(n7079), .ZN(n6770) );
  AOI211_X1 U8484 ( .C1(n6768), .C2(n6767), .A(n6766), .B(n9934), .ZN(n6769)
         );
  AOI211_X1 U8485 ( .C1(n9932), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6770), .B(
        n6769), .ZN(n6775) );
  OAI211_X1 U8486 ( .C1(n6773), .C2(n6772), .A(n9930), .B(n6771), .ZN(n6774)
         );
  OAI211_X1 U8487 ( .C1(n9933), .C2(n6776), .A(n6775), .B(n6774), .ZN(P2_U3251) );
  INV_X1 U8488 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10362) );
  NOR2_X1 U8489 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10362), .ZN(n6780) );
  AOI211_X1 U8490 ( .C1(n4525), .C2(n6778), .A(n6777), .B(n9934), .ZN(n6779)
         );
  AOI211_X1 U8491 ( .C1(n9932), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6780), .B(
        n6779), .ZN(n6785) );
  OAI211_X1 U8492 ( .C1(n6783), .C2(n6782), .A(n9930), .B(n6781), .ZN(n6784)
         );
  OAI211_X1 U8493 ( .C1(n9933), .C2(n6786), .A(n6785), .B(n6784), .ZN(P2_U3252) );
  INV_X1 U8494 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10458) );
  NOR2_X1 U8495 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10458), .ZN(n6791) );
  AOI211_X1 U8496 ( .C1(n6789), .C2(n6788), .A(n6787), .B(n9934), .ZN(n6790)
         );
  AOI211_X1 U8497 ( .C1(n9932), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6791), .B(
        n6790), .ZN(n6796) );
  OAI211_X1 U8498 ( .C1(n6794), .C2(n6793), .A(n9930), .B(n6792), .ZN(n6795)
         );
  OAI211_X1 U8499 ( .C1(n9933), .C2(n6797), .A(n6796), .B(n6795), .ZN(P2_U3253) );
  INV_X1 U8500 ( .A(n6798), .ZN(n6838) );
  AOI22_X1 U8501 ( .A1(n7685), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9545), .ZN(n6799) );
  OAI21_X1 U8502 ( .B1(n6838), .B2(n9548), .A(n6799), .ZN(P1_U3339) );
  INV_X1 U8503 ( .A(n6800), .ZN(n6801) );
  INV_X1 U8504 ( .A(n7451), .ZN(n7137) );
  OAI222_X1 U8505 ( .A1(n9541), .A2(n10387), .B1(n9548), .B2(n6801), .C1(n7137), .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U8506 ( .A(n7426), .ZN(n7321) );
  OAI222_X1 U8507 ( .A1(n7789), .A2(n6802), .B1(n8949), .B2(n6801), .C1(n7321), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  OAI21_X1 U8508 ( .B1(n6805), .B2(n6804), .A(n6803), .ZN(n6811) );
  OAI22_X1 U8509 ( .A1(n9062), .A2(n5294), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6806), .ZN(n6807) );
  AOI21_X1 U8510 ( .B1(n9064), .B2(n9781), .A(n6807), .ZN(n6809) );
  NAND2_X1 U8511 ( .A1(n9076), .A2(n6806), .ZN(n6808) );
  OAI211_X1 U8512 ( .C1(n9840), .C2(n9067), .A(n6809), .B(n6808), .ZN(n6810)
         );
  AOI21_X1 U8513 ( .B1(n6811), .B2(n9056), .A(n6810), .ZN(n6812) );
  INV_X1 U8514 ( .A(n6812), .ZN(P1_U3216) );
  NOR2_X1 U8515 ( .A1(n6813), .A2(P2_U3152), .ZN(n6974) );
  NAND2_X1 U8516 ( .A1(n6981), .A2(n6974), .ZN(n6814) );
  NOR2_X1 U8517 ( .A1(n6972), .A2(n6814), .ZN(n6815) );
  NAND2_X1 U8518 ( .A1(n6976), .A2(n6815), .ZN(n6824) );
  NAND2_X1 U8519 ( .A1(n8784), .A2(n6255), .ZN(n7895) );
  OR2_X1 U8520 ( .A1(n7895), .A2(n7868), .ZN(n6900) );
  INV_X1 U8521 ( .A(n6900), .ZN(n6817) );
  NAND2_X1 U8522 ( .A1(n6892), .A2(n6818), .ZN(n6819) );
  NAND2_X1 U8523 ( .A1(n6820), .A2(n6819), .ZN(n6903) );
  INV_X1 U8524 ( .A(n6915), .ZN(n8550) );
  NAND2_X1 U8525 ( .A1(n8550), .A2(n6821), .ZN(n7940) );
  NAND2_X1 U8526 ( .A1(n6915), .A2(n6941), .ZN(n7938) );
  NAND2_X1 U8527 ( .A1(n6903), .A2(n6902), .ZN(n6823) );
  NAND2_X1 U8528 ( .A1(n6915), .A2(n6821), .ZN(n6822) );
  INV_X1 U8529 ( .A(n6927), .ZN(n8549) );
  NAND2_X1 U8530 ( .A1(n6927), .A2(n8442), .ZN(n7923) );
  XNOR2_X1 U8531 ( .A(n6926), .B(n7873), .ZN(n9971) );
  OR2_X1 U8532 ( .A1(n6824), .A2(n8784), .ZN(n8422) );
  NOR2_X1 U8533 ( .A1(n6917), .A2(n9950), .ZN(n6897) );
  NAND2_X1 U8534 ( .A1(n6897), .A2(n6821), .ZN(n6896) );
  OAI211_X1 U8535 ( .C1(n4667), .C2(n9967), .A(n10014), .B(n6969), .ZN(n9966)
         );
  OAI22_X1 U8536 ( .A1(n8422), .A2(n9966), .B1(n8821), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n6825) );
  AOI21_X1 U8537 ( .B1(n8792), .B2(n9971), .A(n6825), .ZN(n6837) );
  NAND2_X1 U8538 ( .A1(n6914), .A2(n9950), .ZN(n8424) );
  NAND2_X1 U8539 ( .A1(n7937), .A2(n8424), .ZN(n7927) );
  NAND2_X1 U8540 ( .A1(n7927), .A2(n7935), .ZN(n6889) );
  INV_X1 U8541 ( .A(n6889), .ZN(n6826) );
  NAND2_X1 U8542 ( .A1(n6826), .A2(n7869), .ZN(n6891) );
  NAND2_X1 U8543 ( .A1(n6891), .A2(n7938), .ZN(n6827) );
  NAND2_X1 U8544 ( .A1(n6827), .A2(n7930), .ZN(n6921) );
  OAI21_X1 U8545 ( .B1(n7930), .B2(n6827), .A(n6921), .ZN(n6829) );
  NAND2_X1 U8546 ( .A1(n6254), .A2(n8784), .ZN(n8058) );
  NAND2_X1 U8547 ( .A1(n7868), .A2(n6255), .ZN(n7863) );
  OAI22_X1 U8548 ( .A1(n6964), .A2(n8762), .B1(n6915), .B2(n8764), .ZN(n6828)
         );
  AOI21_X1 U8549 ( .B1(n6829), .B2(n8804), .A(n6828), .ZN(n6835) );
  MUX2_X1 U8550 ( .A(n6254), .B(n6830), .S(n8061), .Z(n6833) );
  INV_X1 U8551 ( .A(n6831), .ZN(n6832) );
  NAND2_X1 U8552 ( .A1(n6833), .A2(n6832), .ZN(n7568) );
  INV_X1 U8553 ( .A(n7568), .ZN(n8786) );
  NAND2_X1 U8554 ( .A1(n9971), .A2(n8786), .ZN(n6834) );
  AND2_X1 U8555 ( .A1(n6835), .A2(n6834), .ZN(n9968) );
  MUX2_X1 U8556 ( .A(n6651), .B(n9968), .S(n8696), .Z(n6836) );
  OAI211_X1 U8557 ( .C1(n9967), .C2(n8823), .A(n6837), .B(n6836), .ZN(P2_U3293) );
  INV_X1 U8558 ( .A(n7649), .ZN(n7644) );
  OAI222_X1 U8559 ( .A1(n7789), .A2(n6839), .B1(n8949), .B2(n6838), .C1(n7644), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8560 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6858) );
  OAI21_X1 U8561 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6847), .A(n6840), .ZN(
        n9703) );
  XNOR2_X1 U8562 ( .A(n9707), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n9704) );
  NOR2_X1 U8563 ( .A1(n9703), .A2(n9704), .ZN(n9702) );
  XNOR2_X1 U8564 ( .A(n6850), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9716) );
  MUX2_X1 U8565 ( .A(n9622), .B(P1_REG2_REG_11__SCAN_IN), .S(n6997), .Z(n6841)
         );
  INV_X1 U8566 ( .A(n6841), .ZN(n6842) );
  OAI21_X1 U8567 ( .B1(n6843), .B2(n6842), .A(n6996), .ZN(n6844) );
  NAND2_X1 U8568 ( .A1(n6844), .A2(n9735), .ZN(n6857) );
  INV_X1 U8569 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6845) );
  MUX2_X1 U8570 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6845), .S(n6997), .Z(n6852)
         );
  XOR2_X1 U8571 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9707), .Z(n9710) );
  AOI21_X1 U8572 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6847), .A(n6846), .ZN(
        n9709) );
  AOI22_X1 U8573 ( .A1(n9710), .A2(n9709), .B1(n9926), .B2(n6848), .ZN(n9719)
         );
  INV_X1 U8574 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6849) );
  MUX2_X1 U8575 ( .A(n6849), .B(P1_REG1_REG_10__SCAN_IN), .S(n6850), .Z(n9718)
         );
  OAI21_X1 U8576 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6850), .A(n9722), .ZN(
        n6851) );
  NAND2_X1 U8577 ( .A1(n6851), .A2(n6852), .ZN(n6990) );
  OAI21_X1 U8578 ( .B1(n6852), .B2(n6851), .A(n6990), .ZN(n6855) );
  AND2_X1 U8579 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7546) );
  NOR2_X1 U8580 ( .A1(n9739), .A2(n6853), .ZN(n6854) );
  AOI211_X1 U8581 ( .C1(n9744), .C2(n6855), .A(n7546), .B(n6854), .ZN(n6856)
         );
  OAI211_X1 U8582 ( .C1(n9748), .C2(n6858), .A(n6857), .B(n6856), .ZN(P1_U3252) );
  INV_X1 U8583 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6870) );
  INV_X1 U8584 ( .A(n9739), .ZN(n9708) );
  INV_X1 U8585 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9799) );
  OAI211_X1 U8586 ( .C1(n6861), .C2(n6860), .A(n9744), .B(n6859), .ZN(n6862)
         );
  OAI21_X1 U8587 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9799), .A(n6862), .ZN(n6867) );
  AOI211_X1 U8588 ( .C1(n6865), .C2(n6864), .A(n6863), .B(n9715), .ZN(n6866)
         );
  AOI211_X1 U8589 ( .C1(n9708), .C2(n6868), .A(n6867), .B(n6866), .ZN(n6869)
         );
  OAI21_X1 U8590 ( .B1(n9748), .B2(n6870), .A(n6869), .ZN(P1_U3242) );
  INV_X1 U8591 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10061) );
  INV_X1 U8592 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6876) );
  INV_X1 U8593 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7017) );
  NAND2_X1 U8594 ( .A1(n9098), .A2(n7017), .ZN(n6871) );
  NAND2_X1 U8595 ( .A1(n6872), .A2(n6871), .ZN(n9100) );
  MUX2_X1 U8596 ( .A(n6876), .B(n6873), .S(n8381), .Z(n6874) );
  NOR2_X1 U8597 ( .A1(n6874), .A2(n9100), .ZN(n6875) );
  AOI211_X1 U8598 ( .C1(n6876), .C2(n9100), .A(n9095), .B(n6875), .ZN(n9669)
         );
  INV_X1 U8599 ( .A(n9669), .ZN(n6888) );
  INV_X1 U8600 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7033) );
  OAI211_X1 U8601 ( .C1(n6879), .C2(n6878), .A(n9744), .B(n6877), .ZN(n6880)
         );
  OAI21_X1 U8602 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7033), .A(n6880), .ZN(n6885) );
  AOI211_X1 U8603 ( .C1(n6883), .C2(n6882), .A(n6881), .B(n9715), .ZN(n6884)
         );
  AOI211_X1 U8604 ( .C1(n9708), .C2(n6886), .A(n6885), .B(n6884), .ZN(n6887)
         );
  OAI211_X1 U8605 ( .C1(n10061), .C2(n9748), .A(n6888), .B(n6887), .ZN(
        P1_U3243) );
  NAND2_X1 U8606 ( .A1(n6889), .A2(n6902), .ZN(n6890) );
  INV_X1 U8607 ( .A(n8804), .ZN(n8759) );
  AOI21_X1 U8608 ( .B1(n6891), .B2(n6890), .A(n8759), .ZN(n6894) );
  OAI22_X1 U8609 ( .A1(n6892), .A2(n8764), .B1(n6927), .B2(n8762), .ZN(n6893)
         );
  OR2_X1 U8610 ( .A1(n6894), .A2(n6893), .ZN(n9962) );
  NOR2_X1 U8611 ( .A1(n8696), .A2(n6895), .ZN(n6899) );
  OAI211_X1 U8612 ( .C1(n6897), .C2(n6821), .A(n6896), .B(n10014), .ZN(n9961)
         );
  INV_X1 U8613 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10390) );
  OAI22_X1 U8614 ( .A1(n8422), .A2(n9961), .B1(n10390), .B2(n8821), .ZN(n6898)
         );
  AOI211_X1 U8615 ( .C1(n8696), .C2(n9962), .A(n6899), .B(n6898), .ZN(n6905)
         );
  NAND2_X1 U8616 ( .A1(n7568), .A2(n6900), .ZN(n6901) );
  XNOR2_X1 U8617 ( .A(n6903), .B(n6902), .ZN(n9964) );
  AOI22_X1 U8618 ( .A1(n8826), .A2(n9964), .B1(n8620), .B2(n6941), .ZN(n6904)
         );
  NAND2_X1 U8619 ( .A1(n6905), .A2(n6904), .ZN(P2_U3294) );
  XNOR2_X1 U8620 ( .A(n6907), .B(n6906), .ZN(n6911) );
  INV_X1 U8621 ( .A(n8524), .ZN(n8475) );
  OAI22_X1 U8622 ( .A1(n6964), .A2(n8764), .B1(n7110), .B2(n8762), .ZN(n6967)
         );
  AOI22_X1 U8623 ( .A1(n8475), .A2(n6967), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6910) );
  INV_X1 U8624 ( .A(n8822), .ZN(n7102) );
  AOI22_X1 U8625 ( .A1(n8503), .A2(n7102), .B1(n8526), .B2(n6908), .ZN(n6909)
         );
  OAI211_X1 U8626 ( .C1(n8505), .C2(n6911), .A(n6910), .B(n6909), .ZN(P2_U3229) );
  XOR2_X1 U8627 ( .A(n6938), .B(n6936), .Z(n6913) );
  NOR2_X1 U8628 ( .A1(n6913), .A2(n6912), .ZN(n6937) );
  AOI21_X1 U8629 ( .B1(n6913), .B2(n6912), .A(n6937), .ZN(n6920) );
  OAI22_X1 U8630 ( .A1(n6914), .A2(n8764), .B1(n6915), .B2(n8762), .ZN(n8425)
         );
  NAND2_X1 U8631 ( .A1(n6916), .A2(n6974), .ZN(n7304) );
  AOI22_X1 U8632 ( .A1(n8475), .A2(n8425), .B1(n7304), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6919) );
  NAND2_X1 U8633 ( .A1(n8503), .A2(n6917), .ZN(n6918) );
  OAI211_X1 U8634 ( .C1(n6920), .C2(n8505), .A(n6919), .B(n6918), .ZN(P2_U3224) );
  NAND2_X1 U8635 ( .A1(n6921), .A2(n7923), .ZN(n6966) );
  NAND2_X1 U8636 ( .A1(n6964), .A2(n9973), .ZN(n7922) );
  NAND2_X1 U8637 ( .A1(n7922), .A2(n7918), .ZN(n7872) );
  INV_X1 U8638 ( .A(n7872), .ZN(n6922) );
  XNOR2_X1 U8639 ( .A(n6966), .B(n6922), .ZN(n6925) );
  NAND2_X1 U8640 ( .A1(n8547), .A2(n8810), .ZN(n6923) );
  OAI21_X1 U8641 ( .B1(n6927), .B2(n8764), .A(n6923), .ZN(n6924) );
  AOI21_X1 U8642 ( .B1(n6925), .B2(n8804), .A(n6924), .ZN(n9976) );
  NAND2_X1 U8643 ( .A1(n6927), .A2(n9967), .ZN(n6928) );
  NAND2_X1 U8644 ( .A1(n6929), .A2(n6928), .ZN(n6963) );
  XNOR2_X1 U8645 ( .A(n6963), .B(n7872), .ZN(n9978) );
  AOI22_X1 U8646 ( .A1(n8826), .A2(n9978), .B1(n8620), .B2(n9973), .ZN(n6933)
         );
  NOR2_X2 U8647 ( .A1(n8422), .A2(n10024), .ZN(n8816) );
  XNOR2_X1 U8648 ( .A(n6969), .B(n7070), .ZN(n9974) );
  INV_X1 U8649 ( .A(n6930), .ZN(n7069) );
  OAI22_X1 U8650 ( .A1(n8696), .A2(n6728), .B1(n7069), .B2(n8821), .ZN(n6931)
         );
  AOI21_X1 U8651 ( .B1(n8816), .B2(n9974), .A(n6931), .ZN(n6932) );
  OAI211_X1 U8652 ( .C1(n8788), .C2(n9976), .A(n6933), .B(n6932), .ZN(P2_U3292) );
  NAND2_X1 U8653 ( .A1(n6935), .A2(n6934), .ZN(n6940) );
  AOI21_X1 U8654 ( .B1(n6938), .B2(n4926), .A(n6937), .ZN(n6939) );
  XOR2_X1 U8655 ( .A(n6940), .B(n6939), .Z(n6944) );
  AOI22_X1 U8656 ( .A1(n8510), .A2(n4483), .B1(n8511), .B2(n8549), .ZN(n6943)
         );
  AOI22_X1 U8657 ( .A1(n8503), .A2(n6941), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n7304), .ZN(n6942) );
  OAI211_X1 U8658 ( .C1(n8505), .C2(n6944), .A(n6943), .B(n6942), .ZN(P2_U3239) );
  INV_X1 U8659 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U8660 ( .A1(P2_U3966), .A2(n8402), .ZN(n6945) );
  OAI21_X1 U8661 ( .B1(P2_U3966), .B2(n10181), .A(n6945), .ZN(P2_U3579) );
  NOR2_X1 U8662 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10462), .ZN(n6951) );
  AOI21_X1 U8663 ( .B1(n6952), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6946), .ZN(
        n6949) );
  INV_X1 U8664 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6947) );
  MUX2_X1 U8665 ( .A(n6947), .B(P2_REG1_REG_10__SCAN_IN), .S(n7092), .Z(n6948)
         );
  NOR2_X1 U8666 ( .A1(n6949), .A2(n6948), .ZN(n7091) );
  AOI211_X1 U8667 ( .C1(n6949), .C2(n6948), .A(n7091), .B(n9934), .ZN(n6950)
         );
  AOI211_X1 U8668 ( .C1(n9932), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6951), .B(
        n6950), .ZN(n6960) );
  NAND2_X1 U8669 ( .A1(n6952), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8670 ( .A1(n6954), .A2(n6953), .ZN(n6958) );
  INV_X1 U8671 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6955) );
  MUX2_X1 U8672 ( .A(n6955), .B(P2_REG2_REG_10__SCAN_IN), .S(n7092), .Z(n6956)
         );
  INV_X1 U8673 ( .A(n6956), .ZN(n6957) );
  NAND2_X1 U8674 ( .A1(n6957), .A2(n6958), .ZN(n7085) );
  OAI211_X1 U8675 ( .C1(n6958), .C2(n6957), .A(n9930), .B(n7085), .ZN(n6959)
         );
  OAI211_X1 U8676 ( .C1(n9933), .C2(n6961), .A(n6960), .B(n6959), .ZN(P2_U3255) );
  AND2_X1 U8677 ( .A1(n8061), .A2(n8784), .ZN(n6962) );
  NAND2_X1 U8678 ( .A1(n7786), .A2(n6962), .ZN(n9576) );
  NAND2_X1 U8679 ( .A1(n6964), .A2(n7070), .ZN(n6965) );
  INV_X1 U8680 ( .A(n8547), .ZN(n7104) );
  NAND2_X1 U8681 ( .A1(n7104), .A2(n7102), .ZN(n7924) );
  AND2_X1 U8682 ( .A1(n8822), .A2(n8547), .ZN(n7914) );
  INV_X1 U8683 ( .A(n7914), .ZN(n7919) );
  NAND2_X1 U8684 ( .A1(n7924), .A2(n7919), .ZN(n7871) );
  XNOR2_X1 U8685 ( .A(n7105), .B(n7871), .ZN(n8825) );
  INV_X1 U8686 ( .A(n10013), .ZN(n10022) );
  XNOR2_X1 U8687 ( .A(n7109), .B(n7871), .ZN(n6968) );
  AOI21_X1 U8688 ( .B1(n6968), .B2(n8804), .A(n6967), .ZN(n8819) );
  OAI211_X1 U8689 ( .C1(n6970), .C2(n8822), .A(n10014), .B(n7149), .ZN(n8827)
         );
  OAI211_X1 U8690 ( .C1(n8822), .C2(n10022), .A(n8819), .B(n8827), .ZN(n6971)
         );
  AOI21_X1 U8691 ( .B1(n10029), .B2(n8825), .A(n6971), .ZN(n6985) );
  INV_X1 U8692 ( .A(n6972), .ZN(n6975) );
  NAND3_X1 U8693 ( .A1(n6975), .A2(n6974), .A3(n6973), .ZN(n6977) );
  INV_X1 U8694 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6979) );
  OR2_X1 U8695 ( .A1(n10052), .A2(n6979), .ZN(n6980) );
  OAI21_X1 U8696 ( .B1(n6985), .B2(n10050), .A(n6980), .ZN(P2_U3525) );
  INV_X1 U8697 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6983) );
  OR2_X1 U8698 ( .A1(n10032), .A2(n6983), .ZN(n6984) );
  OAI21_X1 U8699 ( .B1(n6985), .B2(n10030), .A(n6984), .ZN(P2_U3466) );
  INV_X1 U8700 ( .A(n6986), .ZN(n6987) );
  OAI222_X1 U8701 ( .A1(n9541), .A2(n10393), .B1(n9548), .B2(n6987), .C1(
        P1_U3084), .C2(n7697), .ZN(P1_U3338) );
  INV_X1 U8702 ( .A(n8561), .ZN(n8553) );
  OAI222_X1 U8703 ( .A1(n7789), .A2(n6988), .B1(n8949), .B2(n6987), .C1(
        P2_U3152), .C2(n8553), .ZN(P2_U3343) );
  INV_X1 U8704 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6989) );
  MUX2_X1 U8705 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6989), .S(n7139), .Z(n6992)
         );
  OAI21_X1 U8706 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6997), .A(n6990), .ZN(
        n6991) );
  NAND2_X1 U8707 ( .A1(n6991), .A2(n6992), .ZN(n7132) );
  OAI21_X1 U8708 ( .B1(n6992), .B2(n6991), .A(n7132), .ZN(n7003) );
  NAND2_X1 U8709 ( .A1(n9134), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8710 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6993) );
  OAI211_X1 U8711 ( .C1(n9739), .C2(n6995), .A(n6994), .B(n6993), .ZN(n7002)
         );
  OAI21_X1 U8712 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6997), .A(n6996), .ZN(
        n7000) );
  NAND2_X1 U8713 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7139), .ZN(n6998) );
  OAI21_X1 U8714 ( .B1(n7139), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6998), .ZN(
        n6999) );
  AOI211_X1 U8715 ( .C1(n7000), .C2(n6999), .A(n9715), .B(n7138), .ZN(n7001)
         );
  AOI211_X1 U8716 ( .C1(n9744), .C2(n7003), .A(n7002), .B(n7001), .ZN(n7004)
         );
  INV_X1 U8717 ( .A(n7004), .ZN(P1_U3253) );
  NAND2_X1 U8718 ( .A1(n9164), .A2(P1_U4006), .ZN(n7005) );
  OAI21_X1 U8719 ( .B1(P1_U4006), .B2(n5195), .A(n7005), .ZN(P1_U3582) );
  INV_X1 U8720 ( .A(n7006), .ZN(n7007) );
  NAND2_X1 U8721 ( .A1(n7008), .A2(n7007), .ZN(n7032) );
  AND2_X1 U8722 ( .A1(n9816), .A2(n9814), .ZN(n9235) );
  INV_X1 U8723 ( .A(n9235), .ZN(n9326) );
  INV_X1 U8724 ( .A(n9797), .ZN(n9785) );
  OAI21_X1 U8725 ( .B1(n9326), .B2(n7011), .A(n9337), .ZN(n7013) );
  NAND2_X1 U8726 ( .A1(n7013), .A2(n7012), .ZN(n7016) );
  AOI22_X1 U8727 ( .A1(n7014), .A2(n9816), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9787), .ZN(n7015) );
  OAI211_X1 U8728 ( .C1(n9816), .C2(n7017), .A(n7016), .B(n7015), .ZN(P1_U3291) );
  AND2_X1 U8729 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9670) );
  AOI21_X1 U8730 ( .B1(n9074), .B2(n9094), .A(n9670), .ZN(n7019) );
  NAND2_X1 U8731 ( .A1(n9082), .A2(n9847), .ZN(n7018) );
  OAI211_X1 U8732 ( .C1(n9848), .C2(n9079), .A(n7019), .B(n7018), .ZN(n7025)
         );
  INV_X1 U8733 ( .A(n7020), .ZN(n7021) );
  AOI211_X1 U8734 ( .C1(n7023), .C2(n7022), .A(n9085), .B(n7021), .ZN(n7024)
         );
  AOI211_X1 U8735 ( .C1(n7294), .C2(n9076), .A(n7025), .B(n7024), .ZN(n7026)
         );
  INV_X1 U8736 ( .A(n7026), .ZN(P1_U3228) );
  NAND2_X1 U8737 ( .A1(n7027), .A2(n8213), .ZN(n7028) );
  NAND2_X1 U8738 ( .A1(n7029), .A2(n7028), .ZN(n9835) );
  INV_X1 U8739 ( .A(n9835), .ZN(n7042) );
  INV_X2 U8740 ( .A(n9816), .ZN(n9822) );
  OAI211_X1 U8741 ( .C1(n9793), .C2(n9832), .A(n7199), .B(n9794), .ZN(n9831)
         );
  OAI22_X1 U8742 ( .A1(n9361), .A2(n9831), .B1(n7033), .B2(n9800), .ZN(n7035)
         );
  NOR2_X1 U8743 ( .A1(n9337), .A2(n9832), .ZN(n7034) );
  AOI211_X1 U8744 ( .C1(n9822), .C2(P1_REG2_REG_2__SCAN_IN), .A(n7035), .B(
        n7034), .ZN(n7041) );
  INV_X1 U8745 ( .A(n7036), .ZN(n8337) );
  XNOR2_X1 U8746 ( .A(n8213), .B(n8337), .ZN(n7039) );
  INV_X1 U8747 ( .A(n9812), .ZN(n9900) );
  INV_X1 U8748 ( .A(n9866), .ZN(n9886) );
  OAI22_X1 U8749 ( .A1(n8334), .A2(n9886), .B1(n9849), .B2(n9888), .ZN(n7037)
         );
  AOI21_X1 U8750 ( .B1(n9835), .B2(n9900), .A(n7037), .ZN(n7038) );
  OAI21_X1 U8751 ( .B1(n7039), .B2(n9882), .A(n7038), .ZN(n9833) );
  NAND2_X1 U8752 ( .A1(n9833), .A2(n9816), .ZN(n7040) );
  OAI211_X1 U8753 ( .C1(n7042), .C2(n9818), .A(n7041), .B(n7040), .ZN(P1_U3289) );
  INV_X1 U8754 ( .A(n8076), .ZN(n7703) );
  INV_X1 U8755 ( .A(n7043), .ZN(n7044) );
  OAI222_X1 U8756 ( .A1(P1_U3084), .A2(n7703), .B1(n9548), .B2(n7044), .C1(
        n10360), .C2(n9541), .ZN(P1_U3337) );
  INV_X1 U8757 ( .A(n8578), .ZN(n8565) );
  OAI222_X1 U8758 ( .A1(n7789), .A2(n7045), .B1(n8949), .B2(n7044), .C1(n8565), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8759 ( .A(n7046), .ZN(n7131) );
  AOI22_X1 U8760 ( .A1(n9121), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9545), .ZN(n7047) );
  OAI21_X1 U8761 ( .B1(n7131), .B2(n9548), .A(n7047), .ZN(P1_U3336) );
  XNOR2_X1 U8762 ( .A(n7049), .B(n7048), .ZN(n7050) );
  XNOR2_X1 U8763 ( .A(n6338), .B(n7050), .ZN(n7055) );
  AND2_X1 U8764 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9112) );
  AOI21_X1 U8765 ( .B1(n9074), .B2(n9782), .A(n9112), .ZN(n7052) );
  NAND2_X1 U8766 ( .A1(n9076), .A2(n7401), .ZN(n7051) );
  OAI211_X1 U8767 ( .C1(n9875), .C2(n9079), .A(n7052), .B(n7051), .ZN(n7053)
         );
  AOI21_X1 U8768 ( .B1(n9082), .B2(n9879), .A(n7053), .ZN(n7054) );
  OAI21_X1 U8769 ( .B1(n7055), .B2(n9085), .A(n7054), .ZN(P1_U3211) );
  XNOR2_X1 U8770 ( .A(n7057), .B(n7056), .ZN(n7062) );
  INV_X1 U8771 ( .A(n7352), .ZN(n7058) );
  OAI22_X1 U8772 ( .A1(n8498), .A2(n7058), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10458), .ZN(n7060) );
  INV_X1 U8773 ( .A(n7353), .ZN(n9992) );
  OAI22_X1 U8774 ( .A1(n8499), .A2(n7381), .B1(n9992), .B2(n8529), .ZN(n7059)
         );
  AOI211_X1 U8775 ( .C1(n8510), .C2(n5015), .A(n7060), .B(n7059), .ZN(n7061)
         );
  OAI21_X1 U8776 ( .B1(n8505), .B2(n7062), .A(n7061), .ZN(P2_U3223) );
  NAND2_X1 U8777 ( .A1(n7064), .A2(n7063), .ZN(n7066) );
  XOR2_X1 U8778 ( .A(n7066), .B(n7065), .Z(n7074) );
  INV_X1 U8779 ( .A(n7067), .ZN(n7068) );
  OAI21_X1 U8780 ( .B1(n8498), .B2(n7069), .A(n7068), .ZN(n7072) );
  OAI22_X1 U8781 ( .A1(n8499), .A2(n7104), .B1(n7070), .B2(n8529), .ZN(n7071)
         );
  AOI211_X1 U8782 ( .C1(n8510), .C2(n8549), .A(n7072), .B(n7071), .ZN(n7073)
         );
  OAI21_X1 U8783 ( .B1(n7074), .B2(n8505), .A(n7073), .ZN(P2_U3232) );
  INV_X1 U8784 ( .A(n7075), .ZN(n7076) );
  AOI21_X1 U8785 ( .B1(n7078), .B2(n7077), .A(n7076), .ZN(n7084) );
  INV_X1 U8786 ( .A(n7152), .ZN(n7080) );
  OAI21_X1 U8787 ( .B1(n8498), .B2(n7080), .A(n7079), .ZN(n7082) );
  INV_X1 U8788 ( .A(n7155), .ZN(n9980) );
  OAI22_X1 U8789 ( .A1(n8499), .A2(n7358), .B1(n9980), .B2(n8529), .ZN(n7081)
         );
  AOI211_X1 U8790 ( .C1(n8510), .C2(n8547), .A(n7082), .B(n7081), .ZN(n7083)
         );
  OAI21_X1 U8791 ( .B1(n7084), .B2(n8505), .A(n7083), .ZN(P2_U3241) );
  NAND2_X1 U8792 ( .A1(n7092), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7086) );
  NAND2_X1 U8793 ( .A1(n7086), .A2(n7085), .ZN(n7089) );
  INV_X1 U8794 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7087) );
  MUX2_X1 U8795 ( .A(n7087), .B(P2_REG2_REG_11__SCAN_IN), .S(n7174), .Z(n7088)
         );
  NOR2_X1 U8796 ( .A1(n7089), .A2(n7088), .ZN(n7175) );
  AOI21_X1 U8797 ( .B1(n7089), .B2(n7088), .A(n7175), .ZN(n7101) );
  INV_X1 U8798 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7098) );
  INV_X1 U8799 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7090) );
  MUX2_X1 U8800 ( .A(n7090), .B(P2_REG1_REG_11__SCAN_IN), .S(n7174), .Z(n7094)
         );
  AOI21_X1 U8801 ( .B1(n7094), .B2(n7093), .A(n7166), .ZN(n7095) );
  NAND2_X1 U8802 ( .A1(n9929), .A2(n7095), .ZN(n7097) );
  INV_X1 U8803 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10459) );
  OR2_X1 U8804 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10459), .ZN(n7096) );
  OAI211_X1 U8805 ( .C1(n8617), .C2(n7098), .A(n7097), .B(n7096), .ZN(n7099)
         );
  AOI21_X1 U8806 ( .B1(n7174), .B2(n8611), .A(n7099), .ZN(n7100) );
  OAI21_X1 U8807 ( .B1(n7101), .B2(n9935), .A(n7100), .ZN(P2_U3256) );
  NAND2_X1 U8808 ( .A1(n7105), .A2(n7871), .ZN(n7103) );
  NAND2_X1 U8809 ( .A1(n7103), .A2(n7102), .ZN(n7107) );
  INV_X1 U8810 ( .A(n7110), .ZN(n8546) );
  OR2_X1 U8811 ( .A1(n7155), .A2(n8546), .ZN(n7108) );
  NAND2_X1 U8812 ( .A1(n7950), .A2(n7949), .ZN(n7266) );
  INV_X1 U8813 ( .A(n7266), .ZN(n7946) );
  XNOR2_X1 U8814 ( .A(n7267), .B(n7946), .ZN(n9989) );
  OAI21_X1 U8815 ( .B1(n7109), .B2(n7914), .A(n7924), .ZN(n7147) );
  OR2_X1 U8816 ( .A1(n7155), .A2(n7110), .ZN(n7943) );
  NAND2_X1 U8817 ( .A1(n7155), .A2(n7110), .ZN(n7948) );
  NAND2_X1 U8818 ( .A1(n7147), .A2(n7876), .ZN(n7146) );
  NAND2_X1 U8819 ( .A1(n7111), .A2(n7946), .ZN(n7274) );
  OAI211_X1 U8820 ( .C1(n7111), .C2(n7946), .A(n8804), .B(n7274), .ZN(n7113)
         );
  AOI22_X1 U8821 ( .A1(n8809), .A2(n8546), .B1(n8545), .B2(n8810), .ZN(n7112)
         );
  NAND2_X1 U8822 ( .A1(n7113), .A2(n7112), .ZN(n9987) );
  AOI21_X1 U8823 ( .B1(n7114), .B2(n8800), .A(n9987), .ZN(n7115) );
  MUX2_X1 U8824 ( .A(n6722), .B(n7115), .S(n8696), .Z(n7117) );
  INV_X1 U8825 ( .A(n8422), .ZN(n8829) );
  OAI211_X1 U8826 ( .C1(n9989), .C2(n8818), .A(n7117), .B(n7116), .ZN(P2_U3289) );
  INV_X1 U8827 ( .A(n7118), .ZN(n7120) );
  AOI21_X1 U8828 ( .B1(n7394), .B2(n8273), .A(n8223), .ZN(n7119) );
  OR3_X1 U8829 ( .A1(n7120), .A2(n9882), .A3(n7119), .ZN(n9894) );
  OAI21_X1 U8830 ( .B1(n4562), .B2(n5387), .A(n7121), .ZN(n9897) );
  INV_X1 U8831 ( .A(n9897), .ZN(n9899) );
  NAND2_X1 U8832 ( .A1(n9899), .A2(n9350), .ZN(n7129) );
  AOI211_X1 U8833 ( .C1(n9893), .C2(n7398), .A(n9615), .B(n9751), .ZN(n9890)
         );
  INV_X1 U8834 ( .A(n9893), .ZN(n7413) );
  NAND2_X1 U8835 ( .A1(n9816), .A2(n9863), .ZN(n9355) );
  INV_X1 U8836 ( .A(n9355), .ZN(n9322) );
  INV_X1 U8837 ( .A(n7418), .ZN(n7122) );
  OAI22_X1 U8838 ( .A1(n9816), .A2(n7123), .B1(n7122), .B2(n9800), .ZN(n7124)
         );
  AOI21_X1 U8839 ( .B1(n9322), .B2(n9092), .A(n7124), .ZN(n7126) );
  AND2_X1 U8840 ( .A1(n9816), .A2(n9866), .ZN(n9352) );
  NAND2_X1 U8841 ( .A1(n9352), .A2(n9864), .ZN(n7125) );
  OAI211_X1 U8842 ( .C1(n7413), .C2(n9337), .A(n7126), .B(n7125), .ZN(n7127)
         );
  AOI21_X1 U8843 ( .B1(n9890), .B2(n9755), .A(n7127), .ZN(n7128) );
  OAI211_X1 U8844 ( .C1(n9822), .C2(n9894), .A(n7129), .B(n7128), .ZN(P1_U3283) );
  INV_X1 U8845 ( .A(n8592), .ZN(n8585) );
  OAI222_X1 U8846 ( .A1(P2_U3152), .A2(n8585), .B1(n8949), .B2(n7131), .C1(
        n7130), .C2(n7789), .ZN(P2_U3341) );
  OAI21_X1 U8847 ( .B1(n7139), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7132), .ZN(
        n7135) );
  INV_X1 U8848 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7133) );
  MUX2_X1 U8849 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7133), .S(n7451), .Z(n7134)
         );
  NAND2_X1 U8850 ( .A1(n7134), .A2(n7135), .ZN(n7450) );
  OAI21_X1 U8851 ( .B1(n7135), .B2(n7134), .A(n7450), .ZN(n7144) );
  NAND2_X1 U8852 ( .A1(n9134), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7136) );
  NAND2_X1 U8853 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7671) );
  OAI211_X1 U8854 ( .C1(n9739), .C2(n7137), .A(n7136), .B(n7671), .ZN(n7143)
         );
  NAND2_X1 U8855 ( .A1(n7451), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7459) );
  OAI21_X1 U8856 ( .B1(n7451), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7459), .ZN(
        n7140) );
  AOI211_X1 U8857 ( .C1(n7141), .C2(n7140), .A(n7457), .B(n9715), .ZN(n7142)
         );
  AOI211_X1 U8858 ( .C1(n9744), .C2(n7144), .A(n7143), .B(n7142), .ZN(n7145)
         );
  INV_X1 U8859 ( .A(n7145), .ZN(P1_U3254) );
  OAI21_X1 U8860 ( .B1(n7876), .B2(n7147), .A(n7146), .ZN(n7148) );
  AOI222_X1 U8861 ( .A1(n8804), .A2(n7148), .B1(n5015), .B2(n8810), .C1(n8547), 
        .C2(n8809), .ZN(n9982) );
  INV_X1 U8862 ( .A(n7149), .ZN(n7151) );
  OAI21_X1 U8863 ( .B1(n7151), .B2(n9980), .A(n7150), .ZN(n9981) );
  AOI22_X1 U8864 ( .A1(n8788), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7152), .B2(
        n8800), .ZN(n7153) );
  OAI21_X1 U8865 ( .B1(n8629), .B2(n9981), .A(n7153), .ZN(n7154) );
  AOI21_X1 U8866 ( .B1(n8620), .B2(n7155), .A(n7154), .ZN(n7158) );
  XNOR2_X1 U8867 ( .A(n7156), .B(n7876), .ZN(n9985) );
  NAND2_X1 U8868 ( .A1(n9985), .A2(n8826), .ZN(n7157) );
  OAI211_X1 U8869 ( .C1(n9982), .C2(n8788), .A(n7158), .B(n7157), .ZN(P2_U3290) );
  XNOR2_X1 U8870 ( .A(n7160), .B(n7159), .ZN(n7165) );
  INV_X1 U8871 ( .A(n7388), .ZN(n7161) );
  OAI22_X1 U8872 ( .A1(n8498), .A2(n7161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10462), .ZN(n7163) );
  INV_X1 U8873 ( .A(n8542), .ZN(n7478) );
  OAI22_X1 U8874 ( .A1(n7381), .A2(n8500), .B1(n8499), .B2(n7478), .ZN(n7162)
         );
  AOI211_X1 U8875 ( .C1(n10004), .C2(n8503), .A(n7163), .B(n7162), .ZN(n7164)
         );
  OAI21_X1 U8876 ( .B1(n7165), .B2(n8505), .A(n7164), .ZN(P2_U3219) );
  INV_X1 U8877 ( .A(n7323), .ZN(n7183) );
  INV_X1 U8878 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7167) );
  MUX2_X1 U8879 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7167), .S(n7323), .Z(n7168)
         );
  OAI21_X1 U8880 ( .B1(n7169), .B2(n7168), .A(n7322), .ZN(n7173) );
  INV_X1 U8881 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7170) );
  NOR2_X1 U8882 ( .A1(n7170), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7472) );
  INV_X1 U8883 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7171) );
  NOR2_X1 U8884 ( .A1(n8617), .A2(n7171), .ZN(n7172) );
  AOI211_X1 U8885 ( .C1(n9929), .C2(n7173), .A(n7472), .B(n7172), .ZN(n7182)
         );
  INV_X1 U8886 ( .A(n7174), .ZN(n7176) );
  AOI21_X1 U8887 ( .B1(n7176), .B2(n7087), .A(n7175), .ZN(n7180) );
  INV_X1 U8888 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7177) );
  MUX2_X1 U8889 ( .A(n7177), .B(P2_REG2_REG_12__SCAN_IN), .S(n7323), .Z(n7178)
         );
  INV_X1 U8890 ( .A(n7178), .ZN(n7179) );
  NAND2_X1 U8891 ( .A1(n7179), .A2(n7180), .ZN(n7317) );
  OAI211_X1 U8892 ( .C1(n7180), .C2(n7179), .A(n9930), .B(n7317), .ZN(n7181)
         );
  OAI211_X1 U8893 ( .C1(n9933), .C2(n7183), .A(n7182), .B(n7181), .ZN(P2_U3257) );
  INV_X1 U8894 ( .A(n7184), .ZN(n7185) );
  AOI21_X1 U8895 ( .B1(n7187), .B2(n7186), .A(n7185), .ZN(n7194) );
  INV_X1 U8896 ( .A(n7285), .ZN(n7191) );
  INV_X1 U8897 ( .A(n7794), .ZN(n8543) );
  AOI22_X1 U8898 ( .A1(n8510), .A2(n8545), .B1(n8511), .B2(n8543), .ZN(n7190)
         );
  INV_X1 U8899 ( .A(n7188), .ZN(n7189) );
  OAI211_X1 U8900 ( .C1(n7191), .C2(n8498), .A(n7190), .B(n7189), .ZN(n7192)
         );
  AOI21_X1 U8901 ( .B1(n7377), .B2(n8492), .A(n7192), .ZN(n7193) );
  OAI21_X1 U8902 ( .B1(n7194), .B2(n8505), .A(n7193), .ZN(P2_U3233) );
  INV_X1 U8903 ( .A(n7195), .ZN(n8214) );
  XNOR2_X1 U8904 ( .A(n7196), .B(n8214), .ZN(n9844) );
  XNOR2_X1 U8905 ( .A(n8292), .B(n8214), .ZN(n7197) );
  NAND2_X1 U8906 ( .A1(n7197), .A2(n9808), .ZN(n9842) );
  INV_X1 U8907 ( .A(n9842), .ZN(n7205) );
  INV_X1 U8908 ( .A(n9352), .ZN(n9324) );
  INV_X1 U8909 ( .A(n9337), .ZN(n9770) );
  AOI22_X1 U8910 ( .A1(n9770), .A2(n7198), .B1(n9322), .B2(n9781), .ZN(n7203)
         );
  AOI21_X1 U8911 ( .B1(n7199), .B2(n7198), .A(n9615), .ZN(n7200) );
  NAND2_X1 U8912 ( .A1(n7200), .A2(n7295), .ZN(n9839) );
  OAI22_X1 U8913 ( .A1(n9361), .A2(n9839), .B1(n9800), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7201) );
  AOI21_X1 U8914 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n9822), .A(n7201), .ZN(
        n7202) );
  OAI211_X1 U8915 ( .C1(n5294), .C2(n9324), .A(n7203), .B(n7202), .ZN(n7204)
         );
  AOI21_X1 U8916 ( .B1(n7205), .B2(n9816), .A(n7204), .ZN(n7206) );
  OAI21_X1 U8917 ( .B1(n9818), .B2(n9844), .A(n7206), .ZN(P1_U3288) );
  OAI21_X1 U8918 ( .B1(n7208), .B2(n8219), .A(n7207), .ZN(n9873) );
  OAI211_X1 U8919 ( .C1(n9774), .C2(n7209), .A(n9794), .B(n7400), .ZN(n9867)
         );
  AOI22_X1 U8920 ( .A1(n9322), .A2(n9864), .B1(n9787), .B2(n7246), .ZN(n7210)
         );
  OAI21_X1 U8921 ( .B1(n9848), .B2(n9324), .A(n7210), .ZN(n7211) );
  AOI21_X1 U8922 ( .B1(n9770), .B2(n7238), .A(n7211), .ZN(n7212) );
  OAI21_X1 U8923 ( .B1(n9361), .B2(n9867), .A(n7212), .ZN(n7218) );
  INV_X1 U8924 ( .A(n8289), .ZN(n7214) );
  NAND2_X1 U8925 ( .A1(n9778), .A2(n7213), .ZN(n8101) );
  OAI21_X1 U8926 ( .B1(n7214), .B2(n9779), .A(n8101), .ZN(n7215) );
  XNOR2_X1 U8927 ( .A(n7215), .B(n8219), .ZN(n7216) );
  AND2_X1 U8928 ( .A1(n7216), .A2(n9808), .ZN(n9872) );
  MUX2_X1 U8929 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9872), .S(n9816), .Z(n7217)
         );
  AOI211_X1 U8930 ( .C1(n9350), .C2(n9873), .A(n7218), .B(n7217), .ZN(n7219)
         );
  INV_X1 U8931 ( .A(n7219), .ZN(P1_U3285) );
  INV_X1 U8932 ( .A(n8424), .ZN(n7221) );
  OR2_X1 U8933 ( .A1(n6914), .A2(n9950), .ZN(n7936) );
  INV_X1 U8934 ( .A(n7936), .ZN(n7220) );
  NOR2_X1 U8935 ( .A1(n7221), .A2(n7220), .ZN(n7867) );
  INV_X1 U8936 ( .A(n7867), .ZN(n9951) );
  AOI22_X1 U8937 ( .A1(n9951), .A2(n8804), .B1(n8810), .B2(n4483), .ZN(n9953)
         );
  INV_X1 U8938 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7222) );
  OAI22_X1 U8939 ( .A1(n8788), .A2(n9953), .B1(n7222), .B2(n8821), .ZN(n7223)
         );
  AOI21_X1 U8940 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8788), .A(n7223), .ZN(
        n7225) );
  OAI21_X1 U8941 ( .B1(n8816), .B2(n8620), .A(n9950), .ZN(n7224) );
  OAI211_X1 U8942 ( .C1(n7867), .C2(n8818), .A(n7225), .B(n7224), .ZN(P2_U3296) );
  INV_X1 U8943 ( .A(n7226), .ZN(n7228) );
  OAI222_X1 U8944 ( .A1(n7789), .A2(n7227), .B1(n8944), .B2(n7228), .C1(
        P2_U3152), .C2(n8590), .ZN(P2_U3340) );
  INV_X1 U8945 ( .A(n8077), .ZN(n9738) );
  OAI222_X1 U8946 ( .A1(n9541), .A2(n10389), .B1(n9548), .B2(n7228), .C1(
        P1_U3084), .C2(n9738), .ZN(P1_U3335) );
  NOR2_X1 U8947 ( .A1(n7229), .A2(n7230), .ZN(n7231) );
  AOI21_X1 U8948 ( .B1(n7230), .B2(n7229), .A(n7231), .ZN(n7258) );
  NAND2_X1 U8949 ( .A1(n7258), .A2(n7259), .ZN(n7257) );
  INV_X1 U8950 ( .A(n7231), .ZN(n7233) );
  AOI22_X1 U8951 ( .A1(n7257), .A2(n7233), .B1(n7234), .B2(n7232), .ZN(n7249)
         );
  INV_X1 U8952 ( .A(n7234), .ZN(n7235) );
  OAI21_X1 U8953 ( .B1(n7236), .B2(n7235), .A(n9056), .ZN(n7248) );
  INV_X1 U8954 ( .A(n7237), .ZN(n7240) );
  NAND2_X1 U8955 ( .A1(n7238), .A2(n9892), .ZN(n9868) );
  NOR3_X1 U8956 ( .A1(n7240), .A2(n9868), .A3(n7239), .ZN(n7245) );
  NAND2_X1 U8957 ( .A1(n9074), .A2(n9865), .ZN(n7243) );
  NOR2_X1 U8958 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7241), .ZN(n9695) );
  INV_X1 U8959 ( .A(n9695), .ZN(n7242) );
  OAI211_X1 U8960 ( .C1(n9079), .C2(n9887), .A(n7243), .B(n7242), .ZN(n7244)
         );
  AOI211_X1 U8961 ( .C1(n7246), .C2(n9076), .A(n7245), .B(n7244), .ZN(n7247)
         );
  OAI21_X1 U8962 ( .B1(n7249), .B2(n7248), .A(n7247), .ZN(P1_U3237) );
  XNOR2_X1 U8963 ( .A(n7251), .B(n7250), .ZN(n7256) );
  OAI22_X1 U8964 ( .A1(n8498), .A2(n7252), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10362), .ZN(n7253) );
  AOI21_X1 U8965 ( .B1(n8510), .B2(n8546), .A(n7253), .ZN(n7255) );
  OAI211_X1 U8966 ( .C1(n7256), .C2(n8505), .A(n7255), .B(n7254), .ZN(P2_U3215) );
  OAI21_X1 U8967 ( .B1(n7259), .B2(n7258), .A(n7257), .ZN(n7260) );
  NAND2_X1 U8968 ( .A1(n7260), .A2(n9056), .ZN(n7265) );
  AND2_X1 U8969 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9680) );
  AOI21_X1 U8970 ( .B1(n9074), .B2(n9781), .A(n9680), .ZN(n7262) );
  NAND2_X1 U8971 ( .A1(n9082), .A2(n9784), .ZN(n7261) );
  OAI211_X1 U8972 ( .C1(n9876), .C2(n9079), .A(n7262), .B(n7261), .ZN(n7263)
         );
  AOI21_X1 U8973 ( .B1(n9786), .B2(n9076), .A(n7263), .ZN(n7264) );
  NAND2_X1 U8974 ( .A1(n7265), .A2(n7264), .ZN(P1_U3225) );
  OR2_X1 U8975 ( .A1(n7377), .A2(n7381), .ZN(n7909) );
  NAND2_X1 U8976 ( .A1(n7377), .A2(n7381), .ZN(n7956) );
  OR2_X1 U8977 ( .A1(n7353), .A2(n7268), .ZN(n7953) );
  NAND2_X1 U8978 ( .A1(n7353), .A2(n7268), .ZN(n7954) );
  NAND2_X1 U8979 ( .A1(n7953), .A2(n7954), .ZN(n7355) );
  NAND2_X1 U8980 ( .A1(n7353), .A2(n8545), .ZN(n7269) );
  INV_X1 U8981 ( .A(n7379), .ZN(n7272) );
  AOI21_X1 U8982 ( .B1(n7278), .B2(n7273), .A(n7272), .ZN(n7283) );
  AOI22_X1 U8983 ( .A1(n8809), .A2(n8545), .B1(n8543), .B2(n8810), .ZN(n7282)
         );
  NAND2_X1 U8984 ( .A1(n7276), .A2(n7278), .ZN(n7380) );
  INV_X1 U8985 ( .A(n7380), .ZN(n7280) );
  AND3_X1 U8986 ( .A1(n7277), .A2(n7954), .A3(n7271), .ZN(n7279) );
  OAI21_X1 U8987 ( .B1(n7280), .B2(n7279), .A(n8804), .ZN(n7281) );
  OAI211_X1 U8988 ( .C1(n7283), .C2(n7568), .A(n7282), .B(n7281), .ZN(n10000)
         );
  INV_X1 U8989 ( .A(n10000), .ZN(n7290) );
  INV_X1 U8990 ( .A(n7283), .ZN(n10002) );
  INV_X1 U8991 ( .A(n7377), .ZN(n9998) );
  OR2_X1 U8992 ( .A1(n7351), .A2(n9998), .ZN(n7284) );
  NAND2_X1 U8993 ( .A1(n7386), .A2(n7284), .ZN(n9999) );
  AOI22_X1 U8994 ( .A1(n8788), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7285), .B2(
        n8800), .ZN(n7287) );
  NAND2_X1 U8995 ( .A1(n8620), .A2(n7377), .ZN(n7286) );
  OAI211_X1 U8996 ( .C1(n8629), .C2(n9999), .A(n7287), .B(n7286), .ZN(n7288)
         );
  AOI21_X1 U8997 ( .B1(n10002), .B2(n8792), .A(n7288), .ZN(n7289) );
  OAI21_X1 U8998 ( .B1(n7290), .B2(n8788), .A(n7289), .ZN(P2_U3287) );
  XOR2_X1 U8999 ( .A(n7291), .B(n8216), .Z(n9855) );
  INV_X1 U9000 ( .A(n8216), .ZN(n7292) );
  XNOR2_X1 U9001 ( .A(n8110), .B(n7292), .ZN(n7293) );
  AND2_X1 U9002 ( .A1(n7293), .A2(n9808), .ZN(n9853) );
  AOI22_X1 U9003 ( .A1(n9822), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7294), .B2(
        n9787), .ZN(n7299) );
  NAND2_X1 U9004 ( .A1(n7295), .A2(n9847), .ZN(n7296) );
  NAND2_X1 U9005 ( .A1(n7296), .A2(n9794), .ZN(n7297) );
  NOR2_X1 U9006 ( .A1(n9776), .A2(n7297), .ZN(n9852) );
  NAND2_X1 U9007 ( .A1(n9852), .A2(n9755), .ZN(n7298) );
  OAI211_X1 U9008 ( .C1(n7300), .C2(n9337), .A(n7299), .B(n7298), .ZN(n7302)
         );
  OAI22_X1 U9009 ( .A1(n9324), .A2(n9849), .B1(n9848), .B2(n9355), .ZN(n7301)
         );
  AOI211_X1 U9010 ( .C1(n9853), .C2(n9816), .A(n7302), .B(n7301), .ZN(n7303)
         );
  OAI21_X1 U9011 ( .B1(n9818), .B2(n9855), .A(n7303), .ZN(P1_U3287) );
  INV_X1 U9012 ( .A(n7304), .ZN(n7311) );
  OAI21_X1 U9013 ( .B1(n6914), .B2(n7306), .A(n7305), .ZN(n7307) );
  NAND3_X1 U9014 ( .A1(n8517), .A2(n7308), .A3(n7307), .ZN(n7310) );
  NAND2_X1 U9015 ( .A1(n8492), .A2(n9950), .ZN(n7309) );
  OAI211_X1 U9016 ( .C1(n7311), .C2(n7222), .A(n7310), .B(n7309), .ZN(n7312)
         );
  AOI21_X1 U9017 ( .B1(n8511), .B2(n4483), .A(n7312), .ZN(n7313) );
  INV_X1 U9018 ( .A(n7313), .ZN(P2_U3234) );
  INV_X1 U9019 ( .A(n7314), .ZN(n7315) );
  OAI222_X1 U9020 ( .A1(n9541), .A2(n10432), .B1(n9548), .B2(n7315), .C1(
        P1_U3084), .C2(n9814), .ZN(P1_U3334) );
  OAI222_X1 U9021 ( .A1(n7789), .A2(n7316), .B1(n8944), .B2(n7315), .C1(n7892), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U9022 ( .A1(n7323), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7318) );
  NAND2_X1 U9023 ( .A1(n7318), .A2(n7317), .ZN(n7320) );
  INV_X1 U9024 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7570) );
  AOI22_X1 U9025 ( .A1(n7426), .A2(n7570), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7321), .ZN(n7319) );
  NOR2_X1 U9026 ( .A1(n7320), .A2(n7319), .ZN(n7421) );
  AOI21_X1 U9027 ( .B1(n7320), .B2(n7319), .A(n7421), .ZN(n7332) );
  INV_X1 U9028 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9583) );
  AOI22_X1 U9029 ( .A1(n7426), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9583), .B2(
        n7321), .ZN(n7325) );
  OAI21_X1 U9030 ( .B1(n7323), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7322), .ZN(
        n7324) );
  OAI21_X1 U9031 ( .B1(n7325), .B2(n7324), .A(n7425), .ZN(n7326) );
  NAND2_X1 U9032 ( .A1(n7326), .A2(n9929), .ZN(n7331) );
  INV_X1 U9033 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7328) );
  OAI22_X1 U9034 ( .A1(n8617), .A2(n7328), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7327), .ZN(n7329) );
  AOI21_X1 U9035 ( .B1(n8611), .B2(n7426), .A(n7329), .ZN(n7330) );
  OAI211_X1 U9036 ( .C1(n7332), .C2(n9935), .A(n7331), .B(n7330), .ZN(P2_U3258) );
  INV_X1 U9037 ( .A(n8212), .ZN(n7333) );
  OAI21_X1 U9038 ( .B1(n9760), .B2(n7333), .A(n8211), .ZN(n7334) );
  XNOR2_X1 U9039 ( .A(n7334), .B(n4971), .ZN(n7335) );
  NAND2_X1 U9040 ( .A1(n7335), .A2(n9808), .ZN(n7368) );
  OAI21_X1 U9041 ( .B1(n7338), .B2(n7337), .A(n7336), .ZN(n7370) );
  NAND2_X1 U9042 ( .A1(n7370), .A2(n9350), .ZN(n7347) );
  OAI211_X1 U9043 ( .C1(n9752), .C2(n7371), .A(n9794), .B(n9616), .ZN(n7366)
         );
  INV_X1 U9044 ( .A(n7366), .ZN(n7345) );
  INV_X1 U9045 ( .A(n7496), .ZN(n7339) );
  OAI22_X1 U9046 ( .A1(n9816), .A2(n7340), .B1(n7339), .B2(n9800), .ZN(n7341)
         );
  AOI21_X1 U9047 ( .B1(n9322), .B2(n9090), .A(n7341), .ZN(n7343) );
  NAND2_X1 U9048 ( .A1(n9352), .A2(n9092), .ZN(n7342) );
  OAI211_X1 U9049 ( .C1(n7371), .C2(n9337), .A(n7343), .B(n7342), .ZN(n7344)
         );
  AOI21_X1 U9050 ( .B1(n7345), .B2(n9755), .A(n7344), .ZN(n7346) );
  OAI211_X1 U9051 ( .C1(n9822), .C2(n7368), .A(n7347), .B(n7346), .ZN(P1_U3281) );
  XNOR2_X1 U9052 ( .A(n7348), .B(n7275), .ZN(n9996) );
  NOR2_X1 U9053 ( .A1(n7349), .A2(n9992), .ZN(n7350) );
  OR2_X1 U9054 ( .A1(n7351), .A2(n7350), .ZN(n9993) );
  AOI22_X1 U9055 ( .A1(n8620), .A2(n7353), .B1(n8800), .B2(n7352), .ZN(n7354)
         );
  OAI21_X1 U9056 ( .B1(n8629), .B2(n9993), .A(n7354), .ZN(n7364) );
  NAND2_X1 U9057 ( .A1(n7356), .A2(n7355), .ZN(n7357) );
  NAND2_X1 U9058 ( .A1(n7277), .A2(n7357), .ZN(n7360) );
  OAI22_X1 U9059 ( .A1(n7358), .A2(n8764), .B1(n7381), .B2(n8762), .ZN(n7359)
         );
  AOI21_X1 U9060 ( .B1(n7360), .B2(n8804), .A(n7359), .ZN(n7362) );
  NAND2_X1 U9061 ( .A1(n9996), .A2(n8786), .ZN(n7361) );
  NAND2_X1 U9062 ( .A1(n7362), .A2(n7361), .ZN(n9994) );
  MUX2_X1 U9063 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9994), .S(n8696), .Z(n7363)
         );
  AOI211_X1 U9064 ( .C1(n8792), .C2(n9996), .A(n7364), .B(n7363), .ZN(n7365)
         );
  INV_X1 U9065 ( .A(n7365), .ZN(P2_U3288) );
  AOI22_X1 U9066 ( .A1(n9866), .A2(n9092), .B1(n9090), .B2(n9863), .ZN(n7367)
         );
  NAND3_X1 U9067 ( .A1(n7368), .A2(n7367), .A3(n7366), .ZN(n7369) );
  AOI21_X1 U9068 ( .B1(n7370), .B2(n9885), .A(n7369), .ZN(n7376) );
  OAI22_X1 U9069 ( .A1(n7371), .A2(n9532), .B1(n9911), .B2(n5412), .ZN(n7372)
         );
  INV_X1 U9070 ( .A(n7372), .ZN(n7373) );
  OAI21_X1 U9071 ( .B1(n7376), .B2(n9909), .A(n7373), .ZN(P1_U3484) );
  NAND2_X1 U9072 ( .A1(n9928), .A2(n9892), .ZN(n9478) );
  INV_X1 U9073 ( .A(n9478), .ZN(n7374) );
  AOI22_X1 U9074 ( .A1(n7501), .A2(n7374), .B1(n9925), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7375) );
  OAI21_X1 U9075 ( .B1(n7376), .B2(n9925), .A(n7375), .ZN(P1_U3533) );
  INV_X1 U9076 ( .A(n7381), .ZN(n8544) );
  OR2_X1 U9077 ( .A1(n7377), .A2(n8544), .ZN(n7378) );
  NAND2_X1 U9078 ( .A1(n10004), .A2(n7794), .ZN(n7903) );
  NAND2_X1 U9079 ( .A1(n7908), .A2(n7903), .ZN(n7878) );
  XNOR2_X1 U9080 ( .A(n7486), .B(n7485), .ZN(n7385) );
  NAND2_X1 U9081 ( .A1(n7380), .A2(n7956), .ZN(n7477) );
  XNOR2_X1 U9082 ( .A(n7477), .B(n7485), .ZN(n7383) );
  OAI22_X1 U9083 ( .A1(n7478), .A2(n8762), .B1(n7381), .B2(n8764), .ZN(n7382)
         );
  AOI21_X1 U9084 ( .B1(n7383), .B2(n8804), .A(n7382), .ZN(n7384) );
  OAI21_X1 U9085 ( .B1(n7385), .B2(n7568), .A(n7384), .ZN(n10007) );
  INV_X1 U9086 ( .A(n10007), .ZN(n7393) );
  INV_X1 U9087 ( .A(n7385), .ZN(n10009) );
  NAND2_X1 U9088 ( .A1(n7386), .A2(n10004), .ZN(n7387) );
  NAND2_X1 U9089 ( .A1(n7521), .A2(n7387), .ZN(n10006) );
  AOI22_X1 U9090 ( .A1(n8788), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7388), .B2(
        n8800), .ZN(n7390) );
  NAND2_X1 U9091 ( .A1(n8620), .A2(n10004), .ZN(n7389) );
  OAI211_X1 U9092 ( .C1(n8629), .C2(n10006), .A(n7390), .B(n7389), .ZN(n7391)
         );
  AOI21_X1 U9093 ( .B1(n10009), .B2(n8792), .A(n7391), .ZN(n7392) );
  OAI21_X1 U9094 ( .B1(n7393), .B2(n8788), .A(n7392), .ZN(P2_U3286) );
  INV_X1 U9095 ( .A(n7394), .ZN(n7395) );
  AOI21_X1 U9096 ( .B1(n8218), .B2(n7396), .A(n7395), .ZN(n9881) );
  NAND2_X1 U9097 ( .A1(n9816), .A2(n9808), .ZN(n9367) );
  XNOR2_X1 U9098 ( .A(n7397), .B(n8218), .ZN(n9884) );
  NAND2_X1 U9099 ( .A1(n9884), .A2(n9350), .ZN(n7408) );
  INV_X1 U9100 ( .A(n7398), .ZN(n7399) );
  AOI211_X1 U9101 ( .C1(n9879), .C2(n7400), .A(n9615), .B(n7399), .ZN(n9877)
         );
  INV_X1 U9102 ( .A(n9879), .ZN(n7405) );
  AOI22_X1 U9103 ( .A1(n9822), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7401), .B2(
        n9787), .ZN(n7402) );
  OAI21_X1 U9104 ( .B1(n9324), .B2(n9876), .A(n7402), .ZN(n7403) );
  AOI21_X1 U9105 ( .B1(n9322), .B2(n9093), .A(n7403), .ZN(n7404) );
  OAI21_X1 U9106 ( .B1(n7405), .B2(n9337), .A(n7404), .ZN(n7406) );
  AOI21_X1 U9107 ( .B1(n9877), .B2(n9755), .A(n7406), .ZN(n7407) );
  OAI211_X1 U9108 ( .C1(n9881), .C2(n9367), .A(n7408), .B(n7407), .ZN(P1_U3284) );
  NAND2_X1 U9109 ( .A1(n7410), .A2(n7409), .ZN(n7411) );
  XOR2_X1 U9110 ( .A(n7412), .B(n7411), .Z(n7420) );
  NOR2_X1 U9111 ( .A1(n7413), .A2(n9067), .ZN(n7417) );
  NAND2_X1 U9112 ( .A1(n9074), .A2(n9864), .ZN(n7415) );
  OAI211_X1 U9113 ( .C1(n9079), .C2(n9889), .A(n7415), .B(n7414), .ZN(n7416)
         );
  AOI211_X1 U9114 ( .C1(n7418), .C2(n9076), .A(n7417), .B(n7416), .ZN(n7419)
         );
  OAI21_X1 U9115 ( .B1(n7420), .B2(n9085), .A(n7419), .ZN(P1_U3219) );
  NOR2_X1 U9116 ( .A1(n7426), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7422) );
  NOR2_X1 U9117 ( .A1(n7422), .A2(n7421), .ZN(n7424) );
  INV_X1 U9118 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7643) );
  AOI22_X1 U9119 ( .A1(n7649), .A2(n7643), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7644), .ZN(n7423) );
  NOR2_X1 U9120 ( .A1(n7424), .A2(n7423), .ZN(n7642) );
  AOI21_X1 U9121 ( .B1(n7424), .B2(n7423), .A(n7642), .ZN(n7434) );
  INV_X1 U9122 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9575) );
  AOI22_X1 U9123 ( .A1(n7649), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9575), .B2(
        n7644), .ZN(n7428) );
  OAI21_X1 U9124 ( .B1(n7428), .B2(n7427), .A(n7648), .ZN(n7429) );
  NAND2_X1 U9125 ( .A1(n7429), .A2(n9929), .ZN(n7433) );
  INV_X1 U9126 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7430) );
  NAND2_X1 U9127 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7607) );
  OAI21_X1 U9128 ( .B1(n8617), .B2(n7430), .A(n7607), .ZN(n7431) );
  AOI21_X1 U9129 ( .B1(n8611), .B2(n7649), .A(n7431), .ZN(n7432) );
  OAI211_X1 U9130 ( .C1(n7434), .C2(n9935), .A(n7433), .B(n7432), .ZN(P2_U3259) );
  OAI21_X1 U9131 ( .B1(n7437), .B2(n7436), .A(n7435), .ZN(n7442) );
  NOR2_X1 U9132 ( .A1(n9903), .A2(n9067), .ZN(n7441) );
  AND2_X1 U9133 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9706) );
  AOI21_X1 U9134 ( .B1(n9074), .B2(n9093), .A(n9706), .ZN(n7439) );
  NAND2_X1 U9135 ( .A1(n9076), .A2(n9756), .ZN(n7438) );
  OAI211_X1 U9136 ( .C1(n9762), .C2(n9079), .A(n7439), .B(n7438), .ZN(n7440)
         );
  AOI211_X1 U9137 ( .C1(n7442), .C2(n9056), .A(n7441), .B(n7440), .ZN(n7443)
         );
  INV_X1 U9138 ( .A(n7443), .ZN(P1_U3229) );
  INV_X1 U9139 ( .A(n7444), .ZN(n7447) );
  OAI222_X1 U9140 ( .A1(n7446), .A2(P1_U3084), .B1(n9548), .B2(n7447), .C1(
        n7445), .C2(n9541), .ZN(P1_U3333) );
  OAI222_X1 U9141 ( .A1(n7789), .A2(n7448), .B1(P2_U3152), .B2(n8061), .C1(
        n8944), .C2(n7447), .ZN(P2_U3338) );
  INV_X1 U9142 ( .A(n7685), .ZN(n7456) );
  NAND2_X1 U9143 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8955) );
  INV_X1 U9144 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7449) );
  MUX2_X1 U9145 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7449), .S(n7685), .Z(n7453)
         );
  OAI21_X1 U9146 ( .B1(n7451), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7450), .ZN(
        n7452) );
  NAND2_X1 U9147 ( .A1(n7452), .A2(n7453), .ZN(n7684) );
  OAI21_X1 U9148 ( .B1(n7453), .B2(n7452), .A(n7684), .ZN(n7454) );
  NAND2_X1 U9149 ( .A1(n9744), .A2(n7454), .ZN(n7455) );
  OAI211_X1 U9150 ( .C1(n9739), .C2(n7456), .A(n8955), .B(n7455), .ZN(n7465)
         );
  INV_X1 U9151 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U9152 ( .A1(n7459), .A2(n7458), .ZN(n7460) );
  NOR2_X1 U9153 ( .A1(n7460), .A2(n7685), .ZN(n7461) );
  NOR2_X1 U9154 ( .A1(n7462), .A2(n7463), .ZN(n7678) );
  AOI211_X1 U9155 ( .C1(n7463), .C2(n7462), .A(n7678), .B(n9715), .ZN(n7464)
         );
  AOI211_X1 U9156 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9134), .A(n7465), .B(
        n7464), .ZN(n7466) );
  INV_X1 U9157 ( .A(n7466), .ZN(P1_U3255) );
  INV_X1 U9158 ( .A(n7558), .ZN(n10023) );
  OAI21_X1 U9159 ( .B1(n7469), .B2(n7468), .A(n7467), .ZN(n7470) );
  NAND2_X1 U9160 ( .A1(n7470), .A2(n8517), .ZN(n7474) );
  OAI22_X1 U9161 ( .A1(n7478), .A2(n8500), .B1(n8499), .B2(n7581), .ZN(n7471)
         );
  AOI211_X1 U9162 ( .C1(n7524), .C2(n8526), .A(n7472), .B(n7471), .ZN(n7473)
         );
  OAI211_X1 U9163 ( .C1(n10023), .C2(n8529), .A(n7474), .B(n7473), .ZN(
        P2_U3226) );
  INV_X1 U9164 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7476) );
  INV_X1 U9165 ( .A(n7475), .ZN(n7504) );
  OAI222_X1 U9166 ( .A1(n9541), .A2(n7476), .B1(n9548), .B2(n7504), .C1(n8243), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  NAND2_X1 U9167 ( .A1(n10012), .A2(n7478), .ZN(n7959) );
  NAND2_X1 U9168 ( .A1(n4545), .A2(n7959), .ZN(n7879) );
  XNOR2_X1 U9169 ( .A(n7514), .B(n7879), .ZN(n7480) );
  OAI22_X1 U9170 ( .A1(n7794), .A2(n8764), .B1(n7793), .B2(n8762), .ZN(n7479)
         );
  AOI21_X1 U9171 ( .B1(n7480), .B2(n8804), .A(n7479), .ZN(n10017) );
  XNOR2_X1 U9172 ( .A(n7521), .B(n7483), .ZN(n10015) );
  AOI22_X1 U9173 ( .A1(n8788), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7481), .B2(
        n8800), .ZN(n7482) );
  OAI21_X1 U9174 ( .B1(n7483), .B2(n8823), .A(n7482), .ZN(n7489) );
  NAND2_X1 U9175 ( .A1(n10004), .A2(n8543), .ZN(n7484) );
  OAI21_X1 U9176 ( .B1(n7487), .B2(n7879), .A(n7519), .ZN(n10018) );
  NOR2_X1 U9177 ( .A1(n10018), .A2(n8818), .ZN(n7488) );
  AOI211_X1 U9178 ( .C1(n8816), .C2(n10015), .A(n7489), .B(n7488), .ZN(n7490)
         );
  OAI21_X1 U9179 ( .B1(n8788), .B2(n10017), .A(n7490), .ZN(P2_U3285) );
  NAND2_X1 U9180 ( .A1(n7492), .A2(n7491), .ZN(n7493) );
  XNOR2_X1 U9181 ( .A(n7494), .B(n7493), .ZN(n7503) );
  NOR2_X1 U9182 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7495), .ZN(n9724) );
  AOI21_X1 U9183 ( .B1(n9074), .B2(n9092), .A(n9724), .ZN(n7498) );
  NAND2_X1 U9184 ( .A1(n9076), .A2(n7496), .ZN(n7497) );
  OAI211_X1 U9185 ( .C1(n7499), .C2(n9079), .A(n7498), .B(n7497), .ZN(n7500)
         );
  AOI21_X1 U9186 ( .B1(n9082), .B2(n7501), .A(n7500), .ZN(n7502) );
  OAI21_X1 U9187 ( .B1(n7503), .B2(n9085), .A(n7502), .ZN(P1_U3215) );
  INV_X1 U9188 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7506) );
  OAI222_X1 U9189 ( .A1(n7789), .A2(n7506), .B1(P2_U3152), .B2(n7505), .C1(
        n8944), .C2(n7504), .ZN(P2_U3337) );
  XNOR2_X1 U9190 ( .A(n7508), .B(n7507), .ZN(n7513) );
  INV_X1 U9191 ( .A(n7509), .ZN(n7569) );
  OAI22_X1 U9192 ( .A1(n8498), .A2(n7569), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7327), .ZN(n7511) );
  OAI22_X1 U9193 ( .A1(n7793), .A2(n8500), .B1(n8499), .B2(n7709), .ZN(n7510)
         );
  AOI211_X1 U9194 ( .C1(n7586), .C2(n8503), .A(n7511), .B(n7510), .ZN(n7512)
         );
  OAI21_X1 U9195 ( .B1(n7513), .B2(n8505), .A(n7512), .ZN(P2_U3236) );
  OR2_X1 U9196 ( .A1(n7558), .A2(n7793), .ZN(n7968) );
  AND2_X1 U9197 ( .A1(n7558), .A2(n7793), .ZN(n7961) );
  INV_X1 U9198 ( .A(n7961), .ZN(n7967) );
  XNOR2_X1 U9199 ( .A(n7563), .B(n7881), .ZN(n7515) );
  NAND2_X1 U9200 ( .A1(n7515), .A2(n8804), .ZN(n7517) );
  INV_X1 U9201 ( .A(n7581), .ZN(n8540) );
  AOI22_X1 U9202 ( .A1(n8540), .A2(n8810), .B1(n8809), .B2(n8542), .ZN(n7516)
         );
  NAND2_X1 U9203 ( .A1(n7517), .A2(n7516), .ZN(n10026) );
  INV_X1 U9204 ( .A(n10026), .ZN(n7529) );
  NAND2_X1 U9205 ( .A1(n10012), .A2(n8542), .ZN(n7518) );
  INV_X1 U9206 ( .A(n7881), .ZN(n7520) );
  OAI21_X1 U9207 ( .B1(n5078), .B2(n7520), .A(n7560), .ZN(n10028) );
  AND2_X1 U9208 ( .A1(n7523), .A2(n10023), .ZN(n7571) );
  INV_X1 U9209 ( .A(n7571), .ZN(n7522) );
  OAI21_X1 U9210 ( .B1(n10023), .B2(n7523), .A(n7522), .ZN(n10025) );
  AOI22_X1 U9211 ( .A1(n8788), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7524), .B2(
        n8800), .ZN(n7526) );
  NAND2_X1 U9212 ( .A1(n8620), .A2(n7558), .ZN(n7525) );
  OAI211_X1 U9213 ( .C1(n10025), .C2(n8629), .A(n7526), .B(n7525), .ZN(n7527)
         );
  AOI21_X1 U9214 ( .B1(n10028), .B2(n8826), .A(n7527), .ZN(n7528) );
  OAI21_X1 U9215 ( .B1(n7529), .B2(n8788), .A(n7528), .ZN(P2_U3284) );
  NAND2_X1 U9216 ( .A1(n7530), .A2(n8227), .ZN(n7531) );
  XNOR2_X1 U9217 ( .A(n7533), .B(n8227), .ZN(n7535) );
  AOI22_X1 U9218 ( .A1(n9866), .A2(n9090), .B1(n9089), .B2(n9863), .ZN(n7534)
         );
  OAI21_X1 U9219 ( .B1(n7535), .B2(n9882), .A(n7534), .ZN(n7536) );
  AOI21_X1 U9220 ( .B1(n9647), .B2(n9900), .A(n7536), .ZN(n9649) );
  AOI21_X1 U9221 ( .B1(n9617), .B2(n7618), .A(n9615), .ZN(n7537) );
  NAND2_X1 U9222 ( .A1(n7537), .A2(n9593), .ZN(n9644) );
  AOI22_X1 U9223 ( .A1(n9822), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7625), .B2(
        n9787), .ZN(n7539) );
  NAND2_X1 U9224 ( .A1(n7618), .A2(n9770), .ZN(n7538) );
  OAI211_X1 U9225 ( .C1(n9644), .C2(n9361), .A(n7539), .B(n7538), .ZN(n7540)
         );
  AOI21_X1 U9226 ( .B1(n9647), .B2(n9350), .A(n7540), .ZN(n7541) );
  OAI21_X1 U9227 ( .B1(n9649), .B2(n9822), .A(n7541), .ZN(P1_U3279) );
  INV_X1 U9228 ( .A(n9634), .ZN(n9651) );
  AOI21_X1 U9229 ( .B1(n7543), .B2(n7542), .A(n9085), .ZN(n7545) );
  NAND2_X1 U9230 ( .A1(n7545), .A2(n7544), .ZN(n7550) );
  AOI21_X1 U9231 ( .B1(n9074), .B2(n9091), .A(n7546), .ZN(n7547) );
  OAI21_X1 U9232 ( .B1(n9627), .B2(n9079), .A(n7547), .ZN(n7548) );
  AOI21_X1 U9233 ( .B1(n9620), .B2(n9076), .A(n7548), .ZN(n7549) );
  OAI211_X1 U9234 ( .C1(n9651), .C2(n9067), .A(n7550), .B(n7549), .ZN(P1_U3234) );
  INV_X1 U9235 ( .A(n7551), .ZN(n7787) );
  OAI222_X1 U9236 ( .A1(n9541), .A2(n10392), .B1(n9548), .B2(n7787), .C1(
        P1_U3084), .C2(n8386), .ZN(P1_U3331) );
  INV_X1 U9237 ( .A(n7552), .ZN(n7557) );
  AOI21_X1 U9238 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8947), .A(n7553), .ZN(
        n7554) );
  OAI21_X1 U9239 ( .B1(n7557), .B2(n8944), .A(n7554), .ZN(P2_U3335) );
  AND2_X1 U9240 ( .A1(n7555), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8387) );
  AOI21_X1 U9241 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9545), .A(n8387), .ZN(
        n7556) );
  OAI21_X1 U9242 ( .B1(n7557), .B2(n9548), .A(n7556), .ZN(P1_U3330) );
  INV_X1 U9243 ( .A(n7793), .ZN(n8541) );
  OR2_X1 U9244 ( .A1(n7558), .A2(n8541), .ZN(n7559) );
  OR2_X1 U9245 ( .A1(n7586), .A2(n7581), .ZN(n7973) );
  NAND2_X1 U9246 ( .A1(n7586), .A2(n7581), .ZN(n7972) );
  NAND2_X1 U9247 ( .A1(n7561), .A2(n7970), .ZN(n7562) );
  NAND2_X1 U9248 ( .A1(n7588), .A2(n7562), .ZN(n9577) );
  INV_X1 U9249 ( .A(n8792), .ZN(n7577) );
  OAI21_X1 U9250 ( .B1(n7564), .B2(n7970), .A(n7580), .ZN(n7566) );
  OAI22_X1 U9251 ( .A1(n7793), .A2(n8764), .B1(n7709), .B2(n8762), .ZN(n7565)
         );
  AOI21_X1 U9252 ( .B1(n7566), .B2(n8804), .A(n7565), .ZN(n7567) );
  OAI21_X1 U9253 ( .B1(n7568), .B2(n9577), .A(n7567), .ZN(n9580) );
  NAND2_X1 U9254 ( .A1(n9580), .A2(n8696), .ZN(n7576) );
  OAI22_X1 U9255 ( .A1(n8696), .A2(n7570), .B1(n7569), .B2(n8821), .ZN(n7574)
         );
  INV_X1 U9256 ( .A(n7586), .ZN(n9578) );
  OR2_X1 U9257 ( .A1(n7571), .A2(n9578), .ZN(n7572) );
  NAND2_X1 U9258 ( .A1(n7590), .A2(n7572), .ZN(n9579) );
  NOR2_X1 U9259 ( .A1(n9579), .A2(n8629), .ZN(n7573) );
  AOI211_X1 U9260 ( .C1(n8620), .C2(n7586), .A(n7574), .B(n7573), .ZN(n7575)
         );
  OAI211_X1 U9261 ( .C1(n9577), .C2(n7577), .A(n7576), .B(n7575), .ZN(P2_U3283) );
  NAND2_X1 U9262 ( .A1(n7628), .A2(n7709), .ZN(n7978) );
  NAND2_X1 U9263 ( .A1(n7977), .A2(n7978), .ZN(n7883) );
  INV_X1 U9264 ( .A(n7972), .ZN(n7578) );
  NOR2_X1 U9265 ( .A1(n7883), .A2(n7578), .ZN(n7579) );
  NAND2_X1 U9266 ( .A1(n7631), .A2(n8804), .ZN(n7585) );
  INV_X1 U9267 ( .A(n7883), .ZN(n7976) );
  AOI21_X1 U9268 ( .B1(n7580), .B2(n7972), .A(n7976), .ZN(n7584) );
  OR2_X1 U9269 ( .A1(n7743), .A2(n8762), .ZN(n7583) );
  OR2_X1 U9270 ( .A1(n7581), .A2(n8764), .ZN(n7582) );
  AND2_X1 U9271 ( .A1(n7583), .A2(n7582), .ZN(n7609) );
  OAI21_X1 U9272 ( .B1(n7585), .B2(n7584), .A(n7609), .ZN(n9572) );
  AOI21_X1 U9273 ( .B1(n7606), .B2(n8800), .A(n9572), .ZN(n7595) );
  NAND2_X1 U9274 ( .A1(n7586), .A2(n8540), .ZN(n7587) );
  OAI21_X1 U9275 ( .B1(n7589), .B2(n7883), .A(n7630), .ZN(n9574) );
  INV_X1 U9276 ( .A(n7590), .ZN(n7591) );
  INV_X1 U9277 ( .A(n7628), .ZN(n9570) );
  OAI21_X1 U9278 ( .B1(n7591), .B2(n9570), .A(n7635), .ZN(n9571) );
  AOI22_X1 U9279 ( .A1(n7628), .A2(n8620), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8788), .ZN(n7592) );
  OAI21_X1 U9280 ( .B1(n9571), .B2(n8629), .A(n7592), .ZN(n7593) );
  AOI21_X1 U9281 ( .B1(n9574), .B2(n8826), .A(n7593), .ZN(n7594) );
  OAI21_X1 U9282 ( .B1(n7595), .B2(n8788), .A(n7594), .ZN(P2_U3282) );
  XOR2_X1 U9283 ( .A(n8229), .B(n7596), .Z(n7597) );
  AOI22_X1 U9284 ( .A1(n7597), .A2(n9808), .B1(n9863), .B2(n9458), .ZN(n9473)
         );
  XOR2_X1 U9285 ( .A(n8229), .B(n7598), .Z(n9476) );
  NAND2_X1 U9286 ( .A1(n9476), .A2(n9350), .ZN(n7603) );
  AOI22_X1 U9287 ( .A1(n9822), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8957), .B2(
        n9787), .ZN(n7599) );
  OAI21_X1 U9288 ( .B1(n9324), .B2(n9474), .A(n7599), .ZN(n7601) );
  OAI211_X1 U9289 ( .C1(n9533), .C2(n9592), .A(n7661), .B(n9794), .ZN(n9472)
         );
  NOR2_X1 U9290 ( .A1(n9472), .A2(n9361), .ZN(n7600) );
  AOI211_X1 U9291 ( .C1(n9770), .C2(n8962), .A(n7601), .B(n7600), .ZN(n7602)
         );
  OAI211_X1 U9292 ( .C1(n9822), .C2(n9473), .A(n7603), .B(n7602), .ZN(P1_U3277) );
  AOI21_X1 U9293 ( .B1(n7605), .B2(n7604), .A(n4560), .ZN(n7612) );
  NAND2_X1 U9294 ( .A1(n8526), .A2(n7606), .ZN(n7608) );
  OAI211_X1 U9295 ( .C1(n8524), .C2(n7609), .A(n7608), .B(n7607), .ZN(n7610)
         );
  AOI21_X1 U9296 ( .B1(n7628), .B2(n8492), .A(n7610), .ZN(n7611) );
  OAI21_X1 U9297 ( .B1(n7612), .B2(n8505), .A(n7611), .ZN(P2_U3217) );
  INV_X1 U9298 ( .A(n7613), .ZN(n7616) );
  INV_X1 U9299 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7614) );
  OAI222_X1 U9300 ( .A1(P2_U3152), .A2(n7615), .B1(n8944), .B2(n7616), .C1(
        n7614), .C2(n7789), .ZN(P2_U3334) );
  INV_X1 U9301 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10372) );
  OAI222_X1 U9302 ( .A1(n7617), .A2(P1_U3084), .B1(n9548), .B2(n7616), .C1(
        n10372), .C2(n9541), .ZN(P1_U3329) );
  INV_X1 U9303 ( .A(n7618), .ZN(n9645) );
  OAI21_X1 U9304 ( .B1(n7621), .B2(n7620), .A(n7619), .ZN(n7622) );
  NAND2_X1 U9305 ( .A1(n7622), .A2(n9056), .ZN(n7627) );
  AOI22_X1 U9306 ( .A1(n9074), .A2(n9090), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n7623) );
  OAI21_X1 U9307 ( .B1(n9474), .B2(n9079), .A(n7623), .ZN(n7624) );
  AOI21_X1 U9308 ( .B1(n7625), .B2(n9076), .A(n7624), .ZN(n7626) );
  OAI211_X1 U9309 ( .C1(n9645), .C2(n9067), .A(n7627), .B(n7626), .ZN(P1_U3222) );
  INV_X1 U9310 ( .A(n7709), .ZN(n8539) );
  OR2_X1 U9311 ( .A1(n7628), .A2(n8539), .ZN(n7629) );
  NAND2_X1 U9312 ( .A1(n7630), .A2(n7629), .ZN(n7723) );
  NAND2_X1 U9313 ( .A1(n7721), .A2(n7743), .ZN(n7982) );
  XNOR2_X1 U9314 ( .A(n7723), .B(n7884), .ZN(n9568) );
  INV_X1 U9315 ( .A(n9568), .ZN(n7641) );
  NAND2_X1 U9316 ( .A1(n7631), .A2(n7977), .ZN(n7632) );
  NAND2_X1 U9317 ( .A1(n7632), .A2(n7980), .ZN(n7726) );
  OAI211_X1 U9318 ( .C1(n7632), .C2(n7980), .A(n7726), .B(n8804), .ZN(n7634)
         );
  AOI22_X1 U9319 ( .A1(n8539), .A2(n8809), .B1(n8810), .B2(n8537), .ZN(n7633)
         );
  NAND2_X1 U9320 ( .A1(n7634), .A2(n7633), .ZN(n9566) );
  INV_X1 U9321 ( .A(n7635), .ZN(n7636) );
  INV_X1 U9322 ( .A(n7721), .ZN(n9564) );
  OAI21_X1 U9323 ( .B1(n7636), .B2(n9564), .A(n7771), .ZN(n9565) );
  AOI22_X1 U9324 ( .A1(n8788), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7712), .B2(
        n8800), .ZN(n7638) );
  NAND2_X1 U9325 ( .A1(n7721), .A2(n8620), .ZN(n7637) );
  OAI211_X1 U9326 ( .C1(n9565), .C2(n8629), .A(n7638), .B(n7637), .ZN(n7639)
         );
  AOI21_X1 U9327 ( .B1(n9566), .B2(n8696), .A(n7639), .ZN(n7640) );
  OAI21_X1 U9328 ( .B1(n7641), .B2(n8818), .A(n7640), .ZN(P2_U3281) );
  AOI21_X1 U9329 ( .B1(n7644), .B2(n7643), .A(n7642), .ZN(n8560) );
  XNOR2_X1 U9330 ( .A(n8560), .B(n8561), .ZN(n7645) );
  NOR2_X1 U9331 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7645), .ZN(n8562) );
  AOI21_X1 U9332 ( .B1(n7645), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8562), .ZN(
        n7654) );
  INV_X1 U9333 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7647) );
  INV_X1 U9334 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10463) );
  NOR2_X1 U9335 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10463), .ZN(n7711) );
  INV_X1 U9336 ( .A(n7711), .ZN(n7646) );
  OAI21_X1 U9337 ( .B1(n8617), .B2(n7647), .A(n7646), .ZN(n7652) );
  XNOR2_X1 U9338 ( .A(n8552), .B(n8553), .ZN(n7650) );
  INV_X1 U9339 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9569) );
  NOR2_X1 U9340 ( .A1(n9569), .A2(n7650), .ZN(n8554) );
  AOI211_X1 U9341 ( .C1(n7650), .C2(n9569), .A(n8554), .B(n9934), .ZN(n7651)
         );
  AOI211_X1 U9342 ( .C1(n8611), .C2(n8561), .A(n7652), .B(n7651), .ZN(n7653)
         );
  OAI21_X1 U9343 ( .B1(n7654), .B2(n9935), .A(n7653), .ZN(P2_U3260) );
  INV_X1 U9344 ( .A(n8265), .ZN(n8278) );
  XNOR2_X1 U9345 ( .A(n7655), .B(n8230), .ZN(n7656) );
  NAND2_X1 U9346 ( .A1(n7656), .A2(n9808), .ZN(n7658) );
  AOI22_X1 U9347 ( .A1(n9341), .A2(n9863), .B1(n9866), .B2(n9605), .ZN(n7657)
         );
  NAND2_X1 U9348 ( .A1(n7658), .A2(n7657), .ZN(n9467) );
  INV_X1 U9349 ( .A(n9467), .ZN(n7666) );
  XNOR2_X1 U9350 ( .A(n7659), .B(n8230), .ZN(n9469) );
  NAND2_X1 U9351 ( .A1(n9469), .A2(n9350), .ZN(n7665) );
  INV_X1 U9352 ( .A(n9357), .ZN(n7660) );
  AOI211_X1 U9353 ( .C1(n9083), .C2(n7661), .A(n9615), .B(n7660), .ZN(n9468)
         );
  AOI22_X1 U9354 ( .A1(n9822), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9075), .B2(
        n9787), .ZN(n7662) );
  OAI21_X1 U9355 ( .B1(n9528), .B2(n9337), .A(n7662), .ZN(n7663) );
  AOI21_X1 U9356 ( .B1(n9468), .B2(n9755), .A(n7663), .ZN(n7664) );
  OAI211_X1 U9357 ( .C1(n9822), .C2(n7666), .A(n7665), .B(n7664), .ZN(P1_U3276) );
  XNOR2_X1 U9358 ( .A(n7668), .B(n7667), .ZN(n7669) );
  XNOR2_X1 U9359 ( .A(n7670), .B(n7669), .ZN(n7677) );
  INV_X1 U9360 ( .A(n7671), .ZN(n7672) );
  AOI21_X1 U9361 ( .B1(n9074), .B2(n9606), .A(n7672), .ZN(n7674) );
  NAND2_X1 U9362 ( .A1(n9076), .A2(n9597), .ZN(n7673) );
  OAI211_X1 U9363 ( .C1(n8135), .C2(n9079), .A(n7674), .B(n7673), .ZN(n7675)
         );
  AOI21_X1 U9364 ( .B1(n9637), .B2(n9082), .A(n7675), .ZN(n7676) );
  OAI21_X1 U9365 ( .B1(n7677), .B2(n9085), .A(n7676), .ZN(P1_U3232) );
  NOR2_X1 U9366 ( .A1(n7679), .A2(n7678), .ZN(n7690) );
  XNOR2_X1 U9367 ( .A(n7697), .B(n7690), .ZN(n7681) );
  INV_X1 U9368 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7680) );
  NOR2_X1 U9369 ( .A1(n7680), .A2(n7681), .ZN(n7691) );
  AOI21_X1 U9370 ( .B1(n7681), .B2(n7680), .A(n7691), .ZN(n7682) );
  NAND2_X1 U9371 ( .A1(n9735), .A2(n7682), .ZN(n7683) );
  NAND2_X1 U9372 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9072) );
  OAI211_X1 U9373 ( .C1(n9739), .C2(n7697), .A(n7683), .B(n9072), .ZN(n7688)
         );
  INV_X1 U9374 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9470) );
  OAI21_X1 U9375 ( .B1(n7685), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7684), .ZN(
        n7696) );
  XNOR2_X1 U9376 ( .A(n7696), .B(n7697), .ZN(n7686) );
  NOR2_X1 U9377 ( .A1(n9470), .A2(n7686), .ZN(n7698) );
  INV_X1 U9378 ( .A(n9744), .ZN(n9720) );
  AOI211_X1 U9379 ( .C1(n9470), .C2(n7686), .A(n7698), .B(n9720), .ZN(n7687)
         );
  AOI211_X1 U9380 ( .C1(n9134), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7688), .B(
        n7687), .ZN(n7689) );
  INV_X1 U9381 ( .A(n7689), .ZN(P1_U3256) );
  NOR2_X1 U9382 ( .A1(n7690), .A2(n7697), .ZN(n7692) );
  NOR2_X1 U9383 ( .A1(n7692), .A2(n7691), .ZN(n7695) );
  NAND2_X1 U9384 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8076), .ZN(n7693) );
  OAI21_X1 U9385 ( .B1(n8076), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7693), .ZN(
        n7694) );
  NOR2_X1 U9386 ( .A1(n7695), .A2(n7694), .ZN(n8071) );
  AOI211_X1 U9387 ( .C1(n7695), .C2(n7694), .A(n8071), .B(n9715), .ZN(n7706)
         );
  NOR2_X1 U9388 ( .A1(n7697), .A2(n7696), .ZN(n7699) );
  NOR2_X1 U9389 ( .A1(n7699), .A2(n7698), .ZN(n7701) );
  XNOR2_X1 U9390 ( .A(n8076), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7700) );
  NOR2_X1 U9391 ( .A1(n7701), .A2(n7700), .ZN(n8075) );
  AOI211_X1 U9392 ( .C1(n7701), .C2(n7700), .A(n8075), .B(n9720), .ZN(n7705)
         );
  NAND2_X1 U9393 ( .A1(n9134), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U9394 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9006) );
  OAI211_X1 U9395 ( .C1(n9739), .C2(n7703), .A(n7702), .B(n9006), .ZN(n7704)
         );
  OR3_X1 U9396 ( .A1(n7706), .A2(n7705), .A3(n7704), .ZN(P1_U3257) );
  XNOR2_X1 U9397 ( .A(n7708), .B(n7707), .ZN(n7715) );
  INV_X1 U9398 ( .A(n8537), .ZN(n7754) );
  OAI22_X1 U9399 ( .A1(n7709), .A2(n8500), .B1(n8499), .B2(n7754), .ZN(n7710)
         );
  AOI211_X1 U9400 ( .C1(n8526), .C2(n7712), .A(n7711), .B(n7710), .ZN(n7714)
         );
  NAND2_X1 U9401 ( .A1(n7721), .A2(n8492), .ZN(n7713) );
  OAI211_X1 U9402 ( .C1(n7715), .C2(n8505), .A(n7714), .B(n7713), .ZN(P2_U3243) );
  INV_X1 U9403 ( .A(n7716), .ZN(n7720) );
  OAI222_X1 U9404 ( .A1(n7789), .A2(n7718), .B1(n8949), .B2(n7720), .C1(
        P2_U3152), .C2(n7717), .ZN(P2_U3333) );
  OAI222_X1 U9405 ( .A1(n9541), .A2(n10184), .B1(n9548), .B2(n7720), .C1(n7719), .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9406 ( .A(n7743), .ZN(n8538) );
  NOR2_X1 U9407 ( .A1(n7721), .A2(n8538), .ZN(n7722) );
  AOI21_X1 U9408 ( .B1(n7723), .B2(n7884), .A(n7722), .ZN(n7724) );
  NAND2_X1 U9409 ( .A1(n7748), .A2(n8537), .ZN(n7987) );
  NAND2_X1 U9410 ( .A1(n8912), .A2(n7754), .ZN(n7986) );
  NAND2_X1 U9411 ( .A1(n7987), .A2(n7986), .ZN(n7902) );
  NAND2_X1 U9412 ( .A1(n7724), .A2(n7902), .ZN(n7765) );
  OR2_X1 U9413 ( .A1(n7724), .A2(n7902), .ZN(n7725) );
  OAI22_X1 U9414 ( .A1(n7781), .A2(n8762), .B1(n7743), .B2(n8764), .ZN(n7731)
         );
  NAND2_X1 U9415 ( .A1(n7726), .A2(n7983), .ZN(n7728) );
  NAND2_X1 U9416 ( .A1(n7728), .A2(n7902), .ZN(n7729) );
  AOI21_X1 U9417 ( .B1(n7761), .B2(n7729), .A(n8759), .ZN(n7730) );
  AOI211_X1 U9418 ( .C1(n8911), .C2(n8786), .A(n7731), .B(n7730), .ZN(n8915)
         );
  XNOR2_X1 U9419 ( .A(n7748), .B(n7771), .ZN(n8913) );
  NAND2_X1 U9420 ( .A1(n8913), .A2(n8816), .ZN(n7736) );
  INV_X1 U9421 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7733) );
  OAI22_X1 U9422 ( .A1(n8696), .A2(n7733), .B1(n7732), .B2(n8821), .ZN(n7734)
         );
  AOI21_X1 U9423 ( .B1(n8912), .B2(n8620), .A(n7734), .ZN(n7735) );
  NAND2_X1 U9424 ( .A1(n7736), .A2(n7735), .ZN(n7737) );
  AOI21_X1 U9425 ( .B1(n8911), .B2(n8792), .A(n7737), .ZN(n7738) );
  OAI21_X1 U9426 ( .B1(n8915), .B2(n8788), .A(n7738), .ZN(P2_U3280) );
  OAI21_X1 U9427 ( .B1(n7741), .B2(n7740), .A(n7739), .ZN(n7742) );
  NAND2_X1 U9428 ( .A1(n7742), .A2(n8517), .ZN(n7747) );
  AND2_X1 U9429 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8559) );
  OAI22_X1 U9430 ( .A1(n7743), .A2(n8500), .B1(n8499), .B2(n7781), .ZN(n7744)
         );
  AOI211_X1 U9431 ( .C1(n7745), .C2(n8526), .A(n8559), .B(n7744), .ZN(n7746)
         );
  OAI211_X1 U9432 ( .C1(n7748), .C2(n8529), .A(n7747), .B(n7746), .ZN(P2_U3228) );
  INV_X1 U9433 ( .A(n7749), .ZN(n7759) );
  AOI22_X1 U9434 ( .A1(n7750), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8947), .ZN(n7751) );
  OAI21_X1 U9435 ( .B1(n7759), .B2(n8944), .A(n7751), .ZN(P2_U3332) );
  XNOR2_X1 U9436 ( .A(n7753), .B(n7752), .ZN(n7758) );
  INV_X1 U9437 ( .A(n8536), .ZN(n7826) );
  OAI22_X1 U9438 ( .A1(n7826), .A2(n8762), .B1(n7754), .B2(n8764), .ZN(n7762)
         );
  INV_X1 U9439 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10385) );
  NOR2_X1 U9440 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10385), .ZN(n8582) );
  AOI21_X1 U9441 ( .B1(n8475), .B2(n7762), .A(n8582), .ZN(n7755) );
  OAI21_X1 U9442 ( .B1(n7768), .B2(n8498), .A(n7755), .ZN(n7756) );
  AOI21_X1 U9443 ( .B1(n8907), .B2(n8492), .A(n7756), .ZN(n7757) );
  OAI21_X1 U9444 ( .B1(n7758), .B2(n8505), .A(n7757), .ZN(P2_U3230) );
  OAI222_X1 U9445 ( .A1(n7760), .A2(P1_U3084), .B1(n9548), .B2(n7759), .C1(
        n10171), .C2(n9541), .ZN(P1_U3327) );
  NAND2_X1 U9446 ( .A1(n8907), .A2(n7781), .ZN(n7899) );
  NAND2_X1 U9447 ( .A1(n7901), .A2(n7899), .ZN(n7824) );
  XNOR2_X1 U9448 ( .A(n7825), .B(n7990), .ZN(n7763) );
  AOI21_X1 U9449 ( .B1(n7763), .B2(n8804), .A(n7762), .ZN(n8909) );
  NAND2_X1 U9450 ( .A1(n8912), .A2(n8537), .ZN(n7764) );
  NAND2_X1 U9451 ( .A1(n7765), .A2(n7764), .ZN(n7767) );
  INV_X1 U9452 ( .A(n8397), .ZN(n7766) );
  AOI21_X1 U9453 ( .B1(n7990), .B2(n7767), .A(n7766), .ZN(n8910) );
  INV_X1 U9454 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7769) );
  OAI22_X1 U9455 ( .A1(n8696), .A2(n7769), .B1(n7768), .B2(n8821), .ZN(n7770)
         );
  AOI21_X1 U9456 ( .B1(n8907), .B2(n8620), .A(n7770), .ZN(n7776) );
  INV_X1 U9457 ( .A(n8907), .ZN(n7773) );
  OAI21_X1 U9458 ( .B1(n7773), .B2(n7772), .A(n10014), .ZN(n7774) );
  NOR2_X1 U9459 ( .A1(n7774), .A2(n8796), .ZN(n8906) );
  NAND2_X1 U9460 ( .A1(n8906), .A2(n8829), .ZN(n7775) );
  OAI211_X1 U9461 ( .C1(n8910), .C2(n8818), .A(n7776), .B(n7775), .ZN(n7777)
         );
  INV_X1 U9462 ( .A(n7777), .ZN(n7778) );
  OAI21_X1 U9463 ( .B1(n8788), .B2(n8909), .A(n7778), .ZN(P2_U3279) );
  XNOR2_X1 U9464 ( .A(n7779), .B(n7780), .ZN(n7785) );
  INV_X1 U9465 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10222) );
  OAI22_X1 U9466 ( .A1(n8498), .A2(n8799), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10222), .ZN(n7783) );
  OAI22_X1 U9467 ( .A1(n7781), .A2(n8500), .B1(n8499), .B2(n8765), .ZN(n7782)
         );
  AOI211_X1 U9468 ( .C1(n8901), .C2(n8503), .A(n7783), .B(n7782), .ZN(n7784)
         );
  OAI21_X1 U9469 ( .B1(n7785), .B2(n8505), .A(n7784), .ZN(P2_U3240) );
  OAI222_X1 U9470 ( .A1(n7789), .A2(n7788), .B1(n8944), .B2(n7787), .C1(n7786), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  XNOR2_X1 U9471 ( .A(n7791), .B(n7790), .ZN(n7798) );
  OAI22_X1 U9472 ( .A1(n8498), .A2(n7792), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10459), .ZN(n7796) );
  OAI22_X1 U9473 ( .A1(n7794), .A2(n8500), .B1(n8499), .B2(n7793), .ZN(n7795)
         );
  AOI211_X1 U9474 ( .C1(n10012), .C2(n8503), .A(n7796), .B(n7795), .ZN(n7797)
         );
  OAI21_X1 U9475 ( .B1(n7798), .B2(n8505), .A(n7797), .ZN(P2_U3238) );
  INV_X1 U9476 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10147) );
  INV_X1 U9477 ( .A(n7830), .ZN(n8940) );
  OAI222_X1 U9478 ( .A1(n9541), .A2(n10147), .B1(n9548), .B2(n8940), .C1(n7799), .C2(P1_U3084), .ZN(P1_U3324) );
  INV_X1 U9479 ( .A(n7800), .ZN(n7812) );
  NAND2_X1 U9480 ( .A1(n9167), .A2(n7801), .ZN(n7803) );
  NAND2_X1 U9481 ( .A1(n9088), .A2(n7806), .ZN(n7802) );
  NAND2_X1 U9482 ( .A1(n7803), .A2(n7802), .ZN(n7805) );
  XNOR2_X1 U9483 ( .A(n7805), .B(n7804), .ZN(n7810) );
  NAND2_X1 U9484 ( .A1(n9167), .A2(n7806), .ZN(n7807) );
  OAI21_X1 U9485 ( .B1(n9182), .B2(n7808), .A(n7807), .ZN(n7809) );
  XNOR2_X1 U9486 ( .A(n7810), .B(n7809), .ZN(n7817) );
  INV_X1 U9487 ( .A(n7817), .ZN(n7811) );
  NAND2_X1 U9488 ( .A1(n7811), .A2(n9056), .ZN(n7822) );
  NAND2_X1 U9489 ( .A1(n7813), .A2(n7812), .ZN(n7816) );
  NAND4_X1 U9490 ( .A1(n7823), .A2(n9056), .A3(n7817), .A4(n7816), .ZN(n7821)
         );
  AOI22_X1 U9491 ( .A1(n9170), .A2(n9076), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7815) );
  NAND2_X1 U9492 ( .A1(n9163), .A2(n9064), .ZN(n7814) );
  OAI211_X1 U9493 ( .C1(n9199), .C2(n9062), .A(n7815), .B(n7814), .ZN(n7819)
         );
  NOR3_X1 U9494 ( .A1(n7817), .A2(n9085), .A3(n7816), .ZN(n7818) );
  AOI211_X1 U9495 ( .C1(n9082), .C2(n9167), .A(n7819), .B(n7818), .ZN(n7820)
         );
  OAI211_X1 U9496 ( .C1(n7823), .C2(n7822), .A(n7821), .B(n7820), .ZN(P1_U3218) );
  NAND2_X1 U9497 ( .A1(n8901), .A2(n7826), .ZN(n7999) );
  NAND2_X1 U9498 ( .A1(n8807), .A2(n8806), .ZN(n8805) );
  OR2_X1 U9499 ( .A1(n8897), .A2(n8765), .ZN(n7993) );
  NAND2_X1 U9500 ( .A1(n8897), .A2(n8765), .ZN(n8757) );
  NAND2_X1 U9501 ( .A1(n7993), .A2(n8757), .ZN(n7866) );
  INV_X1 U9502 ( .A(n8779), .ZN(n7827) );
  NOR2_X1 U9503 ( .A1(n7866), .A2(n7827), .ZN(n7828) );
  INV_X1 U9504 ( .A(n8757), .ZN(n7994) );
  NAND2_X1 U9505 ( .A1(n8888), .A2(n8464), .ZN(n8001) );
  NAND2_X1 U9506 ( .A1(n8003), .A2(n8001), .ZN(n8400) );
  INV_X1 U9507 ( .A(n8003), .ZN(n7996) );
  XNOR2_X1 U9508 ( .A(n8882), .B(n8535), .ZN(n8749) );
  INV_X1 U9509 ( .A(n8535), .ZN(n8763) );
  NAND2_X1 U9510 ( .A1(n8882), .A2(n8763), .ZN(n8006) );
  NAND2_X1 U9511 ( .A1(n8877), .A2(n8534), .ZN(n8010) );
  NAND2_X1 U9512 ( .A1(n8008), .A2(n8010), .ZN(n8734) );
  INV_X1 U9513 ( .A(n8008), .ZN(n8721) );
  NAND2_X1 U9514 ( .A1(n8872), .A2(n8736), .ZN(n7829) );
  INV_X1 U9515 ( .A(n7829), .ZN(n7896) );
  NAND2_X1 U9516 ( .A1(n8867), .A2(n8472), .ZN(n8017) );
  AND2_X2 U9517 ( .A1(n8020), .A2(n8017), .ZN(n8705) );
  NAND2_X1 U9518 ( .A1(n8706), .A2(n8705), .ZN(n8704) );
  NAND2_X1 U9519 ( .A1(n8704), .A2(n8020), .ZN(n8687) );
  XNOR2_X1 U9520 ( .A(n8864), .B(n8707), .ZN(n8688) );
  NAND2_X1 U9521 ( .A1(n8687), .A2(n8688), .ZN(n8686) );
  OR2_X1 U9522 ( .A1(n8858), .A2(n8657), .ZN(n8025) );
  INV_X1 U9523 ( .A(n8707), .ZN(n8489) );
  OR2_X1 U9524 ( .A1(n8864), .A2(n8489), .ZN(n8673) );
  NAND3_X1 U9525 ( .A1(n8686), .A2(n8675), .A3(n8673), .ZN(n8674) );
  NOR2_X1 U9526 ( .A1(n8852), .A2(n8630), .ZN(n8038) );
  NAND2_X1 U9527 ( .A1(n8847), .A2(n8658), .ZN(n8036) );
  NAND2_X1 U9528 ( .A1(n7830), .A2(n5891), .ZN(n7832) );
  NAND2_X1 U9529 ( .A1(n4487), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7831) );
  NOR2_X1 U9530 ( .A1(n8416), .A2(n8634), .ZN(n8041) );
  INV_X1 U9531 ( .A(n8041), .ZN(n8037) );
  OAI21_X1 U9532 ( .B1(n7833), .B2(n8044), .A(n8037), .ZN(n7849) );
  INV_X1 U9533 ( .A(n7849), .ZN(n7851) );
  NOR2_X1 U9534 ( .A1(n7834), .A2(SI_29_), .ZN(n7836) );
  NAND2_X1 U9535 ( .A1(n7834), .A2(SI_29_), .ZN(n7835) );
  MUX2_X1 U9536 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7856), .Z(n7853) );
  NAND2_X1 U9537 ( .A1(n8935), .A2(n5891), .ZN(n7839) );
  NAND2_X1 U9538 ( .A1(n4487), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7838) );
  INV_X1 U9539 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U9540 ( .A1(n7844), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U9541 ( .A1(n5975), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7840) );
  OAI211_X1 U9542 ( .C1(n7843), .C2(n7842), .A(n7841), .B(n7840), .ZN(n8531)
         );
  INV_X1 U9543 ( .A(n8531), .ZN(n7861) );
  NOR2_X1 U9544 ( .A1(n8837), .A2(n7861), .ZN(n8049) );
  NAND2_X1 U9545 ( .A1(n5975), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U9546 ( .A1(n7844), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7847) );
  NAND2_X1 U9547 ( .A1(n7845), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7846) );
  OAI211_X1 U9548 ( .C1(n7849), .C2(n8837), .A(n6255), .B(n8530), .ZN(n7850)
         );
  OAI21_X1 U9549 ( .B1(n7851), .B2(n8049), .A(n7850), .ZN(n7862) );
  NAND2_X1 U9550 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  MUX2_X1 U9551 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7856), .Z(n7857) );
  XNOR2_X1 U9552 ( .A(n7857), .B(SI_31_), .ZN(n7858) );
  NAND2_X1 U9553 ( .A1(n8194), .A2(n5891), .ZN(n7860) );
  NAND2_X1 U9554 ( .A1(n4487), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7859) );
  OR2_X1 U9555 ( .A1(n8834), .A2(n8530), .ZN(n8054) );
  NAND2_X1 U9556 ( .A1(n8837), .A2(n7861), .ZN(n8048) );
  NAND2_X1 U9557 ( .A1(n8054), .A2(n8048), .ZN(n8052) );
  NAND2_X1 U9558 ( .A1(n8834), .A2(n8530), .ZN(n8055) );
  NAND2_X1 U9559 ( .A1(n7864), .A2(n7863), .ZN(n8066) );
  INV_X1 U9560 ( .A(n8049), .ZN(n7865) );
  NAND2_X1 U9561 ( .A1(n8055), .A2(n7865), .ZN(n8051) );
  INV_X1 U9562 ( .A(n8051), .ZN(n7891) );
  INV_X1 U9563 ( .A(n8052), .ZN(n7890) );
  INV_X1 U9564 ( .A(n7866), .ZN(n8778) );
  NAND4_X1 U9565 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n7874)
         );
  NOR4_X1 U9566 ( .A1(n7874), .A2(n7873), .A3(n7872), .A4(n7871), .ZN(n7875)
         );
  NAND4_X1 U9567 ( .A1(n7876), .A2(n7946), .A3(n7275), .A4(n7875), .ZN(n7877)
         );
  NOR4_X1 U9568 ( .A1(n7879), .A2(n7271), .A3(n7878), .A4(n7877), .ZN(n7880)
         );
  NAND3_X1 U9569 ( .A1(n7970), .A2(n7881), .A3(n7880), .ZN(n7882) );
  NOR4_X1 U9570 ( .A1(n7902), .A2(n7884), .A3(n7883), .A4(n7882), .ZN(n7885)
         );
  NAND4_X1 U9571 ( .A1(n8778), .A2(n7990), .A3(n8806), .A4(n7885), .ZN(n7886)
         );
  NOR4_X1 U9572 ( .A1(n8720), .A2(n8734), .A3(n8400), .A4(n7886), .ZN(n7887)
         );
  NAND4_X1 U9573 ( .A1(n8675), .A2(n8705), .A3(n7887), .A4(n8749), .ZN(n7888)
         );
  INV_X1 U9574 ( .A(n8688), .ZN(n8683) );
  NOR4_X1 U9575 ( .A1(n8643), .A2(n8656), .A3(n7888), .A4(n8683), .ZN(n7889)
         );
  NAND4_X1 U9576 ( .A1(n7891), .A2(n7890), .A3(n8404), .A4(n7889), .ZN(n7893)
         );
  XNOR2_X1 U9577 ( .A(n7893), .B(n7892), .ZN(n8060) );
  INV_X1 U9578 ( .A(n8036), .ZN(n7894) );
  AOI21_X1 U9579 ( .B1(n8630), .B2(n8852), .A(n7894), .ZN(n8035) );
  OR2_X1 U9580 ( .A1(n6254), .A2(n7895), .ZN(n8053) );
  INV_X1 U9581 ( .A(n8053), .ZN(n8034) );
  INV_X1 U9582 ( .A(n8017), .ZN(n7897) );
  OAI21_X1 U9583 ( .B1(n7897), .B2(n7896), .A(n8053), .ZN(n8023) );
  OR2_X1 U9584 ( .A1(n8882), .A2(n8763), .ZN(n8002) );
  INV_X1 U9585 ( .A(n8002), .ZN(n7898) );
  NOR3_X1 U9586 ( .A1(n8721), .A2(n7898), .A3(n8053), .ZN(n8015) );
  AND2_X1 U9587 ( .A1(n7999), .A2(n7899), .ZN(n7900) );
  MUX2_X1 U9588 ( .A(n7901), .B(n7900), .S(n8034), .Z(n7992) );
  NAND2_X1 U9589 ( .A1(n7959), .A2(n7903), .ZN(n7911) );
  INV_X1 U9590 ( .A(n7909), .ZN(n7905) );
  NAND2_X1 U9591 ( .A1(n7903), .A2(n7956), .ZN(n7904) );
  MUX2_X1 U9592 ( .A(n7905), .B(n7904), .S(n8053), .Z(n7907) );
  INV_X1 U9593 ( .A(n7908), .ZN(n7906) );
  OR2_X1 U9594 ( .A1(n7907), .A2(n7906), .ZN(n7912) );
  OAI211_X1 U9595 ( .C1(n7912), .C2(n7909), .A(n4545), .B(n7908), .ZN(n7910)
         );
  MUX2_X1 U9596 ( .A(n7911), .B(n7910), .S(n8053), .Z(n7966) );
  INV_X1 U9597 ( .A(n7912), .ZN(n7958) );
  AND2_X1 U9598 ( .A1(n7924), .A2(n7922), .ZN(n7916) );
  INV_X1 U9599 ( .A(n7918), .ZN(n7913) );
  NOR2_X1 U9600 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  NAND2_X1 U9601 ( .A1(n7918), .A2(n7917), .ZN(n7921) );
  NAND2_X1 U9602 ( .A1(n7919), .A2(n7943), .ZN(n7920) );
  AOI21_X1 U9603 ( .B1(n7931), .B2(n7921), .A(n7920), .ZN(n7945) );
  NAND2_X1 U9604 ( .A1(n7923), .A2(n7922), .ZN(n7926) );
  NAND2_X1 U9605 ( .A1(n7948), .A2(n7924), .ZN(n7925) );
  AOI21_X1 U9606 ( .B1(n7931), .B2(n7926), .A(n7925), .ZN(n7934) );
  AND2_X1 U9607 ( .A1(n7936), .A2(n6255), .ZN(n7928) );
  OAI211_X1 U9608 ( .C1(n7928), .C2(n7927), .A(n7940), .B(n7935), .ZN(n7929)
         );
  NAND3_X1 U9609 ( .A1(n7929), .A2(n7938), .A3(n8053), .ZN(n7932) );
  NAND3_X1 U9610 ( .A1(n7932), .A2(n7931), .A3(n7930), .ZN(n7933) );
  OAI21_X1 U9611 ( .B1(n7934), .B2(n8034), .A(n7933), .ZN(n7944) );
  NAND2_X1 U9612 ( .A1(n7936), .A2(n7935), .ZN(n7939) );
  NAND3_X1 U9613 ( .A1(n7939), .A2(n7938), .A3(n7937), .ZN(n7941) );
  NAND3_X1 U9614 ( .A1(n7941), .A2(n8034), .A3(n7940), .ZN(n7942) );
  OAI211_X1 U9615 ( .C1(n7948), .C2(n8053), .A(n7947), .B(n7946), .ZN(n7952)
         );
  MUX2_X1 U9616 ( .A(n7950), .B(n7949), .S(n8053), .Z(n7951) );
  NAND3_X1 U9617 ( .A1(n7952), .A2(n7275), .A3(n7951), .ZN(n7957) );
  MUX2_X1 U9618 ( .A(n7954), .B(n7953), .S(n8053), .Z(n7955) );
  AND2_X1 U9619 ( .A1(n4545), .A2(n7968), .ZN(n7963) );
  INV_X1 U9620 ( .A(n7959), .ZN(n7960) );
  NOR2_X1 U9621 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  MUX2_X1 U9622 ( .A(n7963), .B(n7962), .S(n8053), .Z(n7964) );
  OAI21_X1 U9623 ( .B1(n7966), .B2(n7965), .A(n7964), .ZN(n7971) );
  MUX2_X1 U9624 ( .A(n7968), .B(n7967), .S(n8034), .Z(n7969) );
  NAND3_X1 U9625 ( .A1(n7971), .A2(n7970), .A3(n7969), .ZN(n7975) );
  MUX2_X1 U9626 ( .A(n7973), .B(n7972), .S(n8053), .Z(n7974) );
  MUX2_X1 U9627 ( .A(n7978), .B(n7977), .S(n8053), .Z(n7979) );
  NAND2_X1 U9628 ( .A1(n7981), .A2(n7980), .ZN(n7985) );
  MUX2_X1 U9629 ( .A(n7983), .B(n7982), .S(n8034), .Z(n7984) );
  NAND3_X1 U9630 ( .A1(n7727), .A2(n7985), .A3(n7984), .ZN(n7989) );
  MUX2_X1 U9631 ( .A(n7987), .B(n7986), .S(n8053), .Z(n7988) );
  NAND3_X1 U9632 ( .A1(n7990), .A2(n7989), .A3(n7988), .ZN(n7991) );
  NAND2_X1 U9633 ( .A1(n7992), .A2(n7991), .ZN(n8000) );
  NAND2_X1 U9634 ( .A1(n7993), .A2(n8779), .ZN(n7998) );
  INV_X1 U9635 ( .A(n7998), .ZN(n7995) );
  AOI21_X1 U9636 ( .B1(n8000), .B2(n7995), .A(n7994), .ZN(n7997) );
  OAI211_X1 U9637 ( .C1(n7997), .C2(n7996), .A(n8006), .B(n8001), .ZN(n8014)
         );
  NAND2_X1 U9638 ( .A1(n8001), .A2(n8757), .ZN(n8004) );
  OAI211_X1 U9639 ( .C1(n8005), .C2(n8004), .A(n8003), .B(n8002), .ZN(n8007)
         );
  NAND2_X1 U9640 ( .A1(n8009), .A2(n8008), .ZN(n8012) );
  INV_X1 U9641 ( .A(n8010), .ZN(n8011) );
  AOI211_X1 U9642 ( .C1(n8015), .C2(n8014), .A(n8720), .B(n8013), .ZN(n8019)
         );
  AOI21_X1 U9643 ( .B1(n8705), .B2(n8016), .A(n8053), .ZN(n8018) );
  OAI21_X1 U9644 ( .B1(n8019), .B2(n8018), .A(n8017), .ZN(n8022) );
  OAI211_X1 U9645 ( .C1(n8034), .C2(n8020), .A(n8675), .B(n8688), .ZN(n8021)
         );
  AOI21_X1 U9646 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n8032) );
  INV_X1 U9647 ( .A(n8028), .ZN(n8024) );
  AOI21_X1 U9648 ( .B1(n8673), .B2(n8025), .A(n8024), .ZN(n8030) );
  NAND2_X1 U9649 ( .A1(n8864), .A2(n8489), .ZN(n8027) );
  INV_X1 U9650 ( .A(n8025), .ZN(n8026) );
  AOI21_X1 U9651 ( .B1(n8028), .B2(n8027), .A(n8026), .ZN(n8029) );
  OAI21_X1 U9652 ( .B1(n8032), .B2(n8031), .A(n5032), .ZN(n8033) );
  OAI211_X1 U9653 ( .C1(n8043), .C2(n8038), .A(n8037), .B(n8036), .ZN(n8040)
         );
  INV_X1 U9654 ( .A(n8044), .ZN(n8039) );
  NAND2_X1 U9655 ( .A1(n8040), .A2(n8039), .ZN(n8047) );
  AOI21_X1 U9656 ( .B1(n8043), .B2(n8042), .A(n8041), .ZN(n8045) );
  NOR2_X1 U9657 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  MUX2_X1 U9658 ( .A(n8047), .B(n8046), .S(n8053), .Z(n8050) );
  MUX2_X1 U9659 ( .A(n8052), .B(n8051), .S(n8053), .Z(n8057) );
  MUX2_X1 U9660 ( .A(n8055), .B(n8054), .S(n8053), .Z(n8056) );
  INV_X1 U9661 ( .A(n8058), .ZN(n8063) );
  OAI21_X1 U9662 ( .B1(n8062), .B2(n8063), .A(n8061), .ZN(n8059) );
  OAI21_X1 U9663 ( .B1(n6255), .B2(n8060), .A(n8059), .ZN(n8065) );
  OAI211_X1 U9664 ( .C1(n4927), .C2(n8063), .A(n8062), .B(n8061), .ZN(n8064)
         );
  NOR2_X1 U9665 ( .A1(n4484), .A2(P2_U3152), .ZN(n8946) );
  NAND3_X1 U9666 ( .A1(n8067), .A2(n8809), .A3(n8946), .ZN(n8068) );
  OAI211_X1 U9667 ( .C1(n6254), .C2(n8070), .A(n8068), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8069) );
  AOI21_X1 U9668 ( .B1(n8076), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8071), .ZN(
        n9131) );
  NAND2_X1 U9669 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9121), .ZN(n8072) );
  OAI21_X1 U9670 ( .B1(n9121), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8072), .ZN(
        n9130) );
  NOR2_X1 U9671 ( .A1(n9131), .A2(n9130), .ZN(n9129) );
  OR2_X1 U9672 ( .A1(n8077), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U9673 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n8077), .ZN(n8073) );
  NAND2_X1 U9674 ( .A1(n8074), .A2(n8073), .ZN(n9733) );
  INV_X1 U9675 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9450) );
  AOI22_X1 U9676 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n8077), .B1(n9738), .B2(
        n9450), .ZN(n9742) );
  AOI21_X1 U9677 ( .B1(n8076), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8075), .ZN(
        n9123) );
  XNOR2_X1 U9678 ( .A(n9121), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9124) );
  NOR2_X1 U9679 ( .A1(n9123), .A2(n9124), .ZN(n9122) );
  AOI21_X1 U9680 ( .B1(n9121), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9122), .ZN(
        n9743) );
  NAND2_X1 U9681 ( .A1(n9742), .A2(n9743), .ZN(n9741) );
  OAI21_X1 U9682 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n8077), .A(n9741), .ZN(
        n8078) );
  XOR2_X1 U9683 ( .A(n8078), .B(n9442), .Z(n8083) );
  INV_X1 U9684 ( .A(n8083), .ZN(n8079) );
  NAND2_X1 U9685 ( .A1(n8079), .A2(n9744), .ZN(n8080) );
  OAI211_X1 U9686 ( .C1(n8084), .C2(n8081), .A(n8080), .B(n9739), .ZN(n8082)
         );
  INV_X1 U9687 ( .A(n8082), .ZN(n8086) );
  AOI22_X1 U9688 ( .A1(n8084), .A2(n9735), .B1(n9744), .B2(n8083), .ZN(n8085)
         );
  MUX2_X1 U9689 ( .A(n8086), .B(n8085), .S(n9814), .Z(n8088) );
  NAND2_X1 U9690 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n8087) );
  OAI211_X1 U9691 ( .C1(n10486), .C2(n9748), .A(n8088), .B(n8087), .ZN(
        P1_U3260) );
  INV_X1 U9692 ( .A(n8165), .ZN(n8089) );
  OAI211_X1 U9693 ( .C1(n8089), .C2(n8091), .A(n8311), .B(n8092), .ZN(n8090)
         );
  INV_X1 U9694 ( .A(n8090), .ZN(n8095) );
  INV_X1 U9695 ( .A(n8166), .ZN(n8094) );
  AND2_X1 U9696 ( .A1(n8092), .A2(n8091), .ZN(n8302) );
  NAND2_X1 U9697 ( .A1(n8178), .A2(n8165), .ZN(n8093) );
  INV_X1 U9698 ( .A(n8200), .ZN(n8198) );
  MUX2_X1 U9699 ( .A(n8095), .B(n8361), .S(n8198), .Z(n8168) );
  INV_X1 U9700 ( .A(n8153), .ZN(n8096) );
  NAND2_X1 U9701 ( .A1(n8298), .A2(n8096), .ZN(n8160) );
  NAND2_X1 U9702 ( .A1(n8161), .A2(n8160), .ZN(n8352) );
  OR3_X1 U9703 ( .A1(n8352), .A2(n8198), .A3(n8298), .ZN(n8163) );
  INV_X1 U9704 ( .A(n8251), .ZN(n8100) );
  NAND2_X1 U9705 ( .A1(n8253), .A2(n8100), .ZN(n8097) );
  NAND2_X1 U9706 ( .A1(n8152), .A2(n8099), .ZN(n8295) );
  MUX2_X1 U9707 ( .A(n8097), .B(n8295), .S(n8200), .Z(n8098) );
  INV_X1 U9708 ( .A(n8098), .ZN(n8151) );
  AND2_X1 U9709 ( .A1(n8284), .A2(n8200), .ZN(n8102) );
  NAND4_X1 U9710 ( .A1(n8101), .A2(n8102), .A3(n8283), .A4(n8108), .ZN(n8117)
         );
  INV_X1 U9711 ( .A(n8102), .ZN(n8106) );
  NOR2_X1 U9712 ( .A1(n9887), .A2(n8200), .ZN(n8104) );
  OAI21_X1 U9713 ( .B1(n8198), .B2(n9864), .A(n9879), .ZN(n8103) );
  OAI21_X1 U9714 ( .B1(n8104), .B2(n9879), .A(n8103), .ZN(n8105) );
  OAI21_X1 U9715 ( .B1(n8106), .B2(n8286), .A(n8105), .ZN(n8107) );
  INV_X1 U9716 ( .A(n8107), .ZN(n8116) );
  INV_X1 U9717 ( .A(n9777), .ZN(n8109) );
  OAI211_X1 U9718 ( .C1(n8110), .C2(n8109), .A(n8108), .B(n8287), .ZN(n8111)
         );
  AND2_X1 U9719 ( .A1(n8273), .A2(n8198), .ZN(n8112) );
  NAND4_X1 U9720 ( .A1(n8111), .A2(n8112), .A3(n8286), .A4(n8289), .ZN(n8115)
         );
  INV_X1 U9721 ( .A(n8112), .ZN(n8113) );
  OR2_X1 U9722 ( .A1(n8113), .A2(n8283), .ZN(n8114) );
  NAND4_X1 U9723 ( .A1(n8117), .A2(n8116), .A3(n8115), .A4(n8114), .ZN(n8122)
         );
  NAND2_X1 U9724 ( .A1(n8211), .A2(n8274), .ZN(n8118) );
  AOI21_X1 U9725 ( .B1(n8122), .B2(n8255), .A(n8118), .ZN(n8120) );
  NAND2_X1 U9726 ( .A1(n8212), .A2(n8255), .ZN(n8121) );
  AOI21_X1 U9727 ( .B1(n8122), .B2(n8274), .A(n8121), .ZN(n8125) );
  INV_X1 U9728 ( .A(n8258), .ZN(n8128) );
  INV_X1 U9729 ( .A(n8129), .ZN(n8131) );
  OAI211_X1 U9730 ( .C1(n8131), .C2(n8130), .A(n8260), .B(n8258), .ZN(n8132)
         );
  INV_X1 U9731 ( .A(n8132), .ZN(n8133) );
  NAND2_X1 U9732 ( .A1(n8137), .A2(n8133), .ZN(n8136) );
  AND2_X1 U9733 ( .A1(n8139), .A2(n8134), .ZN(n8264) );
  AND2_X1 U9734 ( .A1(n8962), .A2(n8135), .ZN(n8138) );
  AOI21_X1 U9735 ( .B1(n8136), .B2(n8264), .A(n8138), .ZN(n8144) );
  INV_X1 U9736 ( .A(n8138), .ZN(n8276) );
  NAND2_X1 U9737 ( .A1(n8276), .A2(n8260), .ZN(n8140) );
  NAND2_X1 U9738 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U9739 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  MUX2_X1 U9740 ( .A(n8144), .B(n8143), .S(n8200), .Z(n8147) );
  MUX2_X1 U9741 ( .A(n8278), .B(n8254), .S(n8200), .Z(n8145) );
  NOR2_X1 U9742 ( .A1(n9346), .A2(n8145), .ZN(n8146) );
  OAI21_X1 U9743 ( .B1(n8147), .B2(n8230), .A(n8146), .ZN(n8149) );
  MUX2_X1 U9744 ( .A(n8270), .B(n8249), .S(n8200), .Z(n8148) );
  NAND3_X1 U9745 ( .A1(n9339), .A2(n8149), .A3(n8148), .ZN(n8150) );
  NAND2_X1 U9746 ( .A1(n8151), .A2(n8150), .ZN(n8157) );
  NAND3_X1 U9747 ( .A1(n8157), .A2(n8156), .A3(n8152), .ZN(n8154) );
  NAND2_X1 U9748 ( .A1(n8303), .A2(n8198), .ZN(n8155) );
  AND2_X1 U9749 ( .A1(n9270), .A2(n8156), .ZN(n8297) );
  AND2_X1 U9750 ( .A1(n8281), .A2(n8253), .ZN(n8296) );
  NAND2_X1 U9751 ( .A1(n8157), .A2(n8296), .ZN(n8158) );
  NAND2_X1 U9752 ( .A1(n8297), .A2(n8158), .ZN(n8159) );
  NAND4_X1 U9753 ( .A1(n8161), .A2(n8200), .A3(n8160), .A4(n8159), .ZN(n8162)
         );
  NAND4_X1 U9754 ( .A1(n8302), .A2(n8166), .A3(n8165), .A4(n8164), .ZN(n8167)
         );
  NAND2_X1 U9755 ( .A1(n8168), .A2(n8167), .ZN(n8175) );
  OAI21_X1 U9756 ( .B1(n8175), .B2(n9216), .A(n8200), .ZN(n8170) );
  AOI21_X1 U9757 ( .B1(n8175), .B2(n8311), .A(n9201), .ZN(n8169) );
  NAND2_X1 U9758 ( .A1(n8170), .A2(n8169), .ZN(n8174) );
  NOR2_X1 U9759 ( .A1(n8178), .A2(n9216), .ZN(n8171) );
  NOR2_X1 U9760 ( .A1(n8171), .A2(n9201), .ZN(n8172) );
  MUX2_X1 U9761 ( .A(n8995), .B(n8172), .S(n8200), .Z(n8173) );
  NAND2_X1 U9762 ( .A1(n8174), .A2(n8173), .ZN(n8185) );
  INV_X1 U9763 ( .A(n8175), .ZN(n8176) );
  NAND2_X1 U9764 ( .A1(n8176), .A2(n9178), .ZN(n8183) );
  NAND2_X1 U9765 ( .A1(n9201), .A2(n8311), .ZN(n8177) );
  NAND2_X1 U9766 ( .A1(n8317), .A2(n8177), .ZN(n8181) );
  NAND2_X1 U9767 ( .A1(n8178), .A2(n9216), .ZN(n8179) );
  NAND2_X1 U9768 ( .A1(n8362), .A2(n8179), .ZN(n8180) );
  MUX2_X1 U9769 ( .A(n8181), .B(n8180), .S(n8200), .Z(n8182) );
  NAND2_X1 U9770 ( .A1(n8183), .A2(n8182), .ZN(n8184) );
  NAND2_X1 U9771 ( .A1(n8185), .A2(n8184), .ZN(n8187) );
  MUX2_X1 U9772 ( .A(n8362), .B(n8317), .S(n8200), .Z(n8186) );
  MUX2_X1 U9773 ( .A(n8318), .B(n8308), .S(n8200), .Z(n8188) );
  INV_X1 U9774 ( .A(n8199), .ZN(n8189) );
  NOR2_X1 U9775 ( .A1(n8189), .A2(n9163), .ZN(n8190) );
  MUX2_X1 U9776 ( .A(n8190), .B(n8198), .S(n8307), .Z(n8204) );
  INV_X1 U9777 ( .A(n9163), .ZN(n8306) );
  NAND2_X1 U9778 ( .A1(n8935), .A2(n8193), .ZN(n8192) );
  NAND2_X1 U9779 ( .A1(n5627), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U9780 ( .A1(n9486), .A2(n9087), .ZN(n8371) );
  NAND2_X1 U9781 ( .A1(n8194), .A2(n8193), .ZN(n8196) );
  NAND2_X1 U9782 ( .A1(n5627), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8195) );
  AOI21_X1 U9783 ( .B1(n9140), .B2(n9087), .A(n9486), .ZN(n8324) );
  INV_X1 U9784 ( .A(n8324), .ZN(n8197) );
  OAI211_X1 U9785 ( .C1(n8306), .C2(n8198), .A(n4582), .B(n8197), .ZN(n8203)
         );
  INV_X1 U9786 ( .A(n9482), .ZN(n8202) );
  INV_X1 U9787 ( .A(n9140), .ZN(n8201) );
  NAND2_X1 U9788 ( .A1(n8202), .A2(n8201), .ZN(n8207) );
  INV_X1 U9789 ( .A(n8246), .ZN(n8395) );
  INV_X1 U9790 ( .A(n8205), .ZN(n8206) );
  NAND4_X1 U9791 ( .A1(n8373), .A2(n8387), .A3(n8206), .A4(n8386), .ZN(n8394)
         );
  INV_X1 U9792 ( .A(n8373), .ZN(n8242) );
  INV_X1 U9793 ( .A(n8207), .ZN(n8374) );
  INV_X1 U9794 ( .A(n8371), .ZN(n8241) );
  INV_X1 U9795 ( .A(n9486), .ZN(n8209) );
  INV_X1 U9796 ( .A(n9087), .ZN(n8208) );
  NAND2_X1 U9797 ( .A1(n8209), .A2(n8208), .ZN(n8369) );
  INV_X1 U9798 ( .A(n9346), .ZN(n9348) );
  NAND2_X1 U9799 ( .A1(n8212), .A2(n8211), .ZN(n9759) );
  NAND4_X1 U9800 ( .A1(n8215), .A2(n8214), .A3(n8213), .A4(n9807), .ZN(n8217)
         );
  NOR3_X1 U9801 ( .A1(n8217), .A2(n5342), .A3(n8216), .ZN(n8222) );
  INV_X1 U9802 ( .A(n8218), .ZN(n8221) );
  INV_X1 U9803 ( .A(n8219), .ZN(n8220) );
  NAND4_X1 U9804 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n8224)
         );
  NOR2_X1 U9805 ( .A1(n9759), .A2(n8224), .ZN(n8226) );
  INV_X1 U9806 ( .A(n9625), .ZN(n8225) );
  NAND4_X1 U9807 ( .A1(n8227), .A2(n4971), .A3(n8226), .A4(n8225), .ZN(n8228)
         );
  NOR4_X1 U9808 ( .A1(n8230), .A2(n8229), .A3(n9600), .A4(n8228), .ZN(n8231)
         );
  NAND3_X1 U9809 ( .A1(n9339), .A2(n9348), .A3(n8231), .ZN(n8232) );
  NOR2_X1 U9810 ( .A1(n8232), .A2(n9317), .ZN(n8233) );
  NAND3_X1 U9811 ( .A1(n9289), .A2(n9304), .A3(n8233), .ZN(n8234) );
  NOR2_X1 U9812 ( .A1(n9274), .A2(n8234), .ZN(n8235) );
  NAND3_X1 U9813 ( .A1(n9240), .A2(n9257), .A3(n8235), .ZN(n8236) );
  NOR2_X1 U9814 ( .A1(n9215), .A2(n8236), .ZN(n8237) );
  INV_X1 U9815 ( .A(n9224), .ZN(n9226) );
  AND4_X1 U9816 ( .A1(n9178), .A2(n9194), .A3(n8237), .A4(n9226), .ZN(n8239)
         );
  NAND4_X1 U9817 ( .A1(n8369), .A2(n9161), .A3(n8239), .A4(n8238), .ZN(n8240)
         );
  NAND2_X1 U9818 ( .A1(n8244), .A2(n8243), .ZN(n8248) );
  OAI21_X1 U9819 ( .B1(n8246), .B2(n8245), .A(n8248), .ZN(n8247) );
  INV_X1 U9820 ( .A(n8248), .ZN(n8329) );
  INV_X1 U9821 ( .A(n8249), .ZN(n8250) );
  NOR2_X1 U9822 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  NAND2_X1 U9823 ( .A1(n8253), .A2(n8252), .ZN(n8279) );
  INV_X1 U9824 ( .A(n8254), .ZN(n8269) );
  NOR2_X1 U9825 ( .A1(n8256), .A2(n4814), .ZN(n8263) );
  AND2_X1 U9826 ( .A1(n8258), .A2(n8257), .ZN(n8259) );
  NAND2_X1 U9827 ( .A1(n8260), .A2(n8259), .ZN(n8272) );
  INV_X1 U9828 ( .A(n8260), .ZN(n8262) );
  OAI22_X1 U9829 ( .A1(n8263), .A2(n8272), .B1(n8262), .B2(n8261), .ZN(n8267)
         );
  INV_X1 U9830 ( .A(n8264), .ZN(n8266) );
  OAI211_X1 U9831 ( .C1(n8267), .C2(n8266), .A(n8265), .B(n8276), .ZN(n8268)
         );
  AND3_X1 U9832 ( .A1(n8270), .A2(n8269), .A3(n8268), .ZN(n8271) );
  OR2_X1 U9833 ( .A1(n8279), .A2(n8271), .ZN(n8355) );
  INV_X1 U9834 ( .A(n8272), .ZN(n8275) );
  NAND4_X1 U9835 ( .A1(n8276), .A2(n8275), .A3(n8274), .A4(n8273), .ZN(n8277)
         );
  OR3_X1 U9836 ( .A1(n8279), .A2(n8278), .A3(n8277), .ZN(n8280) );
  NAND2_X1 U9837 ( .A1(n8355), .A2(n8280), .ZN(n8282) );
  AND2_X1 U9838 ( .A1(n8282), .A2(n8281), .ZN(n8351) );
  INV_X1 U9839 ( .A(n8355), .ZN(n8294) );
  AND2_X1 U9840 ( .A1(n8284), .A2(n8283), .ZN(n8343) );
  AND4_X1 U9841 ( .A1(n8343), .A2(n8287), .A3(n8285), .A4(n8345), .ZN(n8342)
         );
  INV_X1 U9842 ( .A(n8286), .ZN(n8288) );
  OAI21_X1 U9843 ( .B1(n8288), .B2(n8287), .A(n8345), .ZN(n8290) );
  AOI22_X1 U9844 ( .A1(n8344), .A2(n8338), .B1(n8290), .B2(n8289), .ZN(n8291)
         );
  AOI22_X1 U9845 ( .A1(n8342), .A2(n8292), .B1(n8291), .B2(n8343), .ZN(n8293)
         );
  OR2_X1 U9846 ( .A1(n8294), .A2(n8293), .ZN(n8301) );
  INV_X1 U9847 ( .A(n8295), .ZN(n8300) );
  INV_X1 U9848 ( .A(n8296), .ZN(n8299) );
  OAI211_X1 U9849 ( .C1(n8300), .C2(n8299), .A(n8298), .B(n8297), .ZN(n8359)
         );
  AOI21_X1 U9850 ( .B1(n8351), .B2(n8301), .A(n8359), .ZN(n8305) );
  INV_X1 U9851 ( .A(n8302), .ZN(n8304) );
  NOR2_X1 U9852 ( .A1(n8304), .A2(n4595), .ZN(n8356) );
  OAI21_X1 U9853 ( .B1(n8305), .B2(n8352), .A(n8356), .ZN(n8315) );
  INV_X1 U9854 ( .A(n8362), .ZN(n8314) );
  OR2_X1 U9855 ( .A1(n8307), .A2(n8306), .ZN(n8309) );
  NAND2_X1 U9856 ( .A1(n8309), .A2(n8308), .ZN(n8321) );
  INV_X1 U9857 ( .A(n8310), .ZN(n8313) );
  INV_X1 U9858 ( .A(n8311), .ZN(n8312) );
  OR3_X1 U9859 ( .A1(n8321), .A2(n8313), .A3(n8312), .ZN(n8368) );
  AOI211_X1 U9860 ( .C1(n8361), .C2(n8315), .A(n8314), .B(n8368), .ZN(n8323)
         );
  NAND2_X1 U9861 ( .A1(n8317), .A2(n8316), .ZN(n8320) );
  INV_X1 U9862 ( .A(n8318), .ZN(n8319) );
  AOI21_X1 U9863 ( .B1(n8362), .B2(n8320), .A(n8319), .ZN(n8322) );
  OAI22_X1 U9864 ( .A1(n8322), .A2(n8321), .B1(n5690), .B2(n9163), .ZN(n8365)
         );
  NOR3_X1 U9865 ( .A1(n8324), .A2(n8323), .A3(n8365), .ZN(n8326) );
  OAI211_X1 U9866 ( .C1(n8326), .C2(n8325), .A(n8332), .B(n8373), .ZN(n8327)
         );
  NAND4_X1 U9867 ( .A1(n8327), .A2(n8387), .A3(n4481), .A4(n9814), .ZN(n8328)
         );
  NOR2_X1 U9868 ( .A1(n8329), .A2(n8328), .ZN(n8391) );
  INV_X1 U9869 ( .A(n8352), .ZN(n8360) );
  INV_X1 U9870 ( .A(n8330), .ZN(n8331) );
  OAI211_X1 U9871 ( .C1(n8334), .C2(n8333), .A(n8332), .B(n8331), .ZN(n8335)
         );
  NAND3_X1 U9872 ( .A1(n8337), .A2(n8336), .A3(n8335), .ZN(n8341) );
  INV_X1 U9873 ( .A(n8338), .ZN(n8339) );
  AOI21_X1 U9874 ( .B1(n8341), .B2(n8340), .A(n8339), .ZN(n8350) );
  INV_X1 U9875 ( .A(n8342), .ZN(n8349) );
  INV_X1 U9876 ( .A(n8343), .ZN(n8348) );
  INV_X1 U9877 ( .A(n8344), .ZN(n8346) );
  NAND2_X1 U9878 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  OAI22_X1 U9879 ( .A1(n8350), .A2(n8349), .B1(n8348), .B2(n8347), .ZN(n8354)
         );
  INV_X1 U9880 ( .A(n8351), .ZN(n8353) );
  AOI211_X1 U9881 ( .C1(n8355), .C2(n8354), .A(n8353), .B(n8352), .ZN(n8358)
         );
  INV_X1 U9882 ( .A(n8356), .ZN(n8357) );
  AOI211_X1 U9883 ( .C1(n8360), .C2(n8359), .A(n8358), .B(n8357), .ZN(n8364)
         );
  INV_X1 U9884 ( .A(n8361), .ZN(n8363) );
  OAI21_X1 U9885 ( .B1(n8364), .B2(n8363), .A(n8362), .ZN(n8367) );
  INV_X1 U9886 ( .A(n8365), .ZN(n8366) );
  OAI21_X1 U9887 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8372) );
  INV_X1 U9888 ( .A(n8369), .ZN(n8370) );
  AOI21_X1 U9889 ( .B1(n8372), .B2(n8371), .A(n8370), .ZN(n8375) );
  OAI21_X1 U9890 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8377) );
  INV_X1 U9891 ( .A(n8387), .ZN(n8379) );
  NOR4_X1 U9892 ( .A1(n8377), .A2(n4481), .A3(n8379), .A4(n9814), .ZN(n8390)
         );
  INV_X1 U9893 ( .A(n8377), .ZN(n8380) );
  NOR3_X1 U9894 ( .A1(n8380), .A2(n8379), .A3(n8378), .ZN(n8389) );
  NOR3_X1 U9895 ( .A1(n8383), .A2(n8382), .A3(n8381), .ZN(n8384) );
  AOI211_X1 U9896 ( .C1(n8387), .C2(n8386), .A(n8385), .B(n8384), .ZN(n8388)
         );
  NOR4_X1 U9897 ( .A1(n8391), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(n8392)
         );
  OAI211_X1 U9898 ( .C1(n8395), .C2(n8394), .A(n8393), .B(n8392), .ZN(P1_U3240) );
  INV_X1 U9899 ( .A(n8657), .ZN(n8533) );
  INV_X1 U9900 ( .A(n8882), .ZN(n8747) );
  INV_X1 U9901 ( .A(n8464), .ZN(n8751) );
  OR2_X1 U9902 ( .A1(n8907), .A2(n8808), .ZN(n8396) );
  NOR2_X1 U9903 ( .A1(n8901), .A2(n8536), .ZN(n8398) );
  AND2_X1 U9904 ( .A1(n8897), .A2(n8811), .ZN(n8399) );
  NAND2_X1 U9905 ( .A1(n8644), .A2(n8643), .ZN(n8642) );
  XNOR2_X1 U9906 ( .A(n8405), .B(n8404), .ZN(n8412) );
  NAND2_X1 U9907 ( .A1(n8532), .A2(n8809), .ZN(n8410) );
  INV_X1 U9908 ( .A(n4484), .ZN(n8407) );
  AND2_X1 U9909 ( .A1(n8407), .A2(P2_B_REG_SCAN_IN), .ZN(n8408) );
  NOR2_X1 U9910 ( .A1(n8762), .A2(n8408), .ZN(n8618) );
  INV_X1 U9911 ( .A(n8844), .ZN(n8413) );
  NAND2_X1 U9912 ( .A1(n8413), .A2(n8696), .ZN(n8419) );
  INV_X1 U9913 ( .A(n8858), .ZN(n8672) );
  INV_X1 U9914 ( .A(n8901), .ZN(n8803) );
  AOI21_X1 U9915 ( .B1(n8841), .B2(n8635), .A(n8624), .ZN(n8842) );
  AOI22_X1 U9916 ( .A1(n8788), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8414), .B2(
        n8800), .ZN(n8415) );
  OAI21_X1 U9917 ( .B1(n8416), .B2(n8823), .A(n8415), .ZN(n8417) );
  AOI21_X1 U9918 ( .B1(n8842), .B2(n8816), .A(n8417), .ZN(n8418) );
  OAI211_X1 U9919 ( .C1(n8845), .C2(n8818), .A(n8419), .B(n8418), .ZN(P2_U3267) );
  XNOR2_X1 U9920 ( .A(n6818), .B(n9950), .ZN(n8421) );
  NAND2_X1 U9921 ( .A1(n8421), .A2(n10014), .ZN(n9955) );
  OAI22_X1 U9922 ( .A1(n8422), .A2(n9955), .B1(n10338), .B2(n8821), .ZN(n8423)
         );
  AOI21_X1 U9923 ( .B1(n8826), .B2(n9959), .A(n8423), .ZN(n8429) );
  AOI21_X1 U9924 ( .B1(n8426), .B2(n8804), .A(n8425), .ZN(n9956) );
  MUX2_X1 U9925 ( .A(n8427), .B(n9956), .S(n8696), .Z(n8428) );
  OAI211_X1 U9926 ( .C1(n6818), .C2(n8823), .A(n8429), .B(n8428), .ZN(P2_U3295) );
  OAI211_X1 U9927 ( .C1(n8432), .C2(n8431), .A(n8430), .B(n8517), .ZN(n8436)
         );
  AOI22_X1 U9928 ( .A1(n8526), .A2(n8651), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8435) );
  AOI22_X1 U9929 ( .A1(n8511), .A2(n8532), .B1(n8510), .B2(n8533), .ZN(n8434)
         );
  NAND2_X1 U9930 ( .A1(n8852), .A2(n8492), .ZN(n8433) );
  NAND4_X1 U9931 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(
        P2_U3216) );
  XNOR2_X1 U9932 ( .A(n8483), .B(n8482), .ZN(n8441) );
  INV_X1 U9933 ( .A(n8718), .ZN(n8437) );
  OAI22_X1 U9934 ( .A1(n8498), .A2(n8437), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10211), .ZN(n8439) );
  OAI22_X1 U9935 ( .A1(n8472), .A2(n8499), .B1(n8500), .B2(n8534), .ZN(n8438)
         );
  AOI211_X1 U9936 ( .C1(n8872), .C2(n8503), .A(n8439), .B(n8438), .ZN(n8440)
         );
  OAI21_X1 U9937 ( .B1(n8441), .B2(n8505), .A(n8440), .ZN(P2_U3218) );
  AOI22_X1 U9938 ( .A1(n8511), .A2(n8548), .B1(n8510), .B2(n8550), .ZN(n8449)
         );
  MUX2_X1 U9939 ( .A(P2_STATE_REG_SCAN_IN), .B(n8498), .S(n5850), .Z(n8448) );
  NAND2_X1 U9940 ( .A1(n8492), .A2(n8442), .ZN(n8447) );
  OAI211_X1 U9941 ( .C1(n8443), .C2(n8445), .A(n8517), .B(n8444), .ZN(n8446)
         );
  NAND4_X1 U9942 ( .A1(n8449), .A2(n8448), .A3(n8447), .A4(n8446), .ZN(
        P2_U3220) );
  INV_X1 U9943 ( .A(n8450), .ZN(n8451) );
  AOI21_X1 U9944 ( .B1(n8453), .B2(n8452), .A(n8451), .ZN(n8460) );
  INV_X1 U9945 ( .A(n8787), .ZN(n8457) );
  NAND2_X1 U9946 ( .A1(n8536), .A2(n8809), .ZN(n8455) );
  OR2_X1 U9947 ( .A1(n8464), .A2(n8762), .ZN(n8454) );
  NAND2_X1 U9948 ( .A1(n8455), .A2(n8454), .ZN(n8782) );
  AOI22_X1 U9949 ( .A1(n8475), .A2(n8782), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8456) );
  OAI21_X1 U9950 ( .B1(n8457), .B2(n8498), .A(n8456), .ZN(n8458) );
  AOI21_X1 U9951 ( .B1(n8897), .B2(n8492), .A(n8458), .ZN(n8459) );
  OAI21_X1 U9952 ( .B1(n8460), .B2(n8505), .A(n8459), .ZN(P2_U3221) );
  XNOR2_X1 U9953 ( .A(n8461), .B(n8462), .ZN(n8468) );
  INV_X1 U9954 ( .A(n8745), .ZN(n8463) );
  OAI22_X1 U9955 ( .A1(n8498), .A2(n8463), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10483), .ZN(n8466) );
  OAI22_X1 U9956 ( .A1(n8464), .A2(n8500), .B1(n8499), .B2(n8534), .ZN(n8465)
         );
  AOI211_X1 U9957 ( .C1(n8882), .C2(n8492), .A(n8466), .B(n8465), .ZN(n8467)
         );
  OAI21_X1 U9958 ( .B1(n8468), .B2(n8505), .A(n8467), .ZN(P2_U3225) );
  XNOR2_X1 U9959 ( .A(n8470), .B(n8469), .ZN(n8471) );
  XNOR2_X1 U9960 ( .A(n4549), .B(n8471), .ZN(n8480) );
  INV_X1 U9961 ( .A(n8692), .ZN(n8477) );
  OR2_X1 U9962 ( .A1(n8472), .A2(n8764), .ZN(n8474) );
  OR2_X1 U9963 ( .A1(n8657), .A2(n8762), .ZN(n8473) );
  NAND2_X1 U9964 ( .A1(n8474), .A2(n8473), .ZN(n8689) );
  AOI22_X1 U9965 ( .A1(n8475), .A2(n8689), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8476) );
  OAI21_X1 U9966 ( .B1(n8477), .B2(n8498), .A(n8476), .ZN(n8478) );
  AOI21_X1 U9967 ( .B1(n8864), .B2(n8492), .A(n8478), .ZN(n8479) );
  OAI21_X1 U9968 ( .B1(n8480), .B2(n8505), .A(n8479), .ZN(P2_U3227) );
  OAI21_X1 U9969 ( .B1(n8483), .B2(n8482), .A(n8481), .ZN(n8487) );
  XNOR2_X1 U9970 ( .A(n8485), .B(n8484), .ZN(n8486) );
  XNOR2_X1 U9971 ( .A(n8487), .B(n8486), .ZN(n8494) );
  INV_X1 U9972 ( .A(n8701), .ZN(n8488) );
  OAI22_X1 U9973 ( .A1(n8498), .A2(n8488), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10400), .ZN(n8491) );
  OAI22_X1 U9974 ( .A1(n8736), .A2(n8500), .B1(n8499), .B2(n8489), .ZN(n8490)
         );
  AOI211_X1 U9975 ( .C1(n8867), .C2(n8492), .A(n8491), .B(n8490), .ZN(n8493)
         );
  OAI21_X1 U9976 ( .B1(n8494), .B2(n8505), .A(n8493), .ZN(P2_U3231) );
  XNOR2_X1 U9977 ( .A(n8496), .B(n8495), .ZN(n8506) );
  INV_X1 U9978 ( .A(n8769), .ZN(n8497) );
  OAI22_X1 U9979 ( .A1(n8498), .A2(n8497), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10429), .ZN(n8502) );
  OAI22_X1 U9980 ( .A1(n8765), .A2(n8500), .B1(n8499), .B2(n8763), .ZN(n8501)
         );
  AOI211_X1 U9981 ( .C1(n8888), .C2(n8503), .A(n8502), .B(n8501), .ZN(n8504)
         );
  OAI21_X1 U9982 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(P2_U3235) );
  OAI21_X1 U9983 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8515) );
  AOI22_X1 U9984 ( .A1(n8526), .A2(n8730), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8513) );
  AOI22_X1 U9985 ( .A1(n8511), .A2(n5012), .B1(n8510), .B2(n8535), .ZN(n8512)
         );
  OAI211_X1 U9986 ( .C1(n8732), .C2(n8529), .A(n8513), .B(n8512), .ZN(n8514)
         );
  AOI21_X1 U9987 ( .B1(n8515), .B2(n8517), .A(n8514), .ZN(n8516) );
  INV_X1 U9988 ( .A(n8516), .ZN(P2_U3237) );
  OAI211_X1 U9989 ( .C1(n8520), .C2(n8519), .A(n8518), .B(n8517), .ZN(n8528)
         );
  OR2_X1 U9990 ( .A1(n8630), .A2(n8762), .ZN(n8522) );
  NAND2_X1 U9991 ( .A1(n8707), .A2(n8809), .ZN(n8521) );
  NAND2_X1 U9992 ( .A1(n8522), .A2(n8521), .ZN(n8677) );
  INV_X1 U9993 ( .A(n8677), .ZN(n8523) );
  OAI22_X1 U9994 ( .A1(n8524), .A2(n8523), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10182), .ZN(n8525) );
  AOI21_X1 U9995 ( .B1(n8670), .B2(n8526), .A(n8525), .ZN(n8527) );
  OAI211_X1 U9996 ( .C1(n8672), .C2(n8529), .A(n8528), .B(n8527), .ZN(P2_U3242) );
  INV_X1 U9997 ( .A(n8530), .ZN(n8619) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8619), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8531), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8634), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8532), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8533), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8707), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8723), .S(P2_U3966), .Z(
        P2_U3576) );
  INV_X1 U10005 ( .A(n8534), .ZN(n8752) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8752), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10007 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8535), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10008 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8751), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10009 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8811), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10010 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8536), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10011 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8808), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8537), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8538), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8539), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8540), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8541), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8542), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10018 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8543), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10019 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8544), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8545), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n5015), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8546), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8547), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8548), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8549), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10026 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8550), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n4483), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8551), .S(P2_U3966), .Z(
        P2_U3552) );
  NOR2_X1 U10029 ( .A1(n8553), .A2(n8552), .ZN(n8555) );
  NOR2_X1 U10030 ( .A1(n8555), .A2(n8554), .ZN(n8557) );
  XOR2_X1 U10031 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8578), .Z(n8556) );
  NAND2_X1 U10032 ( .A1(n8556), .A2(n8557), .ZN(n8577) );
  OAI21_X1 U10033 ( .B1(n8557), .B2(n8556), .A(n8577), .ZN(n8558) );
  NAND2_X1 U10034 ( .A1(n8558), .A2(n9929), .ZN(n8571) );
  AOI21_X1 U10035 ( .B1(n9932), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8559), .ZN(
        n8570) );
  NOR2_X1 U10036 ( .A1(n8561), .A2(n8560), .ZN(n8563) );
  NOR2_X1 U10037 ( .A1(n8563), .A2(n8562), .ZN(n8567) );
  NAND2_X1 U10038 ( .A1(n8578), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8573) );
  INV_X1 U10039 ( .A(n8573), .ZN(n8564) );
  AOI21_X1 U10040 ( .B1(n7733), .B2(n8565), .A(n8564), .ZN(n8566) );
  NAND2_X1 U10041 ( .A1(n8566), .A2(n8567), .ZN(n8572) );
  OAI211_X1 U10042 ( .C1(n8567), .C2(n8566), .A(n9930), .B(n8572), .ZN(n8569)
         );
  NAND2_X1 U10043 ( .A1(n8611), .A2(n8578), .ZN(n8568) );
  NAND4_X1 U10044 ( .A1(n8571), .A2(n8570), .A3(n8569), .A4(n8568), .ZN(
        P2_U3261) );
  NAND2_X1 U10045 ( .A1(n8573), .A2(n8572), .ZN(n8576) );
  NAND2_X1 U10046 ( .A1(n8592), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8587) );
  INV_X1 U10047 ( .A(n8587), .ZN(n8574) );
  AOI21_X1 U10048 ( .B1(n7769), .B2(n8585), .A(n8574), .ZN(n8575) );
  NAND2_X1 U10049 ( .A1(n8575), .A2(n8576), .ZN(n8586) );
  OAI211_X1 U10050 ( .C1(n8576), .C2(n8575), .A(n9930), .B(n8586), .ZN(n8584)
         );
  OAI21_X1 U10051 ( .B1(n8578), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8577), .ZN(
        n8580) );
  XNOR2_X1 U10052 ( .A(n8592), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8579) );
  NOR2_X1 U10053 ( .A1(n8579), .A2(n8580), .ZN(n8591) );
  AOI211_X1 U10054 ( .C1(n8580), .C2(n8579), .A(n8591), .B(n9934), .ZN(n8581)
         );
  AOI211_X1 U10055 ( .C1(n9932), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8582), .B(
        n8581), .ZN(n8583) );
  OAI211_X1 U10056 ( .C1(n9933), .C2(n8585), .A(n8584), .B(n8583), .ZN(
        P2_U3262) );
  NAND2_X1 U10057 ( .A1(n8587), .A2(n8586), .ZN(n8602) );
  INV_X1 U10058 ( .A(n8590), .ZN(n8607) );
  XNOR2_X1 U10059 ( .A(n8602), .B(n8607), .ZN(n8600) );
  XNOR2_X1 U10060 ( .A(n8600), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10061 ( .A1(n8588), .A2(n9930), .ZN(n8599) );
  NOR2_X1 U10062 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10222), .ZN(n8589) );
  AOI21_X1 U10063 ( .B1(n9932), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8589), .ZN(
        n8598) );
  NAND2_X1 U10064 ( .A1(n8611), .A2(n8607), .ZN(n8597) );
  XNOR2_X1 U10065 ( .A(n8590), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8594) );
  OAI21_X1 U10066 ( .B1(n8594), .B2(n8593), .A(n8606), .ZN(n8595) );
  NAND2_X1 U10067 ( .A1(n9929), .A2(n8595), .ZN(n8596) );
  NAND4_X1 U10068 ( .A1(n8599), .A2(n8598), .A3(n8597), .A4(n8596), .ZN(
        P2_U3263) );
  INV_X1 U10069 ( .A(n8600), .ZN(n8601) );
  NAND2_X1 U10070 ( .A1(n8601), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U10071 ( .A1(n8602), .A2(n8607), .ZN(n8603) );
  NAND2_X1 U10072 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  XOR2_X1 U10073 ( .A(n8605), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8609) );
  INV_X1 U10074 ( .A(n8612), .ZN(n8608) );
  AOI22_X1 U10075 ( .A1(n8609), .A2(n9930), .B1(n8608), .B2(n9929), .ZN(n8614)
         );
  NOR2_X1 U10076 ( .A1(n8609), .A2(n9935), .ZN(n8610) );
  AOI211_X1 U10077 ( .C1(n9929), .C2(n8612), .A(n8611), .B(n8610), .ZN(n8613)
         );
  MUX2_X1 U10078 ( .A(n8614), .B(n8613), .S(n8784), .Z(n8616) );
  NAND2_X1 U10079 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8615) );
  OAI211_X1 U10080 ( .C1(n5036), .C2(n8617), .A(n8616), .B(n8615), .ZN(
        P2_U3264) );
  NAND2_X1 U10081 ( .A1(n8625), .A2(n8624), .ZN(n8623) );
  XNOR2_X1 U10082 ( .A(n8623), .B(n8834), .ZN(n8836) );
  NAND2_X1 U10083 ( .A1(n8619), .A2(n8618), .ZN(n8839) );
  NOR2_X1 U10084 ( .A1(n8788), .A2(n8839), .ZN(n8627) );
  AOI21_X1 U10085 ( .B1(n8788), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8627), .ZN(
        n8622) );
  NAND2_X1 U10086 ( .A1(n8834), .A2(n8620), .ZN(n8621) );
  OAI211_X1 U10087 ( .C1(n8836), .C2(n8629), .A(n8622), .B(n8621), .ZN(
        P2_U3265) );
  OAI21_X1 U10088 ( .B1(n8625), .B2(n8624), .A(n8623), .ZN(n8840) );
  NOR2_X1 U10089 ( .A1(n8625), .A2(n8823), .ZN(n8626) );
  AOI211_X1 U10090 ( .C1(n8788), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8627), .B(
        n8626), .ZN(n8628) );
  OAI21_X1 U10091 ( .B1(n8840), .B2(n8629), .A(n8628), .ZN(P2_U3266) );
  NOR2_X1 U10092 ( .A1(n8630), .A2(n8764), .ZN(n8633) );
  AOI211_X1 U10093 ( .C1(n4528), .C2(n8643), .A(n8759), .B(n8631), .ZN(n8632)
         );
  INV_X1 U10094 ( .A(n8650), .ZN(n8637) );
  INV_X1 U10095 ( .A(n8635), .ZN(n8636) );
  AOI21_X1 U10096 ( .B1(n8847), .B2(n8637), .A(n8636), .ZN(n8848) );
  AOI22_X1 U10097 ( .A1(n8788), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8638), .B2(
        n8800), .ZN(n8639) );
  OAI21_X1 U10098 ( .B1(n8640), .B2(n8823), .A(n8639), .ZN(n8641) );
  AOI21_X1 U10099 ( .B1(n8848), .B2(n8816), .A(n8641), .ZN(n8646) );
  OAI21_X1 U10100 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8846) );
  NAND2_X1 U10101 ( .A1(n8846), .A2(n8826), .ZN(n8645) );
  OAI211_X1 U10102 ( .C1(n8850), .C2(n8788), .A(n8646), .B(n8645), .ZN(
        P2_U3268) );
  OAI21_X1 U10103 ( .B1(n8648), .B2(n8656), .A(n8647), .ZN(n8649) );
  INV_X1 U10104 ( .A(n8649), .ZN(n8856) );
  AOI21_X1 U10105 ( .B1(n8852), .B2(n8668), .A(n8650), .ZN(n8853) );
  INV_X1 U10106 ( .A(n8852), .ZN(n8653) );
  AOI22_X1 U10107 ( .A1(n8788), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8651), .B2(
        n8800), .ZN(n8652) );
  OAI21_X1 U10108 ( .B1(n8653), .B2(n8823), .A(n8652), .ZN(n8662) );
  AOI211_X1 U10109 ( .C1(n8656), .C2(n8655), .A(n8759), .B(n8654), .ZN(n8660)
         );
  OAI22_X1 U10110 ( .A1(n8658), .A2(n8762), .B1(n8657), .B2(n8764), .ZN(n8659)
         );
  NOR2_X1 U10111 ( .A1(n8660), .A2(n8659), .ZN(n8855) );
  NOR2_X1 U10112 ( .A1(n8855), .A2(n8788), .ZN(n8661) );
  AOI211_X1 U10113 ( .C1(n8853), .C2(n8816), .A(n8662), .B(n8661), .ZN(n8663)
         );
  OAI21_X1 U10114 ( .B1(n8856), .B2(n8818), .A(n8663), .ZN(P2_U3269) );
  OAI21_X1 U10115 ( .B1(n8666), .B2(n8665), .A(n8664), .ZN(n8667) );
  INV_X1 U10116 ( .A(n8667), .ZN(n8861) );
  INV_X1 U10117 ( .A(n8668), .ZN(n8669) );
  AOI211_X1 U10118 ( .C1(n8858), .C2(n4899), .A(n10024), .B(n8669), .ZN(n8857)
         );
  AOI22_X1 U10119 ( .A1(n8788), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8670), .B2(
        n8800), .ZN(n8671) );
  OAI21_X1 U10120 ( .B1(n8672), .B2(n8823), .A(n8671), .ZN(n8680) );
  AND2_X1 U10121 ( .A1(n8686), .A2(n8673), .ZN(n8676) );
  OAI21_X1 U10122 ( .B1(n8676), .B2(n8675), .A(n8674), .ZN(n8678) );
  AOI21_X1 U10123 ( .B1(n8678), .B2(n8804), .A(n8677), .ZN(n8860) );
  NOR2_X1 U10124 ( .A1(n8860), .A2(n8788), .ZN(n8679) );
  AOI211_X1 U10125 ( .C1(n8857), .C2(n8829), .A(n8680), .B(n8679), .ZN(n8681)
         );
  OAI21_X1 U10126 ( .B1(n8861), .B2(n8818), .A(n8681), .ZN(P2_U3270) );
  OAI21_X1 U10127 ( .B1(n8684), .B2(n8683), .A(n8682), .ZN(n8685) );
  INV_X1 U10128 ( .A(n8685), .ZN(n8866) );
  OAI211_X1 U10129 ( .C1(n8688), .C2(n8687), .A(n8686), .B(n8804), .ZN(n8691)
         );
  INV_X1 U10130 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U10131 ( .A1(n8691), .A2(n8690), .ZN(n8862) );
  AOI211_X1 U10132 ( .C1(n8864), .C2(n8699), .A(n10024), .B(n4896), .ZN(n8863)
         );
  NAND2_X1 U10133 ( .A1(n8863), .A2(n8829), .ZN(n8694) );
  AOI22_X1 U10134 ( .A1(n8788), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8692), .B2(
        n8800), .ZN(n8693) );
  OAI211_X1 U10135 ( .C1(n4897), .C2(n8823), .A(n8694), .B(n8693), .ZN(n8695)
         );
  AOI21_X1 U10136 ( .B1(n8862), .B2(n8696), .A(n8695), .ZN(n8697) );
  OAI21_X1 U10137 ( .B1(n8866), .B2(n8818), .A(n8697), .ZN(P2_U3271) );
  XOR2_X1 U10138 ( .A(n8698), .B(n8705), .Z(n8871) );
  INV_X1 U10139 ( .A(n8699), .ZN(n8700) );
  AOI21_X1 U10140 ( .B1(n8867), .B2(n8715), .A(n8700), .ZN(n8868) );
  INV_X1 U10141 ( .A(n8867), .ZN(n8703) );
  AOI22_X1 U10142 ( .A1(n8788), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8701), .B2(
        n8800), .ZN(n8702) );
  OAI21_X1 U10143 ( .B1(n8703), .B2(n8823), .A(n8702), .ZN(n8711) );
  OAI211_X1 U10144 ( .C1(n8706), .C2(n8705), .A(n8704), .B(n8804), .ZN(n8709)
         );
  AOI22_X1 U10145 ( .A1(n5012), .A2(n8809), .B1(n8810), .B2(n8707), .ZN(n8708)
         );
  NOR2_X1 U10146 ( .A1(n8870), .A2(n8788), .ZN(n8710) );
  AOI211_X1 U10147 ( .C1(n8868), .C2(n8816), .A(n8711), .B(n8710), .ZN(n8712)
         );
  OAI21_X1 U10148 ( .B1(n8818), .B2(n8871), .A(n8712), .ZN(P2_U3272) );
  OAI21_X1 U10149 ( .B1(n8714), .B2(n8720), .A(n8713), .ZN(n8876) );
  INV_X1 U10150 ( .A(n8728), .ZN(n8717) );
  INV_X1 U10151 ( .A(n8715), .ZN(n8716) );
  AOI21_X1 U10152 ( .B1(n8872), .B2(n8717), .A(n8716), .ZN(n8873) );
  AOI22_X1 U10153 ( .A1(n8788), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8718), .B2(
        n8800), .ZN(n8719) );
  OAI21_X1 U10154 ( .B1(n5009), .B2(n8823), .A(n8719), .ZN(n8726) );
  OAI21_X1 U10155 ( .B1(n8733), .B2(n8721), .A(n8720), .ZN(n8722) );
  NAND2_X1 U10156 ( .A1(n4541), .A2(n8722), .ZN(n8724) );
  AOI222_X1 U10157 ( .A1(n8804), .A2(n8724), .B1(n8752), .B2(n8809), .C1(n8723), .C2(n8810), .ZN(n8875) );
  NOR2_X1 U10158 ( .A1(n8875), .A2(n8788), .ZN(n8725) );
  AOI211_X1 U10159 ( .C1(n8873), .C2(n8816), .A(n8726), .B(n8725), .ZN(n8727)
         );
  OAI21_X1 U10160 ( .B1(n8818), .B2(n8876), .A(n8727), .ZN(P2_U3273) );
  XOR2_X1 U10161 ( .A(n8734), .B(n4510), .Z(n8881) );
  INV_X1 U10162 ( .A(n8743), .ZN(n8729) );
  AOI21_X1 U10163 ( .B1(n8877), .B2(n8729), .A(n8728), .ZN(n8878) );
  AOI22_X1 U10164 ( .A1(n8788), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8730), .B2(
        n8800), .ZN(n8731) );
  OAI21_X1 U10165 ( .B1(n8732), .B2(n8823), .A(n8731), .ZN(n8740) );
  AOI211_X1 U10166 ( .C1(n8735), .C2(n8734), .A(n8759), .B(n8733), .ZN(n8738)
         );
  OAI22_X1 U10167 ( .A1(n8763), .A2(n8764), .B1(n8736), .B2(n8762), .ZN(n8737)
         );
  NOR2_X1 U10168 ( .A1(n8738), .A2(n8737), .ZN(n8880) );
  NOR2_X1 U10169 ( .A1(n8880), .A2(n8788), .ZN(n8739) );
  AOI211_X1 U10170 ( .C1(n8878), .C2(n8816), .A(n8740), .B(n8739), .ZN(n8741)
         );
  OAI21_X1 U10171 ( .B1(n8818), .B2(n8881), .A(n8741), .ZN(P2_U3274) );
  XNOR2_X1 U10172 ( .A(n8742), .B(n8749), .ZN(n8886) );
  INV_X1 U10173 ( .A(n8768), .ZN(n8744) );
  AOI21_X1 U10174 ( .B1(n8882), .B2(n8744), .A(n8743), .ZN(n8883) );
  AOI22_X1 U10175 ( .A1(n8788), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8745), .B2(
        n8800), .ZN(n8746) );
  OAI21_X1 U10176 ( .B1(n8747), .B2(n8823), .A(n8746), .ZN(n8755) );
  OAI21_X1 U10177 ( .B1(n8750), .B2(n8749), .A(n8748), .ZN(n8753) );
  AOI222_X1 U10178 ( .A1(n8804), .A2(n8753), .B1(n8752), .B2(n8810), .C1(n8751), .C2(n8809), .ZN(n8885) );
  NOR2_X1 U10179 ( .A1(n8885), .A2(n8788), .ZN(n8754) );
  AOI211_X1 U10180 ( .C1(n8883), .C2(n8816), .A(n8755), .B(n8754), .ZN(n8756)
         );
  OAI21_X1 U10181 ( .B1(n8886), .B2(n8818), .A(n8756), .ZN(P2_U3275) );
  INV_X1 U10182 ( .A(n8781), .ZN(n8758) );
  AOI21_X1 U10183 ( .B1(n8758), .B2(n8757), .A(n4482), .ZN(n8760) );
  NOR3_X1 U10184 ( .A1(n8761), .A2(n8760), .A3(n8759), .ZN(n8767) );
  OAI22_X1 U10185 ( .A1(n8765), .A2(n8764), .B1(n8763), .B2(n8762), .ZN(n8766)
         );
  NOR2_X1 U10186 ( .A1(n8767), .A2(n8766), .ZN(n8891) );
  AOI21_X1 U10187 ( .B1(n8888), .B2(n8777), .A(n8768), .ZN(n8889) );
  AOI22_X1 U10188 ( .A1(n8788), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8769), .B2(
        n8800), .ZN(n8770) );
  OAI21_X1 U10189 ( .B1(n4673), .B2(n8823), .A(n8770), .ZN(n8771) );
  AOI21_X1 U10190 ( .B1(n8889), .B2(n8816), .A(n8771), .ZN(n8774) );
  NAND2_X1 U10191 ( .A1(n8772), .A2(n4482), .ZN(n8887) );
  NAND3_X1 U10192 ( .A1(n4641), .A2(n8826), .A3(n8887), .ZN(n8773) );
  OAI211_X1 U10193 ( .C1(n8891), .C2(n8788), .A(n8774), .B(n8773), .ZN(
        P2_U3276) );
  XNOR2_X1 U10194 ( .A(n8775), .B(n8778), .ZN(n8894) );
  INV_X1 U10195 ( .A(n8897), .ZN(n8790) );
  INV_X1 U10196 ( .A(n8776), .ZN(n8797) );
  OAI211_X1 U10197 ( .C1(n8790), .C2(n8797), .A(n10014), .B(n8777), .ZN(n8895)
         );
  AOI21_X1 U10198 ( .B1(n8805), .B2(n8779), .A(n8778), .ZN(n8780) );
  OR2_X1 U10199 ( .A1(n8781), .A2(n8780), .ZN(n8783) );
  AOI21_X1 U10200 ( .B1(n8783), .B2(n8804), .A(n8782), .ZN(n8899) );
  OAI21_X1 U10201 ( .B1(n8784), .B2(n8895), .A(n8899), .ZN(n8785) );
  AOI21_X1 U10202 ( .B1(n8786), .B2(n8894), .A(n8785), .ZN(n8794) );
  AOI22_X1 U10203 ( .A1(n8788), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8787), .B2(
        n8800), .ZN(n8789) );
  OAI21_X1 U10204 ( .B1(n8790), .B2(n8823), .A(n8789), .ZN(n8791) );
  AOI21_X1 U10205 ( .B1(n8894), .B2(n8792), .A(n8791), .ZN(n8793) );
  OAI21_X1 U10206 ( .B1(n8794), .B2(n8788), .A(n8793), .ZN(P2_U3277) );
  XNOR2_X1 U10207 ( .A(n8795), .B(n8806), .ZN(n8905) );
  INV_X1 U10208 ( .A(n8796), .ZN(n8798) );
  AOI21_X1 U10209 ( .B1(n8901), .B2(n8798), .A(n8797), .ZN(n8902) );
  INV_X1 U10210 ( .A(n8799), .ZN(n8801) );
  AOI22_X1 U10211 ( .A1(n8788), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8801), .B2(
        n8800), .ZN(n8802) );
  OAI21_X1 U10212 ( .B1(n8803), .B2(n8823), .A(n8802), .ZN(n8815) );
  OAI211_X1 U10213 ( .C1(n8807), .C2(n8806), .A(n8805), .B(n8804), .ZN(n8813)
         );
  AOI22_X1 U10214 ( .A1(n8811), .A2(n8810), .B1(n8809), .B2(n8808), .ZN(n8812)
         );
  NOR2_X1 U10215 ( .A1(n8904), .A2(n8788), .ZN(n8814) );
  AOI211_X1 U10216 ( .C1(n8902), .C2(n8816), .A(n8815), .B(n8814), .ZN(n8817)
         );
  OAI21_X1 U10217 ( .B1(n8905), .B2(n8818), .A(n8817), .ZN(P2_U3278) );
  MUX2_X1 U10218 ( .A(n8819), .B(n6725), .S(n8788), .Z(n8833) );
  OAI22_X1 U10219 ( .A1(n8823), .A2(n8822), .B1(n8821), .B2(n8820), .ZN(n8824)
         );
  INV_X1 U10220 ( .A(n8824), .ZN(n8832) );
  NAND2_X1 U10221 ( .A1(n8826), .A2(n8825), .ZN(n8831) );
  INV_X1 U10222 ( .A(n8827), .ZN(n8828) );
  NAND2_X1 U10223 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  NAND4_X1 U10224 ( .A1(n8833), .A2(n8832), .A3(n8831), .A4(n8830), .ZN(
        P2_U3291) );
  NAND2_X1 U10225 ( .A1(n8834), .A2(n10013), .ZN(n8835) );
  OAI211_X1 U10226 ( .C1(n8836), .C2(n10024), .A(n8839), .B(n8835), .ZN(n8917)
         );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8917), .S(n10052), .Z(
        P2_U3551) );
  NAND2_X1 U10228 ( .A1(n8837), .A2(n10013), .ZN(n8838) );
  OAI211_X1 U10229 ( .C1(n8840), .C2(n10024), .A(n8839), .B(n8838), .ZN(n8918)
         );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8918), .S(n10052), .Z(
        P2_U3550) );
  AOI22_X1 U10231 ( .A1(n8842), .A2(n10014), .B1(n10013), .B2(n8841), .ZN(
        n8843) );
  INV_X1 U10232 ( .A(n8846), .ZN(n8851) );
  AOI22_X1 U10233 ( .A1(n8848), .A2(n10014), .B1(n10013), .B2(n8847), .ZN(
        n8849) );
  OAI211_X1 U10234 ( .C1(n10019), .C2(n8851), .A(n8850), .B(n8849), .ZN(n8919)
         );
  MUX2_X1 U10235 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8919), .S(n10052), .Z(
        P2_U3548) );
  AOI22_X1 U10236 ( .A1(n8853), .A2(n10014), .B1(n10013), .B2(n8852), .ZN(
        n8854) );
  OAI211_X1 U10237 ( .C1(n8856), .C2(n10019), .A(n8855), .B(n8854), .ZN(n8920)
         );
  MUX2_X1 U10238 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8920), .S(n10052), .Z(
        P2_U3547) );
  AOI21_X1 U10239 ( .B1(n10013), .B2(n8858), .A(n8857), .ZN(n8859) );
  OAI211_X1 U10240 ( .C1(n8861), .C2(n10019), .A(n8860), .B(n8859), .ZN(n8921)
         );
  MUX2_X1 U10241 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8921), .S(n10052), .Z(
        P2_U3546) );
  AOI211_X1 U10242 ( .C1(n10013), .C2(n8864), .A(n8863), .B(n8862), .ZN(n8865)
         );
  OAI21_X1 U10243 ( .B1(n8866), .B2(n10019), .A(n8865), .ZN(n8922) );
  MUX2_X1 U10244 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8922), .S(n10052), .Z(
        P2_U3545) );
  AOI22_X1 U10245 ( .A1(n8868), .A2(n10014), .B1(n10013), .B2(n8867), .ZN(
        n8869) );
  OAI211_X1 U10246 ( .C1(n8871), .C2(n10019), .A(n8870), .B(n8869), .ZN(n8923)
         );
  MUX2_X1 U10247 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8923), .S(n10052), .Z(
        P2_U3544) );
  AOI22_X1 U10248 ( .A1(n8873), .A2(n10014), .B1(n10013), .B2(n8872), .ZN(
        n8874) );
  OAI211_X1 U10249 ( .C1(n10019), .C2(n8876), .A(n8875), .B(n8874), .ZN(n8924)
         );
  MUX2_X1 U10250 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8924), .S(n10052), .Z(
        P2_U3543) );
  AOI22_X1 U10251 ( .A1(n8878), .A2(n10014), .B1(n10013), .B2(n8877), .ZN(
        n8879) );
  OAI211_X1 U10252 ( .C1(n8881), .C2(n10019), .A(n8880), .B(n8879), .ZN(n8925)
         );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8925), .S(n10052), .Z(
        P2_U3542) );
  AOI22_X1 U10254 ( .A1(n8883), .A2(n10014), .B1(n10013), .B2(n8882), .ZN(
        n8884) );
  OAI211_X1 U10255 ( .C1(n10019), .C2(n8886), .A(n8885), .B(n8884), .ZN(n8926)
         );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8926), .S(n10052), .Z(
        P2_U3541) );
  NAND2_X1 U10257 ( .A1(n8887), .A2(n10029), .ZN(n8892) );
  AOI22_X1 U10258 ( .A1(n8889), .A2(n10014), .B1(n10013), .B2(n8888), .ZN(
        n8890) );
  OAI211_X1 U10259 ( .C1(n8893), .C2(n8892), .A(n8891), .B(n8890), .ZN(n8927)
         );
  MUX2_X1 U10260 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8927), .S(n10052), .Z(
        P2_U3540) );
  INV_X1 U10261 ( .A(n8894), .ZN(n8900) );
  INV_X1 U10262 ( .A(n8895), .ZN(n8896) );
  AOI21_X1 U10263 ( .B1(n10013), .B2(n8897), .A(n8896), .ZN(n8898) );
  OAI211_X1 U10264 ( .C1(n8900), .C2(n10019), .A(n8899), .B(n8898), .ZN(n8928)
         );
  MUX2_X1 U10265 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8928), .S(n10052), .Z(
        P2_U3539) );
  AOI22_X1 U10266 ( .A1(n8902), .A2(n10014), .B1(n10013), .B2(n8901), .ZN(
        n8903) );
  OAI211_X1 U10267 ( .C1(n8905), .C2(n10019), .A(n8904), .B(n8903), .ZN(n8929)
         );
  MUX2_X1 U10268 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8929), .S(n10052), .Z(
        P2_U3538) );
  AOI21_X1 U10269 ( .B1(n10013), .B2(n8907), .A(n8906), .ZN(n8908) );
  OAI211_X1 U10270 ( .C1(n8910), .C2(n10019), .A(n8909), .B(n8908), .ZN(n8930)
         );
  MUX2_X1 U10271 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8930), .S(n10052), .Z(
        P2_U3537) );
  INV_X1 U10272 ( .A(n8911), .ZN(n8916) );
  AOI22_X1 U10273 ( .A1(n8913), .A2(n10014), .B1(n10013), .B2(n8912), .ZN(
        n8914) );
  OAI211_X1 U10274 ( .C1(n9576), .C2(n8916), .A(n8915), .B(n8914), .ZN(n8931)
         );
  MUX2_X1 U10275 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8931), .S(n10052), .Z(
        P2_U3536) );
  MUX2_X1 U10276 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8917), .S(n10032), .Z(
        P2_U3519) );
  MUX2_X1 U10277 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8918), .S(n10032), .Z(
        P2_U3518) );
  MUX2_X1 U10278 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8919), .S(n10032), .Z(
        P2_U3516) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8920), .S(n10032), .Z(
        P2_U3515) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8921), .S(n10032), .Z(
        P2_U3514) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8922), .S(n10032), .Z(
        P2_U3513) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8923), .S(n10032), .Z(
        P2_U3512) );
  MUX2_X1 U10283 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8924), .S(n10032), .Z(
        P2_U3511) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8925), .S(n10032), .Z(
        P2_U3510) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8926), .S(n10032), .Z(
        P2_U3509) );
  MUX2_X1 U10286 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8927), .S(n10032), .Z(
        P2_U3508) );
  MUX2_X1 U10287 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8928), .S(n10032), .Z(
        P2_U3507) );
  MUX2_X1 U10288 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8929), .S(n10032), .Z(
        P2_U3505) );
  MUX2_X1 U10289 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8930), .S(n10032), .Z(
        P2_U3502) );
  MUX2_X1 U10290 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8931), .S(n10032), .Z(
        P2_U3499) );
  INV_X1 U10291 ( .A(n8194), .ZN(n9537) );
  NOR4_X1 U10292 ( .A1(n8932), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5771), .A4(
        P2_U3152), .ZN(n8933) );
  AOI21_X1 U10293 ( .B1(n8947), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8933), .ZN(
        n8934) );
  OAI21_X1 U10294 ( .B1(n9537), .B2(n8944), .A(n8934), .ZN(P2_U3327) );
  INV_X1 U10295 ( .A(n8935), .ZN(n9540) );
  AOI22_X1 U10296 ( .A1(n8936), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8947), .ZN(n8937) );
  OAI21_X1 U10297 ( .B1(n9540), .B2(n8944), .A(n8937), .ZN(P2_U3328) );
  AOI22_X1 U10298 ( .A1(n8938), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8947), .ZN(n8939) );
  OAI21_X1 U10299 ( .B1(n8940), .B2(n8944), .A(n8939), .ZN(P2_U3329) );
  INV_X1 U10300 ( .A(n8941), .ZN(n9544) );
  AOI22_X1 U10301 ( .A1(n8942), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n8947), .ZN(n8943) );
  OAI21_X1 U10302 ( .B1(n9544), .B2(n8944), .A(n8943), .ZN(P2_U3330) );
  INV_X1 U10303 ( .A(n8945), .ZN(n9549) );
  AOI21_X1 U10304 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8947), .A(n8946), .ZN(
        n8948) );
  OAI21_X1 U10305 ( .B1(n9549), .B2(n8949), .A(n8948), .ZN(P2_U3331) );
  MUX2_X1 U10306 ( .A(n8950), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10307 ( .A(n8952), .B(n8951), .ZN(n8953) );
  XNOR2_X1 U10308 ( .A(n8954), .B(n8953), .ZN(n8964) );
  INV_X1 U10309 ( .A(n8955), .ZN(n8956) );
  AOI21_X1 U10310 ( .B1(n9074), .B2(n9089), .A(n8956), .ZN(n8959) );
  NAND2_X1 U10311 ( .A1(n9076), .A2(n8957), .ZN(n8958) );
  OAI211_X1 U10312 ( .C1(n8960), .C2(n9079), .A(n8959), .B(n8958), .ZN(n8961)
         );
  AOI21_X1 U10313 ( .B1(n8962), .B2(n9082), .A(n8961), .ZN(n8963) );
  OAI21_X1 U10314 ( .B1(n8964), .B2(n9085), .A(n8963), .ZN(P1_U3213) );
  AOI21_X1 U10315 ( .B1(n8968), .B2(n8966), .A(n8965), .ZN(n8967) );
  AOI21_X1 U10316 ( .B1(n4519), .B2(n8968), .A(n8967), .ZN(n8973) );
  INV_X1 U10317 ( .A(n9076), .ZN(n9052) );
  NAND2_X1 U10318 ( .A1(n9242), .A2(n9064), .ZN(n8970) );
  AOI22_X1 U10319 ( .A1(n9421), .A2(n9074), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8969) );
  OAI211_X1 U10320 ( .C1(n9052), .C2(n9247), .A(n8970), .B(n8969), .ZN(n8971)
         );
  AOI21_X1 U10321 ( .B1(n9409), .B2(n9082), .A(n8971), .ZN(n8972) );
  OAI21_X1 U10322 ( .B1(n8973), .B2(n9085), .A(n8972), .ZN(P1_U3214) );
  XOR2_X1 U10323 ( .A(n8975), .B(n8974), .Z(n8980) );
  AOI22_X1 U10324 ( .A1(n9074), .A2(n9435), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n8977) );
  NAND2_X1 U10325 ( .A1(n9076), .A2(n9306), .ZN(n8976) );
  OAI211_X1 U10326 ( .C1(n9309), .C2(n9079), .A(n8977), .B(n8976), .ZN(n8978)
         );
  AOI21_X1 U10327 ( .B1(n9434), .B2(n9082), .A(n8978), .ZN(n8979) );
  OAI21_X1 U10328 ( .B1(n8980), .B2(n9085), .A(n8979), .ZN(P1_U3217) );
  XOR2_X1 U10329 ( .A(n8982), .B(n8981), .Z(n8988) );
  OAI22_X1 U10330 ( .A1(n9309), .A2(n9062), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8983), .ZN(n8984) );
  AOI21_X1 U10331 ( .B1(n9064), .B2(n9421), .A(n8984), .ZN(n8985) );
  OAI21_X1 U10332 ( .B1(n9052), .B2(n9276), .A(n8985), .ZN(n8986) );
  AOI21_X1 U10333 ( .B1(n9284), .B2(n9082), .A(n8986), .ZN(n8987) );
  OAI21_X1 U10334 ( .B1(n8988), .B2(n9085), .A(n8987), .ZN(P1_U3221) );
  XOR2_X1 U10335 ( .A(n8990), .B(n8989), .Z(n8998) );
  OAI22_X1 U10336 ( .A1(n8992), .A2(n9062), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8991), .ZN(n8993) );
  AOI21_X1 U10337 ( .B1(n9211), .B2(n9076), .A(n8993), .ZN(n8994) );
  OAI21_X1 U10338 ( .B1(n8995), .B2(n9079), .A(n8994), .ZN(n8996) );
  AOI21_X1 U10339 ( .B1(n9394), .B2(n9082), .A(n8996), .ZN(n8997) );
  OAI21_X1 U10340 ( .B1(n8998), .B2(n9085), .A(n8997), .ZN(P1_U3223) );
  INV_X1 U10341 ( .A(n8999), .ZN(n9003) );
  OAI21_X1 U10342 ( .B1(n9001), .B2(n9003), .A(n9000), .ZN(n9002) );
  OAI21_X1 U10343 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9005) );
  NAND2_X1 U10344 ( .A1(n9005), .A2(n9056), .ZN(n9011) );
  INV_X1 U10345 ( .A(n9006), .ZN(n9007) );
  AOI21_X1 U10346 ( .B1(n9074), .B2(n9458), .A(n9007), .ZN(n9008) );
  OAI21_X1 U10347 ( .B1(n9356), .B2(n9079), .A(n9008), .ZN(n9009) );
  AOI21_X1 U10348 ( .B1(n9351), .B2(n9076), .A(n9009), .ZN(n9010) );
  OAI211_X1 U10349 ( .C1(n4706), .C2(n9067), .A(n9011), .B(n9010), .ZN(
        P1_U3224) );
  OAI21_X1 U10350 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9015) );
  NAND2_X1 U10351 ( .A1(n9015), .A2(n9056), .ZN(n9020) );
  OAI22_X1 U10352 ( .A1(n9062), .A2(n9080), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9016), .ZN(n9018) );
  NOR2_X1 U10353 ( .A1(n9052), .A2(n9334), .ZN(n9017) );
  AOI211_X1 U10354 ( .C1(n9064), .C2(n9435), .A(n9018), .B(n9017), .ZN(n9019)
         );
  OAI211_X1 U10355 ( .C1(n9338), .C2(n9067), .A(n9020), .B(n9019), .ZN(
        P1_U3226) );
  OAI21_X1 U10356 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(n9024) );
  NAND2_X1 U10357 ( .A1(n9024), .A2(n9056), .ZN(n9028) );
  AOI22_X1 U10358 ( .A1(n9413), .A2(n9074), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9025) );
  OAI21_X1 U10359 ( .B1(n9052), .B2(n9229), .A(n9025), .ZN(n9026) );
  AOI21_X1 U10360 ( .B1(n9196), .B2(n9064), .A(n9026), .ZN(n9027) );
  OAI211_X1 U10361 ( .C1(n9499), .C2(n9067), .A(n9028), .B(n9027), .ZN(
        P1_U3227) );
  XOR2_X1 U10362 ( .A(n9030), .B(n9029), .Z(n9035) );
  NAND2_X1 U10363 ( .A1(n9412), .A2(n9064), .ZN(n9032) );
  AOI22_X1 U10364 ( .A1(n9074), .A2(n9444), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9031) );
  OAI211_X1 U10365 ( .C1(n9052), .C2(n9296), .A(n9032), .B(n9031), .ZN(n9033)
         );
  AOI21_X1 U10366 ( .B1(n9295), .B2(n9082), .A(n9033), .ZN(n9034) );
  OAI21_X1 U10367 ( .B1(n9035), .B2(n9085), .A(n9034), .ZN(P1_U3231) );
  NAND2_X1 U10368 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  XOR2_X1 U10369 ( .A(n9039), .B(n9038), .Z(n9045) );
  OAI22_X1 U10370 ( .A1(n9293), .A2(n9062), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9040), .ZN(n9041) );
  AOI21_X1 U10371 ( .B1(n9413), .B2(n9064), .A(n9041), .ZN(n9042) );
  OAI21_X1 U10372 ( .B1(n9052), .B2(n9259), .A(n9042), .ZN(n9043) );
  AOI21_X1 U10373 ( .B1(n9267), .B2(n9082), .A(n9043), .ZN(n9044) );
  OAI21_X1 U10374 ( .B1(n9045), .B2(n9085), .A(n9044), .ZN(P1_U3233) );
  XNOR2_X1 U10375 ( .A(n9047), .B(n9046), .ZN(n9048) );
  XNOR2_X1 U10376 ( .A(n9049), .B(n9048), .ZN(n9055) );
  NAND2_X1 U10377 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9736) );
  OAI21_X1 U10378 ( .B1(n9062), .B2(n9356), .A(n9736), .ZN(n9050) );
  AOI21_X1 U10379 ( .B1(n9064), .B2(n9444), .A(n9050), .ZN(n9051) );
  OAI21_X1 U10380 ( .B1(n9052), .B2(n9319), .A(n9051), .ZN(n9053) );
  AOI21_X1 U10381 ( .B1(n9329), .B2(n9082), .A(n9053), .ZN(n9054) );
  OAI21_X1 U10382 ( .B1(n9055), .B2(n9085), .A(n9054), .ZN(P1_U3236) );
  OAI211_X1 U10383 ( .C1(n9059), .C2(n9058), .A(n9057), .B(n9056), .ZN(n9066)
         );
  INV_X1 U10384 ( .A(n9060), .ZN(n9202) );
  AOI22_X1 U10385 ( .A1(n9202), .A2(n9076), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9061) );
  OAI21_X1 U10386 ( .B1(n9398), .B2(n9062), .A(n9061), .ZN(n9063) );
  AOI21_X1 U10387 ( .B1(n9164), .B2(n9064), .A(n9063), .ZN(n9065) );
  OAI211_X1 U10388 ( .C1(n9494), .C2(n9067), .A(n9066), .B(n9065), .ZN(
        P1_U3238) );
  NAND2_X1 U10389 ( .A1(n9069), .A2(n9068), .ZN(n9070) );
  XOR2_X1 U10390 ( .A(n9071), .B(n9070), .Z(n9086) );
  INV_X1 U10391 ( .A(n9072), .ZN(n9073) );
  AOI21_X1 U10392 ( .B1(n9074), .B2(n9605), .A(n9073), .ZN(n9078) );
  NAND2_X1 U10393 ( .A1(n9076), .A2(n9075), .ZN(n9077) );
  OAI211_X1 U10394 ( .C1(n9080), .C2(n9079), .A(n9078), .B(n9077), .ZN(n9081)
         );
  AOI21_X1 U10395 ( .B1(n9083), .B2(n9082), .A(n9081), .ZN(n9084) );
  OAI21_X1 U10396 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(P1_U3239) );
  MUX2_X1 U10397 ( .A(n9087), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9095), .Z(
        P1_U3585) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9163), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10399 ( .A(n9088), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9095), .Z(
        P1_U3583) );
  MUX2_X1 U10400 ( .A(n9216), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9095), .Z(
        P1_U3581) );
  MUX2_X1 U10401 ( .A(n9196), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9095), .Z(
        P1_U3580) );
  MUX2_X1 U10402 ( .A(n9242), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9095), .Z(
        P1_U3579) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9421), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10404 ( .A(n9412), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9095), .Z(
        P1_U3576) );
  MUX2_X1 U10405 ( .A(n9436), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9095), .Z(
        P1_U3575) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9444), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9435), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10408 ( .A(n9459), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9095), .Z(
        P1_U3572) );
  MUX2_X1 U10409 ( .A(n9341), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9095), .Z(
        P1_U3571) );
  MUX2_X1 U10410 ( .A(n9458), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9095), .Z(
        P1_U3570) );
  MUX2_X1 U10411 ( .A(n9605), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9095), .Z(
        P1_U3569) );
  MUX2_X1 U10412 ( .A(n9089), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9095), .Z(
        P1_U3568) );
  MUX2_X1 U10413 ( .A(n9606), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9095), .Z(
        P1_U3567) );
  MUX2_X1 U10414 ( .A(n9090), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9095), .Z(
        P1_U3566) );
  MUX2_X1 U10415 ( .A(n9091), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9095), .Z(
        P1_U3565) );
  MUX2_X1 U10416 ( .A(n9092), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9095), .Z(
        P1_U3564) );
  MUX2_X1 U10417 ( .A(n9093), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9095), .Z(
        P1_U3563) );
  MUX2_X1 U10418 ( .A(n9864), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9095), .Z(
        P1_U3562) );
  MUX2_X1 U10419 ( .A(n9782), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9095), .Z(
        P1_U3561) );
  MUX2_X1 U10420 ( .A(n9865), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9095), .Z(
        P1_U3560) );
  MUX2_X1 U10421 ( .A(n9781), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9095), .Z(
        P1_U3559) );
  MUX2_X1 U10422 ( .A(n9094), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9095), .Z(
        P1_U3558) );
  MUX2_X1 U10423 ( .A(n6602), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9095), .Z(
        P1_U3557) );
  MUX2_X1 U10424 ( .A(n9096), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9095), .Z(
        P1_U3556) );
  MUX2_X1 U10425 ( .A(n9804), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9095), .Z(
        P1_U3555) );
  NAND2_X1 U10426 ( .A1(n9134), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n9107) );
  NAND3_X1 U10427 ( .A1(n9744), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6283), .ZN(
        n9106) );
  INV_X1 U10428 ( .A(n9097), .ZN(n9103) );
  NOR2_X1 U10429 ( .A1(n9098), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9099) );
  NOR2_X1 U10430 ( .A1(n9100), .A2(n9099), .ZN(n9101) );
  MUX2_X1 U10431 ( .A(n9101), .B(n9100), .S(P1_IR_REG_0__SCAN_IN), .Z(n9102)
         );
  NAND3_X1 U10432 ( .A1(n9103), .A2(P1_STATE_REG_SCAN_IN), .A3(n9102), .ZN(
        n9105) );
  NAND2_X1 U10433 ( .A1(P1_U3084), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9104) );
  NAND4_X1 U10434 ( .A1(n9107), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(
        P1_U3241) );
  OAI21_X1 U10435 ( .B1(n9110), .B2(n9109), .A(n9108), .ZN(n9111) );
  AOI22_X1 U10436 ( .A1(n9111), .A2(n9744), .B1(n9134), .B2(
        P1_ADDR_REG_7__SCAN_IN), .ZN(n9120) );
  AOI21_X1 U10437 ( .B1(n9708), .B2(n9113), .A(n9112), .ZN(n9119) );
  OAI21_X1 U10438 ( .B1(n9116), .B2(n9115), .A(n9114), .ZN(n9117) );
  NAND2_X1 U10439 ( .A1(n9117), .A2(n9735), .ZN(n9118) );
  NAND3_X1 U10440 ( .A1(n9120), .A2(n9119), .A3(n9118), .ZN(P1_U3248) );
  INV_X1 U10441 ( .A(n9121), .ZN(n9128) );
  NAND2_X1 U10442 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9127) );
  AOI21_X1 U10443 ( .B1(n9124), .B2(n9123), .A(n9122), .ZN(n9125) );
  NAND2_X1 U10444 ( .A1(n9744), .A2(n9125), .ZN(n9126) );
  OAI211_X1 U10445 ( .C1(n9739), .C2(n9128), .A(n9127), .B(n9126), .ZN(n9133)
         );
  AOI211_X1 U10446 ( .C1(n9131), .C2(n9130), .A(n9129), .B(n9715), .ZN(n9132)
         );
  AOI211_X1 U10447 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9134), .A(n9133), .B(
        n9132), .ZN(n9135) );
  INV_X1 U10448 ( .A(n9135), .ZN(P1_U3258) );
  XNOR2_X1 U10449 ( .A(n9482), .B(n9137), .ZN(n9138) );
  NAND2_X1 U10450 ( .A1(n9138), .A2(n9794), .ZN(n9368) );
  NAND2_X1 U10451 ( .A1(n9140), .A2(n9139), .ZN(n9371) );
  NOR2_X1 U10452 ( .A1(n9822), .A2(n9371), .ZN(n9145) );
  NOR2_X1 U10453 ( .A1(n9482), .A2(n9337), .ZN(n9141) );
  AOI211_X1 U10454 ( .C1(n9822), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9145), .B(
        n9141), .ZN(n9142) );
  OAI21_X1 U10455 ( .B1(n9368), .B2(n9361), .A(n9142), .ZN(P1_U3261) );
  XNOR2_X1 U10456 ( .A(n9486), .B(n9143), .ZN(n9144) );
  NAND2_X1 U10457 ( .A1(n9373), .A2(n9755), .ZN(n9147) );
  AOI21_X1 U10458 ( .B1(n9822), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9145), .ZN(
        n9146) );
  OAI211_X1 U10459 ( .C1(n9486), .C2(n9337), .A(n9147), .B(n9146), .ZN(
        P1_U3262) );
  INV_X1 U10460 ( .A(n9148), .ZN(n9156) );
  NAND2_X1 U10461 ( .A1(n9149), .A2(n9755), .ZN(n9152) );
  AOI22_X1 U10462 ( .A1(n9150), .A2(n9787), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9822), .ZN(n9151) );
  OAI211_X1 U10463 ( .C1(n5690), .C2(n9337), .A(n9152), .B(n9151), .ZN(n9153)
         );
  AOI21_X1 U10464 ( .B1(n9154), .B2(n9816), .A(n9153), .ZN(n9155) );
  OAI21_X1 U10465 ( .B1(n9156), .B2(n9818), .A(n9155), .ZN(P1_U3355) );
  AND2_X1 U10466 ( .A1(n9157), .A2(n9161), .ZN(n9158) );
  INV_X1 U10467 ( .A(n9380), .ZN(n9175) );
  OAI211_X1 U10468 ( .C1(n9162), .C2(n9161), .A(n9160), .B(n9808), .ZN(n9166)
         );
  AOI22_X1 U10469 ( .A1(n9164), .A2(n9866), .B1(n9863), .B2(n9163), .ZN(n9165)
         );
  NAND2_X1 U10470 ( .A1(n9166), .A2(n9165), .ZN(n9378) );
  AOI21_X1 U10471 ( .B1(n9167), .B2(n9183), .A(n9615), .ZN(n9169) );
  AND2_X1 U10472 ( .A1(n9169), .A2(n9168), .ZN(n9377) );
  NAND2_X1 U10473 ( .A1(n9377), .A2(n9235), .ZN(n9172) );
  AOI22_X1 U10474 ( .A1(n9170), .A2(n9787), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9822), .ZN(n9171) );
  OAI211_X1 U10475 ( .C1(n4705), .C2(n9337), .A(n9172), .B(n9171), .ZN(n9173)
         );
  AOI21_X1 U10476 ( .B1(n9378), .B2(n9816), .A(n9173), .ZN(n9174) );
  OAI21_X1 U10477 ( .B1(n9175), .B2(n9818), .A(n9174), .ZN(P1_U3263) );
  XOR2_X1 U10478 ( .A(n9178), .B(n4977), .Z(n9387) );
  OAI211_X1 U10479 ( .C1(n9179), .C2(n9178), .A(n9177), .B(n9808), .ZN(n9181)
         );
  NAND2_X1 U10480 ( .A1(n9216), .A2(n9866), .ZN(n9180) );
  OAI211_X1 U10481 ( .C1(n9182), .C2(n9888), .A(n9181), .B(n9180), .ZN(n9383)
         );
  INV_X1 U10482 ( .A(n9200), .ZN(n9185) );
  INV_X1 U10483 ( .A(n9183), .ZN(n9184) );
  AOI211_X1 U10484 ( .C1(n9385), .C2(n9185), .A(n9615), .B(n9184), .ZN(n9384)
         );
  NAND2_X1 U10485 ( .A1(n9384), .A2(n9235), .ZN(n9188) );
  AOI22_X1 U10486 ( .A1(n9186), .A2(n9787), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9822), .ZN(n9187) );
  OAI211_X1 U10487 ( .C1(n9189), .C2(n9337), .A(n9188), .B(n9187), .ZN(n9190)
         );
  AOI21_X1 U10488 ( .B1(n9383), .B2(n9816), .A(n9190), .ZN(n9191) );
  OAI21_X1 U10489 ( .B1(n9387), .B2(n9818), .A(n9191), .ZN(P1_U3264) );
  XOR2_X1 U10490 ( .A(n9192), .B(n9194), .Z(n9390) );
  INV_X1 U10491 ( .A(n9390), .ZN(n9207) );
  OAI211_X1 U10492 ( .C1(n9195), .C2(n9194), .A(n9193), .B(n9808), .ZN(n9198)
         );
  NAND2_X1 U10493 ( .A1(n9196), .A2(n9866), .ZN(n9197) );
  OAI211_X1 U10494 ( .C1(n9199), .C2(n9888), .A(n9198), .B(n9197), .ZN(n9388)
         );
  AOI211_X1 U10495 ( .C1(n9201), .C2(n9209), .A(n9615), .B(n9200), .ZN(n9389)
         );
  NAND2_X1 U10496 ( .A1(n9389), .A2(n9235), .ZN(n9204) );
  AOI22_X1 U10497 ( .A1(n9202), .A2(n9787), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9822), .ZN(n9203) );
  OAI211_X1 U10498 ( .C1(n9494), .C2(n9337), .A(n9204), .B(n9203), .ZN(n9205)
         );
  AOI21_X1 U10499 ( .B1(n9816), .B2(n9388), .A(n9205), .ZN(n9206) );
  OAI21_X1 U10500 ( .B1(n9207), .B2(n9818), .A(n9206), .ZN(P1_U3265) );
  XOR2_X1 U10501 ( .A(n9215), .B(n9208), .Z(n9397) );
  INV_X1 U10502 ( .A(n9209), .ZN(n9210) );
  AOI211_X1 U10503 ( .C1(n9394), .C2(n4714), .A(n9615), .B(n9210), .ZN(n9393)
         );
  AOI22_X1 U10504 ( .A1(n9211), .A2(n9787), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9822), .ZN(n9212) );
  OAI21_X1 U10505 ( .B1(n9213), .B2(n9337), .A(n9212), .ZN(n9219) );
  XOR2_X1 U10506 ( .A(n9215), .B(n9214), .Z(n9217) );
  AOI222_X1 U10507 ( .A1(n9808), .A2(n9217), .B1(n9216), .B2(n9863), .C1(n9242), .C2(n9866), .ZN(n9396) );
  NOR2_X1 U10508 ( .A1(n9396), .A2(n9822), .ZN(n9218) );
  AOI211_X1 U10509 ( .C1(n9393), .C2(n9755), .A(n9219), .B(n9218), .ZN(n9220)
         );
  OAI21_X1 U10510 ( .B1(n9397), .B2(n9818), .A(n9220), .ZN(P1_U3266) );
  INV_X1 U10511 ( .A(n9221), .ZN(n9222) );
  AOI21_X1 U10512 ( .B1(n9224), .B2(n9223), .A(n9222), .ZN(n9402) );
  XNOR2_X1 U10513 ( .A(n9225), .B(n9226), .ZN(n9404) );
  NAND2_X1 U10514 ( .A1(n9404), .A2(n9350), .ZN(n9237) );
  AOI211_X1 U10515 ( .C1(n9228), .C2(n9245), .A(n9615), .B(n9227), .ZN(n9399)
         );
  NOR2_X1 U10516 ( .A1(n9499), .A2(n9337), .ZN(n9234) );
  INV_X1 U10517 ( .A(n9229), .ZN(n9230) );
  AOI22_X1 U10518 ( .A1(n9230), .A2(n9787), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9822), .ZN(n9232) );
  NAND2_X1 U10519 ( .A1(n9413), .A2(n9352), .ZN(n9231) );
  OAI211_X1 U10520 ( .C1(n9398), .C2(n9355), .A(n9232), .B(n9231), .ZN(n9233)
         );
  AOI211_X1 U10521 ( .C1(n9399), .C2(n9235), .A(n9234), .B(n9233), .ZN(n9236)
         );
  OAI211_X1 U10522 ( .C1(n9402), .C2(n9367), .A(n9237), .B(n9236), .ZN(
        P1_U3267) );
  XNOR2_X1 U10523 ( .A(n9238), .B(n9240), .ZN(n9411) );
  OAI211_X1 U10524 ( .C1(n9241), .C2(n9240), .A(n9239), .B(n9808), .ZN(n9244)
         );
  AOI22_X1 U10525 ( .A1(n9242), .A2(n9863), .B1(n9866), .B2(n9421), .ZN(n9243)
         );
  NAND2_X1 U10526 ( .A1(n9244), .A2(n9243), .ZN(n9407) );
  INV_X1 U10527 ( .A(n9409), .ZN(n9251) );
  INV_X1 U10528 ( .A(n9245), .ZN(n9246) );
  AOI211_X1 U10529 ( .C1(n9409), .C2(n9264), .A(n9615), .B(n9246), .ZN(n9408)
         );
  NAND2_X1 U10530 ( .A1(n9408), .A2(n9755), .ZN(n9250) );
  INV_X1 U10531 ( .A(n9247), .ZN(n9248) );
  AOI22_X1 U10532 ( .A1(n9248), .A2(n9787), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9822), .ZN(n9249) );
  OAI211_X1 U10533 ( .C1(n9251), .C2(n9337), .A(n9250), .B(n9249), .ZN(n9252)
         );
  AOI21_X1 U10534 ( .B1(n9816), .B2(n9407), .A(n9252), .ZN(n9253) );
  OAI21_X1 U10535 ( .B1(n9411), .B2(n9818), .A(n9253), .ZN(P1_U3268) );
  NAND2_X1 U10536 ( .A1(n9271), .A2(n9254), .ZN(n9256) );
  INV_X1 U10537 ( .A(n9257), .ZN(n9255) );
  XNOR2_X1 U10538 ( .A(n9256), .B(n9255), .ZN(n9416) );
  XNOR2_X1 U10539 ( .A(n9258), .B(n9257), .ZN(n9418) );
  NAND2_X1 U10540 ( .A1(n9418), .A2(n9350), .ZN(n9269) );
  INV_X1 U10541 ( .A(n9259), .ZN(n9260) );
  AOI22_X1 U10542 ( .A1(n9822), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9260), .B2(
        n9787), .ZN(n9262) );
  NAND2_X1 U10543 ( .A1(n9412), .A2(n9352), .ZN(n9261) );
  OAI211_X1 U10544 ( .C1(n9263), .C2(n9355), .A(n9262), .B(n9261), .ZN(n9266)
         );
  OAI211_X1 U10545 ( .C1(n9504), .C2(n9280), .A(n9794), .B(n9264), .ZN(n9414)
         );
  NOR2_X1 U10546 ( .A1(n9414), .A2(n9361), .ZN(n9265) );
  AOI211_X1 U10547 ( .C1(n9770), .C2(n9267), .A(n9266), .B(n9265), .ZN(n9268)
         );
  OAI211_X1 U10548 ( .C1(n9367), .C2(n9416), .A(n9269), .B(n9268), .ZN(
        P1_U3269) );
  NAND2_X1 U10549 ( .A1(n9288), .A2(n9270), .ZN(n9273) );
  INV_X1 U10550 ( .A(n9271), .ZN(n9272) );
  AOI21_X1 U10551 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9424) );
  XOR2_X1 U10552 ( .A(n9275), .B(n9274), .Z(n9426) );
  NAND2_X1 U10553 ( .A1(n9426), .A2(n9350), .ZN(n9286) );
  INV_X1 U10554 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9277) );
  OAI22_X1 U10555 ( .A1(n9816), .A2(n9277), .B1(n9276), .B2(n9800), .ZN(n9278)
         );
  AOI21_X1 U10556 ( .B1(n9322), .B2(n9421), .A(n9278), .ZN(n9279) );
  OAI21_X1 U10557 ( .B1(n9309), .B2(n9324), .A(n9279), .ZN(n9283) );
  INV_X1 U10558 ( .A(n9280), .ZN(n9281) );
  OAI211_X1 U10559 ( .C1(n9508), .C2(n9294), .A(n9281), .B(n9794), .ZN(n9422)
         );
  NOR2_X1 U10560 ( .A1(n9422), .A2(n9326), .ZN(n9282) );
  AOI211_X1 U10561 ( .C1(n9770), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9285)
         );
  OAI211_X1 U10562 ( .C1(n9424), .C2(n9367), .A(n9286), .B(n9285), .ZN(
        P1_U3270) );
  XOR2_X1 U10563 ( .A(n9287), .B(n9289), .Z(n9431) );
  INV_X1 U10564 ( .A(n9431), .ZN(n9302) );
  OAI211_X1 U10565 ( .C1(n9290), .C2(n9289), .A(n9288), .B(n9808), .ZN(n9292)
         );
  NAND2_X1 U10566 ( .A1(n9444), .A2(n9866), .ZN(n9291) );
  OAI211_X1 U10567 ( .C1(n9293), .C2(n9888), .A(n9292), .B(n9291), .ZN(n9429)
         );
  INV_X1 U10568 ( .A(n9295), .ZN(n9512) );
  AOI211_X1 U10569 ( .C1(n9295), .C2(n9311), .A(n9615), .B(n9294), .ZN(n9430)
         );
  NAND2_X1 U10570 ( .A1(n9430), .A2(n9755), .ZN(n9299) );
  INV_X1 U10571 ( .A(n9296), .ZN(n9297) );
  AOI22_X1 U10572 ( .A1(n9822), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9297), .B2(
        n9787), .ZN(n9298) );
  OAI211_X1 U10573 ( .C1(n9512), .C2(n9337), .A(n9299), .B(n9298), .ZN(n9300)
         );
  AOI21_X1 U10574 ( .B1(n9429), .B2(n9816), .A(n9300), .ZN(n9301) );
  OAI21_X1 U10575 ( .B1(n9302), .B2(n9818), .A(n9301), .ZN(P1_U3271) );
  XOR2_X1 U10576 ( .A(n9304), .B(n9303), .Z(n9439) );
  XNOR2_X1 U10577 ( .A(n9305), .B(n9304), .ZN(n9441) );
  NAND2_X1 U10578 ( .A1(n9441), .A2(n9350), .ZN(n9315) );
  AOI22_X1 U10579 ( .A1(n9822), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9306), .B2(
        n9787), .ZN(n9308) );
  NAND2_X1 U10580 ( .A1(n9352), .A2(n9435), .ZN(n9307) );
  OAI211_X1 U10581 ( .C1(n9309), .C2(n9355), .A(n9308), .B(n9307), .ZN(n9313)
         );
  NAND2_X1 U10582 ( .A1(n9434), .A2(n9325), .ZN(n9310) );
  NAND3_X1 U10583 ( .A1(n9311), .A2(n9794), .A3(n9310), .ZN(n9437) );
  NOR2_X1 U10584 ( .A1(n9437), .A2(n9361), .ZN(n9312) );
  AOI211_X1 U10585 ( .C1(n9770), .C2(n9434), .A(n9313), .B(n9312), .ZN(n9314)
         );
  OAI211_X1 U10586 ( .C1(n9439), .C2(n9367), .A(n9315), .B(n9314), .ZN(
        P1_U3272) );
  AOI21_X1 U10587 ( .B1(n9317), .B2(n9316), .A(n4558), .ZN(n9447) );
  XOR2_X1 U10588 ( .A(n9318), .B(n9317), .Z(n9449) );
  NAND2_X1 U10589 ( .A1(n9449), .A2(n9350), .ZN(n9331) );
  INV_X1 U10590 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9320) );
  OAI22_X1 U10591 ( .A1(n9816), .A2(n9320), .B1(n9319), .B2(n9800), .ZN(n9321)
         );
  AOI21_X1 U10592 ( .B1(n9322), .B2(n9444), .A(n9321), .ZN(n9323) );
  OAI21_X1 U10593 ( .B1(n9356), .B2(n9324), .A(n9323), .ZN(n9328) );
  OAI211_X1 U10594 ( .C1(n9520), .C2(n9333), .A(n9794), .B(n9325), .ZN(n9445)
         );
  NOR2_X1 U10595 ( .A1(n9445), .A2(n9326), .ZN(n9327) );
  AOI211_X1 U10596 ( .C1(n9770), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9330)
         );
  OAI211_X1 U10597 ( .C1(n9447), .C2(n9367), .A(n9331), .B(n9330), .ZN(
        P1_U3273) );
  XOR2_X1 U10598 ( .A(n9332), .B(n9339), .Z(n9457) );
  AOI211_X1 U10599 ( .C1(n9453), .C2(n4708), .A(n9615), .B(n9333), .ZN(n9452)
         );
  INV_X1 U10600 ( .A(n9334), .ZN(n9335) );
  AOI22_X1 U10601 ( .A1(n9822), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9335), .B2(
        n9787), .ZN(n9336) );
  OAI21_X1 U10602 ( .B1(n9338), .B2(n9337), .A(n9336), .ZN(n9344) );
  XNOR2_X1 U10603 ( .A(n9340), .B(n9339), .ZN(n9342) );
  AOI222_X1 U10604 ( .A1(n9808), .A2(n9342), .B1(n9435), .B2(n9863), .C1(n9341), .C2(n9866), .ZN(n9455) );
  NOR2_X1 U10605 ( .A1(n9455), .A2(n9822), .ZN(n9343) );
  AOI211_X1 U10606 ( .C1(n9452), .C2(n9755), .A(n9344), .B(n9343), .ZN(n9345)
         );
  OAI21_X1 U10607 ( .B1(n9457), .B2(n9818), .A(n9345), .ZN(P1_U3274) );
  XNOR2_X1 U10608 ( .A(n9347), .B(n9346), .ZN(n9462) );
  XNOR2_X1 U10609 ( .A(n9349), .B(n9348), .ZN(n9464) );
  NAND2_X1 U10610 ( .A1(n9464), .A2(n9350), .ZN(n9366) );
  AOI22_X1 U10611 ( .A1(n9822), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9351), .B2(
        n9787), .ZN(n9354) );
  NAND2_X1 U10612 ( .A1(n9352), .A2(n9458), .ZN(n9353) );
  OAI211_X1 U10613 ( .C1(n9356), .C2(n9355), .A(n9354), .B(n9353), .ZN(n9363)
         );
  NAND2_X1 U10614 ( .A1(n9357), .A2(n9364), .ZN(n9358) );
  NAND2_X1 U10615 ( .A1(n9358), .A2(n9794), .ZN(n9360) );
  OR2_X1 U10616 ( .A1(n9360), .A2(n9359), .ZN(n9460) );
  NOR2_X1 U10617 ( .A1(n9460), .A2(n9361), .ZN(n9362) );
  AOI211_X1 U10618 ( .C1(n9770), .C2(n9364), .A(n9363), .B(n9362), .ZN(n9365)
         );
  OAI211_X1 U10619 ( .C1(n9462), .C2(n9367), .A(n9366), .B(n9365), .ZN(
        P1_U3275) );
  INV_X1 U10620 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9369) );
  AND2_X1 U10621 ( .A1(n9368), .A2(n9371), .ZN(n9479) );
  MUX2_X1 U10622 ( .A(n9369), .B(n9479), .S(n9928), .Z(n9370) );
  OAI21_X1 U10623 ( .B1(n9482), .B2(n9478), .A(n9370), .ZN(P1_U3554) );
  INV_X1 U10624 ( .A(n9371), .ZN(n9372) );
  NOR2_X1 U10625 ( .A1(n9373), .A2(n9372), .ZN(n9483) );
  MUX2_X1 U10626 ( .A(n9374), .B(n9483), .S(n9928), .Z(n9375) );
  OAI21_X1 U10627 ( .B1(n9486), .B2(n9478), .A(n9375), .ZN(P1_U3553) );
  AOI21_X1 U10628 ( .B1(n9380), .B2(n9885), .A(n9379), .ZN(n9487) );
  MUX2_X1 U10629 ( .A(n9381), .B(n9487), .S(n9928), .Z(n9382) );
  OAI21_X1 U10630 ( .B1(n4705), .B2(n9478), .A(n9382), .ZN(P1_U3551) );
  INV_X1 U10631 ( .A(n9885), .ZN(n9456) );
  AOI211_X1 U10632 ( .C1(n9385), .C2(n9892), .A(n9384), .B(n9383), .ZN(n9386)
         );
  OAI21_X1 U10633 ( .B1(n9387), .B2(n9456), .A(n9386), .ZN(n9490) );
  MUX2_X1 U10634 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9490), .S(n9928), .Z(
        P1_U3550) );
  AOI211_X1 U10635 ( .C1(n9390), .C2(n9885), .A(n9389), .B(n9388), .ZN(n9491)
         );
  MUX2_X1 U10636 ( .A(n9391), .B(n9491), .S(n9928), .Z(n9392) );
  OAI21_X1 U10637 ( .B1(n9494), .B2(n9478), .A(n9392), .ZN(P1_U3549) );
  AOI21_X1 U10638 ( .B1(n9394), .B2(n9892), .A(n9393), .ZN(n9395) );
  OAI211_X1 U10639 ( .C1(n9397), .C2(n9456), .A(n9396), .B(n9395), .ZN(n9495)
         );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9495), .S(n9928), .Z(
        P1_U3548) );
  NOR2_X1 U10641 ( .A1(n9398), .A2(n9888), .ZN(n9400) );
  AOI211_X1 U10642 ( .C1(n9866), .C2(n9413), .A(n9400), .B(n9399), .ZN(n9401)
         );
  OAI21_X1 U10643 ( .B1(n9882), .B2(n9402), .A(n9401), .ZN(n9403) );
  AOI21_X1 U10644 ( .B1(n9404), .B2(n9885), .A(n9403), .ZN(n9497) );
  MUX2_X1 U10645 ( .A(n9497), .B(n9405), .S(n9925), .Z(n9406) );
  OAI21_X1 U10646 ( .B1(n9499), .B2(n9478), .A(n9406), .ZN(P1_U3547) );
  AOI211_X1 U10647 ( .C1(n9409), .C2(n9892), .A(n9408), .B(n9407), .ZN(n9410)
         );
  OAI21_X1 U10648 ( .B1(n9411), .B2(n9456), .A(n9410), .ZN(n9500) );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9500), .S(n9928), .Z(
        P1_U3546) );
  AOI22_X1 U10650 ( .A1(n9413), .A2(n9863), .B1(n9866), .B2(n9412), .ZN(n9415)
         );
  OAI211_X1 U10651 ( .C1(n9416), .C2(n9882), .A(n9415), .B(n9414), .ZN(n9417)
         );
  AOI21_X1 U10652 ( .B1(n9418), .B2(n9885), .A(n9417), .ZN(n9501) );
  MUX2_X1 U10653 ( .A(n9419), .B(n9501), .S(n9928), .Z(n9420) );
  OAI21_X1 U10654 ( .B1(n9504), .B2(n9478), .A(n9420), .ZN(P1_U3545) );
  AOI22_X1 U10655 ( .A1(n9421), .A2(n9863), .B1(n9866), .B2(n9436), .ZN(n9423)
         );
  OAI211_X1 U10656 ( .C1(n9424), .C2(n9882), .A(n9423), .B(n9422), .ZN(n9425)
         );
  AOI21_X1 U10657 ( .B1(n9426), .B2(n9885), .A(n9425), .ZN(n9505) );
  MUX2_X1 U10658 ( .A(n9427), .B(n9505), .S(n9928), .Z(n9428) );
  OAI21_X1 U10659 ( .B1(n9508), .B2(n9478), .A(n9428), .ZN(P1_U3544) );
  AOI211_X1 U10660 ( .C1(n9431), .C2(n9885), .A(n9430), .B(n9429), .ZN(n9509)
         );
  MUX2_X1 U10661 ( .A(n9432), .B(n9509), .S(n9928), .Z(n9433) );
  OAI21_X1 U10662 ( .B1(n9512), .B2(n9478), .A(n9433), .ZN(P1_U3543) );
  INV_X1 U10663 ( .A(n9434), .ZN(n9516) );
  AOI22_X1 U10664 ( .A1(n9436), .A2(n9863), .B1(n9435), .B2(n9866), .ZN(n9438)
         );
  OAI211_X1 U10665 ( .C1(n9439), .C2(n9882), .A(n9438), .B(n9437), .ZN(n9440)
         );
  AOI21_X1 U10666 ( .B1(n9441), .B2(n9885), .A(n9440), .ZN(n9513) );
  MUX2_X1 U10667 ( .A(n9442), .B(n9513), .S(n9928), .Z(n9443) );
  OAI21_X1 U10668 ( .B1(n9516), .B2(n9478), .A(n9443), .ZN(P1_U3542) );
  AOI22_X1 U10669 ( .A1(n9444), .A2(n9863), .B1(n9866), .B2(n9459), .ZN(n9446)
         );
  OAI211_X1 U10670 ( .C1(n9447), .C2(n9882), .A(n9446), .B(n9445), .ZN(n9448)
         );
  AOI21_X1 U10671 ( .B1(n9449), .B2(n9885), .A(n9448), .ZN(n9517) );
  MUX2_X1 U10672 ( .A(n9450), .B(n9517), .S(n9928), .Z(n9451) );
  OAI21_X1 U10673 ( .B1(n9520), .B2(n9478), .A(n9451), .ZN(P1_U3541) );
  AOI21_X1 U10674 ( .B1(n9453), .B2(n9892), .A(n9452), .ZN(n9454) );
  OAI211_X1 U10675 ( .C1(n9457), .C2(n9456), .A(n9455), .B(n9454), .ZN(n9521)
         );
  MUX2_X1 U10676 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9521), .S(n9928), .Z(
        P1_U3540) );
  INV_X1 U10677 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9465) );
  AOI22_X1 U10678 ( .A1(n9459), .A2(n9863), .B1(n9458), .B2(n9866), .ZN(n9461)
         );
  OAI211_X1 U10679 ( .C1(n9462), .C2(n9882), .A(n9461), .B(n9460), .ZN(n9463)
         );
  AOI21_X1 U10680 ( .B1(n9464), .B2(n9885), .A(n9463), .ZN(n9522) );
  MUX2_X1 U10681 ( .A(n9465), .B(n9522), .S(n9928), .Z(n9466) );
  OAI21_X1 U10682 ( .B1(n4706), .B2(n9478), .A(n9466), .ZN(P1_U3539) );
  AOI211_X1 U10683 ( .C1(n9469), .C2(n9885), .A(n9468), .B(n9467), .ZN(n9525)
         );
  MUX2_X1 U10684 ( .A(n9470), .B(n9525), .S(n9928), .Z(n9471) );
  OAI21_X1 U10685 ( .B1(n9528), .B2(n9478), .A(n9471), .ZN(P1_U3538) );
  OAI211_X1 U10686 ( .C1(n9474), .C2(n9886), .A(n9473), .B(n9472), .ZN(n9475)
         );
  AOI21_X1 U10687 ( .B1(n9476), .B2(n9885), .A(n9475), .ZN(n9529) );
  MUX2_X1 U10688 ( .A(n7449), .B(n9529), .S(n9928), .Z(n9477) );
  OAI21_X1 U10689 ( .B1(n9533), .B2(n9478), .A(n9477), .ZN(P1_U3537) );
  INV_X1 U10690 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9480) );
  MUX2_X1 U10691 ( .A(n9480), .B(n9479), .S(n9911), .Z(n9481) );
  OAI21_X1 U10692 ( .B1(n9482), .B2(n9532), .A(n9481), .ZN(P1_U3522) );
  INV_X1 U10693 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9484) );
  MUX2_X1 U10694 ( .A(n9484), .B(n9483), .S(n9911), .Z(n9485) );
  OAI21_X1 U10695 ( .B1(n9486), .B2(n9532), .A(n9485), .ZN(P1_U3521) );
  INV_X1 U10696 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9488) );
  MUX2_X1 U10697 ( .A(n9488), .B(n9487), .S(n9911), .Z(n9489) );
  OAI21_X1 U10698 ( .B1(n4705), .B2(n9532), .A(n9489), .ZN(P1_U3519) );
  MUX2_X1 U10699 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9490), .S(n9911), .Z(
        P1_U3518) );
  INV_X1 U10700 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9492) );
  MUX2_X1 U10701 ( .A(n9492), .B(n9491), .S(n9911), .Z(n9493) );
  OAI21_X1 U10702 ( .B1(n9494), .B2(n9532), .A(n9493), .ZN(P1_U3517) );
  MUX2_X1 U10703 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9495), .S(n9911), .Z(
        P1_U3516) );
  INV_X1 U10704 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9496) );
  MUX2_X1 U10705 ( .A(n9497), .B(n9496), .S(n9909), .Z(n9498) );
  OAI21_X1 U10706 ( .B1(n9499), .B2(n9532), .A(n9498), .ZN(P1_U3515) );
  MUX2_X1 U10707 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9500), .S(n9911), .Z(
        P1_U3514) );
  INV_X1 U10708 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9502) );
  MUX2_X1 U10709 ( .A(n9502), .B(n9501), .S(n9911), .Z(n9503) );
  OAI21_X1 U10710 ( .B1(n9504), .B2(n9532), .A(n9503), .ZN(P1_U3513) );
  INV_X1 U10711 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U10712 ( .A(n9506), .B(n9505), .S(n9911), .Z(n9507) );
  OAI21_X1 U10713 ( .B1(n9508), .B2(n9532), .A(n9507), .ZN(P1_U3512) );
  INV_X1 U10714 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9510) );
  MUX2_X1 U10715 ( .A(n9510), .B(n9509), .S(n9911), .Z(n9511) );
  OAI21_X1 U10716 ( .B1(n9512), .B2(n9532), .A(n9511), .ZN(P1_U3511) );
  INV_X1 U10717 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9514) );
  MUX2_X1 U10718 ( .A(n9514), .B(n9513), .S(n9911), .Z(n9515) );
  OAI21_X1 U10719 ( .B1(n9516), .B2(n9532), .A(n9515), .ZN(P1_U3510) );
  INV_X1 U10720 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9518) );
  MUX2_X1 U10721 ( .A(n9518), .B(n9517), .S(n9911), .Z(n9519) );
  OAI21_X1 U10722 ( .B1(n9520), .B2(n9532), .A(n9519), .ZN(P1_U3508) );
  MUX2_X1 U10723 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9521), .S(n9911), .Z(
        P1_U3505) );
  MUX2_X1 U10724 ( .A(n9523), .B(n9522), .S(n9911), .Z(n9524) );
  OAI21_X1 U10725 ( .B1(n4706), .B2(n9532), .A(n9524), .ZN(P1_U3502) );
  INV_X1 U10726 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9526) );
  MUX2_X1 U10727 ( .A(n9526), .B(n9525), .S(n9911), .Z(n9527) );
  OAI21_X1 U10728 ( .B1(n9528), .B2(n9532), .A(n9527), .ZN(P1_U3499) );
  INV_X1 U10729 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9530) );
  MUX2_X1 U10730 ( .A(n9530), .B(n9529), .S(n9911), .Z(n9531) );
  OAI21_X1 U10731 ( .B1(n9533), .B2(n9532), .A(n9531), .ZN(P1_U3496) );
  NOR4_X1 U10732 ( .A1(n5247), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9534), .A4(
        P1_U3084), .ZN(n9535) );
  AOI21_X1 U10733 ( .B1(n9545), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9535), .ZN(
        n9536) );
  OAI21_X1 U10734 ( .B1(n9537), .B2(n9548), .A(n9536), .ZN(P1_U3322) );
  INV_X1 U10735 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10445) );
  OAI222_X1 U10736 ( .A1(n9541), .A2(n10445), .B1(n9548), .B2(n9540), .C1(
        P1_U3084), .C2(n9538), .ZN(P1_U3323) );
  AOI21_X1 U10737 ( .B1(n9545), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9542), .ZN(
        n9543) );
  OAI21_X1 U10738 ( .B1(n9544), .B2(n9548), .A(n9543), .ZN(P1_U3325) );
  NAND2_X1 U10739 ( .A1(n9545), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9546) );
  OAI211_X1 U10740 ( .C1(n9549), .C2(n9548), .A(n9547), .B(n9546), .ZN(
        P1_U3326) );
  MUX2_X1 U10741 ( .A(n9550), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI211_X1 U10742 ( .C1(n9553), .C2(n9552), .A(n9551), .B(n9720), .ZN(n9558)
         );
  AOI211_X1 U10743 ( .C1(n9556), .C2(n9555), .A(n9554), .B(n9715), .ZN(n9557)
         );
  AOI211_X1 U10744 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(P1_U3084), .A(n9558), 
        .B(n9557), .ZN(n9563) );
  INV_X1 U10745 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9560) );
  OAI22_X1 U10746 ( .A1(n9748), .A2(n9560), .B1(n9559), .B2(n9739), .ZN(n9561)
         );
  INV_X1 U10747 ( .A(n9561), .ZN(n9562) );
  NAND2_X1 U10748 ( .A1(n9563), .A2(n9562), .ZN(P1_U3244) );
  OAI22_X1 U10749 ( .A1(n9565), .A2(n10024), .B1(n9564), .B2(n10022), .ZN(
        n9567) );
  AOI211_X1 U10750 ( .C1(n10029), .C2(n9568), .A(n9567), .B(n9566), .ZN(n9585)
         );
  AOI22_X1 U10751 ( .A1(n10052), .A2(n9585), .B1(n9569), .B2(n10050), .ZN(
        P2_U3535) );
  OAI22_X1 U10752 ( .A1(n9571), .A2(n10024), .B1(n9570), .B2(n10022), .ZN(
        n9573) );
  AOI211_X1 U10753 ( .C1(n10029), .C2(n9574), .A(n9573), .B(n9572), .ZN(n9587)
         );
  AOI22_X1 U10754 ( .A1(n10052), .A2(n9587), .B1(n9575), .B2(n10050), .ZN(
        P2_U3534) );
  INV_X1 U10755 ( .A(n9576), .ZN(n10010) );
  INV_X1 U10756 ( .A(n9577), .ZN(n9582) );
  OAI22_X1 U10757 ( .A1(n9579), .A2(n10024), .B1(n9578), .B2(n10022), .ZN(
        n9581) );
  AOI211_X1 U10758 ( .C1(n10010), .C2(n9582), .A(n9581), .B(n9580), .ZN(n9589)
         );
  AOI22_X1 U10759 ( .A1(n10052), .A2(n9589), .B1(n9583), .B2(n10050), .ZN(
        P2_U3533) );
  INV_X1 U10760 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9584) );
  AOI22_X1 U10761 ( .A1(n10032), .A2(n9585), .B1(n9584), .B2(n10030), .ZN(
        P2_U3496) );
  INV_X1 U10762 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U10763 ( .A1(n10032), .A2(n9587), .B1(n9586), .B2(n10030), .ZN(
        P2_U3493) );
  INV_X1 U10764 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9588) );
  AOI22_X1 U10765 ( .A1(n10032), .A2(n9589), .B1(n9588), .B2(n10030), .ZN(
        P2_U3490) );
  INV_X1 U10766 ( .A(n9600), .ZN(n9590) );
  XNOR2_X1 U10767 ( .A(n9591), .B(n9590), .ZN(n9641) );
  INV_X1 U10768 ( .A(n9592), .ZN(n9595) );
  AOI21_X1 U10769 ( .B1(n9593), .B2(n9637), .A(n9615), .ZN(n9594) );
  NAND2_X1 U10770 ( .A1(n9595), .A2(n9594), .ZN(n9639) );
  INV_X1 U10771 ( .A(n9639), .ZN(n9596) );
  AOI22_X1 U10772 ( .A1(n9641), .A2(n9350), .B1(n9755), .B2(n9596), .ZN(n9613)
         );
  INV_X1 U10773 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9599) );
  INV_X1 U10774 ( .A(n9597), .ZN(n9598) );
  OAI22_X1 U10775 ( .A1(n9816), .A2(n9599), .B1(n9598), .B2(n9800), .ZN(n9611)
         );
  NAND2_X1 U10776 ( .A1(n9601), .A2(n9600), .ZN(n9602) );
  NAND2_X1 U10777 ( .A1(n9603), .A2(n9602), .ZN(n9604) );
  NAND2_X1 U10778 ( .A1(n9604), .A2(n9808), .ZN(n9608) );
  AOI22_X1 U10779 ( .A1(n9606), .A2(n9866), .B1(n9863), .B2(n9605), .ZN(n9607)
         );
  NAND2_X1 U10780 ( .A1(n9608), .A2(n9607), .ZN(n9609) );
  AOI21_X1 U10781 ( .B1(n9641), .B2(n9900), .A(n9609), .ZN(n9643) );
  NOR2_X1 U10782 ( .A1(n9643), .A2(n9822), .ZN(n9610) );
  AOI211_X1 U10783 ( .C1(n9770), .C2(n9637), .A(n9611), .B(n9610), .ZN(n9612)
         );
  NAND2_X1 U10784 ( .A1(n9613), .A2(n9612), .ZN(P1_U3278) );
  XNOR2_X1 U10785 ( .A(n9614), .B(n9625), .ZN(n9653) );
  AOI21_X1 U10786 ( .B1(n9616), .B2(n9634), .A(n9615), .ZN(n9618) );
  NAND2_X1 U10787 ( .A1(n9618), .A2(n9617), .ZN(n9650) );
  INV_X1 U10788 ( .A(n9650), .ZN(n9619) );
  AOI22_X1 U10789 ( .A1(n9653), .A2(n9350), .B1(n9755), .B2(n9619), .ZN(n9636)
         );
  INV_X1 U10790 ( .A(n9620), .ZN(n9621) );
  OAI22_X1 U10791 ( .A1(n9816), .A2(n9622), .B1(n9621), .B2(n9800), .ZN(n9633)
         );
  NAND2_X1 U10792 ( .A1(n9624), .A2(n9623), .ZN(n9626) );
  XNOR2_X1 U10793 ( .A(n9626), .B(n9625), .ZN(n9630) );
  OAI22_X1 U10794 ( .A1(n9762), .A2(n9886), .B1(n9627), .B2(n9888), .ZN(n9628)
         );
  INV_X1 U10795 ( .A(n9628), .ZN(n9629) );
  OAI21_X1 U10796 ( .B1(n9630), .B2(n9882), .A(n9629), .ZN(n9631) );
  AOI21_X1 U10797 ( .B1(n9653), .B2(n9900), .A(n9631), .ZN(n9655) );
  NOR2_X1 U10798 ( .A1(n9655), .A2(n9822), .ZN(n9632) );
  AOI211_X1 U10799 ( .C1(n9770), .C2(n9634), .A(n9633), .B(n9632), .ZN(n9635)
         );
  NAND2_X1 U10800 ( .A1(n9636), .A2(n9635), .ZN(P1_U3280) );
  INV_X1 U10801 ( .A(n9896), .ZN(n9905) );
  NAND2_X1 U10802 ( .A1(n9637), .A2(n9892), .ZN(n9638) );
  NAND2_X1 U10803 ( .A1(n9639), .A2(n9638), .ZN(n9640) );
  AOI21_X1 U10804 ( .B1(n9641), .B2(n9905), .A(n9640), .ZN(n9642) );
  AND2_X1 U10805 ( .A1(n9643), .A2(n9642), .ZN(n9657) );
  AOI22_X1 U10806 ( .A1(n9928), .A2(n9657), .B1(n7133), .B2(n9925), .ZN(
        P1_U3536) );
  OAI21_X1 U10807 ( .B1(n9645), .B2(n9902), .A(n9644), .ZN(n9646) );
  AOI21_X1 U10808 ( .B1(n9647), .B2(n9905), .A(n9646), .ZN(n9648) );
  AND2_X1 U10809 ( .A1(n9649), .A2(n9648), .ZN(n9658) );
  AOI22_X1 U10810 ( .A1(n9928), .A2(n9658), .B1(n6989), .B2(n9925), .ZN(
        P1_U3535) );
  OAI21_X1 U10811 ( .B1(n9651), .B2(n9902), .A(n9650), .ZN(n9652) );
  AOI21_X1 U10812 ( .B1(n9653), .B2(n9905), .A(n9652), .ZN(n9654) );
  AND2_X1 U10813 ( .A1(n9655), .A2(n9654), .ZN(n9660) );
  AOI22_X1 U10814 ( .A1(n9928), .A2(n9660), .B1(n6845), .B2(n9925), .ZN(
        P1_U3534) );
  INV_X1 U10815 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9656) );
  AOI22_X1 U10816 ( .A1(n9911), .A2(n9657), .B1(n9656), .B2(n9909), .ZN(
        P1_U3493) );
  AOI22_X1 U10817 ( .A1(n9911), .A2(n9658), .B1(n5444), .B2(n9909), .ZN(
        P1_U3490) );
  INV_X1 U10818 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U10819 ( .A1(n9911), .A2(n9660), .B1(n9659), .B2(n9909), .ZN(
        P1_U3487) );
  INV_X1 U10820 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10209) );
  XOR2_X1 U10821 ( .A(n10209), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XOR2_X1 U10822 ( .A(P1_RD_REG_SCAN_IN), .B(n5081), .Z(U126) );
  OAI21_X1 U10823 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9668) );
  OAI21_X1 U10824 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9667) );
  AOI22_X1 U10825 ( .A1(n9735), .A2(n9668), .B1(n9744), .B2(n9667), .ZN(n9673)
         );
  AOI211_X1 U10826 ( .C1(n9708), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9672)
         );
  OAI211_X1 U10827 ( .C1(n9748), .C2(n10060), .A(n9673), .B(n9672), .ZN(
        P1_U3245) );
  XNOR2_X1 U10828 ( .A(n9675), .B(n9674), .ZN(n9681) );
  AOI211_X1 U10829 ( .C1(n9678), .C2(n9677), .A(n9676), .B(n9720), .ZN(n9679)
         );
  AOI211_X1 U10830 ( .C1(n9735), .C2(n9681), .A(n9680), .B(n9679), .ZN(n9686)
         );
  INV_X1 U10831 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9683) );
  OAI22_X1 U10832 ( .A1(n9748), .A2(n9683), .B1(n9682), .B2(n9739), .ZN(n9684)
         );
  INV_X1 U10833 ( .A(n9684), .ZN(n9685) );
  NAND2_X1 U10834 ( .A1(n9686), .A2(n9685), .ZN(P1_U3246) );
  OAI21_X1 U10835 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(n9696) );
  NOR2_X1 U10836 ( .A1(n9691), .A2(n9690), .ZN(n9692) );
  NOR3_X1 U10837 ( .A1(n9715), .A2(n9693), .A3(n9692), .ZN(n9694) );
  AOI211_X1 U10838 ( .C1(n9744), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9701)
         );
  INV_X1 U10839 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9698) );
  OAI22_X1 U10840 ( .A1(n9748), .A2(n9698), .B1(n9697), .B2(n9739), .ZN(n9699)
         );
  INV_X1 U10841 ( .A(n9699), .ZN(n9700) );
  NAND2_X1 U10842 ( .A1(n9701), .A2(n9700), .ZN(P1_U3247) );
  INV_X1 U10843 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10492) );
  AOI211_X1 U10844 ( .C1(n9704), .C2(n9703), .A(n9715), .B(n9702), .ZN(n9705)
         );
  AOI211_X1 U10845 ( .C1(n9708), .C2(n9707), .A(n9706), .B(n9705), .ZN(n9713)
         );
  XNOR2_X1 U10846 ( .A(n9710), .B(n9709), .ZN(n9711) );
  NAND2_X1 U10847 ( .A1(n9744), .A2(n9711), .ZN(n9712) );
  OAI211_X1 U10848 ( .C1(n10492), .C2(n9748), .A(n9713), .B(n9712), .ZN(
        P1_U3250) );
  AOI211_X1 U10849 ( .C1(n9717), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9725)
         );
  NAND2_X1 U10850 ( .A1(n9719), .A2(n9718), .ZN(n9721) );
  AOI21_X1 U10851 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9723) );
  NOR3_X1 U10852 ( .A1(n9725), .A2(n9724), .A3(n9723), .ZN(n9730) );
  INV_X1 U10853 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9727) );
  OAI22_X1 U10854 ( .A1(n9748), .A2(n9727), .B1(n9726), .B2(n9739), .ZN(n9728)
         );
  INV_X1 U10855 ( .A(n9728), .ZN(n9729) );
  NAND2_X1 U10856 ( .A1(n9730), .A2(n9729), .ZN(P1_U3251) );
  INV_X1 U10857 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10502) );
  AOI21_X1 U10858 ( .B1(n9733), .B2(n9732), .A(n9731), .ZN(n9734) );
  NAND2_X1 U10859 ( .A1(n9735), .A2(n9734), .ZN(n9737) );
  OAI211_X1 U10860 ( .C1(n9739), .C2(n9738), .A(n9737), .B(n9736), .ZN(n9740)
         );
  INV_X1 U10861 ( .A(n9740), .ZN(n9747) );
  OAI21_X1 U10862 ( .B1(n9743), .B2(n9742), .A(n9741), .ZN(n9745) );
  NAND2_X1 U10863 ( .A1(n9745), .A2(n9744), .ZN(n9746) );
  OAI211_X1 U10864 ( .C1(n10502), .C2(n9748), .A(n9747), .B(n9746), .ZN(
        P1_U3259) );
  INV_X1 U10865 ( .A(n9759), .ZN(n9749) );
  XNOR2_X1 U10866 ( .A(n9750), .B(n9749), .ZN(n9906) );
  OAI21_X1 U10867 ( .B1(n9751), .B2(n9903), .A(n9794), .ZN(n9753) );
  OR2_X1 U10868 ( .A1(n9753), .A2(n9752), .ZN(n9901) );
  INV_X1 U10869 ( .A(n9901), .ZN(n9754) );
  AOI22_X1 U10870 ( .A1(n9906), .A2(n9350), .B1(n9755), .B2(n9754), .ZN(n9772)
         );
  INV_X1 U10871 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9758) );
  INV_X1 U10872 ( .A(n9756), .ZN(n9757) );
  OAI22_X1 U10873 ( .A1(n9816), .A2(n9758), .B1(n9757), .B2(n9800), .ZN(n9768)
         );
  XNOR2_X1 U10874 ( .A(n9760), .B(n9759), .ZN(n9761) );
  NAND2_X1 U10875 ( .A1(n9761), .A2(n9808), .ZN(n9765) );
  OAI22_X1 U10876 ( .A1(n9875), .A2(n9886), .B1(n9762), .B2(n9888), .ZN(n9763)
         );
  INV_X1 U10877 ( .A(n9763), .ZN(n9764) );
  NAND2_X1 U10878 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  AOI21_X1 U10879 ( .B1(n9906), .B2(n9900), .A(n9766), .ZN(n9908) );
  NOR2_X1 U10880 ( .A1(n9908), .A2(n9822), .ZN(n9767) );
  AOI211_X1 U10881 ( .C1(n9770), .C2(n9769), .A(n9768), .B(n9767), .ZN(n9771)
         );
  NAND2_X1 U10882 ( .A1(n9772), .A2(n9771), .ZN(P1_U3282) );
  XNOR2_X1 U10883 ( .A(n9773), .B(n5342), .ZN(n9862) );
  INV_X1 U10884 ( .A(n9774), .ZN(n9775) );
  OAI211_X1 U10885 ( .C1(n9860), .C2(n9776), .A(n9775), .B(n9794), .ZN(n9858)
         );
  NAND2_X1 U10886 ( .A1(n9778), .A2(n9777), .ZN(n9780) );
  XNOR2_X1 U10887 ( .A(n9780), .B(n9779), .ZN(n9783) );
  AOI222_X1 U10888 ( .A1(n9808), .A2(n9783), .B1(n9782), .B2(n9863), .C1(n9781), .C2(n9866), .ZN(n9859) );
  AOI22_X1 U10889 ( .A1(n9787), .A2(n9786), .B1(n9785), .B2(n9784), .ZN(n9788)
         );
  OAI211_X1 U10890 ( .C1(n9789), .C2(n9858), .A(n9859), .B(n9788), .ZN(n9790)
         );
  AOI21_X1 U10891 ( .B1(n9791), .B2(n9862), .A(n9790), .ZN(n9792) );
  AOI22_X1 U10892 ( .A1(n9822), .A2(n6615), .B1(n9792), .B2(n9816), .ZN(
        P1_U3286) );
  INV_X1 U10893 ( .A(n9793), .ZN(n9795) );
  OAI211_X1 U10894 ( .C1(n9798), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9825)
         );
  INV_X1 U10895 ( .A(n9825), .ZN(n9815) );
  OAI22_X1 U10896 ( .A1(n9800), .A2(n9799), .B1(n9798), .B2(n9797), .ZN(n9813)
         );
  OAI21_X1 U10897 ( .B1(n9803), .B2(n9802), .A(n9801), .ZN(n9827) );
  AOI22_X1 U10898 ( .A1(n6602), .A2(n9863), .B1(n9866), .B2(n9804), .ZN(n9811)
         );
  OAI21_X1 U10899 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9809) );
  NAND2_X1 U10900 ( .A1(n9809), .A2(n9808), .ZN(n9810) );
  OAI211_X1 U10901 ( .C1(n9827), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9829)
         );
  AOI211_X1 U10902 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n9829), .ZN(n9821)
         );
  INV_X1 U10903 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9817) );
  OAI22_X1 U10904 ( .A1(n9818), .A2(n9827), .B1(n9817), .B2(n9816), .ZN(n9819)
         );
  INV_X1 U10905 ( .A(n9819), .ZN(n9820) );
  OAI21_X1 U10906 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(P1_U3290) );
  AND2_X1 U10907 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9823), .ZN(P1_U3292) );
  AND2_X1 U10908 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9823), .ZN(P1_U3293) );
  AND2_X1 U10909 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9823), .ZN(P1_U3294) );
  AND2_X1 U10910 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9823), .ZN(P1_U3295) );
  AND2_X1 U10911 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9823), .ZN(P1_U3296) );
  AND2_X1 U10912 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9823), .ZN(P1_U3297) );
  AND2_X1 U10913 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9823), .ZN(P1_U3298) );
  AND2_X1 U10914 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9823), .ZN(P1_U3299) );
  AND2_X1 U10915 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9823), .ZN(P1_U3300) );
  AND2_X1 U10916 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9823), .ZN(P1_U3301) );
  AND2_X1 U10917 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9823), .ZN(P1_U3302) );
  AND2_X1 U10918 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9823), .ZN(P1_U3303) );
  AND2_X1 U10919 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9823), .ZN(P1_U3304) );
  AND2_X1 U10920 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9823), .ZN(P1_U3305) );
  AND2_X1 U10921 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9823), .ZN(P1_U3306) );
  AND2_X1 U10922 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9823), .ZN(P1_U3307) );
  AND2_X1 U10923 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9823), .ZN(P1_U3308) );
  AND2_X1 U10924 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9823), .ZN(P1_U3309) );
  AND2_X1 U10925 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9823), .ZN(P1_U3310) );
  AND2_X1 U10926 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9823), .ZN(P1_U3311) );
  AND2_X1 U10927 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9823), .ZN(P1_U3312) );
  AND2_X1 U10928 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9823), .ZN(P1_U3313) );
  AND2_X1 U10929 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9823), .ZN(P1_U3314) );
  AND2_X1 U10930 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9823), .ZN(P1_U3315) );
  AND2_X1 U10931 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9823), .ZN(P1_U3316) );
  AND2_X1 U10932 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9823), .ZN(P1_U3317) );
  AND2_X1 U10933 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9823), .ZN(P1_U3318) );
  INV_X1 U10934 ( .A(n9823), .ZN(n9824) );
  INV_X1 U10935 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10399) );
  NOR2_X1 U10936 ( .A1(n9824), .A2(n10399), .ZN(P1_U3319) );
  INV_X1 U10937 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U10938 ( .A1(n9824), .A2(n10199), .ZN(P1_U3320) );
  INV_X1 U10939 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U10940 ( .A1(n9824), .A2(n10417), .ZN(P1_U3321) );
  OAI211_X1 U10941 ( .C1(n9827), .C2(n9896), .A(n9826), .B(n9825), .ZN(n9828)
         );
  NOR2_X1 U10942 ( .A1(n9829), .A2(n9828), .ZN(n9912) );
  INV_X1 U10943 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9830) );
  AOI22_X1 U10944 ( .A1(n9911), .A2(n9912), .B1(n9830), .B2(n9909), .ZN(
        P1_U3457) );
  OAI21_X1 U10945 ( .B1(n9832), .B2(n9902), .A(n9831), .ZN(n9834) );
  AOI211_X1 U10946 ( .C1(n9905), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9913)
         );
  AOI22_X1 U10947 ( .A1(n9911), .A2(n9913), .B1(n5268), .B2(n9909), .ZN(
        P1_U3460) );
  INV_X1 U10948 ( .A(n9844), .ZN(n9846) );
  OAI22_X1 U10949 ( .A1(n5294), .A2(n9886), .B1(n9836), .B2(n9888), .ZN(n9837)
         );
  INV_X1 U10950 ( .A(n9837), .ZN(n9838) );
  OAI211_X1 U10951 ( .C1(n9840), .C2(n9902), .A(n9839), .B(n9838), .ZN(n9841)
         );
  INV_X1 U10952 ( .A(n9841), .ZN(n9843) );
  OAI211_X1 U10953 ( .C1(n9844), .C2(n9896), .A(n9843), .B(n9842), .ZN(n9845)
         );
  AOI21_X1 U10954 ( .B1(n9900), .B2(n9846), .A(n9845), .ZN(n9915) );
  AOI22_X1 U10955 ( .A1(n9911), .A2(n9915), .B1(n5297), .B2(n9909), .ZN(
        P1_U3463) );
  INV_X1 U10956 ( .A(n9855), .ZN(n9857) );
  AND2_X1 U10957 ( .A1(n9892), .A2(n9847), .ZN(n9851) );
  OAI22_X1 U10958 ( .A1(n9849), .A2(n9886), .B1(n9848), .B2(n9888), .ZN(n9850)
         );
  NOR4_X1 U10959 ( .A1(n9853), .A2(n9852), .A3(n9851), .A4(n9850), .ZN(n9854)
         );
  OAI21_X1 U10960 ( .B1(n9855), .B2(n9896), .A(n9854), .ZN(n9856) );
  AOI21_X1 U10961 ( .B1(n9900), .B2(n9857), .A(n9856), .ZN(n9917) );
  AOI22_X1 U10962 ( .A1(n9911), .A2(n9917), .B1(n5310), .B2(n9909), .ZN(
        P1_U3466) );
  OAI211_X1 U10963 ( .C1(n9860), .C2(n9902), .A(n9859), .B(n9858), .ZN(n9861)
         );
  AOI21_X1 U10964 ( .B1(n9885), .B2(n9862), .A(n9861), .ZN(n9919) );
  AOI22_X1 U10965 ( .A1(n9911), .A2(n9919), .B1(n5328), .B2(n9909), .ZN(
        P1_U3469) );
  NAND2_X1 U10966 ( .A1(n9873), .A2(n9905), .ZN(n9870) );
  AOI22_X1 U10967 ( .A1(n9866), .A2(n9865), .B1(n9864), .B2(n9863), .ZN(n9869)
         );
  NAND4_X1 U10968 ( .A1(n9870), .A2(n9869), .A3(n9868), .A4(n9867), .ZN(n9871)
         );
  AOI211_X1 U10969 ( .C1(n9900), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9920)
         );
  INV_X1 U10970 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U10971 ( .A1(n9911), .A2(n9920), .B1(n9874), .B2(n9909), .ZN(
        P1_U3472) );
  OAI22_X1 U10972 ( .A1(n9876), .A2(n9886), .B1(n9875), .B2(n9888), .ZN(n9878)
         );
  AOI211_X1 U10973 ( .C1(n9879), .C2(n9892), .A(n9878), .B(n9877), .ZN(n9880)
         );
  OAI21_X1 U10974 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(n9883) );
  AOI21_X1 U10975 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9922) );
  AOI22_X1 U10976 ( .A1(n9911), .A2(n9922), .B1(n5366), .B2(n9909), .ZN(
        P1_U3475) );
  OAI22_X1 U10977 ( .A1(n9889), .A2(n9888), .B1(n9887), .B2(n9886), .ZN(n9891)
         );
  AOI211_X1 U10978 ( .C1(n9893), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9895)
         );
  OAI211_X1 U10979 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9898)
         );
  AOI21_X1 U10980 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(n9924) );
  AOI22_X1 U10981 ( .A1(n9911), .A2(n9924), .B1(n5382), .B2(n9909), .ZN(
        P1_U3478) );
  OAI21_X1 U10982 ( .B1(n9903), .B2(n9902), .A(n9901), .ZN(n9904) );
  AOI21_X1 U10983 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  AND2_X1 U10984 ( .A1(n9908), .A2(n9907), .ZN(n9927) );
  INV_X1 U10985 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U10986 ( .A1(n9911), .A2(n9927), .B1(n9910), .B2(n9909), .ZN(
        P1_U3481) );
  AOI22_X1 U10987 ( .A1(n9928), .A2(n9912), .B1(n6630), .B2(n9925), .ZN(
        P1_U3524) );
  AOI22_X1 U10988 ( .A1(n9928), .A2(n9913), .B1(n6629), .B2(n9925), .ZN(
        P1_U3525) );
  INV_X1 U10989 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9914) );
  AOI22_X1 U10990 ( .A1(n9928), .A2(n9915), .B1(n9914), .B2(n9925), .ZN(
        P1_U3526) );
  INV_X1 U10991 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U10992 ( .A1(n9928), .A2(n9917), .B1(n9916), .B2(n9925), .ZN(
        P1_U3527) );
  INV_X1 U10993 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U10994 ( .A1(n9928), .A2(n9919), .B1(n9918), .B2(n9925), .ZN(
        P1_U3528) );
  AOI22_X1 U10995 ( .A1(n9928), .A2(n9920), .B1(n6636), .B2(n9925), .ZN(
        P1_U3529) );
  INV_X1 U10996 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9921) );
  AOI22_X1 U10997 ( .A1(n9928), .A2(n9922), .B1(n9921), .B2(n9925), .ZN(
        P1_U3530) );
  INV_X1 U10998 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9923) );
  AOI22_X1 U10999 ( .A1(n9928), .A2(n9924), .B1(n9923), .B2(n9925), .ZN(
        P1_U3531) );
  INV_X1 U11000 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U11001 ( .A1(n9928), .A2(n9927), .B1(n9926), .B2(n9925), .ZN(
        P1_U3532) );
  AOI22_X1 U11002 ( .A1(n9930), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9929), .ZN(n9940) );
  AOI22_X1 U11003 ( .A1(n9932), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9939) );
  OAI21_X1 U11004 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9934), .A(n9933), .ZN(
        n9937) );
  NOR2_X1 U11005 ( .A1(n9935), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9936) );
  OAI21_X1 U11006 ( .B1(n9937), .B2(n9936), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9938) );
  OAI211_X1 U11007 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9940), .A(n9939), .B(
        n9938), .ZN(P2_U3245) );
  INV_X1 U11008 ( .A(n9941), .ZN(n9942) );
  AND2_X1 U11009 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9946), .ZN(P2_U3297) );
  AND2_X1 U11010 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9946), .ZN(P2_U3298) );
  AND2_X1 U11011 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9946), .ZN(P2_U3299) );
  AND2_X1 U11012 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9946), .ZN(P2_U3300) );
  AND2_X1 U11013 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9946), .ZN(P2_U3301) );
  AND2_X1 U11014 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9946), .ZN(P2_U3302) );
  AND2_X1 U11015 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9946), .ZN(P2_U3303) );
  AND2_X1 U11016 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9946), .ZN(P2_U3304) );
  AND2_X1 U11017 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9946), .ZN(P2_U3305) );
  AND2_X1 U11018 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9946), .ZN(P2_U3306) );
  AND2_X1 U11019 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9946), .ZN(P2_U3307) );
  AND2_X1 U11020 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9946), .ZN(P2_U3308) );
  AND2_X1 U11021 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9946), .ZN(P2_U3309) );
  AND2_X1 U11022 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9946), .ZN(P2_U3310) );
  AND2_X1 U11023 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9946), .ZN(P2_U3311) );
  AND2_X1 U11024 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9946), .ZN(P2_U3312) );
  AND2_X1 U11025 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9946), .ZN(P2_U3313) );
  AND2_X1 U11026 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9946), .ZN(P2_U3314) );
  AND2_X1 U11027 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9946), .ZN(P2_U3315) );
  AND2_X1 U11028 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9946), .ZN(P2_U3316) );
  AND2_X1 U11029 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9946), .ZN(P2_U3317) );
  AND2_X1 U11030 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9946), .ZN(P2_U3318) );
  AND2_X1 U11031 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9946), .ZN(P2_U3319) );
  AND2_X1 U11032 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9946), .ZN(P2_U3320) );
  AND2_X1 U11033 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9946), .ZN(P2_U3321) );
  AND2_X1 U11034 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9946), .ZN(P2_U3322) );
  AND2_X1 U11035 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9946), .ZN(P2_U3323) );
  AND2_X1 U11036 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9946), .ZN(P2_U3324) );
  AND2_X1 U11037 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9946), .ZN(P2_U3325) );
  AND2_X1 U11038 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9946), .ZN(P2_U3326) );
  AOI22_X1 U11039 ( .A1(n9945), .A2(n9948), .B1(n9944), .B2(n9946), .ZN(
        P2_U3437) );
  AOI22_X1 U11040 ( .A1(n9949), .A2(n9948), .B1(n9947), .B2(n9946), .ZN(
        P2_U3438) );
  AOI22_X1 U11041 ( .A1(n9951), .A2(n10029), .B1(n4927), .B2(n9950), .ZN(n9952) );
  AND2_X1 U11042 ( .A1(n9953), .A2(n9952), .ZN(n10034) );
  INV_X1 U11043 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U11044 ( .A1(n10032), .A2(n10034), .B1(n9954), .B2(n10030), .ZN(
        P2_U3451) );
  OAI21_X1 U11045 ( .B1(n6818), .B2(n10022), .A(n9955), .ZN(n9958) );
  INV_X1 U11046 ( .A(n9956), .ZN(n9957) );
  AOI211_X1 U11047 ( .C1(n10029), .C2(n9959), .A(n9958), .B(n9957), .ZN(n10036) );
  INV_X1 U11048 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11049 ( .A1(n10032), .A2(n10036), .B1(n9960), .B2(n10030), .ZN(
        P2_U3454) );
  OAI21_X1 U11050 ( .B1(n6821), .B2(n10022), .A(n9961), .ZN(n9963) );
  AOI211_X1 U11051 ( .C1(n10029), .C2(n9964), .A(n9963), .B(n9962), .ZN(n10038) );
  INV_X1 U11052 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9965) );
  AOI22_X1 U11053 ( .A1(n10032), .A2(n10038), .B1(n9965), .B2(n10030), .ZN(
        P2_U3457) );
  OAI21_X1 U11054 ( .B1(n9967), .B2(n10022), .A(n9966), .ZN(n9970) );
  INV_X1 U11055 ( .A(n9968), .ZN(n9969) );
  AOI211_X1 U11056 ( .C1(n10010), .C2(n9971), .A(n9970), .B(n9969), .ZN(n10040) );
  INV_X1 U11057 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9972) );
  AOI22_X1 U11058 ( .A1(n10032), .A2(n10040), .B1(n9972), .B2(n10030), .ZN(
        P2_U3460) );
  AOI22_X1 U11059 ( .A1(n9974), .A2(n10014), .B1(n10013), .B2(n9973), .ZN(
        n9975) );
  NAND2_X1 U11060 ( .A1(n9976), .A2(n9975), .ZN(n9977) );
  AOI21_X1 U11061 ( .B1(n10029), .B2(n9978), .A(n9977), .ZN(n10042) );
  INV_X1 U11062 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11063 ( .A1(n10032), .A2(n10042), .B1(n9979), .B2(n10030), .ZN(
        P2_U3463) );
  OAI22_X1 U11064 ( .A1(n9981), .A2(n10024), .B1(n9980), .B2(n10022), .ZN(
        n9984) );
  INV_X1 U11065 ( .A(n9982), .ZN(n9983) );
  AOI211_X1 U11066 ( .C1(n9985), .C2(n10029), .A(n9984), .B(n9983), .ZN(n10043) );
  INV_X1 U11067 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U11068 ( .A1(n10032), .A2(n10043), .B1(n9986), .B2(n10030), .ZN(
        P2_U3469) );
  OAI21_X1 U11069 ( .B1(n10019), .B2(n9989), .A(n9988), .ZN(n9990) );
  INV_X1 U11070 ( .A(n9990), .ZN(n10045) );
  INV_X1 U11071 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11072 ( .A1(n10032), .A2(n10045), .B1(n9991), .B2(n10030), .ZN(
        P2_U3472) );
  OAI22_X1 U11073 ( .A1(n9993), .A2(n10024), .B1(n9992), .B2(n10022), .ZN(
        n9995) );
  AOI211_X1 U11074 ( .C1(n10010), .C2(n9996), .A(n9995), .B(n9994), .ZN(n10046) );
  INV_X1 U11075 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U11076 ( .A1(n10032), .A2(n10046), .B1(n9997), .B2(n10030), .ZN(
        P2_U3475) );
  OAI22_X1 U11077 ( .A1(n9999), .A2(n10024), .B1(n9998), .B2(n10022), .ZN(
        n10001) );
  AOI211_X1 U11078 ( .C1(n10010), .C2(n10002), .A(n10001), .B(n10000), .ZN(
        n10047) );
  INV_X1 U11079 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11080 ( .A1(n10032), .A2(n10047), .B1(n10003), .B2(n10030), .ZN(
        P2_U3478) );
  INV_X1 U11081 ( .A(n10004), .ZN(n10005) );
  OAI22_X1 U11082 ( .A1(n10006), .A2(n10024), .B1(n10005), .B2(n10022), .ZN(
        n10008) );
  AOI211_X1 U11083 ( .C1(n10010), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10048) );
  INV_X1 U11084 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10011) );
  AOI22_X1 U11085 ( .A1(n10032), .A2(n10048), .B1(n10011), .B2(n10030), .ZN(
        P2_U3481) );
  AOI22_X1 U11086 ( .A1(n10015), .A2(n10014), .B1(n10013), .B2(n10012), .ZN(
        n10016) );
  OAI211_X1 U11087 ( .C1(n10019), .C2(n10018), .A(n10017), .B(n10016), .ZN(
        n10020) );
  INV_X1 U11088 ( .A(n10020), .ZN(n10049) );
  INV_X1 U11089 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10021) );
  AOI22_X1 U11090 ( .A1(n10032), .A2(n10049), .B1(n10021), .B2(n10030), .ZN(
        P2_U3484) );
  OAI22_X1 U11091 ( .A1(n10025), .A2(n10024), .B1(n10023), .B2(n10022), .ZN(
        n10027) );
  AOI211_X1 U11092 ( .C1(n10029), .C2(n10028), .A(n10027), .B(n10026), .ZN(
        n10051) );
  INV_X1 U11093 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10031) );
  AOI22_X1 U11094 ( .A1(n10032), .A2(n10051), .B1(n10031), .B2(n10030), .ZN(
        P2_U3487) );
  INV_X1 U11095 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10033) );
  AOI22_X1 U11096 ( .A1(n10052), .A2(n10034), .B1(n10033), .B2(n10050), .ZN(
        P2_U3520) );
  INV_X1 U11097 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10035) );
  AOI22_X1 U11098 ( .A1(n10052), .A2(n10036), .B1(n10035), .B2(n10050), .ZN(
        P2_U3521) );
  INV_X1 U11099 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U11100 ( .A1(n10052), .A2(n10038), .B1(n10037), .B2(n10050), .ZN(
        P2_U3522) );
  INV_X1 U11101 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U11102 ( .A1(n10052), .A2(n10040), .B1(n10039), .B2(n10050), .ZN(
        P2_U3523) );
  INV_X1 U11103 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U11104 ( .A1(n10052), .A2(n10042), .B1(n10041), .B2(n10050), .ZN(
        P2_U3524) );
  AOI22_X1 U11105 ( .A1(n10052), .A2(n10043), .B1(n6710), .B2(n10050), .ZN(
        P2_U3526) );
  INV_X1 U11106 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U11107 ( .A1(n10052), .A2(n10045), .B1(n10044), .B2(n10050), .ZN(
        P2_U3527) );
  AOI22_X1 U11108 ( .A1(n10052), .A2(n10046), .B1(n6713), .B2(n10050), .ZN(
        P2_U3528) );
  AOI22_X1 U11109 ( .A1(n10052), .A2(n10047), .B1(n6714), .B2(n10050), .ZN(
        P2_U3529) );
  AOI22_X1 U11110 ( .A1(n10052), .A2(n10048), .B1(n6947), .B2(n10050), .ZN(
        P2_U3530) );
  AOI22_X1 U11111 ( .A1(n10052), .A2(n10049), .B1(n7090), .B2(n10050), .ZN(
        P2_U3531) );
  AOI22_X1 U11112 ( .A1(n10052), .A2(n10051), .B1(n7167), .B2(n10050), .ZN(
        P2_U3532) );
  NAND3_X1 U11113 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10062) );
  AOI21_X1 U11114 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10064) );
  INV_X1 U11115 ( .A(n10064), .ZN(n10053) );
  NAND2_X1 U11116 ( .A1(n10062), .A2(n10053), .ZN(n10054) );
  XOR2_X1 U11117 ( .A(n10063), .B(n10054), .Z(ADD_1071_U5) );
  XOR2_X1 U11118 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NOR2_X1 U11119 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10055) );
  AOI21_X1 U11120 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10055), .ZN(n10088) );
  NOR2_X1 U11121 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10056) );
  AOI21_X1 U11122 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10056), .ZN(n10091) );
  NOR2_X1 U11123 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10057) );
  AOI21_X1 U11124 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10057), .ZN(n10094) );
  NOR2_X1 U11125 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10058) );
  AOI21_X1 U11126 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10058), .ZN(n10097) );
  NOR2_X1 U11127 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10059) );
  AOI21_X1 U11128 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10059), .ZN(n10100) );
  NOR2_X1 U11129 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10070) );
  XOR2_X1 U11130 ( .A(n10060), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10509) );
  NAND2_X1 U11131 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10068) );
  XOR2_X1 U11132 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10507) );
  NAND2_X1 U11133 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10066) );
  XNOR2_X1 U11134 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n10061), .ZN(n10496) );
  OAI21_X1 U11135 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(n10495) );
  NAND2_X1 U11136 ( .A1(n10496), .A2(n10495), .ZN(n10065) );
  NAND2_X1 U11137 ( .A1(n10066), .A2(n10065), .ZN(n10506) );
  NAND2_X1 U11138 ( .A1(n10507), .A2(n10506), .ZN(n10067) );
  NAND2_X1 U11139 ( .A1(n10068), .A2(n10067), .ZN(n10508) );
  NOR2_X1 U11140 ( .A1(n10509), .A2(n10508), .ZN(n10069) );
  NOR2_X1 U11141 ( .A1(n10070), .A2(n10069), .ZN(n10071) );
  NOR2_X1 U11142 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10071), .ZN(n10498) );
  AND2_X1 U11143 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10071), .ZN(n10497) );
  NOR2_X1 U11144 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10497), .ZN(n10072) );
  NAND2_X1 U11145 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10073), .ZN(n10075) );
  XOR2_X1 U11146 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10073), .Z(n10505) );
  NAND2_X1 U11147 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10505), .ZN(n10074) );
  NAND2_X1 U11148 ( .A1(n10075), .A2(n10074), .ZN(n10076) );
  NAND2_X1 U11149 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10076), .ZN(n10078) );
  XOR2_X1 U11150 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10076), .Z(n10494) );
  NAND2_X1 U11151 ( .A1(n10494), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U11152 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  NAND2_X1 U11153 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10079), .ZN(n10081) );
  XOR2_X1 U11154 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10079), .Z(n10504) );
  NAND2_X1 U11155 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10504), .ZN(n10080) );
  NAND2_X1 U11156 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  AND2_X1 U11157 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10082), .ZN(n10083) );
  XNOR2_X1 U11158 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10082), .ZN(n10493) );
  NOR2_X1 U11159 ( .A1(n10493), .A2(n10492), .ZN(n10491) );
  NAND2_X1 U11160 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10084) );
  OAI21_X1 U11161 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10084), .ZN(n10108) );
  NAND2_X1 U11162 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10085) );
  OAI21_X1 U11163 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10085), .ZN(n10105) );
  NOR2_X1 U11164 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10086) );
  AOI21_X1 U11165 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10086), .ZN(n10102) );
  NAND2_X1 U11166 ( .A1(n10103), .A2(n10102), .ZN(n10101) );
  NAND2_X1 U11167 ( .A1(n10100), .A2(n10099), .ZN(n10098) );
  NAND2_X1 U11168 ( .A1(n10097), .A2(n10096), .ZN(n10095) );
  OAI21_X1 U11169 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10095), .ZN(n10093) );
  NAND2_X1 U11170 ( .A1(n10094), .A2(n10093), .ZN(n10092) );
  OAI21_X1 U11171 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10092), .ZN(n10090) );
  NAND2_X1 U11172 ( .A1(n10091), .A2(n10090), .ZN(n10089) );
  OAI21_X1 U11173 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10089), .ZN(n10087) );
  NAND2_X1 U11174 ( .A1(n10088), .A2(n10087), .ZN(n10484) );
  OAI21_X1 U11175 ( .B1(n10088), .B2(n10087), .A(n10484), .ZN(ADD_1071_U56) );
  OAI21_X1 U11176 ( .B1(n10091), .B2(n10090), .A(n10089), .ZN(ADD_1071_U57) );
  OAI21_X1 U11177 ( .B1(n10094), .B2(n10093), .A(n10092), .ZN(ADD_1071_U58) );
  OAI21_X1 U11178 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(ADD_1071_U59) );
  OAI21_X1 U11179 ( .B1(n10100), .B2(n10099), .A(n10098), .ZN(ADD_1071_U60) );
  OAI21_X1 U11180 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(ADD_1071_U61) );
  AOI21_X1 U11181 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(ADD_1071_U62) );
  AOI21_X1 U11182 ( .B1(n10109), .B2(n10108), .A(n10107), .ZN(ADD_1071_U63) );
  OAI22_X1 U11183 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_g89), .ZN(n10110) );
  AOI221_X1 U11184 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        keyinput_g89), .C2(P2_DATAO_REG_7__SCAN_IN), .A(n10110), .ZN(n10117)
         );
  OAI22_X1 U11185 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        keyinput_g61), .B2(P2_REG3_REG_6__SCAN_IN), .ZN(n10111) );
  AOI221_X1 U11186 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n10111), .ZN(n10116) );
  OAI22_X1 U11187 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_g100), .B1(
        keyinput_g84), .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n10112) );
  AOI221_X1 U11188 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_g100), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_g84), .A(n10112), .ZN(n10115)
         );
  OAI22_X1 U11189 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        keyinput_g28), .B2(SI_4_), .ZN(n10113) );
  AOI221_X1 U11190 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        SI_4_), .C2(keyinput_g28), .A(n10113), .ZN(n10114) );
  NAND4_X1 U11191 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10248) );
  OAI22_X1 U11192 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g30), .B2(SI_2_), .ZN(n10118) );
  AOI221_X1 U11193 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        SI_2_), .C2(keyinput_g30), .A(n10118), .ZN(n10143) );
  OAI22_X1 U11194 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_g119), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .ZN(n10119) );
  AOI221_X1 U11195 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_g119), .C1(
        keyinput_g54), .C2(P2_REG3_REG_0__SCAN_IN), .A(n10119), .ZN(n10122) );
  OAI22_X1 U11196 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        keyinput_g26), .B2(SI_6_), .ZN(n10120) );
  AOI221_X1 U11197 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        SI_6_), .C2(keyinput_g26), .A(n10120), .ZN(n10121) );
  OAI211_X1 U11198 ( .C1(n10375), .C2(keyinput_g10), .A(n10122), .B(n10121), 
        .ZN(n10123) );
  AOI21_X1 U11199 ( .B1(n10375), .B2(keyinput_g10), .A(n10123), .ZN(n10142) );
  AOI22_X1 U11200 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(SI_7_), 
        .B2(keyinput_g25), .ZN(n10124) );
  OAI221_X1 U11201 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(SI_7_), .C2(keyinput_g25), .A(n10124), .ZN(n10131) );
  AOI22_X1 U11202 ( .A1(SI_11_), .A2(keyinput_g21), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n10125) );
  OAI221_X1 U11203 ( .B1(SI_11_), .B2(keyinput_g21), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_g82), .A(n10125), .ZN(n10130)
         );
  AOI22_X1 U11204 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        SI_20_), .B2(keyinput_g12), .ZN(n10126) );
  OAI221_X1 U11205 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        SI_20_), .C2(keyinput_g12), .A(n10126), .ZN(n10129) );
  AOI22_X1 U11206 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        SI_15_), .B2(keyinput_g17), .ZN(n10127) );
  OAI221_X1 U11207 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        SI_15_), .C2(keyinput_g17), .A(n10127), .ZN(n10128) );
  NOR4_X1 U11208 ( .A1(n10131), .A2(n10130), .A3(n10129), .A4(n10128), .ZN(
        n10141) );
  AOI22_X1 U11209 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(SI_19_), .B2(keyinput_g13), .ZN(n10132) );
  OAI221_X1 U11210 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        SI_19_), .C2(keyinput_g13), .A(n10132), .ZN(n10139) );
  AOI22_X1 U11211 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_g120), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_g111), .ZN(n10133) );
  OAI221_X1 U11212 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_g120), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_g111), .A(n10133), .ZN(n10138) );
  AOI22_X1 U11213 ( .A1(SI_31_), .A2(keyinput_g1), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .ZN(n10134) );
  OAI221_X1 U11214 ( .B1(SI_31_), .B2(keyinput_g1), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_g76), .A(n10134), .ZN(n10137)
         );
  AOI22_X1 U11215 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_g66), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_g112), .ZN(n10135) );
  OAI221_X1 U11216 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_g112), .A(n10135), .ZN(n10136) );
  NOR4_X1 U11217 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10140) );
  NAND4_X1 U11218 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n10247) );
  AOI22_X1 U11219 ( .A1(n10145), .A2(keyinput_g23), .B1(keyinput_g36), .B2(
        n6204), .ZN(n10144) );
  OAI221_X1 U11220 ( .B1(n10145), .B2(keyinput_g23), .C1(n6204), .C2(
        keyinput_g36), .A(n10144), .ZN(n10156) );
  AOI22_X1 U11221 ( .A1(n10148), .A2(keyinput_g5), .B1(keyinput_g67), .B2(
        n10147), .ZN(n10146) );
  OAI221_X1 U11222 ( .B1(n10148), .B2(keyinput_g5), .C1(n10147), .C2(
        keyinput_g67), .A(n10146), .ZN(n10155) );
  AOI22_X1 U11223 ( .A1(n10458), .A2(keyinput_g43), .B1(n10150), .B2(
        keyinput_g68), .ZN(n10149) );
  OAI221_X1 U11224 ( .B1(n10458), .B2(keyinput_g43), .C1(n10150), .C2(
        keyinput_g68), .A(n10149), .ZN(n10154) );
  XNOR2_X1 U11225 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_g101), .ZN(n10152)
         );
  XNOR2_X1 U11226 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g91), .ZN(n10151) );
  NAND2_X1 U11227 ( .A1(n10152), .A2(n10151), .ZN(n10153) );
  NOR4_X1 U11228 ( .A1(n10156), .A2(n10155), .A3(n10154), .A4(n10153), .ZN(
        n10195) );
  AOI22_X1 U11229 ( .A1(n10417), .A2(keyinput_g125), .B1(keyinput_g73), .B2(
        n5176), .ZN(n10157) );
  OAI221_X1 U11230 ( .B1(n10417), .B2(keyinput_g125), .C1(n5176), .C2(
        keyinput_g73), .A(n10157), .ZN(n10167) );
  INV_X1 U11231 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U11232 ( .A1(n10159), .A2(keyinput_g109), .B1(keyinput_g74), .B2(
        n10392), .ZN(n10158) );
  OAI221_X1 U11233 ( .B1(n10159), .B2(keyinput_g109), .C1(n10392), .C2(
        keyinput_g74), .A(n10158), .ZN(n10166) );
  INV_X1 U11234 ( .A(SI_17_), .ZN(n10161) );
  AOI22_X1 U11235 ( .A1(n10161), .A2(keyinput_g15), .B1(n10372), .B2(
        keyinput_g72), .ZN(n10160) );
  OAI221_X1 U11236 ( .B1(n10161), .B2(keyinput_g15), .C1(n10372), .C2(
        keyinput_g72), .A(n10160), .ZN(n10165) );
  XNOR2_X1 U11237 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_g115), .ZN(n10163)
         );
  XNOR2_X1 U11238 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g96), .ZN(n10162) );
  NAND2_X1 U11239 ( .A1(n10163), .A2(n10162), .ZN(n10164) );
  NOR4_X1 U11240 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10194) );
  INV_X1 U11241 ( .A(SI_14_), .ZN(n10169) );
  INV_X1 U11242 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U11243 ( .A1(n10169), .A2(keyinput_g18), .B1(keyinput_g41), .B2(
        n10420), .ZN(n10168) );
  OAI221_X1 U11244 ( .B1(n10169), .B2(keyinput_g18), .C1(n10420), .C2(
        keyinput_g41), .A(n10168), .ZN(n10179) );
  AOI22_X1 U11245 ( .A1(n10171), .A2(keyinput_g70), .B1(keyinput_g34), .B2(
        P2_U3152), .ZN(n10170) );
  OAI221_X1 U11246 ( .B1(n10171), .B2(keyinput_g70), .C1(P2_U3152), .C2(
        keyinput_g34), .A(n10170), .ZN(n10178) );
  XNOR2_X1 U11247 ( .A(n10399), .B(keyinput_g127), .ZN(n10177) );
  XOR2_X1 U11248 ( .A(n10172), .B(keyinput_g64), .Z(n10175) );
  XNOR2_X1 U11249 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g116), .ZN(n10174)
         );
  XNOR2_X1 U11250 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_g117), .ZN(n10173)
         );
  NAND3_X1 U11251 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(n10176) );
  NOR4_X1 U11252 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10193) );
  AOI22_X1 U11253 ( .A1(n10182), .A2(keyinput_g62), .B1(n10181), .B2(
        keyinput_g69), .ZN(n10180) );
  OAI221_X1 U11254 ( .B1(n10182), .B2(keyinput_g62), .C1(n10181), .C2(
        keyinput_g69), .A(n10180), .ZN(n10191) );
  AOI22_X1 U11255 ( .A1(n10184), .A2(keyinput_g71), .B1(keyinput_g80), .B2(
        n10360), .ZN(n10183) );
  OAI221_X1 U11256 ( .B1(n10184), .B2(keyinput_g71), .C1(n10360), .C2(
        keyinput_g80), .A(n10183), .ZN(n10190) );
  XOR2_X1 U11257 ( .A(n5203), .B(keyinput_g4), .Z(n10188) );
  XNOR2_X1 U11258 ( .A(SI_3_), .B(keyinput_g29), .ZN(n10187) );
  XNOR2_X1 U11259 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g102), .ZN(n10186)
         );
  XNOR2_X1 U11260 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_g121), .ZN(n10185)
         );
  NAND4_X1 U11261 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10189) );
  NOR3_X1 U11262 ( .A1(n10191), .A2(n10190), .A3(n10189), .ZN(n10192) );
  NAND4_X1 U11263 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n10246) );
  AOI22_X1 U11264 ( .A1(n10430), .A2(keyinput_g108), .B1(keyinput_g123), .B2(
        n10361), .ZN(n10196) );
  OAI221_X1 U11265 ( .B1(n10430), .B2(keyinput_g108), .C1(n10361), .C2(
        keyinput_g123), .A(n10196), .ZN(n10206) );
  AOI22_X1 U11266 ( .A1(n10199), .A2(keyinput_g126), .B1(keyinput_g22), .B2(
        n10198), .ZN(n10197) );
  OAI221_X1 U11267 ( .B1(n10199), .B2(keyinput_g126), .C1(n10198), .C2(
        keyinput_g22), .A(n10197), .ZN(n10205) );
  XOR2_X1 U11268 ( .A(n10463), .B(keyinput_g63), .Z(n10203) );
  XNOR2_X1 U11269 ( .A(SI_16_), .B(keyinput_g16), .ZN(n10202) );
  XNOR2_X1 U11270 ( .A(SI_0_), .B(keyinput_g32), .ZN(n10201) );
  XNOR2_X1 U11271 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g92), .ZN(n10200) );
  NAND4_X1 U11272 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10204) );
  NOR3_X1 U11273 ( .A1(n10206), .A2(n10205), .A3(n10204), .ZN(n10244) );
  AOI22_X1 U11274 ( .A1(n10390), .A2(keyinput_g59), .B1(n5944), .B2(
        keyinput_g53), .ZN(n10207) );
  OAI221_X1 U11275 ( .B1(n10390), .B2(keyinput_g59), .C1(n5944), .C2(
        keyinput_g53), .A(n10207), .ZN(n10218) );
  INV_X1 U11276 ( .A(SI_26_), .ZN(n10373) );
  AOI22_X1 U11277 ( .A1(n10209), .A2(keyinput_g0), .B1(n10373), .B2(
        keyinput_g6), .ZN(n10208) );
  OAI221_X1 U11278 ( .B1(n10209), .B2(keyinput_g0), .C1(n10373), .C2(
        keyinput_g6), .A(n10208), .ZN(n10217) );
  AOI22_X1 U11279 ( .A1(n10212), .A2(keyinput_g20), .B1(keyinput_g38), .B2(
        n10211), .ZN(n10210) );
  OAI221_X1 U11280 ( .B1(n10212), .B2(keyinput_g20), .C1(n10211), .C2(
        keyinput_g38), .A(n10210), .ZN(n10216) );
  XNOR2_X1 U11281 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g122), .ZN(n10214)
         );
  XNOR2_X1 U11282 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_g46), .ZN(n10213)
         );
  NAND2_X1 U11283 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  NOR4_X1 U11284 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10243) );
  AOI22_X1 U11285 ( .A1(n6203), .A2(keyinput_g42), .B1(n10220), .B2(
        keyinput_g9), .ZN(n10219) );
  OAI221_X1 U11286 ( .B1(n6203), .B2(keyinput_g42), .C1(n10220), .C2(
        keyinput_g9), .A(n10219), .ZN(n10229) );
  AOI22_X1 U11287 ( .A1(n10462), .A2(keyinput_g39), .B1(n10222), .B2(
        keyinput_g60), .ZN(n10221) );
  OAI221_X1 U11288 ( .B1(n10462), .B2(keyinput_g39), .C1(n10222), .C2(
        keyinput_g60), .A(n10221), .ZN(n10228) );
  XNOR2_X1 U11289 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10226) );
  XNOR2_X1 U11290 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g98), .ZN(n10225) );
  XNOR2_X1 U11291 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g97), .ZN(n10224) );
  XNOR2_X1 U11292 ( .A(SI_13_), .B(keyinput_g19), .ZN(n10223) );
  NAND4_X1 U11293 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10227) );
  NOR3_X1 U11294 ( .A1(n10229), .A2(n10228), .A3(n10227), .ZN(n10242) );
  INV_X1 U11295 ( .A(SI_5_), .ZN(n10435) );
  AOI22_X1 U11296 ( .A1(n10435), .A2(keyinput_g27), .B1(n10432), .B2(
        keyinput_g77), .ZN(n10230) );
  OAI221_X1 U11297 ( .B1(n10435), .B2(keyinput_g27), .C1(n10432), .C2(
        keyinput_g77), .A(n10230), .ZN(n10240) );
  AOI22_X1 U11298 ( .A1(n10393), .A2(keyinput_g81), .B1(keyinput_g49), .B2(
        n10232), .ZN(n10231) );
  OAI221_X1 U11299 ( .B1(n10393), .B2(keyinput_g81), .C1(n10232), .C2(
        keyinput_g49), .A(n10231), .ZN(n10239) );
  AOI22_X1 U11300 ( .A1(n10429), .A2(keyinput_g55), .B1(n10234), .B2(
        keyinput_g103), .ZN(n10233) );
  OAI221_X1 U11301 ( .B1(n10429), .B2(keyinput_g55), .C1(n10234), .C2(
        keyinput_g103), .A(n10233), .ZN(n10238) );
  XNOR2_X1 U11302 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g118), .ZN(n10236)
         );
  XNOR2_X1 U11303 ( .A(SI_30_), .B(keyinput_g2), .ZN(n10235) );
  NAND2_X1 U11304 ( .A1(n10236), .A2(n10235), .ZN(n10237) );
  NOR4_X1 U11305 ( .A1(n10240), .A2(n10239), .A3(n10238), .A4(n10237), .ZN(
        n10241) );
  NAND4_X1 U11306 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10245) );
  NOR4_X1 U11307 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10287) );
  OAI22_X1 U11308 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g107), .B1(
        keyinput_g90), .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n10249) );
  AOI221_X1 U11309 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g107), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput_g90), .A(n10249), .ZN(n10256)
         );
  OAI22_X1 U11310 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g105), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n10250) );
  AOI221_X1 U11311 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g105), .C1(
        keyinput_g58), .C2(P2_REG3_REG_11__SCAN_IN), .A(n10250), .ZN(n10255)
         );
  OAI22_X1 U11312 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g104), .B1(
        keyinput_g14), .B2(SI_18_), .ZN(n10251) );
  AOI221_X1 U11313 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g104), .C1(
        SI_18_), .C2(keyinput_g14), .A(n10251), .ZN(n10254) );
  OAI22_X1 U11314 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_g106), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .ZN(n10252) );
  AOI221_X1 U11315 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_g106), .C1(
        keyinput_g52), .C2(P2_REG3_REG_4__SCAN_IN), .A(n10252), .ZN(n10253) );
  NAND4_X1 U11316 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n10285) );
  OAI22_X1 U11317 ( .A1(SI_21_), .A2(keyinput_g11), .B1(keyinput_g78), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n10257) );
  AOI221_X1 U11318 ( .B1(SI_21_), .B2(keyinput_g11), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_g78), .A(n10257), .ZN(n10264)
         );
  OAI22_X1 U11319 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n10258) );
  AOI221_X1 U11320 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        keyinput_g56), .C2(P2_REG3_REG_13__SCAN_IN), .A(n10258), .ZN(n10263)
         );
  OAI22_X1 U11321 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_g35), .B1(SI_29_), .B2(keyinput_g3), .ZN(n10259) );
  AOI221_X1 U11322 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_g35), .C1(
        keyinput_g3), .C2(SI_29_), .A(n10259), .ZN(n10262) );
  OAI22_X1 U11323 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g110), .B1(
        keyinput_g95), .B2(P1_IR_REG_4__SCAN_IN), .ZN(n10260) );
  AOI221_X1 U11324 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g110), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_g95), .A(n10260), .ZN(n10261) );
  NAND4_X1 U11325 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10284) );
  OAI22_X1 U11326 ( .A1(SI_25_), .A2(keyinput_g7), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .ZN(n10265) );
  AOI221_X1 U11327 ( .B1(SI_25_), .B2(keyinput_g7), .C1(keyinput_g65), .C2(
        P2_DATAO_REG_31__SCAN_IN), .A(n10265), .ZN(n10272) );
  OAI22_X1 U11328 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_g83), .B1(
        keyinput_g57), .B2(P2_REG3_REG_22__SCAN_IN), .ZN(n10266) );
  AOI221_X1 U11329 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n10266), .ZN(n10271)
         );
  OAI22_X1 U11330 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_g113), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n10267) );
  AOI221_X1 U11331 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_g113), .C1(
        keyinput_g48), .C2(P2_REG3_REG_16__SCAN_IN), .A(n10267), .ZN(n10270)
         );
  OAI22_X1 U11332 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_g114), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n10268) );
  AOI221_X1 U11333 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g33), .C2(P2_RD_REG_SCAN_IN), .A(n10268), .ZN(n10269) );
  NAND4_X1 U11334 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10283) );
  OAI22_X1 U11335 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g93), .B1(
        keyinput_g51), .B2(P2_REG3_REG_24__SCAN_IN), .ZN(n10273) );
  AOI221_X1 U11336 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g93), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n10273), .ZN(n10281)
         );
  OAI22_X1 U11337 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_g124), .B1(
        keyinput_g24), .B2(SI_8_), .ZN(n10274) );
  AOI221_X1 U11338 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_g124), .C1(SI_8_), 
        .C2(keyinput_g24), .A(n10274), .ZN(n10280) );
  OAI22_X1 U11339 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g94), .B1(SI_24_), 
        .B2(keyinput_g8), .ZN(n10275) );
  AOI221_X1 U11340 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g8), .C2(SI_24_), .A(n10275), .ZN(n10279) );
  OAI22_X1 U11341 ( .A1(n10277), .A2(keyinput_g37), .B1(keyinput_g99), .B2(
        P1_IR_REG_8__SCAN_IN), .ZN(n10276) );
  AOI221_X1 U11342 ( .B1(n10277), .B2(keyinput_g37), .C1(P1_IR_REG_8__SCAN_IN), 
        .C2(keyinput_g99), .A(n10276), .ZN(n10278) );
  NAND4_X1 U11343 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  NOR4_X1 U11344 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  AOI22_X1 U11345 ( .A1(n10287), .A2(n10286), .B1(keyinput_g45), .B2(n10483), 
        .ZN(n10482) );
  OAI22_X1 U11346 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_f69), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .ZN(n10288) );
  AOI221_X1 U11347 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .C1(
        keyinput_f87), .C2(P2_DATAO_REG_9__SCAN_IN), .A(n10288), .ZN(n10295)
         );
  OAI22_X1 U11348 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_f70), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .ZN(n10289) );
  AOI221_X1 U11349 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .C1(
        keyinput_f40), .C2(P2_REG3_REG_3__SCAN_IN), .A(n10289), .ZN(n10294) );
  OAI22_X1 U11350 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f126), .B1(
        keyinput_f64), .B2(P2_B_REG_SCAN_IN), .ZN(n10290) );
  AOI221_X1 U11351 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f126), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n10290), .ZN(n10293) );
  OAI22_X1 U11352 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f111), .B1(
        keyinput_f20), .B2(SI_12_), .ZN(n10291) );
  AOI221_X1 U11353 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f111), .C1(
        SI_12_), .C2(keyinput_f20), .A(n10291), .ZN(n10292) );
  NAND4_X1 U11354 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10323) );
  OAI22_X1 U11355 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_f113), .B1(
        keyinput_f11), .B2(SI_21_), .ZN(n10296) );
  AOI221_X1 U11356 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_f113), .C1(
        SI_21_), .C2(keyinput_f11), .A(n10296), .ZN(n10303) );
  OAI22_X1 U11357 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f109), .B1(
        keyinput_f25), .B2(SI_7_), .ZN(n10297) );
  AOI221_X1 U11358 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f109), .C1(SI_7_), .C2(keyinput_f25), .A(n10297), .ZN(n10302) );
  OAI22_X1 U11359 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_f98), .B1(
        keyinput_f49), .B2(P2_REG3_REG_5__SCAN_IN), .ZN(n10298) );
  AOI221_X1 U11360 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_f98), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n10298), .ZN(n10301) );
  OAI22_X1 U11361 ( .A1(SI_18_), .A2(keyinput_f14), .B1(keyinput_f36), .B2(
        P2_REG3_REG_27__SCAN_IN), .ZN(n10299) );
  AOI221_X1 U11362 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10299), .ZN(n10300)
         );
  NAND4_X1 U11363 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10322) );
  OAI22_X1 U11364 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_f91), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput_f116), .ZN(n10304) );
  AOI221_X1 U11365 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_f91), .C1(
        keyinput_f116), .C2(P1_IR_REG_25__SCAN_IN), .A(n10304), .ZN(n10311) );
  OAI22_X1 U11366 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f99), .B1(
        keyinput_f82), .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n10305) );
  AOI221_X1 U11367 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f99), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_f82), .A(n10305), .ZN(n10310)
         );
  OAI22_X1 U11368 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_f37), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n10306) );
  AOI221_X1 U11369 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .C1(
        keyinput_f46), .C2(P2_REG3_REG_12__SCAN_IN), .A(n10306), .ZN(n10309)
         );
  OAI22_X1 U11370 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_f106), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_f71), .ZN(n10307) );
  AOI221_X1 U11371 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_f106), .C1(
        keyinput_f71), .C2(P2_DATAO_REG_25__SCAN_IN), .A(n10307), .ZN(n10308)
         );
  NAND4_X1 U11372 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10321) );
  OAI22_X1 U11373 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_f73), .B1(
        SI_20_), .B2(keyinput_f12), .ZN(n10312) );
  AOI221_X1 U11374 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .C1(
        keyinput_f12), .C2(SI_20_), .A(n10312), .ZN(n10319) );
  OAI22_X1 U11375 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_f107), .B1(
        keyinput_f17), .B2(SI_15_), .ZN(n10313) );
  AOI221_X1 U11376 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_f107), .C1(
        SI_15_), .C2(keyinput_f17), .A(n10313), .ZN(n10318) );
  OAI22_X1 U11377 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f117), .B1(
        keyinput_f67), .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10314) );
  AOI221_X1 U11378 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f117), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_f67), .A(n10314), .ZN(n10317)
         );
  OAI22_X1 U11379 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f102), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10315) );
  AOI221_X1 U11380 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f102), .C1(
        keyinput_f62), .C2(P2_REG3_REG_26__SCAN_IN), .A(n10315), .ZN(n10316)
         );
  NAND4_X1 U11381 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10320) );
  NOR4_X1 U11382 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10479) );
  OAI22_X1 U11383 ( .A1(SI_0_), .A2(keyinput_f32), .B1(keyinput_f65), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n10324) );
  AOI221_X1 U11384 ( .B1(SI_0_), .B2(keyinput_f32), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_f65), .A(n10324), .ZN(n10331)
         );
  OAI22_X1 U11385 ( .A1(SI_8_), .A2(keyinput_f24), .B1(keyinput_f47), .B2(
        P2_REG3_REG_25__SCAN_IN), .ZN(n10325) );
  AOI221_X1 U11386 ( .B1(SI_8_), .B2(keyinput_f24), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n10325), .ZN(n10330)
         );
  OAI22_X1 U11387 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f97), .B1(SI_14_), 
        .B2(keyinput_f18), .ZN(n10326) );
  AOI221_X1 U11388 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f97), .C1(
        keyinput_f18), .C2(SI_14_), .A(n10326), .ZN(n10329) );
  OAI22_X1 U11389 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f120), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n10327) );
  AOI221_X1 U11390 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f120), .C1(
        keyinput_f61), .C2(P2_REG3_REG_6__SCAN_IN), .A(n10327), .ZN(n10328) );
  NAND4_X1 U11391 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10477) );
  OAI22_X1 U11392 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_f76), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n10332) );
  AOI221_X1 U11393 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .C1(
        keyinput_f48), .C2(P2_REG3_REG_16__SCAN_IN), .A(n10332), .ZN(n10358)
         );
  OAI22_X1 U11394 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n10333) );
  AOI221_X1 U11395 ( .B1(SI_11_), .B2(keyinput_f21), .C1(keyinput_f57), .C2(
        P2_REG3_REG_22__SCAN_IN), .A(n10333), .ZN(n10336) );
  OAI22_X1 U11396 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_f114), .B1(
        keyinput_f86), .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n10334) );
  AOI221_X1 U11397 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_f114), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_f86), .A(n10334), .ZN(n10335)
         );
  OAI211_X1 U11398 ( .C1(n10338), .C2(keyinput_f44), .A(n10336), .B(n10335), 
        .ZN(n10337) );
  AOI21_X1 U11399 ( .B1(n10338), .B2(keyinput_f44), .A(n10337), .ZN(n10357) );
  AOI22_X1 U11400 ( .A1(SI_16_), .A2(keyinput_f16), .B1(P1_IR_REG_3__SCAN_IN), 
        .B2(keyinput_f94), .ZN(n10339) );
  OAI221_X1 U11401 ( .B1(SI_16_), .B2(keyinput_f16), .C1(P1_IR_REG_3__SCAN_IN), 
        .C2(keyinput_f94), .A(n10339), .ZN(n10346) );
  AOI22_X1 U11402 ( .A1(SI_9_), .A2(keyinput_f23), .B1(P1_IR_REG_27__SCAN_IN), 
        .B2(keyinput_f118), .ZN(n10340) );
  OAI221_X1 U11403 ( .B1(SI_9_), .B2(keyinput_f23), .C1(P1_IR_REG_27__SCAN_IN), 
        .C2(keyinput_f118), .A(n10340), .ZN(n10345) );
  AOI22_X1 U11404 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_f68), .B1(
        SI_17_), .B2(keyinput_f15), .ZN(n10341) );
  OAI221_X1 U11405 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .C1(
        SI_17_), .C2(keyinput_f15), .A(n10341), .ZN(n10344) );
  AOI22_X1 U11406 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f96), .ZN(n10342) );
  OAI221_X1 U11407 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_f96), .A(n10342), .ZN(n10343) );
  NOR4_X1 U11408 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10356) );
  AOI22_X1 U11409 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P1_IR_REG_4__SCAN_IN), 
        .B2(keyinput_f95), .ZN(n10347) );
  OAI221_X1 U11410 ( .B1(SI_23_), .B2(keyinput_f9), .C1(P1_IR_REG_4__SCAN_IN), 
        .C2(keyinput_f95), .A(n10347), .ZN(n10354) );
  AOI22_X1 U11411 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_f79), .B1(
        SI_19_), .B2(keyinput_f13), .ZN(n10348) );
  OAI221_X1 U11412 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .C1(
        SI_19_), .C2(keyinput_f13), .A(n10348), .ZN(n10353) );
  AOI22_X1 U11413 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .ZN(n10349) );
  OAI221_X1 U11414 ( .B1(SI_31_), .B2(keyinput_f1), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_f88), .A(n10349), .ZN(n10352)
         );
  AOI22_X1 U11415 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n10350) );
  OAI221_X1 U11416 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n10350), .ZN(n10351) );
  NOR4_X1 U11417 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10355) );
  NAND4_X1 U11418 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10476) );
  AOI22_X1 U11419 ( .A1(n10361), .A2(keyinput_f123), .B1(keyinput_f80), .B2(
        n10360), .ZN(n10359) );
  OAI221_X1 U11420 ( .B1(n10361), .B2(keyinput_f123), .C1(n10360), .C2(
        keyinput_f80), .A(n10359), .ZN(n10370) );
  XNOR2_X1 U11421 ( .A(SI_10_), .B(keyinput_f22), .ZN(n10369) );
  XNOR2_X1 U11422 ( .A(keyinput_f35), .B(n10362), .ZN(n10368) );
  XNOR2_X1 U11423 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f92), .ZN(n10366) );
  XNOR2_X1 U11424 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_f121), .ZN(n10365)
         );
  XNOR2_X1 U11425 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_f115), .ZN(n10364)
         );
  XNOR2_X1 U11426 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_f119), .ZN(n10363)
         );
  NAND4_X1 U11427 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10367) );
  NOR4_X1 U11428 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10415) );
  AOI22_X1 U11429 ( .A1(n10373), .A2(keyinput_f6), .B1(keyinput_f72), .B2(
        n10372), .ZN(n10371) );
  OAI221_X1 U11430 ( .B1(n10373), .B2(keyinput_f6), .C1(n10372), .C2(
        keyinput_f72), .A(n10371), .ZN(n10383) );
  INV_X1 U11431 ( .A(SI_6_), .ZN(n10376) );
  AOI22_X1 U11432 ( .A1(n10376), .A2(keyinput_f26), .B1(n10375), .B2(
        keyinput_f10), .ZN(n10374) );
  OAI221_X1 U11433 ( .B1(n10376), .B2(keyinput_f26), .C1(n10375), .C2(
        keyinput_f10), .A(n10374), .ZN(n10382) );
  XNOR2_X1 U11434 ( .A(SI_2_), .B(keyinput_f30), .ZN(n10380) );
  XNOR2_X1 U11435 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_f90), .ZN(n10379)
         );
  XNOR2_X1 U11436 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f105), .ZN(n10378)
         );
  XNOR2_X1 U11437 ( .A(SI_27_), .B(keyinput_f5), .ZN(n10377) );
  NAND4_X1 U11438 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  NOR3_X1 U11439 ( .A1(n10383), .A2(n10382), .A3(n10381), .ZN(n10414) );
  AOI22_X1 U11440 ( .A1(n10385), .A2(keyinput_f50), .B1(keyinput_f54), .B2(
        n7222), .ZN(n10384) );
  OAI221_X1 U11441 ( .B1(n10385), .B2(keyinput_f50), .C1(n7222), .C2(
        keyinput_f54), .A(n10384), .ZN(n10397) );
  AOI22_X1 U11442 ( .A1(n10387), .A2(keyinput_f83), .B1(keyinput_f53), .B2(
        n5944), .ZN(n10386) );
  OAI221_X1 U11443 ( .B1(n10387), .B2(keyinput_f83), .C1(n5944), .C2(
        keyinput_f53), .A(n10386), .ZN(n10396) );
  AOI22_X1 U11444 ( .A1(n10390), .A2(keyinput_f59), .B1(n10389), .B2(
        keyinput_f78), .ZN(n10388) );
  OAI221_X1 U11445 ( .B1(n10390), .B2(keyinput_f59), .C1(n10389), .C2(
        keyinput_f78), .A(n10388), .ZN(n10395) );
  AOI22_X1 U11446 ( .A1(n10393), .A2(keyinput_f81), .B1(n10392), .B2(
        keyinput_f74), .ZN(n10391) );
  OAI221_X1 U11447 ( .B1(n10393), .B2(keyinput_f81), .C1(n10392), .C2(
        keyinput_f74), .A(n10391), .ZN(n10394) );
  NOR4_X1 U11448 ( .A1(n10397), .A2(n10396), .A3(n10395), .A4(n10394), .ZN(
        n10413) );
  AOI22_X1 U11449 ( .A1(n10400), .A2(keyinput_f51), .B1(n10399), .B2(
        keyinput_f127), .ZN(n10398) );
  OAI221_X1 U11450 ( .B1(n10400), .B2(keyinput_f51), .C1(n10399), .C2(
        keyinput_f127), .A(n10398), .ZN(n10411) );
  INV_X1 U11451 ( .A(keyinput_f0), .ZN(n10402) );
  AOI22_X1 U11452 ( .A1(n10403), .A2(keyinput_f52), .B1(P2_WR_REG_SCAN_IN), 
        .B2(n10402), .ZN(n10401) );
  OAI221_X1 U11453 ( .B1(n10403), .B2(keyinput_f52), .C1(n10402), .C2(
        P2_WR_REG_SCAN_IN), .A(n10401), .ZN(n10410) );
  AOI22_X1 U11454 ( .A1(n10405), .A2(keyinput_f89), .B1(keyinput_f34), .B2(
        P2_U3152), .ZN(n10404) );
  OAI221_X1 U11455 ( .B1(n10405), .B2(keyinput_f89), .C1(P2_U3152), .C2(
        keyinput_f34), .A(n10404), .ZN(n10409) );
  XNOR2_X1 U11456 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f101), .ZN(n10407)
         );
  XNOR2_X1 U11457 ( .A(SI_30_), .B(keyinput_f2), .ZN(n10406) );
  NAND2_X1 U11458 ( .A1(n10407), .A2(n10406), .ZN(n10408) );
  NOR4_X1 U11459 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10412) );
  NAND4_X1 U11460 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10475) );
  AOI22_X1 U11461 ( .A1(n5203), .A2(keyinput_f4), .B1(n10417), .B2(
        keyinput_f125), .ZN(n10416) );
  OAI221_X1 U11462 ( .B1(n5203), .B2(keyinput_f4), .C1(n10417), .C2(
        keyinput_f125), .A(n10416), .ZN(n10427) );
  AOI22_X1 U11463 ( .A1(n10420), .A2(keyinput_f41), .B1(n10419), .B2(
        keyinput_f84), .ZN(n10418) );
  OAI221_X1 U11464 ( .B1(n10420), .B2(keyinput_f41), .C1(n10419), .C2(
        keyinput_f84), .A(n10418), .ZN(n10426) );
  XNOR2_X1 U11465 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10424) );
  XNOR2_X1 U11466 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f122), .ZN(n10423)
         );
  XNOR2_X1 U11467 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_f75), .ZN(n10422) );
  XNOR2_X1 U11468 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10421) );
  NAND4_X1 U11469 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10425) );
  NOR3_X1 U11470 ( .A1(n10427), .A2(n10426), .A3(n10425), .ZN(n10473) );
  AOI22_X1 U11471 ( .A1(n10430), .A2(keyinput_f108), .B1(keyinput_f55), .B2(
        n10429), .ZN(n10428) );
  OAI221_X1 U11472 ( .B1(n10430), .B2(keyinput_f108), .C1(n10429), .C2(
        keyinput_f55), .A(n10428), .ZN(n10442) );
  AOI22_X1 U11473 ( .A1(n10432), .A2(keyinput_f77), .B1(n5081), .B2(
        keyinput_f33), .ZN(n10431) );
  OAI221_X1 U11474 ( .B1(n10432), .B2(keyinput_f77), .C1(n5081), .C2(
        keyinput_f33), .A(n10431), .ZN(n10441) );
  AOI22_X1 U11475 ( .A1(n10435), .A2(keyinput_f27), .B1(n10434), .B2(
        keyinput_f112), .ZN(n10433) );
  OAI221_X1 U11476 ( .B1(n10435), .B2(keyinput_f27), .C1(n10434), .C2(
        keyinput_f112), .A(n10433), .ZN(n10440) );
  AOI22_X1 U11477 ( .A1(n10438), .A2(keyinput_f85), .B1(n10437), .B2(
        keyinput_f104), .ZN(n10436) );
  OAI221_X1 U11478 ( .B1(n10438), .B2(keyinput_f85), .C1(n10437), .C2(
        keyinput_f104), .A(n10436), .ZN(n10439) );
  NOR4_X1 U11479 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10472) );
  AOI22_X1 U11480 ( .A1(n5205), .A2(keyinput_f3), .B1(n6553), .B2(
        keyinput_f124), .ZN(n10443) );
  OAI221_X1 U11481 ( .B1(n5205), .B2(keyinput_f3), .C1(n6553), .C2(
        keyinput_f124), .A(n10443), .ZN(n10454) );
  AOI22_X1 U11482 ( .A1(n10446), .A2(keyinput_f8), .B1(keyinput_f66), .B2(
        n10445), .ZN(n10444) );
  OAI221_X1 U11483 ( .B1(n10446), .B2(keyinput_f8), .C1(n10445), .C2(
        keyinput_f66), .A(n10444), .ZN(n10453) );
  INV_X1 U11484 ( .A(SI_4_), .ZN(n10448) );
  AOI22_X1 U11485 ( .A1(n5556), .A2(keyinput_f110), .B1(keyinput_f28), .B2(
        n10448), .ZN(n10447) );
  OAI221_X1 U11486 ( .B1(n5556), .B2(keyinput_f110), .C1(n10448), .C2(
        keyinput_f28), .A(n10447), .ZN(n10452) );
  XNOR2_X1 U11487 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_f100), .ZN(n10450)
         );
  XNOR2_X1 U11488 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_f38), .ZN(n10449)
         );
  NAND2_X1 U11489 ( .A1(n10450), .A2(n10449), .ZN(n10451) );
  NOR4_X1 U11490 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10471) );
  AOI22_X1 U11491 ( .A1(n10456), .A2(keyinput_f19), .B1(keyinput_f56), .B2(
        n7327), .ZN(n10455) );
  OAI221_X1 U11492 ( .B1(n10456), .B2(keyinput_f19), .C1(n7327), .C2(
        keyinput_f56), .A(n10455), .ZN(n10469) );
  AOI22_X1 U11493 ( .A1(n10459), .A2(keyinput_f58), .B1(keyinput_f43), .B2(
        n10458), .ZN(n10457) );
  OAI221_X1 U11494 ( .B1(n10459), .B2(keyinput_f58), .C1(n10458), .C2(
        keyinput_f43), .A(n10457), .ZN(n10468) );
  AOI22_X1 U11495 ( .A1(n10462), .A2(keyinput_f39), .B1(n10461), .B2(
        keyinput_f7), .ZN(n10460) );
  OAI221_X1 U11496 ( .B1(n10462), .B2(keyinput_f39), .C1(n10461), .C2(
        keyinput_f7), .A(n10460), .ZN(n10467) );
  XOR2_X1 U11497 ( .A(n10463), .B(keyinput_f63), .Z(n10465) );
  XNOR2_X1 U11498 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f93), .ZN(n10464) );
  NAND2_X1 U11499 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  NOR4_X1 U11500 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10470) );
  NAND4_X1 U11501 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10474) );
  NOR4_X1 U11502 ( .A1(n10477), .A2(n10476), .A3(n10475), .A4(n10474), .ZN(
        n10478) );
  AOI22_X1 U11503 ( .A1(n10479), .A2(n10478), .B1(keyinput_f45), .B2(
        P2_REG3_REG_21__SCAN_IN), .ZN(n10480) );
  OAI21_X1 U11504 ( .B1(keyinput_f45), .B2(P2_REG3_REG_21__SCAN_IN), .A(n10480), .ZN(n10481) );
  OAI211_X1 U11505 ( .C1(keyinput_g45), .C2(n10483), .A(n10482), .B(n10481), 
        .ZN(n10490) );
  OAI21_X1 U11506 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10484), .ZN(n10501) );
  NOR2_X1 U11507 ( .A1(n10502), .A2(n10501), .ZN(n10485) );
  NAND2_X1 U11508 ( .A1(n10502), .A2(n10501), .ZN(n10500) );
  OAI21_X1 U11509 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10485), .A(n10500), 
        .ZN(n10488) );
  XNOR2_X1 U11510 ( .A(n10486), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n10487) );
  XNOR2_X1 U11511 ( .A(n10488), .B(n10487), .ZN(n10489) );
  XNOR2_X1 U11512 ( .A(n10490), .B(n10489), .ZN(ADD_1071_U4) );
  AOI21_X1 U11513 ( .B1(n10493), .B2(n10492), .A(n10491), .ZN(ADD_1071_U47) );
  XOR2_X1 U11514 ( .A(n10494), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11515 ( .A(n10496), .B(n10495), .Z(ADD_1071_U54) );
  NOR2_X1 U11516 ( .A1(n10498), .A2(n10497), .ZN(n10499) );
  XOR2_X1 U11517 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10499), .Z(ADD_1071_U51) );
  OAI21_X1 U11518 ( .B1(n10502), .B2(n10501), .A(n10500), .ZN(n10503) );
  XNOR2_X1 U11519 ( .A(n10503), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11520 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10504), .Z(ADD_1071_U48) );
  XOR2_X1 U11521 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10505), .Z(ADD_1071_U50) );
  XOR2_X1 U11522 ( .A(n10507), .B(n10506), .Z(ADD_1071_U53) );
  XNOR2_X1 U11523 ( .A(n10509), .B(n10508), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4988 ( .A(n5797), .Z(n6211) );
  CLKBUF_X1 U4989 ( .A(n5851), .Z(n6261) );
  CLKBUF_X1 U4995 ( .A(n8376), .Z(n4481) );
  CLKBUF_X1 U5002 ( .A(n5350), .Z(n6564) );
  CLKBUF_X3 U5022 ( .A(n5285), .Z(n6563) );
  NAND2_X1 U5379 ( .A1(n9777), .A2(n8287), .ZN(n8216) );
  NAND2_X2 U6188 ( .A1(n5035), .A2(n5034), .ZN(n7856) );
endmodule

