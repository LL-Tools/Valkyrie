

module b20_C_AntiSAT_k_128_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188;

  OR2_X1 U4829 ( .A1(n8195), .A2(n8036), .ZN(n5701) );
  AND2_X1 U4830 ( .A1(n5473), .A2(n5472), .ZN(n8036) );
  INV_X1 U4831 ( .A(n7965), .ZN(n8215) );
  AND4_X1 U4832 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n8278)
         );
  INV_X1 U4833 ( .A(n4324), .ZN(n5547) );
  INV_X4 U4834 ( .A(n6626), .ZN(n6895) );
  INV_X2 U4835 ( .A(n6185), .ZN(n6608) );
  AND2_X1 U4836 ( .A1(n5779), .A2(n5855), .ZN(n6718) );
  INV_X2 U4837 ( .A(n5470), .ZN(n5550) );
  BUF_X1 U4838 ( .A(n5023), .Z(n4324) );
  NOR2_X1 U4839 ( .A1(n6047), .A2(n6048), .ZN(n6075) );
  CLKBUF_X3 U4840 ( .A(n5145), .Z(n4325) );
  NAND2_X1 U4841 ( .A1(n6718), .A2(n6726), .ZN(n5781) );
  NAND2_X1 U4842 ( .A1(n5781), .A2(n6724), .ZN(n6586) );
  BUF_X1 U4843 ( .A(n6626), .Z(n8764) );
  INV_X2 U4844 ( .A(n8761), .ZN(n8695) );
  INV_X1 U4846 ( .A(n8074), .ZN(n7261) );
  NAND2_X1 U4847 ( .A1(n8164), .A2(n5500), .ZN(n7865) );
  NAND2_X1 U4848 ( .A1(n5772), .A2(n5771), .ZN(n4997) );
  OR2_X1 U4849 ( .A1(n5499), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8164) );
  OR2_X1 U4850 ( .A1(n8522), .A2(n8325), .ZN(n8289) );
  NAND2_X1 U4851 ( .A1(n5304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5305) );
  INV_X1 U4852 ( .A(n8677), .ZN(n8758) );
  AND2_X1 U4853 ( .A1(n5492), .A2(n5491), .ZN(n7868) );
  NAND2_X1 U4854 ( .A1(n5499), .A2(n5487), .ZN(n8182) );
  AND4_X1 U4855 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n6856)
         );
  NAND2_X1 U4856 ( .A1(n8960), .A2(n8963), .ZN(n9051) );
  INV_X1 U4857 ( .A(n6509), .ZN(n8077) );
  INV_X1 U4858 ( .A(n5971), .ZN(n7877) );
  OAI21_X1 U4859 ( .B1(n9340), .B2(n6367), .A(n6359), .ZN(n9177) );
  OR2_X1 U4860 ( .A1(n9767), .A2(n7072), .ZN(n9760) );
  INV_X2 U4861 ( .A(n9470), .ZN(n9767) );
  INV_X2 U4862 ( .A(n5145), .ZN(n6070) );
  INV_X1 U4863 ( .A(n5015), .ZN(n5470) );
  OAI21_X2 U4864 ( .B1(n7916), .B2(n4920), .A(n4919), .ZN(n4918) );
  NAND2_X2 U4865 ( .A1(n7756), .A2(n5814), .ZN(n7916) );
  NAND2_X2 U4866 ( .A1(n7538), .A2(n4357), .ZN(n7756) );
  INV_X2 U4867 ( .A(n8216), .ZN(n8248) );
  NAND2_X2 U4868 ( .A1(n6160), .A2(n6159), .ZN(n9746) );
  OAI21_X2 U4869 ( .B1(n7124), .B2(n4725), .A(n6427), .ZN(n7237) );
  AND4_X2 U4871 ( .A1(n5004), .A2(n5047), .A3(n4952), .A4(n4951), .ZN(n5067)
         );
  AND2_X2 U4872 ( .A1(n9101), .A2(n9103), .ZN(n9166) );
  NAND2_X2 U4873 ( .A1(n7971), .A2(n7970), .ZN(n7969) );
  NOR2_X2 U4874 ( .A1(n7901), .A2(n4455), .ZN(n7971) );
  NAND2_X2 U4875 ( .A1(n5841), .A2(n7985), .ZN(n7988) );
  OAI21_X2 U4876 ( .B1(n5173), .B2(n5172), .A(n5176), .ZN(n5203) );
  AND2_X1 U4877 ( .A1(n6047), .A2(n6048), .ZN(n6394) );
  XNOR2_X2 U4878 ( .A(n6041), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6047) );
  XNOR2_X2 U4879 ( .A(n5305), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6556) );
  CLKBUF_X1 U4880 ( .A(n5023), .Z(n4323) );
  XNOR2_X2 U4881 ( .A(n6107), .B(n6092), .ZN(n6685) );
  AOI21_X1 U4882 ( .B1(n5719), .B2(n5718), .A(n5717), .ZN(n5751) );
  XNOR2_X1 U4883 ( .A(n6551), .B(n6507), .ZN(n8175) );
  NOR3_X2 U4884 ( .A1(n9390), .A2(n9504), .A3(n4585), .ZN(n4582) );
  OAI21_X1 U4885 ( .B1(n8356), .B2(n5637), .A(n5647), .ZN(n8346) );
  NAND2_X2 U4886 ( .A1(n8289), .A2(n5668), .ZN(n8309) );
  NAND2_X1 U4887 ( .A1(n6434), .A2(n9125), .ZN(n7525) );
  NAND2_X1 U4888 ( .A1(n5322), .A2(n5321), .ZN(n8522) );
  OR2_X1 U4889 ( .A1(n8600), .A2(n8599), .ZN(n4327) );
  NAND2_X1 U4890 ( .A1(n6208), .A2(n6207), .ZN(n9785) );
  NAND2_X1 U4891 ( .A1(n6426), .A2(n9108), .ZN(n7124) );
  AND4_X1 U4892 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n8325)
         );
  AND2_X1 U4893 ( .A1(n4339), .A2(n4326), .ZN(n6893) );
  NAND2_X1 U4894 ( .A1(n6914), .A2(n6913), .ZN(n6912) );
  AND2_X1 U4895 ( .A1(n4454), .A2(n5787), .ZN(n6914) );
  NAND2_X1 U4896 ( .A1(n9110), .A2(n6420), .ZN(n6419) );
  CLKBUF_X2 U4897 ( .A(n5788), .Z(n5850) );
  NOR2_X2 U4898 ( .A1(n6932), .A2(n6926), .ZN(n6940) );
  NAND2_X2 U4899 ( .A1(n7210), .A2(n9865), .ZN(n5592) );
  CLKBUF_X2 U4900 ( .A(n6627), .Z(n8677) );
  INV_X2 U4901 ( .A(n6395), .ZN(n9013) );
  INV_X1 U4902 ( .A(n4344), .ZN(n4345) );
  AND2_X1 U4903 ( .A1(n6154), .A2(n6028), .ZN(n6255) );
  INV_X4 U4904 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9610) );
  AOI211_X1 U4905 ( .C1(n9488), .C2(n9470), .A(n9287), .B(n9286), .ZN(n9288)
         );
  OAI21_X1 U4906 ( .B1(n4843), .B2(n4735), .A(n6499), .ZN(n6503) );
  AOI21_X1 U4907 ( .B1(n4660), .B2(n9158), .A(n4659), .ZN(n4658) );
  OAI21_X1 U4908 ( .B1(n8723), .B2(n8767), .A(n8905), .ZN(n8729) );
  AND2_X1 U4909 ( .A1(n9102), .A2(n4458), .ZN(n4659) );
  OR2_X1 U4910 ( .A1(n8767), .A2(n4451), .ZN(n4450) );
  NAND2_X1 U4911 ( .A1(n4759), .A2(n4757), .ZN(n8767) );
  NAND2_X1 U4912 ( .A1(n8798), .A2(n8704), .ZN(n8904) );
  NAND2_X1 U4913 ( .A1(n8799), .A2(n8800), .ZN(n8798) );
  AOI21_X1 U4914 ( .B1(n7852), .B2(n8392), .A(n7851), .ZN(n8417) );
  NAND2_X1 U4915 ( .A1(n8830), .A2(n8692), .ZN(n8799) );
  OAI21_X1 U4916 ( .B1(n6552), .B2(n4380), .A(n4609), .ZN(n4608) );
  NAND2_X1 U4917 ( .A1(n5474), .A2(n5701), .ZN(n8176) );
  NAND2_X1 U4918 ( .A1(n4334), .A2(n4449), .ZN(n8871) );
  AND2_X1 U4919 ( .A1(n6599), .A2(n6598), .ZN(n9481) );
  NAND2_X1 U4920 ( .A1(n8741), .A2(n8743), .ZN(n8683) );
  OAI22_X1 U4921 ( .A1(n8675), .A2(n4336), .B1(n8674), .B2(n4335), .ZN(n8741)
         );
  NAND2_X1 U4922 ( .A1(n6601), .A2(n6600), .ZN(n9260) );
  INV_X1 U4923 ( .A(n8675), .ZN(n4334) );
  NAND2_X1 U4924 ( .A1(n8675), .A2(n8674), .ZN(n8870) );
  OAI222_X1 U4925 ( .A1(n8389), .A2(n8248), .B1(n8387), .B2(n8279), .C1(n8323), 
        .C2(n8247), .ZN(n8502) );
  NAND2_X1 U4926 ( .A1(n8853), .A2(n8852), .ZN(n8663) );
  OR2_X1 U4927 ( .A1(n8183), .A2(n8191), .ZN(n6548) );
  NAND2_X1 U4928 ( .A1(n8645), .A2(n8644), .ZN(n8647) );
  NAND2_X1 U4929 ( .A1(n6393), .A2(n6392), .ZN(n8773) );
  INV_X1 U4930 ( .A(n4333), .ZN(n4332) );
  NAND2_X1 U4931 ( .A1(n5424), .A2(n5423), .ZN(n8220) );
  OAI21_X1 U4932 ( .B1(n8644), .B2(n4766), .A(n4763), .ZN(n4333) );
  AND2_X1 U4933 ( .A1(n5411), .A2(n5410), .ZN(n8501) );
  NOR2_X1 U4934 ( .A1(n4449), .A2(n8872), .ZN(n4336) );
  NAND2_X1 U4935 ( .A1(n8308), .A2(n4947), .ZN(n8292) );
  NAND2_X1 U4936 ( .A1(n8310), .A2(n8309), .ZN(n8308) );
  INV_X1 U4937 ( .A(n8872), .ZN(n4335) );
  NAND2_X1 U4938 ( .A1(n4328), .A2(n4327), .ZN(n8862) );
  AND2_X1 U4939 ( .A1(n5680), .A2(n5681), .ZN(n8243) );
  NAND2_X1 U4940 ( .A1(n8046), .A2(n4456), .ZN(n7944) );
  NAND2_X1 U4941 ( .A1(n4330), .A2(n4329), .ZN(n4328) );
  OR2_X2 U4942 ( .A1(n9407), .A2(n9530), .ZN(n9390) );
  NAND2_X1 U4943 ( .A1(n4752), .A2(n4331), .ZN(n4330) );
  AND2_X1 U4944 ( .A1(n4753), .A2(n4751), .ZN(n4331) );
  NOR2_X1 U4945 ( .A1(n9459), .A2(n9545), .ZN(n9444) );
  AND2_X1 U4946 ( .A1(n5453), .A2(n5452), .ZN(n7965) );
  NAND2_X1 U4947 ( .A1(n5307), .A2(n5306), .ZN(n8518) );
  INV_X1 U4948 ( .A(n8789), .ZN(n4329) );
  AOI21_X1 U4949 ( .B1(n4744), .B2(n4747), .A(n4400), .ZN(n4741) );
  NOR2_X2 U4950 ( .A1(n9737), .A2(n9785), .ZN(n7530) );
  XNOR2_X1 U4951 ( .A(n5272), .B(n5255), .ZN(n6908) );
  NAND2_X1 U4952 ( .A1(n7313), .A2(n8890), .ZN(n9737) );
  AND2_X1 U4953 ( .A1(n4771), .A2(n7350), .ZN(n4342) );
  NAND2_X1 U4954 ( .A1(n7259), .A2(n5801), .ZN(n8021) );
  INV_X1 U4955 ( .A(n4747), .ZN(n4746) );
  NOR2_X1 U4956 ( .A1(n8843), .A2(n4340), .ZN(n6970) );
  OAI21_X1 U4957 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7710), .A(n7709), .ZN(
        n9678) );
  NAND2_X1 U4958 ( .A1(n8840), .A2(n4375), .ZN(n7350) );
  OR2_X1 U4959 ( .A1(n7285), .A2(n7284), .ZN(n8840) );
  AND2_X1 U4960 ( .A1(n6965), .A2(n4341), .ZN(n4340) );
  AND3_X1 U4961 ( .A1(n5132), .A2(n5131), .A3(n5130), .ZN(n9889) );
  NAND2_X1 U4962 ( .A1(n4496), .A2(n4494), .ZN(n7452) );
  INV_X1 U4963 ( .A(n7364), .ZN(n7354) );
  NAND2_X1 U4964 ( .A1(n6860), .A2(n6861), .ZN(n6902) );
  OAI21_X1 U4965 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6995), .A(n6994), .ZN(
        n9631) );
  OAI21_X1 U4966 ( .B1(n6995), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6984), .ZN(
        n9634) );
  AOI21_X1 U4967 ( .B1(n5591), .B2(n5590), .A(n7267), .ZN(n5600) );
  NOR2_X1 U4968 ( .A1(n6893), .A2(n4338), .ZN(n6860) );
  CLKBUF_X3 U4969 ( .A(n7289), .Z(n8709) );
  AOI21_X1 U4970 ( .B1(n9013), .B2(P1_REG0_REG_4__SCAN_IN), .A(n6104), .ZN(
        n7279) );
  INV_X1 U4971 ( .A(n6852), .ZN(n8761) );
  INV_X1 U4972 ( .A(n6859), .ZN(n4326) );
  NAND2_X1 U4973 ( .A1(n6627), .A2(n6852), .ZN(n7289) );
  AND3_X1 U4974 ( .A1(n6098), .A2(n6097), .A3(n6096), .ZN(n6961) );
  AND4_X1 U4975 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n7676)
         );
  INV_X2 U4976 ( .A(n6561), .ZN(n6584) );
  NAND2_X1 U4977 ( .A1(n6622), .A2(n4761), .ZN(n6852) );
  AND4_X1 U4978 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n7501)
         );
  NAND2_X1 U4979 ( .A1(n4762), .A2(n7071), .ZN(n6627) );
  INV_X1 U4980 ( .A(n6932), .ZN(n7087) );
  AND4_X1 U4981 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n6938)
         );
  NAND2_X1 U4982 ( .A1(n5208), .A2(n7824), .ZN(n5226) );
  AND2_X2 U4983 ( .A1(n6619), .A2(n7557), .ZN(P1_U3973) );
  INV_X2 U4984 ( .A(n6046), .ZN(n9012) );
  NAND2_X1 U4985 ( .A1(n6464), .A2(n6410), .ZN(n9029) );
  NAND2_X1 U4986 ( .A1(n5565), .A2(n5755), .ZN(n7485) );
  NAND2_X1 U4987 ( .A1(n9430), .A2(n6620), .ZN(n7071) );
  AOI21_X1 U4988 ( .B1(n4729), .B2(n4730), .A(n4728), .ZN(n4727) );
  AND2_X1 U4989 ( .A1(n6621), .A2(n6827), .ZN(n4761) );
  OR2_X1 U4990 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  AND2_X2 U4991 ( .A1(n7878), .A2(n4970), .ZN(n5035) );
  INV_X2 U4992 ( .A(n6091), .ZN(n6602) );
  INV_X1 U4993 ( .A(n6394), .ZN(n4344) );
  INV_X1 U4994 ( .A(n4971), .ZN(n7878) );
  INV_X1 U4995 ( .A(n9101), .ZN(n9430) );
  INV_X1 U4997 ( .A(n6556), .ZN(n5770) );
  NAND2_X1 U4998 ( .A1(n5763), .A2(n5759), .ZN(n7700) );
  AOI21_X1 U4999 ( .B1(n4894), .B2(n5202), .A(n4408), .ZN(n4893) );
  INV_X1 U5000 ( .A(n9109), .ZN(n7834) );
  AND2_X1 U5001 ( .A1(n6406), .A2(n6405), .ZN(n6464) );
  NAND2_X1 U5002 ( .A1(n9109), .A2(n9103), .ZN(n6621) );
  NAND2_X1 U5003 ( .A1(n6632), .A2(n4325), .ZN(n6091) );
  NAND2_X1 U5004 ( .A1(n6491), .A2(n6476), .ZN(n6827) );
  XNOR2_X1 U5005 ( .A(n4337), .B(n6298), .ZN(n9101) );
  XNOR2_X1 U5006 ( .A(n6414), .B(n6413), .ZN(n9103) );
  XNOR2_X1 U5007 ( .A(n4966), .B(P2_IR_REG_30__SCAN_IN), .ZN(n4971) );
  NOR2_X1 U5008 ( .A1(n5218), .A2(n4895), .ZN(n4894) );
  NAND2_X4 U5009 ( .A1(n6459), .A2(n6612), .ZN(n6632) );
  NAND2_X1 U5010 ( .A1(n6285), .A2(n6284), .ZN(n6297) );
  NAND2_X1 U5011 ( .A1(n4968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4966) );
  OAI21_X1 U5012 ( .B1(n6283), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4337) );
  NAND2_X1 U5013 ( .A1(n4976), .A2(n4981), .ZN(n5771) );
  NAND2_X1 U5014 ( .A1(n6472), .A2(n6471), .ZN(n7703) );
  OAI21_X2 U5015 ( .B1(n6412), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6416) );
  MUX2_X1 U5016 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5766), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n5768) );
  XNOR2_X1 U5017 ( .A(n4982), .B(n4962), .ZN(n5772) );
  NAND2_X1 U5018 ( .A1(n6283), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6285) );
  INV_X2 U5019 ( .A(n8559), .ZN(n8568) );
  NAND2_X1 U5020 ( .A1(n4647), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U5021 ( .A1(n6403), .A2(n4374), .ZN(n6412) );
  NOR2_X1 U5022 ( .A1(n6060), .A2(n6059), .ZN(n6061) );
  XNOR2_X1 U5023 ( .A(n6475), .B(n6474), .ZN(n7648) );
  NAND2_X1 U5024 ( .A1(n6402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U5025 ( .A1(n4704), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U5026 ( .A1(n6270), .A2(n6269), .ZN(n6402) );
  AND2_X1 U5027 ( .A1(n5301), .A2(n4959), .ZN(n5764) );
  AND2_X1 U5028 ( .A1(n6255), .A2(n4944), .ZN(n6270) );
  NOR2_X1 U5029 ( .A1(n4637), .A2(n4955), .ZN(n4916) );
  NAND3_X1 U5030 ( .A1(n5005), .A2(n4812), .A3(n4810), .ZN(n9800) );
  AND2_X1 U5031 ( .A1(n4858), .A2(n6030), .ZN(n4857) );
  AND2_X1 U5032 ( .A1(n6028), .A2(n6029), .ZN(n4858) );
  INV_X1 U5033 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5204) );
  INV_X1 U5034 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6415) );
  INV_X1 U5035 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5182) );
  INV_X1 U5036 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4569) );
  INV_X1 U5037 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6469) );
  INV_X1 U5038 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5128) );
  INV_X1 U5039 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4953) );
  INV_X1 U5040 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6465) );
  INV_X4 U5041 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5042 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10117) );
  NOR2_X1 U5043 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6028) );
  NOR2_X1 U5044 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4639) );
  NOR2_X1 U5045 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4640) );
  INV_X4 U5046 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  XNOR2_X1 U5047 ( .A(n4330), .B(n8789), .ZN(n8797) );
  OAI21_X2 U5048 ( .B1(n8645), .B2(n4766), .A(n4332), .ZN(n8853) );
  NOR2_X1 U5049 ( .A1(n4339), .A2(n4326), .ZN(n4338) );
  XNOR2_X1 U5050 ( .A(n6857), .B(n8761), .ZN(n4339) );
  NOR2_X1 U5051 ( .A1(n4341), .A2(n6965), .ZN(n7285) );
  NAND2_X1 U5052 ( .A1(n4736), .A2(n4737), .ZN(n4341) );
  AOI21_X1 U5053 ( .B1(n8904), .B2(n8719), .A(n8718), .ZN(n8723) );
  NAND3_X1 U5054 ( .A1(n4771), .A2(n7350), .A3(n7294), .ZN(n7351) );
  OAI21_X1 U5055 ( .B1(n7294), .B2(n4342), .A(n7351), .ZN(n7301) );
  NOR2_X4 U5056 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6082) );
  NAND2_X2 U5057 ( .A1(n5427), .A2(n5413), .ZN(n8226) );
  OR2_X2 U5058 ( .A1(n5412), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5427) );
  NOR2_X4 U5059 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4832) );
  OR2_X1 U5060 ( .A1(n6043), .A2(n9610), .ZN(n6041) );
  NAND2_X2 U5061 ( .A1(n7895), .A2(n8248), .ZN(n8210) );
  INV_X1 U5062 ( .A(n7289), .ZN(n7352) );
  AND2_X4 U5063 ( .A1(n4971), .A2(n7884), .ZN(n5052) );
  AND2_X1 U5064 ( .A1(n7878), .A2(n4970), .ZN(n4343) );
  OR2_X2 U5065 ( .A1(n8183), .A2(n7868), .ZN(n4948) );
  NAND4_X2 U5066 ( .A1(n6082), .A2(n6105), .A3(n4832), .A4(n6027), .ZN(n6138)
         );
  OAI211_X1 U5067 ( .C1(n5695), .C2(n5694), .A(n5693), .B(n5692), .ZN(n5699)
         );
  OR3_X2 U5068 ( .A1(n5684), .A2(n8213), .A3(n5723), .ZN(n5694) );
  AOI21_X1 U5069 ( .B1(n5679), .B2(n5678), .A(n5677), .ZN(n5695) );
  INV_X4 U5070 ( .A(n4344), .ZN(n4346) );
  AND2_X1 U5071 ( .A1(n6047), .A2(n6045), .ZN(n6076) );
  AND2_X1 U5072 ( .A1(n8011), .A2(n4931), .ZN(n4927) );
  NOR2_X1 U5073 ( .A1(n7406), .A2(n4809), .ZN(n5952) );
  NOR2_X1 U5074 ( .A1(n5998), .A2(n7457), .ZN(n4809) );
  AND2_X1 U5075 ( .A1(n4934), .A2(n4959), .ZN(n4624) );
  AND2_X1 U5076 ( .A1(n4376), .A2(n4935), .ZN(n4934) );
  NOR2_X1 U5077 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4935) );
  AND2_X1 U5078 ( .A1(n4916), .A2(n4915), .ZN(n4499) );
  INV_X1 U5079 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4915) );
  INV_X1 U5080 ( .A(n6076), .ZN(n6185) );
  AOI21_X1 U5081 ( .B1(n7183), .B2(n7181), .A(n7182), .ZN(n7180) );
  NAND3_X1 U5082 ( .A1(n4514), .A2(n4350), .A3(n4515), .ZN(n4513) );
  AOI21_X1 U5083 ( .B1(n7466), .B2(n6529), .A(n4941), .ZN(n7627) );
  OAI21_X1 U5084 ( .B1(n9344), .B2(n6350), .A(n4493), .ZN(n9332) );
  OR2_X1 U5085 ( .A1(n9513), .A2(n9178), .ZN(n4493) );
  NAND2_X1 U5086 ( .A1(n4874), .A2(n6552), .ZN(n5714) );
  NOR2_X1 U5087 ( .A1(n5709), .A2(n5710), .ZN(n4874) );
  INV_X1 U5088 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5302) );
  AOI21_X1 U5089 ( .B1(n4746), .B2(n4745), .A(n8571), .ZN(n4744) );
  INV_X1 U5090 ( .A(n4749), .ZN(n4745) );
  AOI21_X1 U5091 ( .B1(n4673), .B2(n9086), .A(n9023), .ZN(n4670) );
  AND2_X1 U5092 ( .A1(n4672), .A2(n4676), .ZN(n4671) );
  NAND2_X1 U5093 ( .A1(n4677), .A2(n9075), .ZN(n4672) );
  INV_X1 U5094 ( .A(n5270), .ZN(n5273) );
  INV_X1 U5095 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4877) );
  OR2_X1 U5096 ( .A1(n5844), .A2(n5845), .ZN(n5848) );
  INV_X1 U5097 ( .A(n7884), .ZN(n4970) );
  AOI21_X1 U5098 ( .B1(n4803), .B2(n4801), .A(n4533), .ZN(n5919) );
  NAND2_X1 U5099 ( .A1(n7180), .A2(n6678), .ZN(n4521) );
  AND2_X1 U5100 ( .A1(n6764), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4819) );
  AOI21_X1 U5101 ( .B1(n4369), .B2(n4614), .A(n4613), .ZN(n4612) );
  NOR2_X1 U5102 ( .A1(n6549), .A2(n8418), .ZN(n4613) );
  AND2_X1 U5103 ( .A1(n7226), .A2(n5593), .ZN(n4627) );
  OR2_X1 U5104 ( .A1(n8437), .A2(n8279), .ZN(n5725) );
  NAND2_X1 U5105 ( .A1(n7665), .A2(n6533), .ZN(n8386) );
  OR2_X1 U5106 ( .A1(n7521), .A2(n5770), .ZN(n6554) );
  INV_X1 U5107 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4961) );
  INV_X1 U5108 ( .A(n8880), .ZN(n4755) );
  OR2_X1 U5109 ( .A1(n9029), .A2(n7834), .ZN(n9099) );
  INV_X1 U5110 ( .A(n4854), .ZN(n4852) );
  OR2_X1 U5111 ( .A1(n9499), .A2(n6449), .ZN(n9071) );
  NOR2_X1 U5112 ( .A1(n9048), .A2(n4720), .ZN(n4719) );
  INV_X1 U5113 ( .A(n8956), .ZN(n4720) );
  INV_X1 U5114 ( .A(n6075), .ZN(n6395) );
  AND2_X1 U5115 ( .A1(n9029), .A2(n7834), .ZN(n6836) );
  NAND2_X1 U5116 ( .A1(n5513), .A2(n5512), .ZN(n5524) );
  NAND2_X1 U5117 ( .A1(n5509), .A2(n5508), .ZN(n5513) );
  XNOR2_X1 U5118 ( .A(n5524), .B(n5525), .ZN(n5523) );
  AND2_X1 U5119 ( .A1(n5495), .A2(n5481), .ZN(n5493) );
  AND2_X1 U5120 ( .A1(n5477), .A2(n5462), .ZN(n5475) );
  INV_X1 U5121 ( .A(n4886), .ZN(n4885) );
  AND2_X1 U5122 ( .A1(n5457), .A2(n5442), .ZN(n5455) );
  AND2_X1 U5123 ( .A1(n5437), .A2(n5422), .ZN(n5435) );
  NAND2_X1 U5124 ( .A1(n4907), .A2(n5350), .ZN(n5366) );
  NAND2_X1 U5125 ( .A1(n5250), .A2(n4940), .ZN(n5254) );
  INV_X1 U5126 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U5127 ( .A1(n5160), .A2(n5159), .ZN(n5173) );
  INV_X1 U5128 ( .A(n7759), .ZN(n4914) );
  OR2_X1 U5129 ( .A1(n7180), .A2(n4787), .ZN(n4784) );
  OR2_X1 U5130 ( .A1(n4946), .A2(n6678), .ZN(n4787) );
  AND2_X1 U5131 ( .A1(n4373), .A2(n6678), .ZN(n4783) );
  NAND2_X1 U5132 ( .A1(n4535), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4808) );
  AND2_X1 U5133 ( .A1(n4807), .A2(n4553), .ZN(n7614) );
  INV_X1 U5134 ( .A(n7615), .ZN(n4553) );
  NAND2_X1 U5135 ( .A1(n4816), .A2(n4815), .ZN(n4813) );
  INV_X1 U5136 ( .A(n7822), .ZN(n4815) );
  INV_X1 U5137 ( .A(n5930), .ZN(n4782) );
  OR2_X1 U5138 ( .A1(n5220), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5221) );
  AND2_X1 U5139 ( .A1(n5855), .A2(n5769), .ZN(n5972) );
  OR2_X1 U5140 ( .A1(n8129), .A2(n5939), .ZN(n4792) );
  OAI21_X1 U5141 ( .B1(n4566), .B2(n9805), .A(n7902), .ZN(n5975) );
  NAND2_X1 U5142 ( .A1(n5225), .A2(n5224), .ZN(n5242) );
  INV_X1 U5143 ( .A(n5226), .ZN(n5225) );
  AOI21_X1 U5144 ( .B1(n7626), .B2(n4646), .A(n4645), .ZN(n4644) );
  AND2_X1 U5145 ( .A1(n4416), .A2(n5616), .ZN(n4646) );
  OAI21_X1 U5146 ( .B1(n7321), .B2(n6523), .A(n6522), .ZN(n7439) );
  INV_X1 U5147 ( .A(n4604), .ZN(n4603) );
  OAI21_X1 U5148 ( .B1(n6542), .B2(n6543), .A(n4396), .ZN(n4604) );
  NAND2_X1 U5149 ( .A1(n8238), .A2(n5681), .ZN(n4642) );
  OR2_X1 U5150 ( .A1(n8252), .A2(n8264), .ZN(n5680) );
  AND2_X1 U5151 ( .A1(n4624), .A2(n4963), .ZN(n4623) );
  AOI21_X1 U5152 ( .B1(n9164), .B2(n4459), .A(n4371), .ZN(n4654) );
  INV_X1 U5153 ( .A(n4658), .ZN(n4459) );
  AND4_X1 U5154 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n7570)
         );
  NAND2_X1 U5155 ( .A1(n6443), .A2(n9105), .ZN(n9396) );
  AOI21_X1 U5156 ( .B1(n4470), .B2(n4472), .A(n4394), .ZN(n4468) );
  OR2_X1 U5157 ( .A1(n9499), .A2(n9176), .ZN(n4854) );
  NOR2_X1 U5158 ( .A1(n6373), .A2(n4856), .ZN(n4855) );
  INV_X1 U5159 ( .A(n6361), .ZN(n4856) );
  OR2_X1 U5160 ( .A1(n9332), .A2(n6360), .ZN(n6362) );
  OR2_X1 U5161 ( .A1(n9389), .A2(n6321), .ZN(n4841) );
  NOR2_X1 U5162 ( .A1(n4381), .A2(n4834), .ZN(n4833) );
  INV_X1 U5163 ( .A(n4479), .ZN(n4478) );
  OAI21_X1 U5164 ( .B1(n9047), .B2(n4480), .A(n6239), .ZN(n4479) );
  AND2_X1 U5165 ( .A1(n9156), .A2(n6836), .ZN(n9546) );
  XNOR2_X1 U5166 ( .A(n6468), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U5167 ( .A1(n6472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6468) );
  XNOR2_X1 U5168 ( .A(n5476), .B(n5475), .ZN(n8564) );
  NAND2_X1 U5169 ( .A1(n6470), .A2(n6469), .ZN(n6472) );
  NAND2_X1 U5170 ( .A1(n6412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6414) );
  AND2_X1 U5171 ( .A1(n4923), .A2(n4922), .ZN(n4921) );
  INV_X1 U5172 ( .A(n7899), .ZN(n4922) );
  NAND2_X1 U5173 ( .A1(n4918), .A2(n7918), .ZN(n7977) );
  OR2_X1 U5174 ( .A1(n7996), .A2(n4410), .ZN(n4920) );
  INV_X1 U5175 ( .A(n5823), .ZN(n4919) );
  OR2_X1 U5176 ( .A1(n7783), .A2(n7782), .ZN(n4538) );
  NAND2_X1 U5177 ( .A1(n6900), .A2(n6959), .ZN(n4737) );
  OAI21_X1 U5178 ( .B1(n6839), .B2(n7072), .A(n9401), .ZN(n9650) );
  NAND2_X1 U5179 ( .A1(n4567), .A2(n4566), .ZN(n4570) );
  INV_X1 U5180 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U5181 ( .A1(n9360), .A2(n4690), .ZN(n4689) );
  INV_X1 U5182 ( .A(n9079), .ZN(n4690) );
  NAND2_X1 U5183 ( .A1(n4692), .A2(n4691), .ZN(n8994) );
  NAND2_X1 U5184 ( .A1(n4422), .A2(n9161), .ZN(n4691) );
  NAND2_X1 U5185 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  AOI21_X1 U5186 ( .B1(n8978), .B2(n9023), .A(n4695), .ZN(n4694) );
  NOR2_X1 U5187 ( .A1(n4871), .A2(n4866), .ZN(n4865) );
  INV_X1 U5188 ( .A(n5475), .ZN(n4866) );
  INV_X1 U5189 ( .A(n5495), .ZN(n4868) );
  AND2_X1 U5190 ( .A1(n4900), .A2(n5289), .ZN(n4557) );
  INV_X1 U5191 ( .A(n5286), .ZN(n5288) );
  INV_X1 U5192 ( .A(SI_16_), .ZN(n5287) );
  INV_X1 U5193 ( .A(n5249), .ZN(n5252) );
  INV_X1 U5194 ( .A(SI_14_), .ZN(n5251) );
  AOI21_X1 U5195 ( .B1(n4891), .B2(n4893), .A(n5233), .ZN(n4890) );
  INV_X1 U5196 ( .A(n4894), .ZN(n4891) );
  INV_X1 U5197 ( .A(n4893), .ZN(n4892) );
  AND2_X1 U5198 ( .A1(n4881), .A2(n4379), .ZN(n4729) );
  NOR2_X1 U5199 ( .A1(n5143), .A2(n4882), .ZN(n4881) );
  INV_X1 U5200 ( .A(n5121), .ZN(n4882) );
  INV_X1 U5201 ( .A(n5117), .ZN(n4730) );
  NAND2_X1 U5202 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U5203 ( .A1(n4880), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4878) );
  AOI21_X1 U5204 ( .B1(n7200), .B2(n7390), .A(n5892), .ZN(n5782) );
  CLKBUF_X1 U5205 ( .A(n5812), .Z(n5817) );
  NAND2_X1 U5206 ( .A1(n4930), .A2(n5831), .ZN(n4929) );
  INV_X1 U5207 ( .A(n4932), .ZN(n4930) );
  NAND2_X1 U5208 ( .A1(n4909), .A2(n4908), .ZN(n5853) );
  AOI21_X1 U5209 ( .B1(n4910), .B2(n4912), .A(n4423), .ZN(n4908) );
  NAND2_X1 U5210 ( .A1(n4806), .A2(n5947), .ZN(n5948) );
  NAND2_X1 U5211 ( .A1(n4534), .A2(n4533), .ZN(n5949) );
  INV_X1 U5212 ( .A(n5948), .ZN(n4534) );
  INV_X1 U5213 ( .A(n7172), .ZN(n4823) );
  NAND2_X1 U5214 ( .A1(n7174), .A2(n5951), .ZN(n4541) );
  NAND2_X1 U5215 ( .A1(n8132), .A2(n4444), .ZN(n6015) );
  NAND2_X1 U5216 ( .A1(n8220), .A2(n8232), .ZN(n4605) );
  AND2_X1 U5217 ( .A1(n4603), .A2(n4605), .ZN(n4600) );
  OR2_X1 U5218 ( .A1(n8220), .A2(n7938), .ZN(n5688) );
  AND2_X1 U5219 ( .A1(n8501), .A2(n8216), .ZN(n5723) );
  AND2_X1 U5220 ( .A1(n5650), .A2(n5651), .ZN(n6538) );
  OR2_X1 U5221 ( .A1(n8549), .A2(n8390), .ZN(n5641) );
  OAI21_X1 U5222 ( .B1(n7627), .B2(n4594), .A(n4592), .ZN(n7663) );
  INV_X1 U5223 ( .A(n4595), .ZN(n4594) );
  AOI21_X1 U5224 ( .B1(n4595), .B2(n4593), .A(n4401), .ZN(n4592) );
  AOI21_X1 U5225 ( .B1(n6530), .B2(n4596), .A(n4395), .ZN(n4595) );
  NOR2_X1 U5226 ( .A1(n5609), .A2(n4636), .ZN(n4635) );
  INV_X1 U5227 ( .A(n5615), .ZN(n4636) );
  NAND2_X1 U5228 ( .A1(n5764), .A2(n4933), .ZN(n4647) );
  NAND2_X1 U5229 ( .A1(n5561), .A2(n5560), .ZN(n5567) );
  NOR2_X1 U5230 ( .A1(n5185), .A2(n5184), .ZN(n5189) );
  NOR2_X1 U5231 ( .A1(n7566), .A2(n4750), .ZN(n4749) );
  INV_X1 U5232 ( .A(n7443), .ZN(n4750) );
  OAI22_X1 U5233 ( .A1(n7566), .A2(n4748), .B1(n7564), .B2(n7565), .ZN(n4747)
         );
  AND2_X1 U5234 ( .A1(n9031), .A2(n4563), .ZN(n4562) );
  NOR2_X1 U5235 ( .A1(n9271), .A2(n4564), .ZN(n4563) );
  NAND2_X1 U5236 ( .A1(n4671), .A2(n9086), .ZN(n4668) );
  INV_X1 U5237 ( .A(n4670), .ZN(n4669) );
  AOI21_X1 U5238 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9637), .A(n9629), .ZN(
        n9662) );
  AOI21_X1 U5239 ( .B1(n9637), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9632), .ZN(
        n9657) );
  AND2_X1 U5240 ( .A1(n4487), .A2(n4849), .ZN(n4486) );
  INV_X1 U5241 ( .A(n9290), .ZN(n4487) );
  AND2_X1 U5242 ( .A1(n4710), .A2(n9373), .ZN(n4709) );
  NAND2_X1 U5243 ( .A1(n4711), .A2(n8988), .ZN(n4710) );
  INV_X1 U5244 ( .A(n9397), .ZN(n4711) );
  NAND2_X1 U5245 ( .A1(n4722), .A2(n9124), .ZN(n4721) );
  INV_X1 U5246 ( .A(n7525), .ZN(n4722) );
  INV_X1 U5247 ( .A(n9746), .ZN(n4574) );
  OAI21_X1 U5248 ( .B1(n7237), .B2(n7236), .A(n7238), .ZN(n7371) );
  NOR2_X1 U5249 ( .A1(n9390), .A2(n4584), .ZN(n9364) );
  INV_X1 U5250 ( .A(n4586), .ZN(n4584) );
  INV_X1 U5251 ( .A(n6322), .ZN(n4840) );
  NAND2_X1 U5252 ( .A1(n7372), .A2(n7502), .ZN(n7235) );
  NAND2_X1 U5253 ( .A1(n4939), .A2(n6474), .ZN(n4861) );
  NOR2_X1 U5254 ( .A1(n5400), .A2(n5399), .ZN(n4555) );
  NAND2_X1 U5255 ( .A1(n5295), .A2(n4905), .ZN(n4904) );
  NOR2_X1 U5256 ( .A1(n5317), .A2(n4906), .ZN(n4905) );
  INV_X1 U5257 ( .A(n5294), .ZN(n4906) );
  NAND2_X1 U5258 ( .A1(n4556), .A2(n4559), .ZN(n5295) );
  INV_X1 U5259 ( .A(n4560), .ZN(n4559) );
  NAND2_X1 U5260 ( .A1(n5254), .A2(n4557), .ZN(n4556) );
  OAI21_X1 U5261 ( .B1(n4897), .B2(n4561), .A(n5330), .ZN(n4560) );
  AND2_X2 U5262 ( .A1(n5773), .A2(n7200), .ZN(n6561) );
  AND2_X1 U5263 ( .A1(n5805), .A2(n5804), .ZN(n4913) );
  XNOR2_X1 U5264 ( .A(n5812), .B(n5783), .ZN(n5785) );
  AND2_X1 U5265 ( .A1(n7909), .A2(n7910), .ZN(n5838) );
  XNOR2_X1 U5266 ( .A(n8501), .B(n5850), .ZN(n7928) );
  NAND2_X1 U5267 ( .A1(n5830), .A2(n8312), .ZN(n4931) );
  OR2_X1 U5268 ( .A1(n7943), .A2(n4929), .ZN(n4928) );
  NAND2_X1 U5269 ( .A1(n4928), .A2(n4927), .ZN(n8009) );
  NAND2_X1 U5270 ( .A1(n4876), .A2(n4873), .ZN(n5719) );
  NOR2_X1 U5271 ( .A1(n4368), .A2(n5919), .ZN(n4773) );
  NOR2_X1 U5272 ( .A1(n4804), .A2(n6979), .ZN(n4802) );
  NAND2_X1 U5273 ( .A1(n4773), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7183) );
  NAND2_X1 U5274 ( .A1(n4519), .A2(n4522), .ZN(n7403) );
  NOR2_X1 U5275 ( .A1(n4351), .A2(n7333), .ZN(n4520) );
  AND2_X1 U5276 ( .A1(n4447), .A2(n4364), .ZN(n7331) );
  NOR2_X1 U5277 ( .A1(n7343), .A2(n4500), .ZN(n7400) );
  NOR2_X1 U5278 ( .A1(n4501), .A2(n7348), .ZN(n4500) );
  INV_X1 U5279 ( .A(n5997), .ZN(n4501) );
  NAND2_X1 U5280 ( .A1(n7400), .A2(n7399), .ZN(n7398) );
  NAND2_X1 U5281 ( .A1(n4808), .A2(n4378), .ZN(n4807) );
  NOR2_X1 U5282 ( .A1(n7735), .A2(n4778), .ZN(n4777) );
  OAI21_X1 U5283 ( .B1(n7604), .B2(n5988), .A(n4776), .ZN(n4518) );
  NAND2_X1 U5284 ( .A1(n7735), .A2(n4778), .ZN(n4776) );
  NAND2_X1 U5285 ( .A1(n4514), .A2(n4350), .ZN(n4517) );
  INV_X1 U5286 ( .A(n7817), .ZN(n4781) );
  OR2_X1 U5287 ( .A1(n7784), .A2(n5928), .ZN(n5930) );
  NAND2_X1 U5288 ( .A1(n9836), .A2(n4551), .ZN(n4550) );
  NOR2_X1 U5289 ( .A1(n9839), .A2(n9840), .ZN(n9838) );
  OAI21_X1 U5290 ( .B1(n4510), .B2(n4509), .A(n4508), .ZN(n5935) );
  INV_X1 U5291 ( .A(n4805), .ZN(n4509) );
  XNOR2_X1 U5292 ( .A(n5935), .B(n8100), .ZN(n8105) );
  OR2_X1 U5293 ( .A1(n8096), .A2(n8454), .ZN(n4827) );
  INV_X1 U5294 ( .A(n5964), .ZN(n4826) );
  OR2_X1 U5295 ( .A1(n8096), .A2(n4365), .ZN(n4543) );
  NAND2_X1 U5296 ( .A1(n5937), .A2(n8138), .ZN(n5938) );
  NAND2_X1 U5297 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  NAND2_X1 U5298 ( .A1(n6552), .A2(n4612), .ZN(n4609) );
  INV_X1 U5299 ( .A(n4614), .ZN(n4610) );
  NAND2_X1 U5300 ( .A1(n6551), .A2(n4612), .ZN(n4611) );
  OAI21_X1 U5301 ( .B1(n8176), .B2(n4626), .A(n5700), .ZN(n7854) );
  INV_X1 U5302 ( .A(n4948), .ZN(n4626) );
  XNOR2_X1 U5303 ( .A(n7872), .B(n8179), .ZN(n7862) );
  INV_X1 U5304 ( .A(n7862), .ZN(n7847) );
  NAND2_X1 U5305 ( .A1(n5426), .A2(n5425), .ZN(n5446) );
  INV_X1 U5306 ( .A(n5427), .ZN(n5426) );
  OR2_X1 U5307 ( .A1(n8533), .A2(n8326), .ZN(n8318) );
  INV_X1 U5308 ( .A(n5209), .ZN(n5208) );
  OR2_X1 U5309 ( .A1(n7625), .A2(n7626), .ZN(n7623) );
  OR2_X1 U5310 ( .A1(n8068), .A2(n7762), .ZN(n4596) );
  AND2_X1 U5311 ( .A1(n5612), .A2(n5615), .ZN(n7415) );
  OAI21_X1 U5312 ( .B1(n7439), .B2(n6526), .A(n6525), .ZN(n7466) );
  NAND2_X1 U5313 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  NOR2_X1 U5314 ( .A1(n4942), .A2(n7271), .ZN(n6517) );
  NOR2_X1 U5315 ( .A1(n4386), .A2(n4630), .ZN(n4629) );
  AND2_X1 U5316 ( .A1(n7390), .A2(n6556), .ZN(n7201) );
  NAND2_X1 U5317 ( .A1(n7224), .A2(n7226), .ZN(n7223) );
  NAND2_X1 U5318 ( .A1(n6511), .A2(n6510), .ZN(n7209) );
  OAI21_X1 U5319 ( .B1(n8036), .B2(n8483), .A(n6547), .ZN(n8178) );
  AOI21_X1 U5320 ( .B1(n4603), .B2(n6542), .A(n4405), .ZN(n4602) );
  NAND2_X1 U5321 ( .A1(n5373), .A2(n5372), .ZN(n8437) );
  NAND2_X1 U5322 ( .A1(n8292), .A2(n4950), .ZN(n8258) );
  AOI21_X1 U5323 ( .B1(n8322), .B2(n8321), .A(n4591), .ZN(n8310) );
  AND2_X1 U5324 ( .A1(n7955), .A2(n8312), .ZN(n4591) );
  OAI21_X1 U5325 ( .B1(n8386), .B2(n4619), .A(n4616), .ZN(n8360) );
  INV_X1 U5326 ( .A(n4620), .ZN(n4619) );
  AND2_X1 U5327 ( .A1(n4617), .A2(n6537), .ZN(n4616) );
  NAND2_X1 U5328 ( .A1(n6563), .A2(n6561), .ZN(n8389) );
  INV_X1 U5329 ( .A(n8377), .ZN(n8387) );
  INV_X1 U5330 ( .A(n5046), .ZN(n5335) );
  INV_X1 U5331 ( .A(n6562), .ZN(n5334) );
  INV_X1 U5332 ( .A(n8389), .ZN(n8375) );
  NOR2_X2 U5333 ( .A1(n6563), .A2(n6584), .ZN(n8377) );
  AND2_X1 U5334 ( .A1(n7485), .A2(n7521), .ZN(n9914) );
  NOR2_X1 U5335 ( .A1(n5902), .A2(n6581), .ZN(n6570) );
  AND2_X1 U5336 ( .A1(n5875), .A2(n5874), .ZN(n6571) );
  NAND2_X1 U5337 ( .A1(n6555), .A2(n6554), .ZN(n8392) );
  NAND2_X1 U5338 ( .A1(n4980), .A2(n4979), .ZN(n4981) );
  NAND2_X1 U5339 ( .A1(n4963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4979) );
  INV_X1 U5340 ( .A(n5772), .ZN(n5971) );
  XNOR2_X1 U5341 ( .A(n5760), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5855) );
  INV_X1 U5342 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5756) );
  OAI21_X1 U5343 ( .B1(n5755), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  INV_X1 U5344 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U5345 ( .A1(n5566), .A2(n5562), .ZN(n5564) );
  INV_X1 U5346 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5562) );
  INV_X1 U5347 ( .A(n5567), .ZN(n5566) );
  OR2_X1 U5348 ( .A1(n5564), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U5349 ( .A1(n5087), .A2(n4916), .ZN(n5276) );
  NAND2_X1 U5350 ( .A1(n8892), .A2(n8891), .ZN(n4768) );
  INV_X1 U5351 ( .A(n4766), .ZN(n4765) );
  OAI21_X1 U5352 ( .B1(n4769), .B2(n4767), .A(n8750), .ZN(n4766) );
  INV_X1 U5353 ( .A(n4768), .ZN(n4767) );
  NAND2_X1 U5354 ( .A1(n4448), .A2(n4389), .ZN(n4752) );
  INV_X1 U5355 ( .A(n9644), .ZN(n4448) );
  INV_X1 U5356 ( .A(n9645), .ZN(n4754) );
  NAND2_X1 U5357 ( .A1(n8587), .A2(n4755), .ZN(n4753) );
  AND4_X1 U5358 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n7355)
         );
  AND4_X1 U5359 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n7097)
         );
  AND2_X1 U5360 ( .A1(n7743), .A2(n7715), .ZN(n7716) );
  AND2_X1 U5361 ( .A1(n9071), .A2(n9083), .ZN(n9323) );
  OR2_X1 U5362 ( .A1(n9594), .A2(n6439), .ZN(n9408) );
  NAND2_X1 U5363 ( .A1(n6302), .A2(n6301), .ZN(n8648) );
  AND2_X1 U5364 ( .A1(n6438), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U5365 ( .A1(n4719), .A2(n6435), .ZN(n4717) );
  NAND2_X1 U5366 ( .A1(n7525), .A2(n4719), .ZN(n4712) );
  NAND2_X1 U5367 ( .A1(n4721), .A2(n4719), .ZN(n7652) );
  AND2_X1 U5368 ( .A1(n9118), .A2(n4724), .ZN(n4723) );
  INV_X1 U5369 ( .A(n6174), .ZN(n4472) );
  INV_X1 U5370 ( .A(n4471), .ZN(n4470) );
  OAI21_X1 U5371 ( .B1(n7379), .B2(n4472), .A(n9032), .ZN(n4471) );
  NAND2_X1 U5372 ( .A1(n7499), .A2(n6161), .ZN(n7380) );
  NAND2_X1 U5373 ( .A1(n7380), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U5374 ( .A1(n6364), .A2(n6363), .ZN(n9499) );
  NAND2_X1 U5375 ( .A1(n6352), .A2(n6351), .ZN(n9504) );
  OAI21_X1 U5376 ( .B1(n9357), .B2(n6337), .A(n6338), .ZN(n9344) );
  NOR2_X1 U5377 ( .A1(n4398), .A2(n4491), .ZN(n4490) );
  INV_X1 U5378 ( .A(n6267), .ZN(n4491) );
  INV_X1 U5379 ( .A(n6227), .ZN(n4481) );
  NAND2_X1 U5380 ( .A1(n7524), .A2(n9047), .ZN(n7523) );
  NAND2_X1 U5381 ( .A1(n6195), .A2(n6194), .ZN(n8592) );
  INV_X1 U5382 ( .A(n6112), .ZN(n6300) );
  NAND2_X1 U5383 ( .A1(n6452), .A2(n9158), .ZN(n9729) );
  NAND2_X1 U5384 ( .A1(n6488), .A2(n6491), .ZN(n9768) );
  INV_X1 U5385 ( .A(n9768), .ZN(n6494) );
  NAND2_X1 U5386 ( .A1(n5528), .A2(n5527), .ZN(n5546) );
  XNOR2_X1 U5387 ( .A(n5546), .B(n5545), .ZN(n7844) );
  INV_X1 U5388 ( .A(n6058), .ZN(n6060) );
  AND2_X1 U5389 ( .A1(n6037), .A2(n4701), .ZN(n4700) );
  AND2_X1 U5390 ( .A1(n4702), .A2(n6474), .ZN(n4701) );
  INV_X1 U5391 ( .A(n6063), .ZN(n4702) );
  XNOR2_X1 U5392 ( .A(n5494), .B(n5493), .ZN(n7875) );
  NAND2_X1 U5393 ( .A1(n6467), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6470) );
  AND2_X1 U5394 ( .A1(n6037), .A2(n6474), .ZN(n4703) );
  NAND2_X1 U5395 ( .A1(n5408), .A2(n5407), .ZN(n5418) );
  INV_X1 U5396 ( .A(n4558), .ZN(n5331) );
  AOI21_X1 U5397 ( .B1(n4899), .B2(n4897), .A(n4561), .ZN(n4558) );
  NAND2_X1 U5398 ( .A1(n4899), .A2(n5274), .ZN(n5291) );
  NAND2_X1 U5399 ( .A1(n4889), .A2(n4893), .ZN(n5234) );
  NAND2_X1 U5400 ( .A1(n5203), .A2(n4894), .ZN(n4889) );
  NAND2_X1 U5401 ( .A1(n4896), .A2(n5201), .ZN(n5219) );
  INV_X1 U5402 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6030) );
  AND3_X1 U5403 ( .A1(n5398), .A2(n5397), .A3(n5396), .ZN(n8264) );
  INV_X1 U5404 ( .A(n8501), .ZN(n7895) );
  AND4_X1 U5405 ( .A1(n5199), .A2(n5198), .A3(n5197), .A4(n5196), .ZN(n8388)
         );
  AND4_X1 U5406 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n7599)
         );
  NAND2_X1 U5407 ( .A1(n5828), .A2(n4457), .ZN(n4456) );
  INV_X1 U5408 ( .A(n8362), .ZN(n4457) );
  AND4_X1 U5409 ( .A1(n5247), .A2(n5246), .A3(n5245), .A4(n5244), .ZN(n8050)
         );
  INV_X1 U5410 ( .A(n7521), .ZN(n5773) );
  INV_X1 U5411 ( .A(n8264), .ZN(n8231) );
  NAND4_X1 U5412 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n8067)
         );
  INV_X1 U5413 ( .A(n7599), .ZN(n8068) );
  INV_X1 U5414 ( .A(n4803), .ZN(n9801) );
  AND2_X1 U5415 ( .A1(n4498), .A2(n4497), .ZN(n6973) );
  NAND2_X1 U5416 ( .A1(n5994), .A2(n9800), .ZN(n4497) );
  INV_X1 U5417 ( .A(n9806), .ZN(n4498) );
  OR2_X1 U5418 ( .A1(n7607), .A2(n7606), .ZN(n7604) );
  NOR2_X1 U5419 ( .A1(n7723), .A2(n4539), .ZN(n7783) );
  AND2_X1 U5420 ( .A1(n5954), .A2(n7735), .ZN(n4539) );
  NAND2_X1 U5421 ( .A1(n8153), .A2(n8152), .ZN(n4532) );
  NOR2_X1 U5422 ( .A1(n4830), .A2(n8158), .ZN(n4829) );
  NOR2_X1 U5423 ( .A1(n4383), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U5424 ( .A1(n6025), .A2(n4545), .ZN(n4503) );
  INV_X1 U5425 ( .A(n5975), .ZN(n4545) );
  NAND2_X1 U5426 ( .A1(n5393), .A2(n5392), .ZN(n8252) );
  INV_X1 U5427 ( .A(n6531), .ZN(n9905) );
  NOR2_X1 U5428 ( .A1(n7703), .A2(n7648), .ZN(n6476) );
  XNOR2_X1 U5429 ( .A(n6466), .B(n6465), .ZN(n7557) );
  NAND2_X1 U5430 ( .A1(n6464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U5431 ( .A1(n6324), .A2(n6323), .ZN(n9382) );
  NAND2_X1 U5432 ( .A1(n6314), .A2(n6313), .ZN(n9530) );
  NAND2_X1 U5433 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  INV_X1 U5434 ( .A(n6898), .ZN(n4739) );
  NOR2_X2 U5435 ( .A1(n6839), .A2(n6832), .ZN(n8905) );
  NAND2_X1 U5436 ( .A1(n6375), .A2(n6374), .ZN(n8913) );
  NAND2_X1 U5437 ( .A1(n4654), .A2(n4655), .ZN(n4653) );
  INV_X1 U5438 ( .A(n9163), .ZN(n4655) );
  AOI21_X1 U5439 ( .B1(n4654), .B2(n4652), .A(n9170), .ZN(n4650) );
  INV_X1 U5440 ( .A(n4656), .ZN(n4652) );
  NAND2_X1 U5441 ( .A1(n6372), .A2(n6371), .ZN(n9176) );
  OAI21_X1 U5442 ( .B1(n9724), .B2(n4569), .A(n9254), .ZN(n4462) );
  NAND2_X1 U5443 ( .A1(n6838), .A2(n9771), .ZN(n9401) );
  NOR2_X1 U5444 ( .A1(n9509), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U5445 ( .A1(n4846), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4848) );
  NAND2_X1 U5446 ( .A1(n7836), .A2(n7837), .ZN(n4843) );
  NOR2_X1 U5447 ( .A1(n4382), .A2(n4495), .ZN(n4494) );
  OR2_X1 U5448 ( .A1(n6698), .A2(n6091), .ZN(n4496) );
  NOR2_X1 U5449 ( .A1(n6632), .A2(n6747), .ZN(n4495) );
  NAND2_X1 U5450 ( .A1(n6632), .A2(n4683), .ZN(n4682) );
  AND2_X1 U5451 ( .A1(n6459), .A2(n9206), .ZN(n4685) );
  MUX2_X1 U5452 ( .A(n8952), .B(n8951), .S(n9023), .Z(n8957) );
  NOR2_X1 U5453 ( .A1(n9438), .A2(n9133), .ZN(n4681) );
  NOR2_X1 U5454 ( .A1(n9438), .A2(n4680), .ZN(n4679) );
  NOR2_X1 U5455 ( .A1(n9135), .A2(n9023), .ZN(n4680) );
  INV_X1 U5456 ( .A(n9304), .ZN(n4565) );
  AND2_X1 U5457 ( .A1(n9408), .A2(n9422), .ZN(n8970) );
  NAND2_X1 U5458 ( .A1(n8990), .A2(n4696), .ZN(n4695) );
  INV_X1 U5459 ( .A(n8981), .ZN(n4696) );
  INV_X1 U5460 ( .A(n4596), .ZN(n4593) );
  INV_X1 U5461 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4936) );
  AND2_X1 U5462 ( .A1(n4376), .A2(n4960), .ZN(n4933) );
  INV_X1 U5463 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5183) );
  AOI21_X1 U5464 ( .B1(n9166), .B2(n9029), .A(n6631), .ZN(n4762) );
  NOR2_X1 U5465 ( .A1(n9516), .A2(n9382), .ZN(n4586) );
  OAI21_X1 U5466 ( .B1(n5407), .B2(n4887), .A(n5435), .ZN(n4886) );
  INV_X1 U5467 ( .A(n5417), .ZN(n4887) );
  INV_X1 U5468 ( .A(n5401), .ZN(n4884) );
  NOR2_X1 U5469 ( .A1(n4864), .A2(n4428), .ZN(n4863) );
  INV_X1 U5470 ( .A(n5369), .ZN(n4864) );
  NOR2_X1 U5471 ( .A1(n5351), .A2(n4903), .ZN(n4902) );
  INV_X1 U5472 ( .A(n5300), .ZN(n4903) );
  NOR2_X1 U5473 ( .A1(n5271), .A2(n4901), .ZN(n4900) );
  INV_X1 U5474 ( .A(n5253), .ZN(n4901) );
  NAND2_X1 U5475 ( .A1(n5715), .A2(n6584), .ZN(n4876) );
  OAI211_X1 U5476 ( .C1(n5713), .C2(n4875), .A(n4393), .B(n5714), .ZN(n4873)
         );
  NAND2_X1 U5477 ( .A1(n6552), .A2(n8418), .ZN(n4875) );
  AND2_X1 U5478 ( .A1(n5770), .A2(n7390), .ZN(n5892) );
  INV_X1 U5479 ( .A(n5924), .ZN(n4778) );
  NAND2_X1 U5480 ( .A1(n4538), .A2(n5956), .ZN(n5957) );
  NOR2_X1 U5481 ( .A1(n7822), .A2(n4818), .ZN(n4817) );
  INV_X1 U5482 ( .A(n5958), .ZN(n4816) );
  INV_X1 U5483 ( .A(n4819), .ZN(n4551) );
  NAND2_X1 U5484 ( .A1(n8085), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4805) );
  INV_X1 U5485 ( .A(n8122), .ZN(n4828) );
  INV_X1 U5486 ( .A(n5940), .ZN(n4789) );
  OR2_X1 U5487 ( .A1(n6576), .A2(n7869), .ZN(n5721) );
  NOR2_X1 U5488 ( .A1(n4615), .A2(n6550), .ZN(n4614) );
  INV_X1 U5489 ( .A(n6548), .ZN(n4615) );
  AND2_X1 U5490 ( .A1(n4937), .A2(n8305), .ZN(n6541) );
  INV_X1 U5491 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7824) );
  INV_X1 U5492 ( .A(n5624), .ZN(n4645) );
  NAND2_X1 U5493 ( .A1(n5135), .A2(n5134), .ZN(n5165) );
  INV_X1 U5494 ( .A(n5136), .ZN(n5135) );
  OR2_X1 U5495 ( .A1(n6514), .A2(n7261), .ZN(n6515) );
  INV_X1 U5496 ( .A(n5592), .ZN(n4631) );
  NAND2_X1 U5497 ( .A1(n4620), .A2(n4618), .ZN(n4617) );
  INV_X1 U5498 ( .A(n6534), .ZN(n4618) );
  INV_X1 U5499 ( .A(n5640), .ZN(n4634) );
  NOR2_X1 U5500 ( .A1(n8372), .A2(n4621), .ZN(n4620) );
  INV_X1 U5501 ( .A(n6535), .ZN(n4621) );
  AND4_X1 U5502 ( .A1(n4958), .A2(n4957), .A3(n4956), .A4(n5573), .ZN(n4959)
         );
  INV_X1 U5503 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4954) );
  NAND2_X1 U5504 ( .A1(n5087), .A2(n4953), .ZN(n5100) );
  NAND2_X1 U5505 ( .A1(n4742), .A2(n4741), .ZN(n8583) );
  AND2_X1 U5506 ( .A1(n9481), .A2(n9094), .ZN(n9159) );
  INV_X1 U5507 ( .A(n9162), .ZN(n4662) );
  AOI21_X1 U5508 ( .B1(n8994), .B2(n8991), .A(n8993), .ZN(n8985) );
  NOR2_X1 U5509 ( .A1(n8994), .A2(n4689), .ZN(n8996) );
  NOR2_X1 U5510 ( .A1(n9295), .A2(n8773), .ZN(n6606) );
  OR2_X1 U5511 ( .A1(n9504), .A2(n6447), .ZN(n9068) );
  NAND2_X1 U5512 ( .A1(n9354), .A2(n4586), .ZN(n4585) );
  NOR2_X1 U5513 ( .A1(n8609), .A2(n4578), .ZN(n4577) );
  INV_X1 U5514 ( .A(n4579), .ZN(n4578) );
  NOR2_X1 U5515 ( .A1(n8867), .A2(n8738), .ZN(n4579) );
  AND2_X1 U5516 ( .A1(n7314), .A2(n9780), .ZN(n7313) );
  AND2_X1 U5517 ( .A1(n7235), .A2(n7096), .ZN(n4492) );
  AND2_X1 U5518 ( .A1(n6117), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U5519 ( .A1(n9197), .A2(n7087), .ZN(n9111) );
  NAND2_X1 U5520 ( .A1(n4688), .A2(n4687), .ZN(n6883) );
  INV_X1 U5521 ( .A(n6881), .ZN(n4687) );
  INV_X1 U5522 ( .A(n6419), .ZN(n4688) );
  NAND2_X1 U5523 ( .A1(n6856), .A2(n6890), .ZN(n6420) );
  OR2_X1 U5524 ( .A1(n9011), .A2(n9010), .ZN(n9065) );
  NAND2_X1 U5525 ( .A1(n9327), .A2(n9071), .ZN(n9305) );
  INV_X1 U5526 ( .A(n6280), .ZN(n4834) );
  NAND2_X1 U5527 ( .A1(n7530), .A2(n7535), .ZN(n7589) );
  NOR2_X1 U5528 ( .A1(n7509), .A2(n7687), .ZN(n7314) );
  NAND2_X1 U5529 ( .A1(n6883), .A2(n6420), .ZN(n6927) );
  INV_X1 U5530 ( .A(n9166), .ZN(n9156) );
  INV_X1 U5531 ( .A(SI_17_), .ZN(n10129) );
  NAND2_X1 U5532 ( .A1(n4870), .A2(n4867), .ZN(n5509) );
  AOI21_X1 U5533 ( .B1(n5493), .B2(n4869), .A(n4868), .ZN(n4867) );
  INV_X1 U5534 ( .A(n5477), .ZN(n4869) );
  INV_X1 U5535 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6039) );
  NOR2_X1 U5536 ( .A1(n5290), .A2(n4898), .ZN(n4897) );
  INV_X1 U5537 ( .A(n5274), .ZN(n4898) );
  NAND2_X1 U5538 ( .A1(n5254), .A2(n4900), .ZN(n4899) );
  AOI21_X1 U5539 ( .B1(n4890), .B2(n4892), .A(n4404), .ZN(n4888) );
  INV_X1 U5540 ( .A(n5201), .ZN(n4895) );
  INV_X1 U5541 ( .A(n5144), .ZN(n4728) );
  OAI21_X1 U5542 ( .B1(n4325), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n4466), .ZN(
        n5105) );
  NAND2_X1 U5543 ( .A1(n4325), .A2(n6683), .ZN(n4466) );
  OAI21_X1 U5544 ( .B1(n4733), .B2(n4732), .A(n4731), .ZN(n5009) );
  NAND2_X1 U5545 ( .A1(n4733), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5546 ( .A1(n4734), .A2(n4879), .ZN(n4733) );
  OAI21_X1 U5547 ( .B1(n5145), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5012), .ZN(
        n5026) );
  NAND2_X1 U5548 ( .A1(n4926), .A2(n7898), .ZN(n4925) );
  INV_X1 U5549 ( .A(n4929), .ZN(n4926) );
  OR2_X1 U5550 ( .A1(n4927), .A2(n5833), .ZN(n4923) );
  XNOR2_X1 U5551 ( .A(n5810), .B(n5808), .ZN(n7539) );
  OR2_X1 U5552 ( .A1(n5111), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5136) );
  INV_X1 U5553 ( .A(n5812), .ZN(n5788) );
  AOI21_X1 U5554 ( .B1(n4943), .B2(n4384), .A(n4911), .ZN(n4910) );
  INV_X1 U5555 ( .A(n7932), .ZN(n4911) );
  INV_X1 U5556 ( .A(n4943), .ZN(n4912) );
  NAND2_X1 U5557 ( .A1(n5799), .A2(n7256), .ZN(n7259) );
  OR2_X1 U5558 ( .A1(n5165), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U5559 ( .A1(n6561), .A2(n5892), .ZN(n6559) );
  XNOR2_X1 U5560 ( .A(n5993), .B(n4504), .ZN(n6662) );
  NOR2_X1 U5561 ( .A1(n7051), .A2(n7057), .ZN(n7050) );
  NOR2_X1 U5562 ( .A1(n6662), .A2(n7050), .ZN(n6661) );
  NAND2_X1 U5563 ( .A1(n4801), .A2(n4798), .ZN(n9802) );
  NAND2_X1 U5564 ( .A1(n4800), .A2(n4799), .ZN(n4798) );
  NAND2_X1 U5565 ( .A1(n4797), .A2(n4796), .ZN(n4803) );
  INV_X1 U5566 ( .A(n9802), .ZN(n4797) );
  INV_X1 U5567 ( .A(n9803), .ZN(n4796) );
  NAND2_X1 U5568 ( .A1(n4441), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U5569 ( .A1(n4822), .A2(n4821), .ZN(n7174) );
  AOI21_X1 U5570 ( .B1(n7171), .B2(n4824), .A(n4823), .ZN(n4822) );
  NAND2_X1 U5571 ( .A1(n6971), .A2(n4372), .ZN(n7168) );
  NOR2_X1 U5572 ( .A1(n7168), .A2(n7169), .ZN(n7167) );
  XNOR2_X1 U5573 ( .A(n4541), .B(n7348), .ZN(n7337) );
  AND2_X1 U5574 ( .A1(n7337), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7339) );
  NOR2_X1 U5575 ( .A1(n7339), .A2(n4540), .ZN(n7408) );
  AND2_X1 U5576 ( .A1(n4541), .A2(n6678), .ZN(n4540) );
  XNOR2_X1 U5577 ( .A(n5922), .B(n9825), .ZN(n9820) );
  NAND2_X1 U5578 ( .A1(n7398), .A2(n6000), .ZN(n9830) );
  NAND2_X1 U5579 ( .A1(n9830), .A2(n9831), .ZN(n9829) );
  NOR2_X1 U5580 ( .A1(n7403), .A2(n5921), .ZN(n5922) );
  NOR2_X1 U5581 ( .A1(n5998), .A2(n5920), .ZN(n5921) );
  NAND2_X1 U5582 ( .A1(n7604), .A2(n5924), .ZN(n4775) );
  NOR2_X1 U5583 ( .A1(n7614), .A2(n4552), .ZN(n5953) );
  AND2_X1 U5584 ( .A1(n6701), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4552) );
  XNOR2_X1 U5585 ( .A(n5957), .B(n5984), .ZN(n7803) );
  NAND2_X1 U5586 ( .A1(n7803), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7802) );
  AND2_X1 U5587 ( .A1(n4361), .A2(n4780), .ZN(n7808) );
  NOR2_X1 U5588 ( .A1(n9838), .A2(n5961), .ZN(n8088) );
  AOI21_X1 U5589 ( .B1(n4349), .B2(n9843), .A(n8079), .ZN(n4510) );
  NAND2_X1 U5590 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  NOR2_X1 U5591 ( .A1(n8113), .A2(n8352), .ZN(n4526) );
  NAND2_X1 U5592 ( .A1(n4525), .A2(n4524), .ZN(n5937) );
  AND2_X1 U5593 ( .A1(n4528), .A2(n4442), .ZN(n4524) );
  NAND2_X1 U5594 ( .A1(n8133), .A2(n8134), .ZN(n8132) );
  INV_X1 U5595 ( .A(n8152), .ZN(n4791) );
  INV_X1 U5596 ( .A(n6016), .ZN(n8148) );
  NOR2_X1 U5597 ( .A1(n5967), .A2(n8140), .ZN(n8157) );
  AOI21_X1 U5598 ( .B1(n5939), .B2(n4791), .A(n4789), .ZN(n4788) );
  NAND2_X1 U5599 ( .A1(n5445), .A2(n7937), .ZN(n5465) );
  NAND2_X1 U5600 ( .A1(n5375), .A2(n5374), .ZN(n5394) );
  INV_X1 U5601 ( .A(n5376), .ZN(n5375) );
  NAND2_X1 U5602 ( .A1(n5311), .A2(n5310), .ZN(n5355) );
  INV_X1 U5603 ( .A(n5325), .ZN(n5311) );
  NAND2_X1 U5604 ( .A1(n5309), .A2(n5308), .ZN(n5323) );
  INV_X1 U5605 ( .A(n5338), .ZN(n5309) );
  OR2_X1 U5606 ( .A1(n5323), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5325) );
  OR2_X1 U5607 ( .A1(n5280), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5608 ( .A1(n5263), .A2(n5262), .ZN(n5280) );
  INV_X1 U5609 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5262) );
  INV_X1 U5610 ( .A(n5264), .ZN(n5263) );
  OR2_X1 U5611 ( .A1(n5242), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5264) );
  OR2_X1 U5612 ( .A1(n5194), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5209) );
  AND2_X1 U5613 ( .A1(n5627), .A2(n5628), .ZN(n7662) );
  AND2_X1 U5614 ( .A1(n5164), .A2(n5163), .ZN(n6531) );
  INV_X1 U5615 ( .A(n8069), .ZN(n7629) );
  AND4_X1 U5616 ( .A1(n5099), .A2(n5098), .A3(n5097), .A4(n5096), .ZN(n8026)
         );
  INV_X1 U5617 ( .A(n7415), .ZN(n7465) );
  OR2_X1 U5618 ( .A1(n5075), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5094) );
  NOR2_X1 U5619 ( .A1(n6514), .A2(n4589), .ZN(n4588) );
  INV_X1 U5620 ( .A(n6512), .ZN(n4589) );
  AND2_X1 U5621 ( .A1(n5586), .A2(n5585), .ZN(n7206) );
  INV_X1 U5622 ( .A(n7206), .ZN(n7208) );
  INV_X1 U5623 ( .A(n6508), .ZN(n4999) );
  NAND2_X1 U5624 ( .A1(n6589), .A2(n6588), .ZN(n7027) );
  AND2_X1 U5625 ( .A1(n6583), .A2(n6582), .ZN(n7029) );
  AND2_X1 U5626 ( .A1(n4948), .A2(n5700), .ZN(n8177) );
  NAND2_X1 U5627 ( .A1(n4599), .A2(n4597), .ZN(n8201) );
  OR2_X1 U5628 ( .A1(n4411), .A2(n4598), .ZN(n4597) );
  INV_X1 U5629 ( .A(n4605), .ZN(n4598) );
  AND2_X1 U5630 ( .A1(n6544), .A2(n6546), .ZN(n8200) );
  NAND2_X1 U5631 ( .A1(n4642), .A2(n4641), .ZN(n8211) );
  AND2_X1 U5632 ( .A1(n5416), .A2(n5680), .ZN(n4641) );
  AND4_X1 U5633 ( .A1(n5381), .A2(n5380), .A3(n5379), .A4(n5378), .ZN(n8279)
         );
  OR2_X1 U5634 ( .A1(n5363), .A2(n5362), .ZN(n8270) );
  AND2_X1 U5635 ( .A1(n8318), .A2(n8286), .ZN(n8332) );
  AND2_X1 U5636 ( .A1(n8348), .A2(n8347), .ZN(n6539) );
  NAND2_X1 U5637 ( .A1(n8386), .A2(n6534), .ZN(n4622) );
  NAND2_X1 U5638 ( .A1(n4622), .A2(n4620), .ZN(n8373) );
  OR2_X1 U5639 ( .A1(n8399), .A2(n8400), .ZN(n8397) );
  AND3_X1 U5640 ( .A1(n5072), .A2(n5071), .A3(n5070), .ZN(n9876) );
  AND3_X1 U5641 ( .A1(n5051), .A2(n5050), .A3(n5049), .ZN(n9872) );
  INV_X1 U5642 ( .A(n9914), .ZN(n9893) );
  OR2_X1 U5643 ( .A1(n6723), .A2(n5972), .ZN(n6581) );
  NAND2_X1 U5644 ( .A1(n5973), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6723) );
  XNOR2_X1 U5645 ( .A(n5568), .B(P2_IR_REG_20__SCAN_IN), .ZN(n5746) );
  INV_X1 U5646 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5237) );
  INV_X1 U5647 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5188) );
  INV_X1 U5648 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U5649 ( .A1(n8584), .A2(n8586), .ZN(n9644) );
  OR2_X1 U5650 ( .A1(n8583), .A2(n8582), .ZN(n8584) );
  OR2_X1 U5651 ( .A1(n8892), .A2(n8891), .ZN(n4769) );
  AND2_X1 U5652 ( .A1(n8715), .A2(n8714), .ZN(n8774) );
  AND2_X1 U5653 ( .A1(n6325), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6333) );
  OR2_X1 U5654 ( .A1(n8622), .A2(n8918), .ZN(n8625) );
  NAND2_X1 U5655 ( .A1(n7444), .A2(n4749), .ZN(n4743) );
  INV_X1 U5656 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6312) );
  AND2_X1 U5657 ( .A1(n6221), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6233) );
  INV_X1 U5658 ( .A(n8674), .ZN(n4449) );
  OR2_X1 U5659 ( .A1(n9644), .A2(n9645), .ZN(n4756) );
  INV_X1 U5660 ( .A(n9099), .ZN(n6831) );
  AND2_X1 U5661 ( .A1(n9162), .A2(n9101), .ZN(n4458) );
  AND2_X1 U5662 ( .A1(n9022), .A2(n4665), .ZN(n4664) );
  AND2_X1 U5663 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  NAND2_X1 U5664 ( .A1(n4666), .A2(n4392), .ZN(n4665) );
  AND2_X1 U5665 ( .A1(n6648), .A2(n6831), .ZN(n9167) );
  AND4_X1 U5666 ( .A1(n6266), .A2(n6265), .A3(n6264), .A4(n6263), .ZN(n8821)
         );
  AND4_X1 U5667 ( .A1(n6216), .A2(n6215), .A3(n6214), .A4(n6213), .ZN(n7527)
         );
  AND4_X1 U5668 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6186), .ZN(n8585)
         );
  NAND2_X1 U5669 ( .A1(n9201), .A2(n9200), .ZN(n9199) );
  AOI21_X1 U5670 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6813), .A(n6810), .ZN(
        n6758) );
  AOI21_X1 U5671 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6813), .A(n6807), .ZN(
        n6748) );
  AOI21_X1 U5672 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9681), .A(n9676), .ZN(
        n9687) );
  AOI21_X1 U5673 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9681), .A(n9673), .ZN(
        n9690) );
  AOI21_X1 U5674 ( .B1(n9693), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9685), .ZN(
        n7712) );
  AOI21_X1 U5675 ( .B1(n9693), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9688), .ZN(
        n7705) );
  OR2_X1 U5676 ( .A1(n7746), .A2(n7745), .ZN(n7743) );
  OR2_X1 U5677 ( .A1(n9711), .A2(n9710), .ZN(n9714) );
  NOR2_X1 U5678 ( .A1(n9260), .A2(n9282), .ZN(n9259) );
  NAND2_X1 U5679 ( .A1(n6606), .A2(n6605), .ZN(n9282) );
  INV_X1 U5680 ( .A(n6606), .ZN(n9281) );
  AOI21_X1 U5681 ( .B1(n4486), .B2(n4488), .A(n4348), .ZN(n4485) );
  AOI21_X1 U5682 ( .B1(n4850), .B2(n4851), .A(n4387), .ZN(n4849) );
  INV_X1 U5683 ( .A(n4855), .ZN(n4850) );
  INV_X1 U5684 ( .A(n4851), .ZN(n4488) );
  OAI21_X1 U5685 ( .B1(n9305), .B2(n9304), .A(n9146), .ZN(n9291) );
  AND2_X1 U5686 ( .A1(n9008), .A2(n9007), .ZN(n9290) );
  NAND2_X1 U5687 ( .A1(n9322), .A2(n9323), .ZN(n9327) );
  NOR2_X1 U5688 ( .A1(n9499), .A2(n4949), .ZN(n9317) );
  NAND2_X1 U5689 ( .A1(n6333), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6343) );
  AOI21_X1 U5690 ( .B1(n4709), .B2(n8989), .A(n4707), .ZN(n4706) );
  INV_X1 U5691 ( .A(n8991), .ZN(n4707) );
  NOR2_X1 U5692 ( .A1(n9390), .A2(n9382), .ZN(n9380) );
  NAND2_X1 U5693 ( .A1(n9395), .A2(n8988), .ZN(n9374) );
  NAND2_X1 U5694 ( .A1(n9396), .A2(n9397), .ZN(n9395) );
  AND2_X1 U5695 ( .A1(n9444), .A2(n9433), .ZN(n9420) );
  NOR2_X1 U5696 ( .A1(n6274), .A2(n6273), .ZN(n6289) );
  AOI21_X1 U5697 ( .B1(n4716), .B2(n4718), .A(n4714), .ZN(n4713) );
  INV_X1 U5698 ( .A(n8960), .ZN(n4714) );
  NAND2_X1 U5699 ( .A1(n7530), .A2(n4577), .ZN(n9458) );
  OR2_X1 U5700 ( .A1(n6246), .A2(n8922), .ZN(n6261) );
  NAND2_X1 U5701 ( .A1(n4721), .A2(n8956), .ZN(n7582) );
  OR2_X1 U5702 ( .A1(n6196), .A2(n8884), .ZN(n6210) );
  NAND2_X1 U5703 ( .A1(n9114), .A2(n9118), .ZN(n7303) );
  AOI21_X1 U5704 ( .B1(n4705), .B2(n7376), .A(n7375), .ZN(n8935) );
  NAND2_X1 U5705 ( .A1(n7371), .A2(n7370), .ZN(n4705) );
  NAND3_X1 U5706 ( .A1(n7510), .A2(n7243), .A3(n7247), .ZN(n7509) );
  NAND2_X1 U5707 ( .A1(n4836), .A2(n4837), .ZN(n7500) );
  AOI21_X1 U5708 ( .B1(n7235), .B2(n4838), .A(n4402), .ZN(n4837) );
  NAND2_X1 U5709 ( .A1(n7093), .A2(n4492), .ZN(n4836) );
  INV_X1 U5710 ( .A(n6142), .ZN(n4838) );
  INV_X1 U5711 ( .A(n9115), .ZN(n4725) );
  NOR2_X1 U5712 ( .A1(n4575), .A2(n7123), .ZN(n7243) );
  NAND2_X1 U5713 ( .A1(n7354), .A2(n9761), .ZN(n4575) );
  NOR2_X1 U5714 ( .A1(n7123), .A2(n7290), .ZN(n7122) );
  INV_X1 U5715 ( .A(n9729), .ZN(n9425) );
  XNOR2_X1 U5716 ( .A(n9196), .B(n6961), .ZN(n9034) );
  NAND2_X1 U5717 ( .A1(n6421), .A2(n9111), .ZN(n9033) );
  NAND2_X1 U5718 ( .A1(n7078), .A2(n6872), .ZN(n6926) );
  INV_X1 U5719 ( .A(n8874), .ZN(n8907) );
  NAND2_X1 U5720 ( .A1(n4484), .A2(n4482), .ZN(n9265) );
  AND2_X1 U5721 ( .A1(n4485), .A2(n4483), .ZN(n4482) );
  INV_X1 U5722 ( .A(n9267), .ZN(n4483) );
  AND4_X1 U5723 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(n9277)
         );
  AND2_X1 U5724 ( .A1(n6836), .A2(n9103), .ZN(n9505) );
  AND2_X1 U5725 ( .A1(n8984), .A2(n9077), .ZN(n9346) );
  NOR2_X1 U5726 ( .A1(n4397), .A2(n4840), .ZN(n4839) );
  AND2_X1 U5727 ( .A1(n8980), .A2(n8988), .ZN(n9397) );
  AND2_X1 U5728 ( .A1(n9408), .A2(n8974), .ZN(n9424) );
  AOI21_X1 U5729 ( .B1(n4347), .B2(n4480), .A(n4390), .ZN(n4474) );
  INV_X1 U5730 ( .A(n9546), .ZN(n9787) );
  NAND2_X1 U5731 ( .A1(n7095), .A2(n6142), .ZN(n7234) );
  NAND2_X1 U5732 ( .A1(n7093), .A2(n7096), .ZN(n7095) );
  NAND2_X1 U5733 ( .A1(n4409), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U5734 ( .A1(n6070), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4684) );
  AND3_X1 U5735 ( .A1(n6825), .A2(P1_STATE_REG_SCAN_IN), .A3(n6824), .ZN(n7068) );
  XNOR2_X1 U5736 ( .A(n5523), .B(n5514), .ZN(n7882) );
  XNOR2_X1 U5737 ( .A(n5509), .B(n5508), .ZN(n6391) );
  NAND2_X1 U5738 ( .A1(n5418), .A2(n5417), .ZN(n5436) );
  INV_X1 U5739 ( .A(n4555), .ZN(n5402) );
  INV_X1 U5740 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U5741 ( .A1(n5370), .A2(n5369), .ZN(n5383) );
  NAND2_X1 U5742 ( .A1(n4904), .A2(n5300), .ZN(n5352) );
  INV_X1 U5743 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U5744 ( .A1(n5254), .A2(n5253), .ZN(n5272) );
  AND2_X1 U5745 ( .A1(n6206), .A2(n6228), .ZN(n7710) );
  INV_X1 U5746 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6027) );
  XNOR2_X1 U5747 ( .A(n5026), .B(SI_2_), .ZN(n5024) );
  NAND2_X1 U5748 ( .A1(n8021), .A2(n5804), .ZN(n7428) );
  NAND2_X1 U5749 ( .A1(n6949), .A2(n5792), .ZN(n7043) );
  AND4_X1 U5750 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n8297)
         );
  AND4_X1 U5751 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n8390)
         );
  NAND2_X1 U5752 ( .A1(n5207), .A2(n5206), .ZN(n9913) );
  NAND2_X1 U5753 ( .A1(n7538), .A2(n5811), .ZN(n7758) );
  AND2_X1 U5754 ( .A1(n5834), .A2(n8278), .ZN(n4455) );
  AND4_X1 U5755 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n8003)
         );
  AND4_X1 U5756 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n8340)
         );
  AND2_X1 U5757 ( .A1(n4928), .A2(n4931), .ZN(n8010) );
  NAND2_X1 U5758 ( .A1(n5889), .A2(n8227), .ZN(n8030) );
  AND4_X1 U5759 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n8326)
         );
  NAND2_X1 U5760 ( .A1(n6570), .A2(n5891), .ZN(n8052) );
  AND2_X1 U5761 ( .A1(n5827), .A2(n8050), .ZN(n4917) );
  INV_X1 U5762 ( .A(n8040), .ZN(n8055) );
  AND2_X1 U5763 ( .A1(n5557), .A2(n5544), .ZN(n8163) );
  INV_X1 U5764 ( .A(n8036), .ZN(n8202) );
  INV_X1 U5765 ( .A(n8279), .ZN(n8062) );
  INV_X1 U5766 ( .A(n8340), .ZN(n8312) );
  INV_X1 U5767 ( .A(n8050), .ZN(n8376) );
  INV_X1 U5768 ( .A(n8003), .ZN(n8378) );
  NAND2_X1 U5769 ( .A1(n9813), .A2(n9812), .ZN(n4806) );
  NAND2_X1 U5770 ( .A1(n7183), .A2(n4772), .ZN(n6974) );
  OR2_X1 U5771 ( .A1(n4773), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4772) );
  NAND2_X1 U5772 ( .A1(n6973), .A2(n6972), .ZN(n6971) );
  NAND2_X1 U5773 ( .A1(n4364), .A2(n4784), .ZN(n7332) );
  NOR2_X1 U5774 ( .A1(n7331), .A2(n4783), .ZN(n7405) );
  NOR2_X1 U5775 ( .A1(n9818), .A2(n4536), .ZN(n9827) );
  INV_X1 U5776 ( .A(n4808), .ZN(n9818) );
  INV_X1 U5777 ( .A(n4807), .ZN(n7616) );
  OR2_X1 U5778 ( .A1(n4518), .A2(n4516), .ZN(n7727) );
  INV_X1 U5779 ( .A(n7808), .ZN(n4779) );
  NAND2_X1 U5780 ( .A1(n4505), .A2(n4506), .ZN(n7816) );
  NAND2_X1 U5781 ( .A1(n5930), .A2(n4426), .ZN(n4506) );
  OR2_X1 U5782 ( .A1(n9842), .A2(n9843), .ZN(n4511) );
  OR2_X1 U5783 ( .A1(P2_U3150), .A2(n5974), .ZN(n9805) );
  INV_X1 U5784 ( .A(n4827), .ZN(n8095) );
  NOR2_X1 U5785 ( .A1(n8105), .A2(n8352), .ZN(n8104) );
  NAND2_X1 U5786 ( .A1(n4543), .A2(n4825), .ZN(n8121) );
  NAND2_X1 U5787 ( .A1(n4525), .A2(n4528), .ZN(n8112) );
  NAND2_X1 U5788 ( .A1(n4608), .A2(n4611), .ZN(n4607) );
  XNOR2_X1 U5789 ( .A(n7848), .B(n7847), .ZN(n7852) );
  NAND2_X1 U5790 ( .A1(n5483), .A2(n5482), .ZN(n8183) );
  NAND2_X1 U5791 ( .A1(n5464), .A2(n5463), .ZN(n8195) );
  NAND2_X1 U5792 ( .A1(n5444), .A2(n5443), .ZN(n8206) );
  NAND2_X1 U5793 ( .A1(n7623), .A2(n5616), .ZN(n7595) );
  OAI21_X1 U5794 ( .B1(n7627), .B2(n6530), .A(n4596), .ZN(n7597) );
  AND2_X1 U5795 ( .A1(n7204), .A2(n8401), .ZN(n8406) );
  NAND2_X1 U5796 ( .A1(n7418), .A2(n5615), .ZN(n7480) );
  NAND2_X1 U5797 ( .A1(n7223), .A2(n5592), .ZN(n7266) );
  INV_X1 U5798 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7229) );
  NAND2_X1 U5799 ( .A1(n7203), .A2(n8219), .ZN(n8403) );
  AND2_X1 U5800 ( .A1(n7036), .A2(n8227), .ZN(n8408) );
  INV_X1 U5801 ( .A(n8227), .ZN(n8396) );
  INV_X2 U5802 ( .A(n8408), .ZN(n8401) );
  NAND2_X1 U5803 ( .A1(n5549), .A2(n5548), .ZN(n8412) );
  OR2_X1 U5804 ( .A1(n5046), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4625) );
  AND4_X2 U5805 ( .A1(n7029), .A2(n6591), .A3(n6590), .A4(n7027), .ZN(n9938)
         );
  INV_X1 U5806 ( .A(n8412), .ZN(n8469) );
  INV_X1 U5807 ( .A(n8183), .ZN(n8477) );
  INV_X1 U5808 ( .A(n8195), .ZN(n8483) );
  NAND2_X1 U5809 ( .A1(n4601), .A2(n4602), .ZN(n8214) );
  NAND2_X1 U5810 ( .A1(n8241), .A2(n4603), .ZN(n4601) );
  AOI21_X1 U5811 ( .B1(n8241), .B2(n6543), .A(n6542), .ZN(n8230) );
  NAND2_X1 U5812 ( .A1(n4642), .A2(n5680), .ZN(n8225) );
  NAND2_X1 U5813 ( .A1(n5354), .A2(n5353), .ZN(n8513) );
  NAND2_X1 U5814 ( .A1(n5279), .A2(n5278), .ZN(n8533) );
  NAND2_X1 U5815 ( .A1(n5223), .A2(n5222), .ZN(n8549) );
  AND3_X1 U5816 ( .A1(n5091), .A2(n5090), .A3(n5089), .ZN(n7461) );
  INV_X1 U5817 ( .A(n5783), .ZN(n7011) );
  INV_X2 U5818 ( .A(n9921), .ZN(n9919) );
  OR2_X1 U5819 ( .A1(n5855), .A2(n5780), .ZN(n6724) );
  NAND2_X1 U5820 ( .A1(n6720), .A2(n6719), .ZN(n6729) );
  NAND2_X1 U5821 ( .A1(n4969), .A2(n4968), .ZN(n7884) );
  MUX2_X1 U5822 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5762), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5763) );
  INV_X1 U5823 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10114) );
  INV_X1 U5824 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7522) );
  XNOR2_X1 U5825 ( .A(n5574), .B(n5573), .ZN(n7521) );
  INV_X1 U5826 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7484) );
  INV_X1 U5827 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7389) );
  INV_X1 U5828 ( .A(n5746), .ZN(n7390) );
  INV_X1 U5829 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6909) );
  XNOR2_X1 U5830 ( .A(n5257), .B(n5256), .ZN(n8085) );
  INV_X1 U5831 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10105) );
  INV_X1 U5832 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6712) );
  INV_X1 U5833 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6706) );
  INV_X1 U5834 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6703) );
  INV_X1 U5835 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6699) );
  INV_X1 U5836 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U5837 ( .A1(n4977), .A2(n4951), .ZN(n4812) );
  OR2_X1 U5838 ( .A1(n5004), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U5839 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4811) );
  AOI21_X1 U5840 ( .B1(n7444), .B2(n7443), .A(n4353), .ZN(n7567) );
  AND2_X1 U5841 ( .A1(n6386), .A2(n6454), .ZN(n9297) );
  NAND2_X1 U5842 ( .A1(n7875), .A2(n6602), .ZN(n4554) );
  NAND2_X1 U5843 ( .A1(n6341), .A2(n6340), .ZN(n9513) );
  CLKBUF_X1 U5844 ( .A(n7285), .Z(n8843) );
  NAND2_X1 U5845 ( .A1(n4764), .A2(n4768), .ZN(n8751) );
  NAND2_X1 U5846 ( .A1(n8647), .A2(n4769), .ZN(n4764) );
  NAND2_X1 U5847 ( .A1(n4453), .A2(n4452), .ZN(n4451) );
  NOR2_X1 U5848 ( .A1(n8774), .A2(n9646), .ZN(n4453) );
  INV_X1 U5849 ( .A(n8775), .ZN(n4452) );
  NAND2_X1 U5850 ( .A1(n8722), .A2(n4758), .ZN(n4757) );
  INV_X1 U5851 ( .A(n8704), .ZN(n4758) );
  NAND2_X1 U5852 ( .A1(n8663), .A2(n8662), .ZN(n8784) );
  INV_X1 U5853 ( .A(n8882), .ZN(n4751) );
  NAND2_X1 U5854 ( .A1(n6272), .A2(n6271), .ZN(n9545) );
  INV_X1 U5855 ( .A(n8842), .ZN(n7283) );
  INV_X1 U5856 ( .A(n8841), .ZN(n7282) );
  AOI21_X1 U5857 ( .B1(n4765), .B2(n4767), .A(n4407), .ZN(n4763) );
  INV_X1 U5858 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8884) );
  INV_X1 U5859 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U5860 ( .A1(n6834), .A2(n9166), .ZN(n9641) );
  INV_X1 U5861 ( .A(n9653), .ZN(n8929) );
  INV_X1 U5862 ( .A(n8585), .ZN(n9189) );
  AOI21_X1 U5863 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6757), .A(n6756), .ZN(
        n6793) );
  AOI21_X1 U5864 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6757), .A(n6744), .ZN(
        n6796) );
  AOI21_X1 U5865 ( .B1(n6771), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6765), .ZN(
        n6780) );
  AOI21_X1 U5866 ( .B1(n6771), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6768), .ZN(
        n6783) );
  AND2_X1 U5867 ( .A1(n9239), .A2(n9238), .ZN(n9719) );
  NAND2_X1 U5868 ( .A1(n6362), .A2(n6361), .ZN(n9316) );
  NAND2_X1 U5869 ( .A1(n4712), .A2(n4716), .ZN(n7650) );
  NAND2_X1 U5870 ( .A1(n7523), .A2(n6227), .ZN(n7581) );
  NAND2_X1 U5871 ( .A1(n6204), .A2(n6203), .ZN(n9733) );
  NAND2_X1 U5872 ( .A1(n7378), .A2(n6174), .ZN(n7311) );
  NAND2_X1 U5873 ( .A1(n4467), .A2(n4470), .ZN(n7310) );
  OR2_X1 U5874 ( .A1(n7380), .A2(n4472), .ZN(n4467) );
  INV_X1 U5875 ( .A(n7452), .ZN(n7247) );
  INV_X1 U5876 ( .A(n9740), .ZN(n9754) );
  INV_X1 U5877 ( .A(n9260), .ZN(n9559) );
  OAI21_X1 U5878 ( .B1(n7835), .B2(n9509), .A(n9793), .ZN(n4735) );
  INV_X1 U5879 ( .A(n8913), .ZN(n9566) );
  NAND2_X1 U5880 ( .A1(n6362), .A2(n4855), .ZN(n4853) );
  OR3_X1 U5881 ( .A1(n9519), .A2(n9518), .A3(n9517), .ZN(n9577) );
  NAND2_X1 U5882 ( .A1(n4841), .A2(n6322), .ZN(n9372) );
  NAND2_X1 U5883 ( .A1(n6288), .A2(n6287), .ZN(n9594) );
  NAND2_X1 U5884 ( .A1(n4475), .A2(n4478), .ZN(n7649) );
  NAND2_X1 U5885 ( .A1(n4477), .A2(n4476), .ZN(n4475) );
  INV_X1 U5886 ( .A(n8592), .ZN(n8890) );
  AND2_X1 U5887 ( .A1(n6828), .A2(n7557), .ZN(n9771) );
  AND2_X1 U5888 ( .A1(n6496), .A2(n6495), .ZN(n9608) );
  XNOR2_X1 U5889 ( .A(n5537), .B(n5536), .ZN(n9609) );
  OAI21_X1 U5890 ( .B1(n5546), .B2(n5545), .A(n5533), .ZN(n5537) );
  NOR2_X1 U5891 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6059) );
  INV_X1 U5892 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6064) );
  OR2_X1 U5893 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  INV_X1 U5894 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10146) );
  INV_X1 U5895 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7832) );
  INV_X1 U5896 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6922) );
  INV_X1 U5897 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10120) );
  AND2_X1 U5898 ( .A1(n6179), .A2(n6178), .ZN(n9637) );
  NOR2_X1 U5899 ( .A1(n4325), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9613) );
  INV_X1 U5900 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6696) );
  INV_X1 U5901 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6683) );
  INV_X1 U5902 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6688) );
  INV_X1 U5903 ( .A(n4538), .ZN(n7781) );
  NAND2_X1 U5904 ( .A1(n4531), .A2(n6975), .ZN(n4530) );
  NAND2_X1 U5905 ( .A1(n4532), .A2(n4795), .ZN(n4531) );
  OR2_X1 U5906 ( .A1(n6021), .A2(n9807), .ZN(n6026) );
  NOR2_X1 U5907 ( .A1(n4445), .A2(n6900), .ZN(n6960) );
  OR2_X1 U5908 ( .A1(n9160), .A2(n4651), .ZN(n4649) );
  INV_X1 U5909 ( .A(n4462), .ZN(n4461) );
  OR2_X1 U5910 ( .A1(n9252), .A2(n9101), .ZN(n4463) );
  OR2_X1 U5911 ( .A1(n9562), .A2(n9555), .ZN(n4464) );
  NAND2_X1 U5912 ( .A1(n4843), .A2(n9799), .ZN(n4847) );
  OAI22_X1 U5913 ( .A1(n9481), .A2(n6501), .B1(n9793), .B2(n6615), .ZN(n6616)
         );
  OR2_X1 U5914 ( .A1(n9562), .A2(n9606), .ZN(n4465) );
  AND2_X1 U5915 ( .A1(n4478), .A2(n4377), .ZN(n4347) );
  AND2_X1 U5916 ( .A1(n8908), .A2(n4489), .ZN(n4348) );
  OR2_X1 U5917 ( .A1(n9836), .A2(n5933), .ZN(n4349) );
  INV_X1 U5918 ( .A(n5193), .ZN(n5053) );
  NAND2_X1 U5919 ( .A1(n5004), .A2(n4951), .ZN(n5005) );
  AND4_X2 U5920 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n5789)
         );
  INV_X1 U5921 ( .A(n6979), .ZN(n4533) );
  AND2_X1 U5922 ( .A1(n4774), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4350) );
  NOR2_X1 U5923 ( .A1(n6473), .A2(n4406), .ZN(n6043) );
  INV_X1 U5924 ( .A(n5598), .ZN(n4630) );
  INV_X1 U5925 ( .A(n7404), .ZN(n4523) );
  INV_X1 U5926 ( .A(n4480), .ZN(n4476) );
  OR2_X1 U5927 ( .A1(n4481), .A2(n6240), .ZN(n4480) );
  OR2_X1 U5928 ( .A1(n7404), .A2(n4785), .ZN(n4351) );
  AND2_X1 U5929 ( .A1(n8157), .A2(n8156), .ZN(n4352) );
  AND4_X1 U5930 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n8908)
         );
  NOR2_X1 U5931 ( .A1(n7357), .A2(n7356), .ZN(n4353) );
  AND2_X1 U5932 ( .A1(n4662), .A2(n9023), .ZN(n4354) );
  NAND2_X1 U5933 ( .A1(n9065), .A2(n9090), .ZN(n9271) );
  INV_X1 U5934 ( .A(n9271), .ZN(n4675) );
  AND2_X1 U5935 ( .A1(n4825), .A2(n4440), .ZN(n4355) );
  AND2_X1 U5936 ( .A1(n4577), .A2(n4576), .ZN(n4356) );
  AND2_X1 U5937 ( .A1(n5811), .A2(n4914), .ZN(n4357) );
  AND2_X1 U5938 ( .A1(n4464), .A2(n4443), .ZN(n4358) );
  AND2_X1 U5939 ( .A1(n4465), .A2(n4439), .ZN(n4359) );
  AND2_X1 U5940 ( .A1(n4510), .A2(n4507), .ZN(n4360) );
  AND2_X1 U5941 ( .A1(n5929), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4361) );
  AND2_X1 U5942 ( .A1(n4781), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4362) );
  AND2_X1 U5943 ( .A1(n4517), .A2(n5925), .ZN(n4363) );
  NAND2_X1 U5944 ( .A1(n4946), .A2(n6678), .ZN(n4786) );
  AND2_X1 U5945 ( .A1(n4521), .A2(n4786), .ZN(n4364) );
  NAND2_X1 U5946 ( .A1(n4828), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4365) );
  INV_X1 U5947 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n4799) );
  INV_X1 U5948 ( .A(n6046), .ZN(n6116) );
  NAND2_X1 U5949 ( .A1(n5761), .A2(n4961), .ZN(n5759) );
  AND4_X1 U5950 ( .A1(n4975), .A2(n4974), .A3(n4973), .A4(n4972), .ZN(n6509)
         );
  AND4_X1 U5951 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n4989), .ZN(n4366)
         );
  AND2_X1 U5952 ( .A1(n4587), .A2(n6516), .ZN(n4367) );
  INV_X1 U5953 ( .A(n5053), .ZN(n5467) );
  AND2_X1 U5954 ( .A1(n4803), .A2(n4802), .ZN(n4368) );
  NAND2_X1 U5955 ( .A1(n6038), .A2(n4703), .ZN(n6467) );
  AND2_X1 U5956 ( .A1(n8949), .A2(n9125), .ZN(n9732) );
  NAND2_X1 U5957 ( .A1(n4853), .A2(n4854), .ZN(n9303) );
  NOR2_X1 U5958 ( .A1(n6382), .A2(n4852), .ZN(n4851) );
  NOR2_X1 U5959 ( .A1(n8477), .A2(n7868), .ZN(n4369) );
  AND3_X1 U5960 ( .A1(n4988), .A2(n4987), .A3(n4625), .ZN(n5783) );
  OR2_X1 U5961 ( .A1(n9095), .A2(n9161), .ZN(n4370) );
  AND2_X1 U5962 ( .A1(n4354), .A2(n9163), .ZN(n4371) );
  NAND2_X1 U5963 ( .A1(n4686), .A2(n4682), .ZN(n6890) );
  INV_X1 U5964 ( .A(n6890), .ZN(n7078) );
  OAI21_X1 U5965 ( .B1(n7927), .B2(n4912), .A(n4910), .ZN(n7934) );
  INV_X1 U5966 ( .A(n9032), .ZN(n4724) );
  INV_X1 U5967 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6474) );
  OR2_X1 U5968 ( .A1(n5995), .A2(n6979), .ZN(n4372) );
  INV_X1 U5969 ( .A(n9064), .ZN(n4674) );
  OR2_X1 U5970 ( .A1(n7180), .A2(n4946), .ZN(n4373) );
  AND3_X1 U5971 ( .A1(n6298), .A2(n6281), .A3(n6284), .ZN(n4374) );
  AND2_X1 U5972 ( .A1(n7293), .A2(n7288), .ZN(n4375) );
  AND2_X1 U5973 ( .A1(n4961), .A2(n4936), .ZN(n4376) );
  OR2_X1 U5974 ( .A1(n8609), .A2(n9184), .ZN(n4377) );
  OR2_X1 U5975 ( .A1(n9825), .A2(n5952), .ZN(n4378) );
  OR2_X1 U5976 ( .A1(n5107), .A2(n4730), .ZN(n4379) );
  AND2_X1 U5977 ( .A1(n4612), .A2(n4610), .ZN(n4380) );
  OR2_X1 U5978 ( .A1(n9296), .A2(n8908), .ZN(n9008) );
  NOR2_X1 U5979 ( .A1(n9594), .A2(n8822), .ZN(n4381) );
  NOR2_X1 U5980 ( .A1(n6112), .A2(n6696), .ZN(n4382) );
  NAND2_X1 U5981 ( .A1(n6332), .A2(n6331), .ZN(n9516) );
  AND2_X1 U5982 ( .A1(n5941), .A2(n6975), .ZN(n4383) );
  OR2_X1 U5983 ( .A1(n5844), .A2(n5843), .ZN(n4384) );
  INV_X1 U5984 ( .A(n8609), .ZN(n8925) );
  NOR2_X1 U5985 ( .A1(n7821), .A2(n4819), .ZN(n4385) );
  INV_X1 U5986 ( .A(n9086), .ZN(n4677) );
  AND2_X1 U5987 ( .A1(n6044), .A2(n9611), .ZN(n6048) );
  INV_X1 U5988 ( .A(n4573), .ZN(n9295) );
  NOR2_X1 U5989 ( .A1(n9309), .A2(n9296), .ZN(n4573) );
  AND2_X1 U5990 ( .A1(n4631), .A2(n5593), .ZN(n4386) );
  AND2_X1 U5991 ( .A1(n8913), .A2(n9175), .ZN(n4387) );
  AND2_X1 U5992 ( .A1(n5433), .A2(n5432), .ZN(n7938) );
  INV_X1 U5993 ( .A(n7938), .ZN(n8232) );
  AND2_X1 U5994 ( .A1(n4827), .A2(n4826), .ZN(n4388) );
  AND2_X1 U5995 ( .A1(n4755), .A2(n4754), .ZN(n4389) );
  AND2_X1 U5996 ( .A1(n8609), .A2(n9184), .ZN(n4390) );
  INV_X1 U5997 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U5998 ( .A1(n6552), .A2(n4614), .ZN(n4391) );
  NOR2_X1 U5999 ( .A1(n4670), .A2(n4671), .ZN(n4392) );
  AND2_X1 U6000 ( .A1(n5721), .A2(n6561), .ZN(n4393) );
  NOR2_X1 U6001 ( .A1(n9651), .A2(n9189), .ZN(n4394) );
  NOR2_X1 U6002 ( .A1(n7630), .A2(n6531), .ZN(n4395) );
  OR2_X1 U6003 ( .A1(n8501), .A2(n8248), .ZN(n4396) );
  AND2_X1 U6004 ( .A1(n9382), .A2(n9180), .ZN(n4397) );
  AND2_X1 U6005 ( .A1(n9545), .A2(n9182), .ZN(n4398) );
  OR2_X1 U6006 ( .A1(n8220), .A2(n8232), .ZN(n4399) );
  NAND2_X1 U6007 ( .A1(n8579), .A2(n8578), .ZN(n4400) );
  INV_X1 U6008 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4960) );
  AND2_X1 U6009 ( .A1(n6531), .A2(n7630), .ZN(n4401) );
  AND2_X1 U6010 ( .A1(n7501), .A2(n7247), .ZN(n4402) );
  OR2_X1 U6011 ( .A1(n5826), .A2(n8065), .ZN(n4403) );
  AND2_X1 U6012 ( .A1(n5235), .A2(SI_13_), .ZN(n4404) );
  NOR2_X1 U6013 ( .A1(n7895), .A2(n8216), .ZN(n4405) );
  OR2_X1 U6014 ( .A1(n4859), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4406) );
  AOI21_X1 U6015 ( .B1(n4677), .B2(n9075), .A(n4674), .ZN(n4673) );
  INV_X1 U6016 ( .A(n6551), .ZN(n6552) );
  NAND2_X1 U6017 ( .A1(n5721), .A2(n5572), .ZN(n6551) );
  AND2_X1 U6018 ( .A1(n8655), .A2(n8654), .ZN(n4407) );
  AND2_X1 U6019 ( .A1(n5217), .A2(SI_12_), .ZN(n4408) );
  INV_X1 U6020 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6682) );
  OR2_X1 U6021 ( .A1(n6691), .A2(n6070), .ZN(n4409) );
  AND2_X1 U6022 ( .A1(n7773), .A2(n8067), .ZN(n4410) );
  AND2_X1 U6023 ( .A1(n4602), .A2(n4399), .ZN(n4411) );
  AND2_X1 U6024 ( .A1(n4349), .A2(n4805), .ZN(n4412) );
  AND2_X1 U6025 ( .A1(n9336), .A2(n8984), .ZN(n4413) );
  AND2_X1 U6026 ( .A1(n4608), .A2(n4391), .ZN(n4414) );
  AND2_X1 U6027 ( .A1(n4831), .A2(n4829), .ZN(n4415) );
  NAND2_X1 U6028 ( .A1(n6531), .A2(n8067), .ZN(n4416) );
  INV_X1 U6029 ( .A(n4572), .ZN(n4660) );
  OAI21_X1 U6030 ( .B1(n9063), .B2(n9103), .A(n4446), .ZN(n4572) );
  INV_X1 U6031 ( .A(n5289), .ZN(n4561) );
  AND2_X1 U6032 ( .A1(n9323), .A2(n4565), .ZN(n4417) );
  AND2_X1 U6033 ( .A1(n8671), .A2(n8662), .ZN(n4418) );
  AND2_X1 U6034 ( .A1(n4546), .A2(n4502), .ZN(n4419) );
  AND2_X1 U6035 ( .A1(n9725), .A2(n6203), .ZN(n4420) );
  INV_X1 U6036 ( .A(n4860), .ZN(n4859) );
  NOR2_X1 U6037 ( .A1(n4861), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4860) );
  AND2_X1 U6038 ( .A1(n9064), .A2(n9269), .ZN(n9267) );
  INV_X1 U6039 ( .A(n9164), .ZN(n4657) );
  INV_X1 U6040 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4952) );
  INV_X1 U6041 ( .A(n4667), .ZN(n4666) );
  OAI211_X1 U6042 ( .C1(n4669), .C2(n4673), .A(n4675), .B(n4668), .ZN(n4667)
         );
  NAND2_X1 U6043 ( .A1(n4554), .A2(n6383), .ZN(n9296) );
  INV_X1 U6044 ( .A(n9296), .ZN(n4489) );
  NAND2_X1 U6045 ( .A1(n7539), .A2(n7629), .ZN(n7538) );
  NAND2_X1 U6046 ( .A1(n4743), .A2(n4746), .ZN(n8580) );
  OAI21_X1 U6047 ( .B1(n8346), .B2(n5645), .A(n5650), .ZN(n8285) );
  AND2_X1 U6048 ( .A1(n6154), .A2(n4858), .ZN(n6177) );
  INV_X1 U6049 ( .A(n5998), .ZN(n7402) );
  NAND2_X1 U6050 ( .A1(n6604), .A2(n6603), .ZN(n9011) );
  AND2_X1 U6051 ( .A1(n7530), .A2(n4579), .ZN(n4421) );
  NAND2_X1 U6052 ( .A1(n8360), .A2(n6539), .ZN(n8333) );
  INV_X1 U6053 ( .A(n5988), .ZN(n7735) );
  AND2_X1 U6054 ( .A1(n5154), .A2(n5161), .ZN(n5988) );
  XNOR2_X1 U6055 ( .A(n4986), .B(P2_IR_REG_1__SCAN_IN), .ZN(n5992) );
  INV_X1 U6056 ( .A(n5992), .ZN(n4504) );
  NAND2_X1 U6057 ( .A1(n4469), .A2(n4468), .ZN(n7486) );
  NAND2_X1 U6058 ( .A1(n4835), .A2(n6280), .ZN(n9419) );
  NAND2_X1 U6059 ( .A1(n6330), .A2(n6329), .ZN(n9357) );
  NAND2_X1 U6060 ( .A1(n6268), .A2(n6267), .ZN(n9437) );
  OR2_X1 U6061 ( .A1(n8987), .A2(n8933), .ZN(n4422) );
  NAND2_X1 U6062 ( .A1(n5516), .A2(n5515), .ZN(n6576) );
  NAND2_X1 U6063 ( .A1(n5498), .A2(n5497), .ZN(n7872) );
  INV_X1 U6064 ( .A(n7872), .ZN(n8418) );
  INV_X1 U6065 ( .A(n4719), .ZN(n4718) );
  AND2_X1 U6066 ( .A1(n5849), .A2(n7965), .ZN(n4423) );
  NOR2_X1 U6067 ( .A1(n8104), .A2(n5936), .ZN(n4424) );
  OR2_X1 U6068 ( .A1(n9603), .A2(n8821), .ZN(n8966) );
  AND2_X1 U6069 ( .A1(n4622), .A2(n6535), .ZN(n4425) );
  AND2_X1 U6070 ( .A1(n4781), .A2(n7807), .ZN(n4426) );
  NAND2_X1 U6071 ( .A1(n8648), .A2(n8854), .ZN(n4427) );
  AND2_X1 U6072 ( .A1(n5385), .A2(n5384), .ZN(n4428) );
  AND2_X1 U6073 ( .A1(n4752), .A2(n4753), .ZN(n4429) );
  INV_X1 U6074 ( .A(n4583), .ZN(n9349) );
  NOR2_X1 U6075 ( .A1(n9390), .A2(n4585), .ZN(n4583) );
  INV_X1 U6076 ( .A(n7785), .ZN(n4515) );
  AND2_X1 U6077 ( .A1(n8982), .A2(n9078), .ZN(n9360) );
  NOR2_X1 U6078 ( .A1(n7943), .A2(n4932), .ZN(n4430) );
  INV_X1 U6079 ( .A(n5984), .ZN(n7807) );
  AND2_X1 U6080 ( .A1(n5190), .A2(n5220), .ZN(n5984) );
  AND2_X1 U6081 ( .A1(n8776), .A2(n8777), .ZN(n4431) );
  AND2_X1 U6082 ( .A1(n4511), .A2(n4349), .ZN(n4432) );
  AND2_X1 U6083 ( .A1(n7802), .A2(n5958), .ZN(n4433) );
  AND2_X1 U6084 ( .A1(n6506), .A2(n4848), .ZN(n4434) );
  AND2_X1 U6085 ( .A1(n4756), .A2(n8586), .ZN(n4435) );
  OR2_X1 U6086 ( .A1(n4884), .A2(n4887), .ZN(n4436) );
  AND2_X1 U6087 ( .A1(n7243), .A2(n7247), .ZN(n4437) );
  NAND2_X1 U6088 ( .A1(n8397), .A2(n5632), .ZN(n8371) );
  NAND2_X1 U6089 ( .A1(n6259), .A2(n6258), .ZN(n9603) );
  INV_X1 U6090 ( .A(n9603), .ZN(n4576) );
  NAND2_X1 U6091 ( .A1(n7234), .A2(n7235), .ZN(n7233) );
  INV_X1 U6092 ( .A(n5052), .ZN(n5074) );
  NAND2_X1 U6093 ( .A1(n5930), .A2(n7807), .ZN(n5929) );
  AND2_X1 U6094 ( .A1(n4779), .A2(n5929), .ZN(n4438) );
  INV_X1 U6095 ( .A(n5925), .ZN(n5926) );
  NAND2_X1 U6096 ( .A1(n4775), .A2(n7735), .ZN(n5925) );
  AND3_X2 U6097 ( .A1(n7068), .A2(n6504), .A3(n9608), .ZN(n9799) );
  INV_X1 U6098 ( .A(n9799), .ZN(n4846) );
  AND2_X1 U6099 ( .A1(n7491), .A2(n7511), .ZN(n9509) );
  INV_X1 U6100 ( .A(n9509), .ZN(n9791) );
  OR2_X1 U6101 ( .A1(n7053), .A2(n7877), .ZN(n9844) );
  OR2_X1 U6102 ( .A1(n9793), .A2(n9561), .ZN(n4439) );
  OR2_X1 U6103 ( .A1(n5977), .A2(n5965), .ZN(n4440) );
  AND2_X1 U6104 ( .A1(n5949), .A2(n7171), .ZN(n4441) );
  INV_X1 U6105 ( .A(n4353), .ZN(n4748) );
  OR2_X1 U6106 ( .A1(n5977), .A2(n8342), .ZN(n4442) );
  OR2_X1 U6107 ( .A1(n9799), .A2(n9489), .ZN(n4443) );
  INV_X1 U6108 ( .A(n8113), .ZN(n4529) );
  OR2_X1 U6109 ( .A1(n6013), .A2(n8138), .ZN(n4444) );
  AND2_X1 U6110 ( .A1(n6902), .A2(n6901), .ZN(n4445) );
  OR2_X1 U6111 ( .A1(n9158), .A2(n6411), .ZN(n4446) );
  INV_X1 U6112 ( .A(n9170), .ZN(n4661) );
  INV_X1 U6113 ( .A(n5976), .ZN(n8138) );
  AND2_X1 U6114 ( .A1(n4784), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4447) );
  INV_X1 U6115 ( .A(n9800), .ZN(n4800) );
  INV_X1 U6116 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4732) );
  INV_X1 U6117 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n4824) );
  INV_X1 U6118 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n4818) );
  INV_X1 U6119 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4566) );
  OAI21_X1 U6120 ( .B1(n8985), .B2(n8995), .A(n4413), .ZN(n8986) );
  INV_X1 U6121 ( .A(n4580), .ZN(n6473) );
  NAND2_X1 U6122 ( .A1(n8977), .A2(n9161), .ZN(n4693) );
  NAND2_X1 U6123 ( .A1(n6937), .A2(n6423), .ZN(n6424) );
  NOR2_X1 U6124 ( .A1(n8975), .A2(n9137), .ZN(n8976) );
  AOI21_X1 U6125 ( .B1(n8967), .B2(n4681), .A(n4679), .ZN(n4678) );
  NOR3_X1 U6126 ( .A1(n9006), .A2(n9005), .A3(n9004), .ZN(n9009) );
  OR2_X1 U6127 ( .A1(n9253), .A2(n9430), .ZN(n4460) );
  NAND2_X1 U6128 ( .A1(n9114), .A2(n4723), .ZN(n7305) );
  NAND2_X1 U6129 ( .A1(n4883), .A2(n5121), .ZN(n5142) );
  NAND3_X1 U6130 ( .A1(n8778), .A2(n4431), .A3(n4450), .ZN(P1_U3220) );
  INV_X1 U6131 ( .A(n5949), .ZN(n4820) );
  OAI211_X1 U6132 ( .C1(n9836), .C2(n4551), .A(n4549), .B(n4548), .ZN(n9839)
         );
  NAND2_X1 U6133 ( .A1(n4542), .A2(n8138), .ZN(n5966) );
  NAND2_X1 U6134 ( .A1(n6026), .A2(n4419), .ZN(P2_U3201) );
  XNOR2_X1 U6135 ( .A(n5953), .B(n5988), .ZN(n7724) );
  XNOR2_X1 U6136 ( .A(n5970), .B(n6017), .ZN(n4547) );
  NAND2_X1 U6137 ( .A1(n4547), .A2(n9815), .ZN(n4546) );
  NAND2_X1 U6138 ( .A1(n7426), .A2(n5807), .ZN(n5810) );
  NAND2_X1 U6139 ( .A1(n5784), .A2(n8077), .ZN(n4454) );
  AND2_X2 U6140 ( .A1(n4924), .A2(n4921), .ZN(n7901) );
  NAND2_X1 U6141 ( .A1(n6950), .A2(n6951), .ZN(n6949) );
  NAND3_X1 U6142 ( .A1(n6949), .A2(n5792), .A3(n5793), .ZN(n7044) );
  NOR2_X2 U6143 ( .A1(n7944), .A2(n7945), .ZN(n7943) );
  NAND2_X1 U6144 ( .A1(n4862), .A2(n5387), .ZN(n5400) );
  NAND2_X1 U6145 ( .A1(n5476), .A2(n4865), .ZN(n4870) );
  NAND2_X1 U6146 ( .A1(n4571), .A2(n4888), .ZN(n5248) );
  NAND2_X1 U6147 ( .A1(n5086), .A2(n5085), .ZN(n5104) );
  NAND2_X1 U6148 ( .A1(n4653), .A2(n4661), .ZN(n4651) );
  INV_X1 U6149 ( .A(n9030), .ZN(n9091) );
  NAND2_X1 U6150 ( .A1(n4983), .A2(n4569), .ZN(n4734) );
  OAI21_X1 U6151 ( .B1(n4555), .B2(n4436), .A(n4885), .ZN(n5438) );
  OR2_X2 U6152 ( .A1(n9337), .A2(n9057), .ZN(n6448) );
  AOI211_X2 U6153 ( .C1(n9492), .C2(n9791), .A(n9491), .B(n9490), .ZN(n9563)
         );
  OAI21_X2 U6154 ( .B1(n7525), .B2(n4715), .A(n4713), .ZN(n9455) );
  OR2_X1 U6155 ( .A1(n9726), .A2(n9725), .ZN(n6434) );
  NAND2_X1 U6156 ( .A1(n5118), .A2(n5117), .ZN(n4883) );
  NAND3_X1 U6157 ( .A1(n4463), .A2(n4461), .A3(n4460), .ZN(P1_U3262) );
  NAND2_X1 U6158 ( .A1(n4857), .A2(n6154), .ZN(n6192) );
  NOR2_X2 U6159 ( .A1(n6138), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U6160 ( .A1(n8782), .A2(n8672), .ZN(n8675) );
  NAND2_X1 U6161 ( .A1(n5158), .A2(n4945), .ZN(n5160) );
  NAND2_X1 U6162 ( .A1(n4727), .A2(n4726), .ZN(n5158) );
  INV_X1 U6163 ( .A(n4716), .ZN(n4715) );
  NAND2_X1 U6164 ( .A1(n5203), .A2(n4890), .ZN(n4571) );
  NAND2_X1 U6165 ( .A1(n4708), .A2(n4706), .ZN(n9359) );
  OAI21_X1 U6166 ( .B1(n9560), .B2(n4846), .A(n4358), .ZN(P1_U3551) );
  OAI21_X1 U6167 ( .B1(n9560), .B2(n6614), .A(n4359), .ZN(P1_U3519) );
  NAND2_X1 U6168 ( .A1(n7380), .A2(n4470), .ZN(n4469) );
  INV_X1 U6169 ( .A(n7524), .ZN(n4477) );
  NAND2_X1 U6170 ( .A1(n4473), .A2(n4474), .ZN(n9451) );
  NAND2_X1 U6171 ( .A1(n7524), .A2(n4347), .ZN(n4473) );
  NAND2_X1 U6172 ( .A1(n6362), .A2(n4486), .ZN(n4484) );
  NAND2_X1 U6173 ( .A1(n4484), .A2(n4485), .ZN(n6400) );
  OAI21_X1 U6174 ( .B1(n6362), .B2(n4488), .A(n4849), .ZN(n9289) );
  NAND2_X1 U6175 ( .A1(n6268), .A2(n4490), .ZN(n4835) );
  NAND2_X1 U6176 ( .A1(n4835), .A2(n4833), .ZN(n6296) );
  XNOR2_X1 U6177 ( .A(n5118), .B(n5117), .ZN(n6698) );
  MUX2_X1 U6178 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5145), .Z(n5042) );
  AND2_X2 U6179 ( .A1(n4568), .A2(n4878), .ZN(n5145) );
  AND2_X2 U6180 ( .A1(n5087), .A2(n4499), .ZN(n5301) );
  AND2_X2 U6181 ( .A1(n5067), .A2(n5068), .ZN(n5087) );
  MUX2_X1 U6182 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n5971), .Z(n7051) );
  MUX2_X1 U6183 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n5971), .Z(n5993) );
  NOR2_X1 U6184 ( .A1(n7816), .A2(n5932), .ZN(n5933) );
  NAND3_X1 U6185 ( .A1(n4780), .A2(n4362), .A3(n5929), .ZN(n4505) );
  NAND2_X1 U6186 ( .A1(n9842), .A2(n4349), .ZN(n4507) );
  NAND2_X1 U6187 ( .A1(n9842), .A2(n4412), .ZN(n4508) );
  INV_X1 U6188 ( .A(n4511), .ZN(n9841) );
  NAND2_X1 U6189 ( .A1(n4513), .A2(n4512), .ZN(n7784) );
  NAND2_X1 U6190 ( .A1(n5926), .A2(n4515), .ZN(n4512) );
  INV_X1 U6191 ( .A(n4518), .ZN(n4514) );
  INV_X1 U6192 ( .A(n4774), .ZN(n4516) );
  INV_X1 U6193 ( .A(n4517), .ZN(n7725) );
  NAND2_X1 U6194 ( .A1(n4783), .A2(n4523), .ZN(n4519) );
  NAND3_X1 U6195 ( .A1(n4784), .A2(n4520), .A3(n4521), .ZN(n4522) );
  INV_X1 U6196 ( .A(n8105), .ZN(n4527) );
  NAND2_X1 U6197 ( .A1(n5936), .A2(n4529), .ZN(n4528) );
  NAND3_X1 U6198 ( .A1(n4415), .A2(n8154), .A3(n4530), .ZN(P2_U3200) );
  INV_X1 U6199 ( .A(n4537), .ZN(n4535) );
  AND2_X1 U6200 ( .A1(n4537), .A2(n9928), .ZN(n4536) );
  XNOR2_X1 U6201 ( .A(n5952), .B(n9825), .ZN(n4537) );
  NAND3_X1 U6202 ( .A1(n4543), .A2(n4825), .A3(n4440), .ZN(n4542) );
  NAND2_X1 U6203 ( .A1(n4544), .A2(n5966), .ZN(n8141) );
  NAND3_X1 U6204 ( .A1(n4355), .A2(n4543), .A3(n5976), .ZN(n4544) );
  NOR2_X1 U6205 ( .A1(n8141), .A2(n8450), .ZN(n8140) );
  NAND2_X1 U6206 ( .A1(n7821), .A2(n6821), .ZN(n4548) );
  OR2_X1 U6207 ( .A1(n7821), .A2(n4550), .ZN(n4549) );
  NAND3_X1 U6208 ( .A1(n9059), .A2(n9091), .A3(n4562), .ZN(n9098) );
  NAND4_X1 U6209 ( .A1(n9267), .A2(n9058), .A3(n4417), .A4(n9290), .ZN(n4564)
         );
  INV_X1 U6210 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4567) );
  INV_X1 U6211 ( .A(n4570), .ZN(n4983) );
  NAND3_X1 U6212 ( .A1(n4568), .A2(n4878), .A3(n6687), .ZN(n5012) );
  AOI21_X1 U6213 ( .B1(n4658), .B2(n4572), .A(n4657), .ZN(n4656) );
  MUX2_X1 U6214 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9628), .S(n6632), .Z(n9473) );
  NAND2_X1 U6215 ( .A1(n4356), .A2(n7530), .ZN(n9459) );
  INV_X1 U6216 ( .A(n6192), .ZN(n6038) );
  NAND2_X1 U6217 ( .A1(n4580), .A2(n4860), .ZN(n6058) );
  NOR2_X2 U6218 ( .A1(n6192), .A2(n4581), .ZN(n4580) );
  INV_X1 U6219 ( .A(n6037), .ZN(n4581) );
  INV_X1 U6220 ( .A(n4582), .ZN(n4949) );
  NAND2_X1 U6221 ( .A1(n7209), .A2(n7208), .ZN(n4590) );
  NAND2_X1 U6222 ( .A1(n4590), .A2(n4588), .ZN(n4587) );
  NAND2_X1 U6223 ( .A1(n4590), .A2(n6512), .ZN(n7225) );
  INV_X1 U6224 ( .A(n7663), .ZN(n6532) );
  NAND2_X1 U6225 ( .A1(n8241), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U6226 ( .A1(n8178), .A2(n4414), .ZN(n4606) );
  OAI211_X1 U6227 ( .C1(n8178), .C2(n4607), .A(n8392), .B(n4606), .ZN(n6567)
         );
  OAI21_X1 U6228 ( .B1(n8178), .B2(n4369), .A(n6548), .ZN(n7848) );
  NAND2_X1 U6229 ( .A1(n5301), .A2(n4623), .ZN(n4976) );
  AND2_X1 U6230 ( .A1(n5301), .A2(n4624), .ZN(n4978) );
  INV_X1 U6231 ( .A(n4976), .ZN(n4965) );
  NAND2_X4 U6232 ( .A1(n4997), .A2(n4325), .ZN(n5046) );
  NAND2_X1 U6233 ( .A1(n7224), .A2(n4627), .ZN(n4628) );
  NAND2_X1 U6234 ( .A1(n4628), .A2(n4629), .ZN(n7319) );
  NAND2_X1 U6235 ( .A1(n8399), .A2(n5632), .ZN(n4632) );
  NAND2_X1 U6236 ( .A1(n4632), .A2(n4633), .ZN(n5232) );
  AOI21_X1 U6237 ( .B1(n8400), .B2(n5632), .A(n4634), .ZN(n4633) );
  NAND2_X1 U6238 ( .A1(n7416), .A2(n7415), .ZN(n7418) );
  NAND2_X1 U6239 ( .A1(n7418), .A2(n4635), .ZN(n5133) );
  NAND4_X1 U6240 ( .A1(n4640), .A2(n4639), .A3(n4953), .A4(n4638), .ZN(n4637)
         );
  NAND2_X1 U6241 ( .A1(n7625), .A2(n4646), .ZN(n4643) );
  NAND2_X1 U6242 ( .A1(n4643), .A2(n4644), .ZN(n7661) );
  NAND2_X1 U6243 ( .A1(n5576), .A2(n5578), .ZN(n6508) );
  NAND3_X1 U6244 ( .A1(n5576), .A2(n5578), .A3(n4998), .ZN(n7007) );
  NAND2_X1 U6245 ( .A1(n7007), .A2(n5578), .ZN(n7207) );
  NAND3_X1 U6246 ( .A1(n4649), .A2(n4648), .A3(n9169), .ZN(P1_U3242) );
  NAND2_X1 U6247 ( .A1(n9160), .A2(n4650), .ZN(n4648) );
  OR2_X1 U6248 ( .A1(n9009), .A2(n4667), .ZN(n4663) );
  NAND2_X1 U6249 ( .A1(n4663), .A2(n4664), .ZN(n9028) );
  NOR2_X1 U6250 ( .A1(n4674), .A2(n9161), .ZN(n4676) );
  AOI21_X1 U6251 ( .B1(n8968), .B2(n9023), .A(n4678), .ZN(n8975) );
  NAND2_X2 U6252 ( .A1(n6632), .A2(n6070), .ZN(n6112) );
  NAND2_X1 U6253 ( .A1(n4685), .A2(n6612), .ZN(n4686) );
  OAI21_X2 U6254 ( .B1(n6927), .B2(n6422), .A(n9111), .ZN(n6937) );
  NAND2_X1 U6255 ( .A1(n4697), .A2(n8943), .ZN(n8946) );
  NAND2_X1 U6256 ( .A1(n8942), .A2(n8941), .ZN(n4697) );
  NAND2_X1 U6257 ( .A1(n4699), .A2(n4698), .ZN(n8942) );
  OR2_X1 U6258 ( .A1(n8937), .A2(n9023), .ZN(n4698) );
  INV_X1 U6259 ( .A(n8936), .ZN(n4699) );
  NAND2_X1 U6260 ( .A1(n6038), .A2(n4700), .ZN(n4704) );
  NAND2_X1 U6261 ( .A1(n9028), .A2(n4938), .ZN(n9160) );
  XNOR2_X2 U6262 ( .A(n6065), .B(n6064), .ZN(n6612) );
  NAND2_X1 U6263 ( .A1(n9396), .A2(n4709), .ZN(n4708) );
  OR2_X2 U6264 ( .A1(n7237), .A2(n9043), .ZN(n9114) );
  OR2_X1 U6265 ( .A1(n6432), .A2(n7236), .ZN(n9043) );
  NAND2_X1 U6266 ( .A1(n5108), .A2(n4729), .ZN(n4726) );
  NAND2_X1 U6267 ( .A1(n5108), .A2(n5107), .ZN(n5118) );
  NAND3_X1 U6268 ( .A1(n6902), .A2(n6901), .A3(n6959), .ZN(n4736) );
  NAND2_X1 U6269 ( .A1(n6959), .A2(n4738), .ZN(n6900) );
  INV_X1 U6270 ( .A(n6899), .ZN(n4740) );
  AOI22_X1 U6271 ( .A1(n6854), .A2(n6855), .B1(n6853), .B2(n8761), .ZN(n6861)
         );
  NAND2_X1 U6272 ( .A1(n7444), .A2(n4744), .ZN(n4742) );
  INV_X1 U6273 ( .A(n4756), .ZN(n9643) );
  NAND2_X1 U6274 ( .A1(n8799), .A2(n4760), .ZN(n4759) );
  AND2_X1 U6275 ( .A1(n8722), .A2(n8800), .ZN(n4760) );
  NAND2_X1 U6276 ( .A1(n8663), .A2(n4418), .ZN(n8782) );
  NAND2_X1 U6277 ( .A1(n6411), .A2(n9101), .ZN(n6622) );
  NAND2_X1 U6278 ( .A1(n8840), .A2(n7288), .ZN(n4770) );
  NAND2_X1 U6279 ( .A1(n4770), .A2(n7292), .ZN(n4771) );
  NAND2_X1 U6280 ( .A1(n7604), .A2(n4777), .ZN(n4774) );
  NAND2_X1 U6281 ( .A1(n4780), .A2(n5929), .ZN(n7810) );
  NAND2_X1 U6282 ( .A1(n4782), .A2(n5984), .ZN(n4780) );
  INV_X1 U6283 ( .A(n4786), .ZN(n4785) );
  INV_X1 U6284 ( .A(n4792), .ZN(n8153) );
  NAND2_X1 U6285 ( .A1(n4790), .A2(n4788), .ZN(n4794) );
  NAND2_X1 U6286 ( .A1(n8129), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U6287 ( .A1(n4792), .A2(n4791), .ZN(n4795) );
  XNOR2_X1 U6288 ( .A(n4794), .B(n4793), .ZN(n5941) );
  INV_X1 U6289 ( .A(n6018), .ZN(n4793) );
  NAND2_X1 U6290 ( .A1(n9800), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4801) );
  AND2_X1 U6291 ( .A1(n9800), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4804) );
  OAI21_X1 U6292 ( .B1(n9813), .B2(n9812), .A(n4806), .ZN(n9814) );
  NAND2_X1 U6293 ( .A1(n4814), .A2(n4813), .ZN(n7821) );
  NAND2_X1 U6294 ( .A1(n7803), .A2(n4817), .ZN(n4814) );
  NAND2_X1 U6295 ( .A1(n4820), .A2(n7171), .ZN(n4821) );
  NAND2_X1 U6296 ( .A1(n5964), .A2(n4828), .ZN(n4825) );
  XNOR2_X1 U6297 ( .A(n5963), .B(n8100), .ZN(n8096) );
  OAI22_X1 U6298 ( .A1(n8160), .A2(n8159), .B1(n9805), .B2(n9946), .ZN(n4830)
         );
  OAI21_X1 U6299 ( .B1(n8155), .B2(n4352), .A(n9815), .ZN(n4831) );
  NOR2_X4 U6300 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6105) );
  NAND3_X1 U6301 ( .A1(n4832), .A2(n6105), .A3(n6082), .ZN(n6136) );
  NAND2_X1 U6302 ( .A1(n4841), .A2(n4839), .ZN(n6330) );
  NAND2_X1 U6303 ( .A1(n9735), .A2(n6217), .ZN(n7524) );
  NAND2_X1 U6304 ( .A1(n6204), .A2(n4420), .ZN(n9735) );
  INV_X1 U6305 ( .A(n7835), .ZN(n4842) );
  NAND2_X1 U6306 ( .A1(n4842), .A2(n4845), .ZN(n4844) );
  NAND3_X1 U6307 ( .A1(n4847), .A2(n4844), .A3(n4434), .ZN(P1_U3550) );
  NOR2_X1 U6308 ( .A1(n6473), .A2(n4861), .ZN(n6057) );
  NAND2_X1 U6309 ( .A1(n5370), .A2(n4863), .ZN(n4862) );
  NAND2_X1 U6310 ( .A1(n5476), .A2(n5475), .ZN(n4872) );
  NAND2_X1 U6311 ( .A1(n4872), .A2(n5477), .ZN(n5494) );
  INV_X1 U6312 ( .A(n5493), .ZN(n4871) );
  NOR2_X2 U6313 ( .A1(n5707), .A2(n5708), .ZN(n5713) );
  NAND2_X1 U6314 ( .A1(n4877), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4880) );
  NAND3_X1 U6315 ( .A1(n4877), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U6316 ( .A1(n5402), .A2(n5401), .ZN(n5408) );
  OR2_X1 U6317 ( .A1(n5203), .A2(n5202), .ZN(n4896) );
  NAND2_X1 U6318 ( .A1(n4904), .A2(n4902), .ZN(n4907) );
  NAND2_X1 U6319 ( .A1(n5295), .A2(n5294), .ZN(n5319) );
  AND2_X1 U6320 ( .A1(n7044), .A2(n5795), .ZN(n7159) );
  NAND2_X1 U6321 ( .A1(n7927), .A2(n4910), .ZN(n4909) );
  NAND2_X1 U6322 ( .A1(n8021), .A2(n4913), .ZN(n7426) );
  NAND3_X1 U6323 ( .A1(n4952), .A2(n5004), .A3(n4951), .ZN(n5021) );
  AOI21_X2 U6324 ( .B1(n7885), .B2(n7886), .A(n4917), .ZN(n8048) );
  OAI21_X2 U6325 ( .B1(n7977), .B2(n7978), .A(n4403), .ZN(n7885) );
  OR2_X1 U6326 ( .A1(n7943), .A2(n4925), .ZN(n4924) );
  AND2_X1 U6327 ( .A1(n5829), .A2(n8326), .ZN(n4932) );
  AND2_X1 U6328 ( .A1(n5764), .A2(n4960), .ZN(n5761) );
  NAND2_X1 U6329 ( .A1(n7351), .A2(n7350), .ZN(n7444) );
  NAND2_X1 U6330 ( .A1(n6935), .A2(n6099), .ZN(n7015) );
  NAND2_X1 U6331 ( .A1(n4997), .A2(n6070), .ZN(n5023) );
  NAND2_X1 U6332 ( .A1(n7853), .A2(n5507), .ZN(n6507) );
  OAI21_X1 U6333 ( .B1(n4978), .B2(n4977), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n4980) );
  NAND2_X1 U6334 ( .A1(n5073), .A2(n5602), .ZN(n7437) );
  NAND2_X1 U6335 ( .A1(n8077), .A2(n7011), .ZN(n5576) );
  INV_X1 U6336 ( .A(n5035), .ZN(n5553) );
  OR2_X1 U6337 ( .A1(n7955), .A2(n8340), .ZN(n4937) );
  INV_X1 U6338 ( .A(n8543), .ZN(n6577) );
  INV_X1 U6339 ( .A(n7983), .ZN(n5886) );
  AND2_X1 U6340 ( .A1(n9793), .A2(n9546), .ZN(n9604) );
  INV_X1 U6341 ( .A(n9793), .ZN(n6614) );
  AND2_X1 U6342 ( .A1(n9027), .A2(n4370), .ZN(n4938) );
  INV_X1 U6343 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6498) );
  INV_X1 U6344 ( .A(n9825), .ZN(n6697) );
  INV_X1 U6345 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4963) );
  NOR2_X1 U6346 ( .A1(n6063), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4939) );
  OR2_X1 U6347 ( .A1(n5252), .A2(n5251), .ZN(n4940) );
  NOR2_X1 U6348 ( .A1(n6528), .A2(n7470), .ZN(n4941) );
  NOR2_X1 U6349 ( .A1(n7261), .A2(n6516), .ZN(n4942) );
  AND2_X1 U6350 ( .A1(n5848), .A2(n7931), .ZN(n4943) );
  AND4_X1 U6351 ( .A1(n6254), .A2(n6253), .A3(n6252), .A4(n10117), .ZN(n4944)
         );
  AND2_X1 U6352 ( .A1(n5159), .A2(n5150), .ZN(n4945) );
  AND2_X1 U6353 ( .A1(n7190), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4946) );
  INV_X1 U6354 ( .A(n9103), .ZN(n6835) );
  INV_X1 U6355 ( .A(n7006), .ZN(n4998) );
  INV_X1 U6356 ( .A(n7626), .ZN(n5157) );
  INV_X1 U6357 ( .A(n6576), .ZN(n8169) );
  AND2_X1 U6358 ( .A1(n8293), .A2(n8294), .ZN(n4947) );
  AND2_X1 U6359 ( .A1(n8273), .A2(n8274), .ZN(n4950) );
  NAND2_X2 U6360 ( .A1(n7074), .A2(n9401), .ZN(n9470) );
  AND2_X1 U6361 ( .A1(n8944), .A2(n9117), .ZN(n8945) );
  AND2_X1 U6362 ( .A1(n8960), .A2(n9129), .ZN(n8961) );
  NAND2_X1 U6363 ( .A1(n9105), .A2(n8974), .ZN(n8969) );
  AOI21_X1 U6364 ( .B1(n8971), .B2(n8970), .A(n8969), .ZN(n8978) );
  OR2_X1 U6365 ( .A1(n8574), .A2(n8573), .ZN(n8579) );
  INV_X1 U6366 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6252) );
  INV_X1 U6367 ( .A(n9029), .ZN(n6411) );
  INV_X1 U6368 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5134) );
  AND2_X1 U6369 ( .A1(n8336), .A2(n8334), .ZN(n6540) );
  OAI22_X1 U6370 ( .A1(n7078), .A2(n7352), .B1(n6856), .B2(n8764), .ZN(n6857)
         );
  OAI22_X1 U6371 ( .A1(n6938), .A2(n8764), .B1(n7087), .B2(n7352), .ZN(n6894)
         );
  INV_X1 U6372 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6040) );
  INV_X1 U6373 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6374 ( .A1(n5569), .A2(n6553), .ZN(n5571) );
  OR2_X1 U6375 ( .A1(n5046), .A2(n6680), .ZN(n5014) );
  INV_X1 U6376 ( .A(n5723), .ZN(n5416) );
  OR2_X1 U6377 ( .A1(n5151), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5185) );
  OAI21_X1 U6378 ( .B1(n6856), .B2(n8677), .A(n6858), .ZN(n6859) );
  OR2_X1 U6379 ( .A1(n6261), .A2(n6260), .ZN(n6274) );
  INV_X1 U6380 ( .A(n7371), .ZN(n7239) );
  AND2_X1 U6381 ( .A1(n5417), .A2(n5406), .ZN(n5407) );
  INV_X1 U6382 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6269) );
  INV_X1 U6383 ( .A(n7429), .ZN(n5805) );
  INV_X1 U6384 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6385 ( .A1(n5571), .A2(n5570), .ZN(n5720) );
  NOR2_X1 U6386 ( .A1(n6666), .A2(n5918), .ZN(n9803) );
  INV_X1 U6387 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5033) );
  AND2_X1 U6388 ( .A1(n6561), .A2(n6557), .ZN(n6580) );
  INV_X1 U6389 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4964) );
  AND2_X1 U6390 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NOR2_X1 U6391 ( .A1(n6377), .A2(n6376), .ZN(n6385) );
  OR2_X1 U6392 ( .A1(n6343), .A2(n6342), .ZN(n6353) );
  INV_X1 U6393 ( .A(n9011), .ZN(n6605) );
  INV_X1 U6394 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6209) );
  AND2_X1 U6395 ( .A1(n6129), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6143) );
  AND2_X1 U6396 ( .A1(n6831), .A2(n6459), .ZN(n8874) );
  INV_X1 U6397 ( .A(n7530), .ZN(n9738) );
  INV_X1 U6398 ( .A(n6632), .ZN(n6299) );
  INV_X1 U6399 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6413) );
  INV_X1 U6400 ( .A(n5215), .ZN(n5218) );
  AOI21_X1 U6401 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8085), .A(n8086), .ZN(
        n5963) );
  INV_X1 U6402 ( .A(n6541), .ZN(n8321) );
  INV_X1 U6403 ( .A(n7485), .ZN(n7200) );
  AND2_X1 U6404 ( .A1(n5592), .A2(n5599), .ZN(n7226) );
  INV_X1 U6405 ( .A(n8067), .ZN(n7630) );
  INV_X1 U6406 ( .A(n8392), .ZN(n8323) );
  XNOR2_X1 U6407 ( .A(n5757), .B(n5756), .ZN(n5973) );
  OR2_X1 U6408 ( .A1(n6303), .A2(n8752), .ZN(n6315) );
  AND2_X1 U6409 ( .A1(n7572), .A2(n7571), .ZN(n8575) );
  AND2_X1 U6410 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6117) );
  INV_X1 U6411 ( .A(n8620), .ZN(n8917) );
  NOR2_X1 U6412 ( .A1(n6353), .A2(n8836), .ZN(n6365) );
  NOR2_X1 U6413 ( .A1(n6315), .A2(n8856), .ZN(n6325) );
  INV_X1 U6414 ( .A(n8648), .ZN(n9535) );
  NOR2_X1 U6415 ( .A1(n6210), .A2(n6209), .ZN(n6221) );
  INV_X1 U6416 ( .A(n9167), .ZN(n9276) );
  OR2_X1 U6417 ( .A1(n7074), .A2(n9430), .ZN(n9740) );
  INV_X1 U6418 ( .A(n9505), .ZN(n9736) );
  OR2_X1 U6419 ( .A1(n9161), .A2(n6835), .ZN(n7511) );
  OAI21_X1 U6420 ( .B1(n9768), .B2(P1_D_REG_1__SCAN_IN), .A(n6492), .ZN(n7066)
         );
  NAND2_X1 U6421 ( .A1(n5458), .A2(n5457), .ZN(n5476) );
  OR2_X1 U6422 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6405) );
  OAI21_X1 U6423 ( .B1(n8477), .B2(n8058), .A(n5909), .ZN(n5910) );
  AND2_X1 U6424 ( .A1(n5904), .A2(n5903), .ZN(n6844) );
  INV_X1 U6425 ( .A(n8049), .ZN(n8038) );
  INV_X1 U6426 ( .A(n8052), .ZN(n8043) );
  AND2_X1 U6427 ( .A1(n5557), .A2(n5522), .ZN(n7869) );
  INV_X1 U6428 ( .A(n9849), .ZN(n9807) );
  NOR2_X1 U6429 ( .A1(n9819), .A2(n5923), .ZN(n7607) );
  INV_X1 U6430 ( .A(n9805), .ZN(n9835) );
  AND2_X1 U6431 ( .A1(P2_U3893), .A2(n5771), .ZN(n9849) );
  INV_X1 U6432 ( .A(n8139), .ZN(n9837) );
  NAND2_X1 U6433 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  NAND2_X1 U6434 ( .A1(n6720), .A2(n5888), .ZN(n8227) );
  INV_X1 U6435 ( .A(n8403), .ZN(n8381) );
  INV_X1 U6436 ( .A(n8457), .ZN(n6594) );
  AND2_X1 U6437 ( .A1(n9938), .A2(n9915), .ZN(n8445) );
  AND2_X1 U6438 ( .A1(n5725), .A2(n5724), .ZN(n8260) );
  INV_X1 U6439 ( .A(n8552), .ZN(n8523) );
  INV_X1 U6440 ( .A(n6538), .ZN(n8348) );
  NAND2_X1 U6441 ( .A1(n9901), .A2(n9902), .ZN(n9915) );
  AND2_X1 U6442 ( .A1(n5857), .A2(n5856), .ZN(n6708) );
  INV_X1 U6443 ( .A(n9641), .ZN(n8895) );
  INV_X1 U6444 ( .A(n8924), .ZN(n8912) );
  AND3_X1 U6445 ( .A1(n9016), .A2(n9015), .A3(n9014), .ZN(n9275) );
  OR2_X1 U6446 ( .A1(n9318), .A2(n6367), .ZN(n6372) );
  INV_X1 U6447 ( .A(n4345), .ZN(n6367) );
  AND4_X1 U6448 ( .A1(n6226), .A2(n6225), .A3(n6224), .A4(n6223), .ZN(n8790)
         );
  OR2_X1 U6449 ( .A1(n6649), .A2(n6648), .ZN(n9668) );
  INV_X1 U6450 ( .A(n9716), .ZN(n9700) );
  INV_X1 U6451 ( .A(n9709), .ZN(n9660) );
  AND2_X1 U6452 ( .A1(n6739), .A2(n6643), .ZN(n9716) );
  INV_X1 U6453 ( .A(n9057), .ZN(n9336) );
  INV_X1 U6454 ( .A(n9466), .ZN(n9764) );
  INV_X1 U6455 ( .A(n9760), .ZN(n9745) );
  AND2_X1 U6456 ( .A1(n9799), .A2(n9546), .ZN(n9553) );
  INV_X1 U6457 ( .A(n6961), .ZN(n7191) );
  AND2_X1 U6458 ( .A1(n7066), .A2(n6837), .ZN(n6504) );
  INV_X1 U6459 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6298) );
  AND2_X1 U6460 ( .A1(n6241), .A2(n6230), .ZN(n9693) );
  INV_X1 U6461 ( .A(n5910), .ZN(n5911) );
  AND2_X1 U6462 ( .A1(n6844), .A2(n7560), .ZN(n8040) );
  AND2_X1 U6463 ( .A1(n5880), .A2(n5879), .ZN(n7983) );
  INV_X1 U6464 ( .A(n8030), .ZN(n8058) );
  AND4_X1 U6465 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n8362)
         );
  OR2_X1 U6466 ( .A1(n6723), .A2(n5914), .ZN(n8073) );
  OR2_X1 U6467 ( .A1(n7053), .A2(n5971), .ZN(n9853) );
  INV_X1 U6468 ( .A(n8406), .ZN(n8384) );
  NAND2_X1 U6469 ( .A1(n9938), .A2(n9914), .ZN(n8457) );
  INV_X1 U6470 ( .A(n9938), .ZN(n9935) );
  INV_X1 U6471 ( .A(n8410), .ZN(n8466) );
  OR2_X1 U6472 ( .A1(n9921), .A2(n9893), .ZN(n8543) );
  OR2_X1 U6473 ( .A1(n9921), .A2(n8473), .ZN(n8552) );
  AND2_X1 U6474 ( .A1(n6574), .A2(n6573), .ZN(n9921) );
  INV_X1 U6475 ( .A(n6729), .ZN(n6731) );
  INV_X1 U6476 ( .A(n6581), .ZN(n6720) );
  INV_X1 U6477 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8566) );
  INV_X1 U6478 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U6479 ( .A1(n6966), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9653) );
  INV_X1 U6480 ( .A(n9650), .ZN(n8924) );
  INV_X1 U6481 ( .A(n8905), .ZN(n9646) );
  INV_X1 U6482 ( .A(n7527), .ZN(n9187) );
  OR2_X1 U6483 ( .A1(n6649), .A2(n9165), .ZN(n9709) );
  NAND2_X1 U6484 ( .A1(n6642), .A2(n6640), .ZN(n9724) );
  OR2_X1 U6485 ( .A1(n9767), .A2(n7071), .ZN(n7498) );
  AND2_X1 U6486 ( .A1(n7498), .A2(n7083), .ZN(n9466) );
  NAND2_X1 U6487 ( .A1(n9799), .A2(n9791), .ZN(n9555) );
  NAND2_X1 U6488 ( .A1(n8773), .A2(n9604), .ZN(n6502) );
  NAND2_X1 U6489 ( .A1(n9793), .A2(n9791), .ZN(n9606) );
  AND3_X2 U6490 ( .A1(n7068), .A2(n6504), .A3(n6497), .ZN(n9793) );
  NAND2_X1 U6491 ( .A1(n9771), .A2(n9768), .ZN(n9972) );
  INV_X1 U6492 ( .A(n6047), .ZN(n7846) );
  INV_X1 U6493 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U6494 ( .A1(n4325), .A2(P1_U3086), .ZN(n9626) );
  INV_X2 U6495 ( .A(n8073), .ZN(P2_U3893) );
  NOR2_X4 U6496 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5004) );
  NAND4_X1 U6497 ( .A1(n5128), .A2(n5182), .A3(n4954), .A4(n5204), .ZN(n4955)
         );
  NOR2_X1 U6498 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4958) );
  NOR2_X1 U6499 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4957) );
  NOR2_X1 U6500 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4956) );
  INV_X1 U6501 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U6502 ( .A1(n4965), .A2(n4964), .ZN(n4968) );
  NAND2_X1 U6503 ( .A1(n4976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4967) );
  MUX2_X1 U6504 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4967), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4969) );
  NAND2_X1 U6505 ( .A1(n5035), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4975) );
  AND2_X2 U6506 ( .A1(n7878), .A2(n7884), .ZN(n5015) );
  NAND2_X1 U6507 ( .A1(n5015), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4974) );
  AND2_X2 U6508 ( .A1(n4971), .A2(n4970), .ZN(n5193) );
  NAND2_X1 U6509 ( .A1(n5193), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6510 ( .A1(n5052), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4972) );
  INV_X1 U6511 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4977) );
  XNOR2_X1 U6512 ( .A(n5009), .B(SI_1_), .ZN(n5006) );
  AND2_X1 U6513 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6514 ( .A1(n5145), .A2(n4984), .ZN(n6055) );
  AND2_X1 U6515 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6516 ( .A1(n6070), .A2(n4985), .ZN(n4995) );
  NAND2_X1 U6517 ( .A1(n6055), .A2(n4995), .ZN(n5007) );
  XNOR2_X1 U6518 ( .A(n5006), .B(n5007), .ZN(n6071) );
  OR2_X1 U6519 ( .A1(n4323), .A2(n6071), .ZN(n4988) );
  NAND2_X1 U6520 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4986) );
  OR2_X1 U6521 ( .A1(n4997), .A2(n5992), .ZN(n4987) );
  NAND2_X1 U6522 ( .A1(n6509), .A2(n5783), .ZN(n5578) );
  NAND2_X1 U6523 ( .A1(n4343), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6524 ( .A1(n5193), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6525 ( .A1(n5052), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U6526 ( .A1(n5015), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6527 ( .A1(n6070), .A2(SI_0_), .ZN(n4994) );
  INV_X1 U6528 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6529 ( .A1(n4994), .A2(n4993), .ZN(n4996) );
  AND2_X1 U6530 ( .A1(n4996), .A2(n4995), .ZN(n8569) );
  MUX2_X1 U6531 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8569), .S(n6562), .Z(n6845) );
  NAND2_X1 U6532 ( .A1(n4366), .A2(n6845), .ZN(n7006) );
  NAND2_X1 U6533 ( .A1(n5035), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6534 ( .A1(n5052), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U6535 ( .A1(n5015), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U6536 ( .A1(n5193), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5000) );
  INV_X1 U6537 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6680) );
  INV_X1 U6538 ( .A(n5006), .ZN(n5008) );
  NAND2_X1 U6539 ( .A1(n5008), .A2(n5007), .ZN(n5011) );
  NAND2_X1 U6540 ( .A1(n5009), .A2(SI_1_), .ZN(n5010) );
  NAND2_X1 U6541 ( .A1(n5011), .A2(n5010), .ZN(n5025) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6687) );
  XNOR2_X1 U6543 ( .A(n5025), .B(n5024), .ZN(n6686) );
  OR2_X1 U6544 ( .A1(n4324), .A2(n6686), .ZN(n5013) );
  OAI211_X1 U6545 ( .C1(n6562), .C2(n9800), .A(n5014), .B(n5013), .ZN(n9858)
         );
  NAND2_X1 U6546 ( .A1(n5789), .A2(n9858), .ZN(n5586) );
  INV_X1 U6547 ( .A(n5789), .ZN(n8076) );
  INV_X1 U6548 ( .A(n9858), .ZN(n6953) );
  NAND2_X1 U6549 ( .A1(n8076), .A2(n6953), .ZN(n5585) );
  NAND2_X1 U6550 ( .A1(n7207), .A2(n7206), .ZN(n7205) );
  NAND2_X1 U6551 ( .A1(n7205), .A2(n5586), .ZN(n7224) );
  INV_X1 U6552 ( .A(n5053), .ZN(n5448) );
  NAND2_X1 U6553 ( .A1(n5448), .A2(n7229), .ZN(n5019) );
  NAND2_X1 U6554 ( .A1(n5052), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U6555 ( .A1(n5035), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6556 ( .A1(n5015), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5016) );
  AND4_X2 U6557 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n7210)
         );
  NAND2_X1 U6558 ( .A1(n5005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5020) );
  MUX2_X1 U6559 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5020), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5022) );
  NAND2_X1 U6560 ( .A1(n5022), .A2(n5021), .ZN(n6979) );
  INV_X1 U6561 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6681) );
  OR2_X1 U6562 ( .A1(n5046), .A2(n6681), .ZN(n5032) );
  NAND2_X1 U6563 ( .A1(n5025), .A2(n5024), .ZN(n5029) );
  INV_X1 U6564 ( .A(n5026), .ZN(n5027) );
  NAND2_X1 U6565 ( .A1(n5027), .A2(SI_2_), .ZN(n5028) );
  NAND2_X1 U6566 ( .A1(n5029), .A2(n5028), .ZN(n5041) );
  INV_X1 U6567 ( .A(SI_3_), .ZN(n5030) );
  XNOR2_X1 U6568 ( .A(n5042), .B(n5030), .ZN(n5040) );
  XNOR2_X1 U6569 ( .A(n5041), .B(n5040), .ZN(n6694) );
  OR2_X1 U6570 ( .A1(n4324), .A2(n6694), .ZN(n5031) );
  OAI211_X1 U6571 ( .C1(n6562), .C2(n6979), .A(n5032), .B(n5031), .ZN(n9865)
         );
  INV_X1 U6572 ( .A(n7210), .ZN(n8075) );
  INV_X1 U6573 ( .A(n9865), .ZN(n6513) );
  NAND2_X1 U6574 ( .A1(n8075), .A2(n6513), .ZN(n5599) );
  NAND2_X1 U6575 ( .A1(n5550), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U6576 ( .A1(n5052), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6577 ( .A1(n5033), .A2(n7229), .ZN(n5056) );
  NAND2_X1 U6578 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5034) );
  NAND2_X1 U6579 ( .A1(n5056), .A2(n5034), .ZN(n7270) );
  NAND2_X1 U6580 ( .A1(n5467), .A2(n7270), .ZN(n5037) );
  NAND2_X1 U6581 ( .A1(n5035), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5036) );
  NAND4_X1 U6582 ( .A1(n5039), .A2(n5038), .A3(n5037), .A4(n5036), .ZN(n8074)
         );
  NAND2_X1 U6583 ( .A1(n5041), .A2(n5040), .ZN(n5044) );
  NAND2_X1 U6584 ( .A1(n5042), .A2(SI_3_), .ZN(n5043) );
  NAND2_X1 U6585 ( .A1(n5044), .A2(n5043), .ZN(n5063) );
  MUX2_X1 U6586 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5145), .Z(n5064) );
  INV_X1 U6587 ( .A(SI_4_), .ZN(n5045) );
  XNOR2_X1 U6588 ( .A(n5064), .B(n5045), .ZN(n5062) );
  XNOR2_X1 U6589 ( .A(n5063), .B(n5062), .ZN(n6676) );
  OR2_X1 U6590 ( .A1(n4324), .A2(n6676), .ZN(n5051) );
  INV_X1 U6591 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6677) );
  OR2_X1 U6592 ( .A1(n5046), .A2(n6677), .ZN(n5050) );
  NAND2_X1 U6593 ( .A1(n5021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5048) );
  INV_X1 U6594 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5047) );
  XNOR2_X1 U6595 ( .A(n5048), .B(n5047), .ZN(n7190) );
  OR2_X1 U6596 ( .A1(n6562), .A2(n7190), .ZN(n5049) );
  NAND2_X1 U6597 ( .A1(n8074), .A2(n9872), .ZN(n5593) );
  INV_X1 U6598 ( .A(n9872), .ZN(n7271) );
  NAND2_X1 U6599 ( .A1(n7261), .A2(n7271), .ZN(n5598) );
  NAND2_X1 U6600 ( .A1(n5550), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6601 ( .A1(n5052), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5060) );
  INV_X1 U6602 ( .A(n5056), .ZN(n5055) );
  NAND2_X1 U6603 ( .A1(n5055), .A2(n5054), .ZN(n5075) );
  NAND2_X1 U6604 ( .A1(n5056), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6605 ( .A1(n5075), .A2(n5057), .ZN(n7254) );
  NAND2_X1 U6606 ( .A1(n5448), .A2(n7254), .ZN(n5059) );
  NAND2_X1 U6607 ( .A1(n5035), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5058) );
  NAND4_X1 U6608 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n8072)
         );
  NAND2_X1 U6609 ( .A1(n5063), .A2(n5062), .ZN(n5066) );
  NAND2_X1 U6610 ( .A1(n5064), .A2(SI_4_), .ZN(n5065) );
  NAND2_X1 U6611 ( .A1(n5066), .A2(n5065), .ZN(n5082) );
  MUX2_X1 U6612 ( .A(n6679), .B(n6688), .S(n5145), .Z(n5083) );
  XNOR2_X1 U6613 ( .A(n5083), .B(SI_5_), .ZN(n5081) );
  XNOR2_X1 U6614 ( .A(n5082), .B(n5081), .ZN(n6689) );
  OR2_X1 U6615 ( .A1(n4324), .A2(n6689), .ZN(n5072) );
  OR2_X1 U6616 ( .A1(n5046), .A2(n6679), .ZN(n5071) );
  OR2_X1 U6617 ( .A1(n5067), .A2(n4977), .ZN(n5069) );
  XNOR2_X1 U6618 ( .A(n5069), .B(n5068), .ZN(n6678) );
  OR2_X1 U6619 ( .A1(n6562), .A2(n6678), .ZN(n5070) );
  NAND2_X1 U6620 ( .A1(n8072), .A2(n9876), .ZN(n5601) );
  NAND2_X1 U6621 ( .A1(n7319), .A2(n5601), .ZN(n5073) );
  INV_X1 U6622 ( .A(n8072), .ZN(n7161) );
  INV_X1 U6623 ( .A(n9876), .ZN(n7327) );
  NAND2_X1 U6624 ( .A1(n7161), .A2(n7327), .ZN(n5602) );
  NAND2_X1 U6625 ( .A1(n5550), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6626 ( .A1(n5052), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6627 ( .A1(n5075), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6628 ( .A1(n5094), .A2(n5076), .ZN(n8028) );
  NAND2_X1 U6629 ( .A1(n5448), .A2(n8028), .ZN(n5078) );
  NAND2_X1 U6630 ( .A1(n5035), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5077) );
  NAND4_X1 U6631 ( .A1(n5080), .A2(n5079), .A3(n5078), .A4(n5077), .ZN(n8071)
         );
  NAND2_X1 U6632 ( .A1(n5082), .A2(n5081), .ZN(n5086) );
  INV_X1 U6633 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6634 ( .A1(n5084), .A2(SI_5_), .ZN(n5085) );
  XNOR2_X1 U6635 ( .A(n5105), .B(SI_6_), .ZN(n5103) );
  XNOR2_X1 U6636 ( .A(n5104), .B(n5103), .ZN(n6684) );
  OR2_X1 U6637 ( .A1(n4324), .A2(n6684), .ZN(n5091) );
  OR2_X1 U6638 ( .A1(n5046), .A2(n6682), .ZN(n5090) );
  OR2_X1 U6639 ( .A1(n5087), .A2(n4977), .ZN(n5088) );
  XNOR2_X1 U6640 ( .A(n5088), .B(P2_IR_REG_6__SCAN_IN), .ZN(n5998) );
  OR2_X1 U6641 ( .A1(n6562), .A2(n7402), .ZN(n5089) );
  NOR2_X1 U6642 ( .A1(n8071), .A2(n7461), .ZN(n5605) );
  NAND2_X1 U6643 ( .A1(n8071), .A2(n7461), .ZN(n5732) );
  OAI21_X1 U6644 ( .B1(n7437), .B2(n5605), .A(n5732), .ZN(n7416) );
  NAND2_X1 U6645 ( .A1(n5550), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6646 ( .A1(n5052), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5098) );
  INV_X1 U6647 ( .A(n5094), .ZN(n5093) );
  NAND2_X1 U6648 ( .A1(n5093), .A2(n5092), .ZN(n5111) );
  NAND2_X1 U6649 ( .A1(n5094), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6650 ( .A1(n5111), .A2(n5095), .ZN(n7422) );
  NAND2_X1 U6651 ( .A1(n5448), .A2(n7422), .ZN(n5097) );
  NAND2_X1 U6652 ( .A1(n5035), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6653 ( .A1(n5100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5101) );
  MUX2_X1 U6654 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5101), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5102) );
  OR2_X1 U6655 ( .A1(n5100), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5151) );
  AND2_X1 U6656 ( .A1(n5102), .A2(n5151), .ZN(n9825) );
  NAND2_X1 U6657 ( .A1(n5104), .A2(n5103), .ZN(n5108) );
  INV_X1 U6658 ( .A(n5105), .ZN(n5106) );
  NAND2_X1 U6659 ( .A1(n5106), .A2(SI_6_), .ZN(n5107) );
  MUX2_X1 U6660 ( .A(n6699), .B(n6696), .S(n5145), .Z(n5119) );
  XNOR2_X1 U6661 ( .A(n5119), .B(SI_7_), .ZN(n5117) );
  OR2_X1 U6662 ( .A1(n4324), .A2(n6698), .ZN(n5110) );
  OR2_X1 U6663 ( .A1(n5046), .A2(n6699), .ZN(n5109) );
  OAI211_X1 U6664 ( .C1(n6562), .C2(n6697), .A(n5110), .B(n5109), .ZN(n7434)
         );
  NAND2_X1 U6665 ( .A1(n8026), .A2(n7434), .ZN(n5612) );
  INV_X1 U6666 ( .A(n8026), .ZN(n8070) );
  INV_X1 U6667 ( .A(n7434), .ZN(n9882) );
  NAND2_X1 U6668 ( .A1(n8070), .A2(n9882), .ZN(n5615) );
  NAND2_X1 U6669 ( .A1(n5550), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6670 ( .A1(n5052), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6671 ( .A1(n5111), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6672 ( .A1(n5136), .A2(n5112), .ZN(n7544) );
  NAND2_X1 U6673 ( .A1(n5467), .A2(n7544), .ZN(n5114) );
  NAND2_X1 U6674 ( .A1(n5035), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5113) );
  NAND4_X1 U6675 ( .A1(n5116), .A2(n5115), .A3(n5114), .A4(n5113), .ZN(n8069)
         );
  INV_X1 U6676 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6677 ( .A1(n5120), .A2(SI_7_), .ZN(n5121) );
  INV_X1 U6678 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5122) );
  MUX2_X1 U6679 ( .A(n6703), .B(n5122), .S(n5145), .Z(n5124) );
  INV_X1 U6680 ( .A(SI_8_), .ZN(n5123) );
  NAND2_X1 U6681 ( .A1(n5124), .A2(n5123), .ZN(n5144) );
  INV_X1 U6682 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6683 ( .A1(n5125), .A2(SI_8_), .ZN(n5126) );
  NAND2_X1 U6684 ( .A1(n5144), .A2(n5126), .ZN(n5143) );
  INV_X1 U6685 ( .A(n5143), .ZN(n5127) );
  XNOR2_X1 U6686 ( .A(n5142), .B(n5127), .ZN(n6702) );
  OR2_X1 U6687 ( .A1(n6702), .A2(n4324), .ZN(n5132) );
  OR2_X1 U6688 ( .A1(n5046), .A2(n6703), .ZN(n5131) );
  NAND2_X1 U6689 ( .A1(n5151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5129) );
  XNOR2_X1 U6690 ( .A(n5129), .B(n5128), .ZN(n6701) );
  OR2_X1 U6691 ( .A1(n6562), .A2(n6701), .ZN(n5130) );
  AND2_X1 U6692 ( .A1(n8069), .A2(n9889), .ZN(n5609) );
  INV_X1 U6693 ( .A(n9889), .ZN(n7478) );
  NAND2_X1 U6694 ( .A1(n7629), .A2(n7478), .ZN(n5729) );
  NAND2_X1 U6695 ( .A1(n5133), .A2(n5729), .ZN(n7625) );
  NAND2_X1 U6696 ( .A1(n5550), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6697 ( .A1(n5052), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6698 ( .A1(n5136), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6699 ( .A1(n5165), .A2(n5137), .ZN(n7631) );
  NAND2_X1 U6700 ( .A1(n5448), .A2(n7631), .ZN(n5139) );
  NAND2_X1 U6701 ( .A1(n5035), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5138) );
  INV_X1 U6702 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5146) );
  MUX2_X1 U6703 ( .A(n6706), .B(n5146), .S(n5145), .Z(n5148) );
  INV_X1 U6704 ( .A(SI_9_), .ZN(n5147) );
  NAND2_X1 U6705 ( .A1(n5148), .A2(n5147), .ZN(n5159) );
  INV_X1 U6706 ( .A(n5148), .ZN(n5149) );
  NAND2_X1 U6707 ( .A1(n5149), .A2(SI_9_), .ZN(n5150) );
  XNOR2_X1 U6708 ( .A(n5158), .B(n4945), .ZN(n6704) );
  NAND2_X1 U6709 ( .A1(n6704), .A2(n5547), .ZN(n5156) );
  NAND2_X1 U6710 ( .A1(n5185), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5153) );
  INV_X1 U6711 ( .A(n5153), .ZN(n5152) );
  NAND2_X1 U6712 ( .A1(n5152), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6713 ( .A1(n5153), .A2(n5183), .ZN(n5161) );
  AOI22_X1 U6714 ( .A1(n5335), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5334), .B2(
        n5988), .ZN(n5155) );
  NAND2_X1 U6715 ( .A1(n5156), .A2(n5155), .ZN(n7762) );
  NAND2_X1 U6716 ( .A1(n7599), .A2(n7762), .ZN(n5613) );
  INV_X1 U6717 ( .A(n7762), .ZN(n9894) );
  NAND2_X1 U6718 ( .A1(n8068), .A2(n9894), .ZN(n5616) );
  NAND2_X1 U6719 ( .A1(n5613), .A2(n5616), .ZN(n7626) );
  MUX2_X1 U6720 ( .A(n6712), .B(n10120), .S(n4325), .Z(n5174) );
  XNOR2_X1 U6721 ( .A(n5174), .B(SI_10_), .ZN(n5171) );
  XNOR2_X1 U6722 ( .A(n5173), .B(n5171), .ZN(n6711) );
  NAND2_X1 U6723 ( .A1(n6711), .A2(n5547), .ZN(n5164) );
  NAND2_X1 U6724 ( .A1(n5161), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5162) );
  XNOR2_X1 U6725 ( .A(n5162), .B(P2_IR_REG_10__SCAN_IN), .ZN(n5986) );
  AOI22_X1 U6726 ( .A1(n5335), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5334), .B2(
        n5986), .ZN(n5163) );
  NAND2_X1 U6727 ( .A1(n5550), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6728 ( .A1(n5052), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6729 ( .A1(n5165), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6730 ( .A1(n5194), .A2(n5166), .ZN(n7774) );
  NAND2_X1 U6731 ( .A1(n5467), .A2(n7774), .ZN(n5168) );
  NAND2_X1 U6732 ( .A1(n5035), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6733 ( .A1(n7630), .A2(n9905), .ZN(n5624) );
  INV_X1 U6734 ( .A(n5171), .ZN(n5172) );
  INV_X1 U6735 ( .A(n5174), .ZN(n5175) );
  NAND2_X1 U6736 ( .A1(n5175), .A2(SI_10_), .ZN(n5176) );
  INV_X1 U6737 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5177) );
  MUX2_X1 U6738 ( .A(n6728), .B(n5177), .S(n4325), .Z(n5179) );
  INV_X1 U6739 ( .A(SI_11_), .ZN(n5178) );
  NAND2_X1 U6740 ( .A1(n5179), .A2(n5178), .ZN(n5201) );
  INV_X1 U6741 ( .A(n5179), .ZN(n5180) );
  NAND2_X1 U6742 ( .A1(n5180), .A2(SI_11_), .ZN(n5181) );
  NAND2_X1 U6743 ( .A1(n5201), .A2(n5181), .ZN(n5202) );
  XNOR2_X1 U6744 ( .A(n5203), .B(n5202), .ZN(n6721) );
  NAND2_X1 U6745 ( .A1(n6721), .A2(n5547), .ZN(n5192) );
  NAND2_X1 U6746 ( .A1(n5183), .A2(n5182), .ZN(n5184) );
  INV_X1 U6747 ( .A(n5189), .ZN(n5186) );
  NAND2_X1 U6748 ( .A1(n5186), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5187) );
  MUX2_X1 U6749 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5187), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5190) );
  NAND2_X1 U6750 ( .A1(n5189), .A2(n5188), .ZN(n5220) );
  AOI22_X1 U6751 ( .A1(n5335), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5334), .B2(
        n5984), .ZN(n5191) );
  NAND2_X1 U6752 ( .A1(n5192), .A2(n5191), .ZN(n9908) );
  NAND2_X1 U6753 ( .A1(n5052), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6754 ( .A1(n5035), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6755 ( .A1(n5194), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6756 ( .A1(n5209), .A2(n5195), .ZN(n8005) );
  NAND2_X1 U6757 ( .A1(n5448), .A2(n8005), .ZN(n5197) );
  NAND2_X1 U6758 ( .A1(n5550), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5196) );
  OR2_X1 U6759 ( .A1(n9908), .A2(n8388), .ZN(n5627) );
  NAND2_X1 U6760 ( .A1(n9908), .A2(n8388), .ZN(n5628) );
  NAND2_X1 U6761 ( .A1(n7661), .A2(n7662), .ZN(n5200) );
  NAND2_X1 U6762 ( .A1(n5200), .A2(n5628), .ZN(n8399) );
  MUX2_X1 U6763 ( .A(n10105), .B(n6803), .S(n4325), .Z(n5216) );
  XNOR2_X1 U6764 ( .A(n5216), .B(SI_12_), .ZN(n5215) );
  XNOR2_X1 U6765 ( .A(n5219), .B(n5215), .ZN(n6763) );
  NAND2_X1 U6766 ( .A1(n6763), .A2(n5547), .ZN(n5207) );
  NAND2_X1 U6767 ( .A1(n5220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  XNOR2_X1 U6768 ( .A(n5205), .B(n5204), .ZN(n6764) );
  INV_X1 U6769 ( .A(n6764), .ZN(n7823) );
  AOI22_X1 U6770 ( .A1(n5335), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5334), .B2(
        n7823), .ZN(n5206) );
  NAND2_X1 U6771 ( .A1(n5052), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6772 ( .A1(n5035), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6773 ( .A1(n5209), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6774 ( .A1(n5226), .A2(n5210), .ZN(n8395) );
  NAND2_X1 U6775 ( .A1(n5193), .A2(n8395), .ZN(n5212) );
  NAND2_X1 U6776 ( .A1(n5550), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5211) );
  XNOR2_X1 U6777 ( .A(n9913), .B(n8003), .ZN(n8400) );
  OR2_X1 U6778 ( .A1(n9913), .A2(n8003), .ZN(n5632) );
  INV_X1 U6779 ( .A(n5216), .ZN(n5217) );
  MUX2_X1 U6780 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4325), .Z(n5235) );
  XNOR2_X1 U6781 ( .A(n5235), .B(SI_13_), .ZN(n5233) );
  XNOR2_X1 U6782 ( .A(n5234), .B(n5233), .ZN(n6805) );
  NAND2_X1 U6783 ( .A1(n6805), .A2(n5547), .ZN(n5223) );
  NAND2_X1 U6784 ( .A1(n5221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5238) );
  XNOR2_X1 U6785 ( .A(n5238), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U6786 ( .A1(n5335), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5334), .B2(
        n9836), .ZN(n5222) );
  NAND2_X1 U6787 ( .A1(n5550), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6788 ( .A1(n5052), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5230) );
  INV_X1 U6789 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6790 ( .A1(n5226), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6791 ( .A1(n5242), .A2(n5227), .ZN(n8380) );
  NAND2_X1 U6792 ( .A1(n5193), .A2(n8380), .ZN(n5229) );
  NAND2_X1 U6793 ( .A1(n5035), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6794 ( .A1(n8549), .A2(n8390), .ZN(n5640) );
  NAND2_X1 U6795 ( .A1(n5232), .A2(n5641), .ZN(n8356) );
  MUX2_X1 U6796 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4325), .Z(n5249) );
  XNOR2_X1 U6797 ( .A(n5249), .B(SI_14_), .ZN(n5236) );
  XNOR2_X1 U6798 ( .A(n5248), .B(n5236), .ZN(n6850) );
  NAND2_X1 U6799 ( .A1(n6850), .A2(n5547), .ZN(n5241) );
  NAND2_X1 U6800 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  NAND2_X1 U6801 ( .A1(n5239), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5257) );
  INV_X1 U6802 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5256) );
  INV_X1 U6803 ( .A(n8085), .ZN(n5980) );
  AOI22_X1 U6804 ( .A1(n5335), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5334), .B2(
        n5980), .ZN(n5240) );
  NAND2_X1 U6805 ( .A1(n5241), .A2(n5240), .ZN(n8368) );
  NAND2_X1 U6806 ( .A1(n5052), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6807 ( .A1(n5550), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6808 ( .A1(n5242), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6809 ( .A1(n5264), .A2(n5243), .ZN(n8367) );
  NAND2_X1 U6810 ( .A1(n5193), .A2(n8367), .ZN(n5245) );
  NAND2_X1 U6811 ( .A1(n5035), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5244) );
  NOR2_X1 U6812 ( .A1(n8368), .A2(n8050), .ZN(n5637) );
  NAND2_X1 U6813 ( .A1(n8368), .A2(n8050), .ZN(n5647) );
  INV_X1 U6814 ( .A(n5248), .ZN(n5250) );
  NAND2_X1 U6815 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  MUX2_X1 U6816 ( .A(n6909), .B(n6922), .S(n4325), .Z(n5270) );
  XNOR2_X1 U6817 ( .A(n5270), .B(SI_15_), .ZN(n5255) );
  NAND2_X1 U6818 ( .A1(n6908), .A2(n5547), .ZN(n5261) );
  NAND2_X1 U6819 ( .A1(n5257), .A2(n5256), .ZN(n5258) );
  NAND2_X1 U6820 ( .A1(n5258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5259) );
  XNOR2_X1 U6821 ( .A(n5259), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8100) );
  AOI22_X1 U6822 ( .A1(n5335), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5334), .B2(
        n8100), .ZN(n5260) );
  NAND2_X1 U6823 ( .A1(n5261), .A2(n5260), .ZN(n8538) );
  NAND2_X1 U6824 ( .A1(n5550), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6825 ( .A1(n5052), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6826 ( .A1(n5264), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6827 ( .A1(n5280), .A2(n5265), .ZN(n8353) );
  NAND2_X1 U6828 ( .A1(n5467), .A2(n8353), .ZN(n5267) );
  NAND2_X1 U6829 ( .A1(n5035), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5266) );
  AND2_X1 U6830 ( .A1(n8538), .A2(n8362), .ZN(n5645) );
  OR2_X1 U6831 ( .A1(n8538), .A2(n8362), .ZN(n5650) );
  NOR2_X1 U6832 ( .A1(n5273), .A2(SI_15_), .ZN(n5271) );
  NAND2_X1 U6833 ( .A1(n5273), .A2(SI_15_), .ZN(n5274) );
  MUX2_X1 U6834 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4325), .Z(n5286) );
  XNOR2_X1 U6835 ( .A(n5286), .B(SI_16_), .ZN(n5275) );
  XNOR2_X1 U6836 ( .A(n5291), .B(n5275), .ZN(n7002) );
  NAND2_X1 U6837 ( .A1(n7002), .A2(n5547), .ZN(n5279) );
  NAND2_X1 U6838 ( .A1(n5276), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5277) );
  XNOR2_X1 U6839 ( .A(n5277), .B(P2_IR_REG_16__SCAN_IN), .ZN(n5977) );
  AOI22_X1 U6840 ( .A1(n5335), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5334), .B2(
        n5977), .ZN(n5278) );
  NAND2_X1 U6841 ( .A1(n5052), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6842 ( .A1(n5550), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6843 ( .A1(n5280), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6844 ( .A1(n5338), .A2(n5281), .ZN(n8343) );
  NAND2_X1 U6845 ( .A1(n5193), .A2(n8343), .ZN(n5283) );
  NAND2_X1 U6846 ( .A1(n5035), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6847 ( .A1(n8533), .A2(n8326), .ZN(n8286) );
  NOR2_X1 U6848 ( .A1(n5288), .A2(n5287), .ZN(n5290) );
  NAND2_X1 U6849 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  MUX2_X1 U6850 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4325), .Z(n5292) );
  XNOR2_X1 U6851 ( .A(n5292), .B(n10129), .ZN(n5330) );
  INV_X1 U6852 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6853 ( .A1(n5293), .A2(n10129), .ZN(n5294) );
  MUX2_X1 U6854 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4325), .Z(n5296) );
  NAND2_X1 U6855 ( .A1(n5296), .A2(SI_18_), .ZN(n5300) );
  INV_X1 U6856 ( .A(n5296), .ZN(n5298) );
  INV_X1 U6857 ( .A(SI_18_), .ZN(n5297) );
  NAND2_X1 U6858 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6859 ( .A1(n5300), .A2(n5299), .ZN(n5317) );
  MUX2_X1 U6860 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4325), .Z(n5347) );
  XNOR2_X1 U6861 ( .A(n5347), .B(SI_19_), .ZN(n5351) );
  XNOR2_X1 U6862 ( .A(n5352), .B(n5351), .ZN(n7252) );
  NAND2_X1 U6863 ( .A1(n7252), .A2(n5547), .ZN(n5307) );
  NAND2_X1 U6864 ( .A1(n5301), .A2(n5302), .ZN(n5559) );
  NAND2_X1 U6865 ( .A1(n5559), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5320) );
  INV_X1 U6866 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6867 ( .A1(n5320), .A2(n5303), .ZN(n5304) );
  AOI22_X1 U6868 ( .A1(n5335), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6556), .B2(
        n5334), .ZN(n5306) );
  NAND2_X1 U6869 ( .A1(n5052), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6870 ( .A1(n5550), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5315) );
  INV_X1 U6871 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5308) );
  INV_X1 U6872 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6873 ( .A1(n5325), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6874 ( .A1(n5355), .A2(n5312), .ZN(n8302) );
  NAND2_X1 U6875 ( .A1(n5193), .A2(n8302), .ZN(n5314) );
  NAND2_X1 U6876 ( .A1(n5035), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6877 ( .A1(n8518), .A2(n8278), .ZN(n5726) );
  OR2_X1 U6878 ( .A1(n8518), .A2(n8278), .ZN(n5727) );
  INV_X1 U6879 ( .A(n5317), .ZN(n5318) );
  XNOR2_X1 U6880 ( .A(n5319), .B(n5318), .ZN(n7064) );
  NAND2_X1 U6881 ( .A1(n7064), .A2(n5547), .ZN(n5322) );
  XNOR2_X1 U6882 ( .A(n5320), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8150) );
  AOI22_X1 U6883 ( .A1(n5335), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5334), .B2(
        n8150), .ZN(n5321) );
  NAND2_X1 U6884 ( .A1(n5052), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6885 ( .A1(n5035), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6886 ( .A1(n5323), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6887 ( .A1(n5325), .A2(n5324), .ZN(n8314) );
  NAND2_X1 U6888 ( .A1(n5448), .A2(n8314), .ZN(n5327) );
  NAND2_X1 U6889 ( .A1(n5550), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5326) );
  AND2_X1 U6890 ( .A1(n5727), .A2(n8289), .ZN(n5663) );
  INV_X1 U6891 ( .A(n5663), .ZN(n5344) );
  NAND2_X1 U6892 ( .A1(n8522), .A2(n8325), .ZN(n5668) );
  INV_X1 U6893 ( .A(n8309), .ZN(n5343) );
  XNOR2_X1 U6894 ( .A(n5331), .B(n5330), .ZN(n7060) );
  NAND2_X1 U6895 ( .A1(n7060), .A2(n5547), .ZN(n5337) );
  INV_X1 U6896 ( .A(n5301), .ZN(n5332) );
  NAND2_X1 U6897 ( .A1(n5332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5333) );
  XNOR2_X1 U6898 ( .A(n5333), .B(P2_IR_REG_17__SCAN_IN), .ZN(n5976) );
  AOI22_X1 U6899 ( .A1(n5335), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5334), .B2(
        n5976), .ZN(n5336) );
  NAND2_X1 U6900 ( .A1(n5337), .A2(n5336), .ZN(n7955) );
  NAND2_X1 U6901 ( .A1(n5550), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6902 ( .A1(n5052), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5341) );
  XNOR2_X1 U6903 ( .A(n5338), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U6904 ( .A1(n5193), .A2(n8327), .ZN(n5340) );
  NAND2_X1 U6905 ( .A1(n5035), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6906 ( .A1(n7955), .A2(n8340), .ZN(n8305) );
  AND2_X1 U6907 ( .A1(n5343), .A2(n8305), .ZN(n8288) );
  OR2_X1 U6908 ( .A1(n5344), .A2(n8288), .ZN(n5345) );
  AND2_X1 U6909 ( .A1(n5726), .A2(n5345), .ZN(n5361) );
  AND2_X1 U6910 ( .A1(n8286), .A2(n5361), .ZN(n5346) );
  NAND2_X1 U6911 ( .A1(n8285), .A2(n5346), .ZN(n8271) );
  INV_X1 U6912 ( .A(n5347), .ZN(n5349) );
  INV_X1 U6913 ( .A(SI_19_), .ZN(n5348) );
  NAND2_X1 U6914 ( .A1(n5349), .A2(n5348), .ZN(n5350) );
  MUX2_X1 U6915 ( .A(n7389), .B(n6312), .S(n4325), .Z(n5368) );
  XNOR2_X1 U6916 ( .A(n5368), .B(SI_20_), .ZN(n5365) );
  XNOR2_X1 U6917 ( .A(n5366), .B(n5365), .ZN(n7367) );
  NAND2_X1 U6918 ( .A1(n7367), .A2(n5547), .ZN(n5354) );
  OR2_X1 U6919 ( .A1(n5046), .A2(n7389), .ZN(n5353) );
  NAND2_X1 U6920 ( .A1(n5550), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6921 ( .A1(n5052), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5359) );
  OR2_X2 U6922 ( .A1(n5355), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6923 ( .A1(n5355), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6924 ( .A1(n5376), .A2(n5356), .ZN(n8282) );
  NAND2_X1 U6925 ( .A1(n5467), .A2(n8282), .ZN(n5358) );
  NAND2_X1 U6926 ( .A1(n5035), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5357) );
  OR2_X1 U6927 ( .A1(n8513), .A2(n8297), .ZN(n5670) );
  INV_X1 U6928 ( .A(n5361), .ZN(n5363) );
  AND2_X1 U6929 ( .A1(n8318), .A2(n4937), .ZN(n8287) );
  AND2_X1 U6930 ( .A1(n8287), .A2(n5663), .ZN(n5362) );
  AND2_X1 U6931 ( .A1(n5670), .A2(n8270), .ZN(n5364) );
  NAND2_X1 U6932 ( .A1(n8271), .A2(n5364), .ZN(n8256) );
  NAND2_X1 U6933 ( .A1(n5366), .A2(n5365), .ZN(n5370) );
  INV_X1 U6934 ( .A(SI_20_), .ZN(n5367) );
  NAND2_X1 U6935 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  MUX2_X1 U6936 ( .A(n7484), .B(n7832), .S(n4325), .Z(n5385) );
  XNOR2_X1 U6937 ( .A(n5385), .B(SI_21_), .ZN(n5371) );
  XNOR2_X1 U6938 ( .A(n5383), .B(n5371), .ZN(n7483) );
  NAND2_X1 U6939 ( .A1(n7483), .A2(n5547), .ZN(n5373) );
  OR2_X1 U6940 ( .A1(n5046), .A2(n7484), .ZN(n5372) );
  INV_X1 U6941 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6942 ( .A1(n5376), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6943 ( .A1(n5394), .A2(n5377), .ZN(n8265) );
  NAND2_X1 U6944 ( .A1(n8265), .A2(n5193), .ZN(n5381) );
  NAND2_X1 U6945 ( .A1(n5052), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6946 ( .A1(n5550), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6947 ( .A1(n5035), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6948 ( .A1(n8437), .A2(n8279), .ZN(n5724) );
  NAND2_X1 U6949 ( .A1(n8513), .A2(n8297), .ZN(n8255) );
  AND2_X1 U6950 ( .A1(n5724), .A2(n8255), .ZN(n5673) );
  NAND2_X1 U6951 ( .A1(n8256), .A2(n5673), .ZN(n5382) );
  NAND2_X1 U6952 ( .A1(n5382), .A2(n5725), .ZN(n8238) );
  INV_X1 U6953 ( .A(SI_21_), .ZN(n5384) );
  INV_X1 U6954 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U6955 ( .A1(n5386), .A2(SI_21_), .ZN(n5387) );
  MUX2_X1 U6956 ( .A(n7522), .B(n10146), .S(n4325), .Z(n5389) );
  INV_X1 U6957 ( .A(SI_22_), .ZN(n5388) );
  NAND2_X1 U6958 ( .A1(n5389), .A2(n5388), .ZN(n5401) );
  INV_X1 U6959 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6960 ( .A1(n5390), .A2(SI_22_), .ZN(n5391) );
  NAND2_X1 U6961 ( .A1(n5401), .A2(n5391), .ZN(n5399) );
  XNOR2_X1 U6962 ( .A(n5400), .B(n5399), .ZN(n7520) );
  NAND2_X1 U6963 ( .A1(n7520), .A2(n5547), .ZN(n5393) );
  OR2_X1 U6964 ( .A1(n5046), .A2(n7522), .ZN(n5392) );
  OR2_X2 U6965 ( .A1(n5394), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6966 ( .A1(n5394), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6967 ( .A1(n5412), .A2(n5395), .ZN(n8251) );
  NAND2_X1 U6968 ( .A1(n8251), .A2(n5193), .ZN(n5398) );
  AOI22_X1 U6969 ( .A1(n5550), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n5052), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6970 ( .A1(n5035), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6971 ( .A1(n8252), .A2(n8264), .ZN(n5681) );
  INV_X1 U6972 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7562) );
  INV_X1 U6973 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7559) );
  MUX2_X1 U6974 ( .A(n7562), .B(n7559), .S(n4325), .Z(n5404) );
  INV_X1 U6975 ( .A(SI_23_), .ZN(n5403) );
  NAND2_X1 U6976 ( .A1(n5404), .A2(n5403), .ZN(n5417) );
  INV_X1 U6977 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U6978 ( .A1(n5405), .A2(SI_23_), .ZN(n5406) );
  OR2_X1 U6979 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  NAND2_X1 U6980 ( .A1(n5418), .A2(n5409), .ZN(n6339) );
  NAND2_X1 U6981 ( .A1(n6339), .A2(n5547), .ZN(n5411) );
  OR2_X1 U6982 ( .A1(n5046), .A2(n7562), .ZN(n5410) );
  INV_X1 U6983 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U6984 ( .A1(n5412), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6985 ( .A1(n8226), .A2(n5467), .ZN(n5415) );
  AOI22_X1 U6986 ( .A1(n5550), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n5052), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5414) );
  OAI211_X2 U6987 ( .C1(n5553), .C2(n8431), .A(n5415), .B(n5414), .ZN(n8216)
         );
  INV_X1 U6988 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7644) );
  INV_X1 U6989 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7646) );
  MUX2_X1 U6990 ( .A(n7644), .B(n7646), .S(n4325), .Z(n5420) );
  INV_X1 U6991 ( .A(SI_24_), .ZN(n5419) );
  NAND2_X1 U6992 ( .A1(n5420), .A2(n5419), .ZN(n5437) );
  INV_X1 U6993 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6994 ( .A1(n5421), .A2(SI_24_), .ZN(n5422) );
  XNOR2_X1 U6995 ( .A(n5436), .B(n5435), .ZN(n7643) );
  NAND2_X1 U6996 ( .A1(n7643), .A2(n5547), .ZN(n5424) );
  OR2_X1 U6997 ( .A1(n5046), .A2(n7644), .ZN(n5423) );
  INV_X1 U6998 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6999 ( .A1(n5427), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U7000 ( .A1(n5446), .A2(n5428), .ZN(n8218) );
  NAND2_X1 U7001 ( .A1(n8218), .A2(n5193), .ZN(n5433) );
  INV_X1 U7002 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U7003 ( .A1(n5550), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7004 ( .A1(n5052), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5429) );
  OAI211_X1 U7005 ( .C1(n8428), .C2(n5553), .A(n5430), .B(n5429), .ZN(n5431)
         );
  INV_X1 U7006 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U7007 ( .A1(n8220), .A2(n7938), .ZN(n5685) );
  AND2_X1 U7008 ( .A1(n5685), .A2(n8210), .ZN(n5687) );
  NAND2_X1 U7009 ( .A1(n8211), .A2(n5687), .ZN(n5434) );
  NAND2_X1 U7010 ( .A1(n5434), .A2(n5688), .ZN(n8199) );
  NAND2_X1 U7011 ( .A1(n5438), .A2(n5437), .ZN(n5456) );
  INV_X1 U7012 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7701) );
  MUX2_X1 U7013 ( .A(n10114), .B(n7701), .S(n4325), .Z(n5440) );
  INV_X1 U7014 ( .A(SI_25_), .ZN(n5439) );
  NAND2_X1 U7015 ( .A1(n5440), .A2(n5439), .ZN(n5457) );
  INV_X1 U7016 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U7017 ( .A1(n5441), .A2(SI_25_), .ZN(n5442) );
  XNOR2_X1 U7018 ( .A(n5456), .B(n5455), .ZN(n7699) );
  NAND2_X1 U7019 ( .A1(n7699), .A2(n5547), .ZN(n5444) );
  OR2_X1 U7020 ( .A1(n5046), .A2(n10114), .ZN(n5443) );
  INV_X1 U7021 ( .A(n5446), .ZN(n5445) );
  INV_X1 U7022 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U7023 ( .A1(n5446), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7024 ( .A1(n5465), .A2(n5447), .ZN(n8205) );
  NAND2_X1 U7025 ( .A1(n8205), .A2(n5448), .ZN(n5453) );
  INV_X1 U7026 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U7027 ( .A1(n5550), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U7028 ( .A1(n5052), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U7029 ( .C1(n8425), .C2(n5553), .A(n5450), .B(n5449), .ZN(n5451)
         );
  INV_X1 U7030 ( .A(n5451), .ZN(n5452) );
  NAND2_X1 U7031 ( .A1(n8206), .A2(n7965), .ZN(n5697) );
  NAND2_X1 U7032 ( .A1(n8199), .A2(n5697), .ZN(n5454) );
  OR2_X1 U7033 ( .A1(n8206), .A2(n7965), .ZN(n5696) );
  NAND2_X1 U7034 ( .A1(n5454), .A2(n5696), .ZN(n8187) );
  NAND2_X1 U7035 ( .A1(n5456), .A2(n5455), .ZN(n5458) );
  INV_X1 U7036 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U7037 ( .A(n8566), .B(n9624), .S(n4325), .Z(n5460) );
  INV_X1 U7038 ( .A(SI_26_), .ZN(n5459) );
  NAND2_X1 U7039 ( .A1(n5460), .A2(n5459), .ZN(n5477) );
  INV_X1 U7040 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U7041 ( .A1(n5461), .A2(SI_26_), .ZN(n5462) );
  NAND2_X1 U7042 ( .A1(n8564), .A2(n5547), .ZN(n5464) );
  OR2_X1 U7043 ( .A1(n5046), .A2(n8566), .ZN(n5463) );
  OR2_X2 U7044 ( .A1(n5465), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U7045 ( .A1(n5465), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7046 ( .A1(n5486), .A2(n5466), .ZN(n8194) );
  NAND2_X1 U7047 ( .A1(n8194), .A2(n5467), .ZN(n5473) );
  INV_X1 U7048 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U7049 ( .A1(n5052), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7050 ( .A1(n5035), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5468) );
  OAI211_X1 U7051 ( .C1(n5470), .C2(n8479), .A(n5469), .B(n5468), .ZN(n5471)
         );
  INV_X1 U7052 ( .A(n5471), .ZN(n5472) );
  NAND2_X1 U7053 ( .A1(n8195), .A2(n8036), .ZN(n5702) );
  NAND2_X1 U7054 ( .A1(n8187), .A2(n5702), .ZN(n5474) );
  INV_X1 U7055 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7876) );
  INV_X1 U7056 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9621) );
  MUX2_X1 U7057 ( .A(n7876), .B(n9621), .S(n4325), .Z(n5479) );
  INV_X1 U7058 ( .A(SI_27_), .ZN(n5478) );
  NAND2_X1 U7059 ( .A1(n5479), .A2(n5478), .ZN(n5495) );
  INV_X1 U7060 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U7061 ( .A1(n5480), .A2(SI_27_), .ZN(n5481) );
  NAND2_X1 U7062 ( .A1(n7875), .A2(n5547), .ZN(n5483) );
  OR2_X1 U7063 ( .A1(n5046), .A2(n7876), .ZN(n5482) );
  INV_X1 U7064 ( .A(n5486), .ZN(n5485) );
  INV_X1 U7065 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7066 ( .A1(n5485), .A2(n5484), .ZN(n5499) );
  NAND2_X1 U7067 ( .A1(n5486), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7068 ( .A1(n8182), .A2(n5193), .ZN(n5492) );
  INV_X1 U7069 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U7070 ( .A1(n5550), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7071 ( .A1(n5052), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5488) );
  OAI211_X1 U7072 ( .C1(n8419), .C2(n5553), .A(n5489), .B(n5488), .ZN(n5490)
         );
  INV_X1 U7073 ( .A(n5490), .ZN(n5491) );
  NAND2_X1 U7074 ( .A1(n8183), .A2(n7868), .ZN(n5700) );
  INV_X1 U7075 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5496) );
  INV_X1 U7076 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9618) );
  MUX2_X1 U7077 ( .A(n5496), .B(n9618), .S(n4325), .Z(n5511) );
  XNOR2_X1 U7078 ( .A(n5511), .B(SI_28_), .ZN(n5508) );
  NAND2_X1 U7079 ( .A1(n6391), .A2(n5547), .ZN(n5498) );
  OR2_X1 U7080 ( .A1(n5046), .A2(n5496), .ZN(n5497) );
  NAND2_X1 U7081 ( .A1(n5499), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7082 ( .A1(n7865), .A2(n5467), .ZN(n5506) );
  INV_X1 U7083 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7084 ( .A1(n5550), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7085 ( .A1(n5052), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5501) );
  OAI211_X1 U7086 ( .C1(n5503), .C2(n5553), .A(n5502), .B(n5501), .ZN(n5504)
         );
  INV_X1 U7087 ( .A(n5504), .ZN(n5505) );
  NAND2_X2 U7088 ( .A1(n5506), .A2(n5505), .ZN(n8179) );
  NAND2_X1 U7089 ( .A1(n7854), .A2(n7862), .ZN(n7853) );
  INV_X1 U7090 ( .A(n8179), .ZN(n6549) );
  NAND2_X1 U7091 ( .A1(n7872), .A2(n6549), .ZN(n5507) );
  INV_X1 U7092 ( .A(SI_28_), .ZN(n5510) );
  NAND2_X1 U7093 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  MUX2_X1 U7094 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4325), .Z(n5525) );
  INV_X1 U7095 ( .A(SI_29_), .ZN(n5514) );
  NAND2_X1 U7096 ( .A1(n7882), .A2(n5547), .ZN(n5516) );
  INV_X1 U7097 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7883) );
  OR2_X1 U7098 ( .A1(n5046), .A2(n7883), .ZN(n5515) );
  INV_X1 U7099 ( .A(n8164), .ZN(n5517) );
  NAND2_X1 U7100 ( .A1(n5517), .A2(n5448), .ZN(n5557) );
  INV_X1 U7101 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7102 ( .A1(n5550), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7103 ( .A1(n5035), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5518) );
  OAI211_X1 U7104 ( .C1(n5074), .C2(n5520), .A(n5519), .B(n5518), .ZN(n5521)
         );
  INV_X1 U7105 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U7106 ( .A1(n5523), .A2(SI_29_), .ZN(n5528) );
  INV_X1 U7107 ( .A(n5524), .ZN(n5526) );
  NAND2_X1 U7108 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  INV_X1 U7109 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7880) );
  INV_X1 U7110 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7845) );
  MUX2_X1 U7111 ( .A(n7880), .B(n7845), .S(n4325), .Z(n5530) );
  INV_X1 U7112 ( .A(SI_30_), .ZN(n5529) );
  NAND2_X1 U7113 ( .A1(n5530), .A2(n5529), .ZN(n5533) );
  INV_X1 U7114 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7115 ( .A1(n5531), .A2(SI_30_), .ZN(n5532) );
  NAND2_X1 U7116 ( .A1(n5533), .A2(n5532), .ZN(n5545) );
  MUX2_X1 U7117 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4325), .Z(n5535) );
  INV_X1 U7118 ( .A(SI_31_), .ZN(n5534) );
  XNOR2_X1 U7119 ( .A(n5535), .B(n5534), .ZN(n5536) );
  NAND2_X1 U7120 ( .A1(n9609), .A2(n5547), .ZN(n5539) );
  INV_X1 U7121 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8556) );
  OR2_X1 U7122 ( .A1(n5046), .A2(n8556), .ZN(n5538) );
  NAND2_X1 U7123 ( .A1(n5539), .A2(n5538), .ZN(n8410) );
  INV_X1 U7124 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7125 ( .A1(n5550), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7126 ( .A1(n5052), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5540) );
  OAI211_X1 U7127 ( .C1(n5542), .C2(n5553), .A(n5541), .B(n5540), .ZN(n5543)
         );
  INV_X1 U7128 ( .A(n5543), .ZN(n5544) );
  OR2_X1 U7129 ( .A1(n8410), .A2(n8163), .ZN(n5558) );
  NAND2_X1 U7130 ( .A1(n7844), .A2(n5547), .ZN(n5549) );
  OR2_X1 U7131 ( .A1(n5046), .A2(n7880), .ZN(n5548) );
  INV_X1 U7132 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7133 ( .A1(n5550), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7134 ( .A1(n5052), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5551) );
  OAI211_X1 U7135 ( .C1(n5554), .C2(n5553), .A(n5552), .B(n5551), .ZN(n5555)
         );
  INV_X1 U7136 ( .A(n5555), .ZN(n5556) );
  AND2_X1 U7137 ( .A1(n5557), .A2(n5556), .ZN(n6560) );
  NAND2_X1 U7138 ( .A1(n8412), .A2(n6560), .ZN(n5716) );
  NAND2_X1 U7139 ( .A1(n6576), .A2(n7869), .ZN(n5572) );
  AND2_X1 U7140 ( .A1(n5716), .A2(n5572), .ZN(n5712) );
  NAND2_X1 U7141 ( .A1(n5558), .A2(n5712), .ZN(n5745) );
  AOI21_X1 U7142 ( .B1(n6507), .B2(n5721), .A(n5745), .ZN(n5747) );
  NOR2_X1 U7143 ( .A1(n8412), .A2(n6560), .ZN(n5744) );
  OR2_X1 U7144 ( .A1(n5747), .A2(n5744), .ZN(n5569) );
  INV_X1 U7145 ( .A(n5559), .ZN(n5561) );
  NOR2_X1 U7146 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5560) );
  NAND2_X1 U7147 ( .A1(n5564), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5563) );
  MUX2_X1 U7148 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5563), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5565) );
  NAND2_X1 U7149 ( .A1(n5567), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5568) );
  AND2_X1 U7150 ( .A1(n7200), .A2(n5746), .ZN(n6553) );
  INV_X1 U7151 ( .A(n8163), .ZN(n5570) );
  NAND2_X1 U7152 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5574) );
  MUX2_X1 U7153 ( .A(n5700), .B(n4948), .S(n6561), .Z(n5706) );
  INV_X1 U7154 ( .A(n4366), .ZN(n8078) );
  INV_X1 U7155 ( .A(n6845), .ZN(n7041) );
  NAND2_X1 U7156 ( .A1(n8078), .A2(n7041), .ZN(n5730) );
  NAND2_X1 U7157 ( .A1(n5730), .A2(n7521), .ZN(n5575) );
  MUX2_X1 U7158 ( .A(n5575), .B(n7006), .S(n7485), .Z(n5581) );
  INV_X1 U7159 ( .A(n5576), .ZN(n5577) );
  OAI21_X1 U7160 ( .B1(n5581), .B2(n5577), .A(n5578), .ZN(n5579) );
  MUX2_X1 U7161 ( .A(n5579), .B(n5578), .S(n6561), .Z(n5584) );
  INV_X1 U7162 ( .A(n5730), .ZN(n5580) );
  NOR2_X1 U7163 ( .A1(n6508), .A2(n5580), .ZN(n5582) );
  AOI21_X1 U7164 ( .B1(n5582), .B2(n5581), .A(n7208), .ZN(n5583) );
  NAND2_X1 U7165 ( .A1(n5584), .A2(n5583), .ZN(n5591) );
  NAND2_X1 U7166 ( .A1(n5599), .A2(n5585), .ZN(n5588) );
  NAND2_X1 U7167 ( .A1(n5592), .A2(n5586), .ZN(n5587) );
  MUX2_X1 U7168 ( .A(n5588), .B(n5587), .S(n6584), .Z(n5589) );
  INV_X1 U7169 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7170 ( .A1(n5598), .A2(n5593), .ZN(n7267) );
  NAND2_X1 U7171 ( .A1(n5600), .A2(n5592), .ZN(n5594) );
  NAND3_X1 U7172 ( .A1(n5594), .A2(n5601), .A3(n5593), .ZN(n5597) );
  INV_X1 U7173 ( .A(n5605), .ZN(n5733) );
  AND2_X1 U7174 ( .A1(n5733), .A2(n5602), .ZN(n5596) );
  INV_X1 U7175 ( .A(n5732), .ZN(n5595) );
  AOI21_X1 U7176 ( .B1(n5597), .B2(n5596), .A(n5595), .ZN(n5608) );
  AOI21_X1 U7177 ( .B1(n5600), .B2(n5599), .A(n4630), .ZN(n5604) );
  INV_X1 U7178 ( .A(n5601), .ZN(n5603) );
  OAI21_X1 U7179 ( .B1(n5604), .B2(n5603), .A(n5602), .ZN(n5606) );
  AOI21_X1 U7180 ( .B1(n5606), .B2(n5732), .A(n5605), .ZN(n5607) );
  MUX2_X1 U7181 ( .A(n5608), .B(n5607), .S(n6584), .Z(n5623) );
  INV_X1 U7182 ( .A(n5609), .ZN(n5728) );
  NAND2_X1 U7183 ( .A1(n5616), .A2(n5728), .ZN(n5611) );
  NAND2_X1 U7184 ( .A1(n5729), .A2(n5613), .ZN(n5610) );
  MUX2_X1 U7185 ( .A(n5611), .B(n5610), .S(n6584), .Z(n5618) );
  NOR2_X1 U7186 ( .A1(n5618), .A2(n7465), .ZN(n5622) );
  AND2_X1 U7187 ( .A1(n5729), .A2(n5612), .ZN(n5614) );
  OAI211_X1 U7188 ( .C1(n5618), .C2(n5614), .A(n5624), .B(n5613), .ZN(n5620)
         );
  AND2_X1 U7189 ( .A1(n5728), .A2(n5615), .ZN(n5617) );
  OAI211_X1 U7190 ( .C1(n5618), .C2(n5617), .A(n4416), .B(n5616), .ZN(n5619)
         );
  MUX2_X1 U7191 ( .A(n5620), .B(n5619), .S(n6584), .Z(n5621) );
  AOI21_X1 U7192 ( .B1(n5623), .B2(n5622), .A(n5621), .ZN(n5631) );
  NAND2_X1 U7193 ( .A1(n5627), .A2(n4416), .ZN(n5626) );
  NAND2_X1 U7194 ( .A1(n5628), .A2(n5624), .ZN(n5625) );
  MUX2_X1 U7195 ( .A(n5626), .B(n5625), .S(n6584), .Z(n5630) );
  MUX2_X1 U7196 ( .A(n5628), .B(n5627), .S(n6584), .Z(n5629) );
  INV_X1 U7197 ( .A(n8400), .ZN(n8385) );
  OAI211_X1 U7198 ( .C1(n5631), .C2(n5630), .A(n5629), .B(n8385), .ZN(n5636)
         );
  NAND2_X1 U7199 ( .A1(n5641), .A2(n6561), .ZN(n5639) );
  NAND3_X1 U7200 ( .A1(n5639), .A2(n8003), .A3(n9913), .ZN(n5635) );
  INV_X1 U7201 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U7202 ( .A1(n5640), .A2(n6584), .ZN(n5638) );
  OAI21_X1 U7203 ( .B1(n5639), .B2(n5633), .A(n5638), .ZN(n5634) );
  NAND3_X1 U7204 ( .A1(n5636), .A2(n5635), .A3(n5634), .ZN(n5644) );
  INV_X1 U7205 ( .A(n5637), .ZN(n5646) );
  NAND2_X1 U7206 ( .A1(n5646), .A2(n5647), .ZN(n6536) );
  INV_X1 U7207 ( .A(n6536), .ZN(n8358) );
  NAND2_X1 U7208 ( .A1(n5639), .A2(n5638), .ZN(n5642) );
  NAND2_X1 U7209 ( .A1(n5641), .A2(n5640), .ZN(n8374) );
  NAND2_X1 U7210 ( .A1(n5642), .A2(n8374), .ZN(n5643) );
  NAND3_X1 U7211 ( .A1(n5644), .A2(n8358), .A3(n5643), .ZN(n5649) );
  INV_X1 U7212 ( .A(n5645), .ZN(n5651) );
  MUX2_X1 U7213 ( .A(n5647), .B(n5646), .S(n6561), .Z(n5648) );
  NAND3_X1 U7214 ( .A1(n5649), .A2(n6538), .A3(n5648), .ZN(n5656) );
  INV_X1 U7215 ( .A(n5650), .ZN(n5653) );
  NAND2_X1 U7216 ( .A1(n8286), .A2(n5651), .ZN(n5652) );
  MUX2_X1 U7217 ( .A(n5653), .B(n5652), .S(n6561), .Z(n5654) );
  INV_X1 U7218 ( .A(n8318), .ZN(n5658) );
  NOR2_X1 U7219 ( .A1(n5654), .A2(n5658), .ZN(n5655) );
  NAND2_X1 U7220 ( .A1(n5656), .A2(n5655), .ZN(n5657) );
  NAND2_X1 U7221 ( .A1(n5657), .A2(n6541), .ZN(n5660) );
  NOR2_X1 U7222 ( .A1(n5660), .A2(n5658), .ZN(n5662) );
  INV_X1 U7223 ( .A(n8286), .ZN(n5659) );
  OAI211_X1 U7224 ( .C1(n5660), .C2(n5659), .A(n8289), .B(n4937), .ZN(n5661)
         );
  MUX2_X1 U7225 ( .A(n5662), .B(n5661), .S(n6584), .Z(n5669) );
  NAND2_X1 U7226 ( .A1(n5668), .A2(n8305), .ZN(n5664) );
  OAI21_X1 U7227 ( .B1(n5669), .B2(n5664), .A(n5663), .ZN(n5665) );
  NAND3_X1 U7228 ( .A1(n5665), .A2(n8255), .A3(n5726), .ZN(n5666) );
  NAND3_X1 U7229 ( .A1(n5666), .A2(n5670), .A3(n5725), .ZN(n5667) );
  NAND2_X1 U7230 ( .A1(n5667), .A2(n6561), .ZN(n5679) );
  NAND3_X1 U7231 ( .A1(n5669), .A2(n5726), .A3(n5668), .ZN(n5672) );
  NAND2_X1 U7232 ( .A1(n5670), .A2(n8255), .ZN(n8273) );
  INV_X1 U7233 ( .A(n8273), .ZN(n5671) );
  NAND3_X1 U7234 ( .A1(n5672), .A2(n5671), .A3(n5727), .ZN(n5674) );
  NAND2_X1 U7235 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND3_X1 U7236 ( .A1(n5675), .A2(n6584), .A3(n5725), .ZN(n5678) );
  NAND3_X1 U7237 ( .A1(n8437), .A2(n8279), .A3(n6561), .ZN(n5676) );
  NAND2_X1 U7238 ( .A1(n8243), .A2(n5676), .ZN(n5677) );
  INV_X1 U7239 ( .A(n5680), .ZN(n5683) );
  NAND2_X1 U7240 ( .A1(n8210), .A2(n5681), .ZN(n5682) );
  MUX2_X1 U7241 ( .A(n5683), .B(n5682), .S(n6584), .Z(n5684) );
  NAND2_X1 U7242 ( .A1(n5688), .A2(n5685), .ZN(n8213) );
  NAND2_X1 U7243 ( .A1(n5688), .A2(n5416), .ZN(n5686) );
  NAND2_X1 U7244 ( .A1(n5686), .A2(n5685), .ZN(n5691) );
  INV_X1 U7245 ( .A(n5687), .ZN(n5689) );
  NAND2_X1 U7246 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  MUX2_X1 U7247 ( .A(n5691), .B(n5690), .S(n6561), .Z(n5693) );
  OR2_X1 U7248 ( .A1(n8206), .A2(n8215), .ZN(n6544) );
  NAND2_X1 U7249 ( .A1(n8206), .A2(n8215), .ZN(n6546) );
  INV_X1 U7250 ( .A(n8200), .ZN(n5692) );
  NAND2_X1 U7251 ( .A1(n5701), .A2(n5702), .ZN(n8188) );
  INV_X1 U7252 ( .A(n8188), .ZN(n8189) );
  MUX2_X1 U7253 ( .A(n5697), .B(n5696), .S(n6561), .Z(n5698) );
  NAND3_X1 U7254 ( .A1(n5699), .A2(n8189), .A3(n5698), .ZN(n5704) );
  MUX2_X1 U7255 ( .A(n5702), .B(n5701), .S(n6584), .Z(n5703) );
  NAND3_X1 U7256 ( .A1(n5704), .A2(n8177), .A3(n5703), .ZN(n5705) );
  AND2_X2 U7257 ( .A1(n5706), .A2(n5705), .ZN(n5709) );
  INV_X1 U7258 ( .A(n5709), .ZN(n5708) );
  MUX2_X1 U7259 ( .A(n6549), .B(n8418), .S(n6584), .Z(n5710) );
  INV_X1 U7260 ( .A(n5710), .ZN(n5707) );
  OR3_X2 U7261 ( .A1(n6551), .A2(n5713), .A3(n8179), .ZN(n5711) );
  NAND3_X1 U7262 ( .A1(n5712), .A2(n5711), .A3(n5714), .ZN(n5715) );
  INV_X1 U7263 ( .A(n5744), .ZN(n5718) );
  NAND2_X1 U7264 ( .A1(n5716), .A2(n7390), .ZN(n5717) );
  NOR2_X1 U7265 ( .A1(n5720), .A2(n5751), .ZN(n5753) );
  INV_X1 U7266 ( .A(n5721), .ZN(n5743) );
  INV_X1 U7267 ( .A(n8210), .ZN(n5722) );
  NOR2_X1 U7268 ( .A1(n5723), .A2(n5722), .ZN(n8229) );
  NAND2_X1 U7269 ( .A1(n5727), .A2(n5726), .ZN(n8293) );
  NAND2_X1 U7270 ( .A1(n5729), .A2(n5728), .ZN(n7479) );
  NAND2_X1 U7271 ( .A1(n5730), .A2(n7006), .ZN(n7032) );
  NOR3_X1 U7272 ( .A1(n7267), .A2(n7208), .A3(n7032), .ZN(n5731) );
  NAND2_X1 U7273 ( .A1(n7161), .A2(n9876), .ZN(n6521) );
  NAND2_X1 U7274 ( .A1(n8072), .A2(n7327), .ZN(n6522) );
  NAND2_X1 U7275 ( .A1(n6521), .A2(n6522), .ZN(n7320) );
  NAND4_X1 U7276 ( .A1(n7226), .A2(n4999), .A3(n5731), .A4(n7320), .ZN(n5734)
         );
  NAND2_X1 U7277 ( .A1(n5733), .A2(n5732), .ZN(n7438) );
  NOR4_X1 U7278 ( .A1(n7465), .A2(n7479), .A3(n5734), .A4(n7438), .ZN(n5735)
         );
  XNOR2_X1 U7279 ( .A(n9905), .B(n8067), .ZN(n7596) );
  NAND4_X1 U7280 ( .A1(n5735), .A2(n7662), .A3(n5157), .A4(n7596), .ZN(n5736)
         );
  NOR4_X1 U7281 ( .A1(n6536), .A2(n8400), .A3(n8374), .A4(n5736), .ZN(n5737)
         );
  NAND4_X1 U7282 ( .A1(n6541), .A2(n6538), .A3(n8332), .A4(n5737), .ZN(n5738)
         );
  NOR4_X1 U7283 ( .A1(n8273), .A2(n8309), .A3(n8293), .A4(n5738), .ZN(n5739)
         );
  NAND4_X1 U7284 ( .A1(n8229), .A2(n8243), .A3(n8260), .A4(n5739), .ZN(n5740)
         );
  NOR4_X1 U7285 ( .A1(n8188), .A2(n8200), .A3(n8213), .A4(n5740), .ZN(n5741)
         );
  NAND3_X1 U7286 ( .A1(n8177), .A2(n5741), .A3(n7862), .ZN(n5742) );
  NOR4_X1 U7287 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5749)
         );
  NAND2_X1 U7288 ( .A1(n7485), .A2(n5746), .ZN(n5870) );
  NAND3_X1 U7289 ( .A1(n5747), .A2(n8469), .A3(n6553), .ZN(n5748) );
  OAI21_X1 U7290 ( .B1(n5749), .B2(n5870), .A(n5748), .ZN(n5750) );
  AOI21_X1 U7291 ( .B1(n5751), .B2(n8163), .A(n5750), .ZN(n5752) );
  OAI21_X1 U7292 ( .B1(n5753), .B2(n8466), .A(n5752), .ZN(n5754) );
  XNOR2_X1 U7293 ( .A(n5754), .B(n5770), .ZN(n5777) );
  INV_X1 U7294 ( .A(n5973), .ZN(n5758) );
  NAND2_X1 U7295 ( .A1(n5758), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7560) );
  NAND2_X1 U7296 ( .A1(n5759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5760) );
  INV_X1 U7297 ( .A(n5761), .ZN(n5767) );
  NAND2_X1 U7298 ( .A1(n5767), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5762) );
  INV_X1 U7299 ( .A(n5764), .ZN(n5765) );
  NAND2_X1 U7300 ( .A1(n5765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5766) );
  NAND2_X2 U7301 ( .A1(n5768), .A2(n5767), .ZN(n7645) );
  NOR2_X1 U7302 ( .A1(n7700), .A2(n7645), .ZN(n5769) );
  NOR4_X1 U7303 ( .A1(n6581), .A2(n6559), .A3(n5771), .A4(n5971), .ZN(n5775)
         );
  OAI21_X1 U7304 ( .B1(n7560), .B2(n5773), .A(P2_B_REG_SCAN_IN), .ZN(n5774) );
  OR2_X1 U7305 ( .A1(n5775), .A2(n5774), .ZN(n5776) );
  OAI21_X1 U7306 ( .B1(n5777), .B2(n7560), .A(n5776), .ZN(P2_U3296) );
  XNOR2_X1 U7307 ( .A(n7645), .B(P2_B_REG_SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7308 ( .A1(n5778), .A2(n7700), .ZN(n5779) );
  INV_X1 U7309 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6726) );
  INV_X1 U7310 ( .A(n7645), .ZN(n5780) );
  OAI21_X2 U7311 ( .B1(n6586), .B2(n5870), .A(n5782), .ZN(n5812) );
  XNOR2_X1 U7312 ( .A(n8252), .B(n5824), .ZN(n5840) );
  INV_X1 U7313 ( .A(n5840), .ZN(n5842) );
  XNOR2_X1 U7314 ( .A(n8518), .B(n5817), .ZN(n5834) );
  XNOR2_X1 U7315 ( .A(n8533), .B(n5824), .ZN(n5829) );
  INV_X1 U7316 ( .A(n8538), .ZN(n8059) );
  XNOR2_X1 U7317 ( .A(n8059), .B(n5824), .ZN(n5828) );
  XNOR2_X1 U7318 ( .A(n6531), .B(n5824), .ZN(n7773) );
  XNOR2_X1 U7319 ( .A(n7662), .B(n5850), .ZN(n7996) );
  XNOR2_X1 U7320 ( .A(n9865), .B(n5817), .ZN(n5794) );
  XNOR2_X1 U7321 ( .A(n7210), .B(n5794), .ZN(n7042) );
  INV_X1 U7322 ( .A(n7042), .ZN(n5793) );
  INV_X1 U7323 ( .A(n5785), .ZN(n5784) );
  NAND2_X1 U7324 ( .A1(n6509), .A2(n5785), .ZN(n5787) );
  NAND2_X1 U7325 ( .A1(n7041), .A2(n5788), .ZN(n5786) );
  NAND2_X1 U7326 ( .A1(n7006), .A2(n5786), .ZN(n6913) );
  NAND2_X1 U7327 ( .A1(n6912), .A2(n5787), .ZN(n6950) );
  XNOR2_X1 U7328 ( .A(n9858), .B(n5788), .ZN(n5790) );
  XNOR2_X1 U7329 ( .A(n5790), .B(n5789), .ZN(n6951) );
  INV_X1 U7330 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7331 ( .A1(n5789), .A2(n5791), .ZN(n5792) );
  OR2_X1 U7332 ( .A1(n7210), .A2(n5794), .ZN(n5795) );
  XNOR2_X1 U7333 ( .A(n9872), .B(n5850), .ZN(n5796) );
  NAND2_X1 U7334 ( .A1(n7261), .A2(n5796), .ZN(n7255) );
  INV_X1 U7335 ( .A(n5796), .ZN(n5797) );
  NAND2_X1 U7336 ( .A1(n5797), .A2(n8074), .ZN(n5798) );
  AND2_X1 U7337 ( .A1(n7255), .A2(n5798), .ZN(n7158) );
  NAND2_X1 U7338 ( .A1(n7159), .A2(n7158), .ZN(n7157) );
  NAND2_X1 U7339 ( .A1(n7157), .A2(n7255), .ZN(n5799) );
  XNOR2_X1 U7340 ( .A(n9876), .B(n5850), .ZN(n5800) );
  XNOR2_X1 U7341 ( .A(n5800), .B(n8072), .ZN(n7256) );
  XNOR2_X1 U7342 ( .A(n7461), .B(n5850), .ZN(n5802) );
  XNOR2_X1 U7343 ( .A(n5802), .B(n8071), .ZN(n8022) );
  NAND2_X1 U7344 ( .A1(n7161), .A2(n5800), .ZN(n8018) );
  AND2_X1 U7345 ( .A1(n8022), .A2(n8018), .ZN(n5801) );
  INV_X1 U7346 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U7347 ( .A1(n5803), .A2(n8071), .ZN(n5804) );
  XNOR2_X1 U7348 ( .A(n7434), .B(n5824), .ZN(n5806) );
  XNOR2_X1 U7349 ( .A(n8026), .B(n5806), .ZN(n7429) );
  NAND2_X1 U7350 ( .A1(n8026), .A2(n5806), .ZN(n5807) );
  XNOR2_X1 U7351 ( .A(n9889), .B(n5824), .ZN(n5808) );
  INV_X1 U7352 ( .A(n5808), .ZN(n5809) );
  NAND2_X1 U7353 ( .A1(n5810), .A2(n5809), .ZN(n5811) );
  XNOR2_X1 U7354 ( .A(n7762), .B(n5824), .ZN(n5813) );
  XNOR2_X1 U7355 ( .A(n5813), .B(n7599), .ZN(n7759) );
  OR2_X1 U7356 ( .A1(n7599), .A2(n5813), .ZN(n5814) );
  NOR3_X1 U7357 ( .A1(n6531), .A2(n5850), .A3(n8067), .ZN(n5816) );
  INV_X1 U7358 ( .A(n7662), .ZN(n5815) );
  AOI211_X1 U7359 ( .C1(n8388), .C2(n5850), .A(n5816), .B(n5815), .ZN(n5820)
         );
  NOR3_X1 U7360 ( .A1(n9905), .A2(n8067), .A3(n5817), .ZN(n5818) );
  AOI211_X1 U7361 ( .C1(n8388), .C2(n5824), .A(n5818), .B(n7662), .ZN(n5819)
         );
  XNOR2_X1 U7362 ( .A(n9913), .B(n5824), .ZN(n5821) );
  NAND2_X1 U7363 ( .A1(n5821), .A2(n8003), .ZN(n7917) );
  OAI21_X1 U7364 ( .B1(n5820), .B2(n5819), .A(n7917), .ZN(n5823) );
  INV_X1 U7365 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U7366 ( .A1(n5822), .A2(n8378), .ZN(n7918) );
  XNOR2_X1 U7367 ( .A(n8549), .B(n5824), .ZN(n5825) );
  XNOR2_X1 U7368 ( .A(n5825), .B(n8390), .ZN(n7978) );
  INV_X1 U7369 ( .A(n5825), .ZN(n5826) );
  INV_X1 U7370 ( .A(n8390), .ZN(n8065) );
  XNOR2_X1 U7371 ( .A(n8368), .B(n5824), .ZN(n5827) );
  XNOR2_X1 U7372 ( .A(n5827), .B(n8376), .ZN(n7886) );
  XNOR2_X1 U7373 ( .A(n5828), .B(n8362), .ZN(n8047) );
  NAND2_X1 U7374 ( .A1(n8048), .A2(n8047), .ZN(n8046) );
  XNOR2_X1 U7375 ( .A(n5829), .B(n8326), .ZN(n7945) );
  XNOR2_X1 U7376 ( .A(n7955), .B(n5824), .ZN(n7952) );
  NAND2_X1 U7377 ( .A1(n7952), .A2(n8340), .ZN(n5831) );
  INV_X1 U7378 ( .A(n7952), .ZN(n5830) );
  XNOR2_X1 U7379 ( .A(n8522), .B(n5850), .ZN(n5832) );
  INV_X1 U7380 ( .A(n8325), .ZN(n8064) );
  NOR2_X1 U7381 ( .A1(n5832), .A2(n8064), .ZN(n5833) );
  AOI21_X1 U7382 ( .B1(n5832), .B2(n8064), .A(n5833), .ZN(n8011) );
  INV_X1 U7383 ( .A(n5833), .ZN(n7898) );
  XNOR2_X1 U7384 ( .A(n5834), .B(n8278), .ZN(n7899) );
  XNOR2_X1 U7385 ( .A(n8513), .B(n5824), .ZN(n5836) );
  XOR2_X1 U7386 ( .A(n8297), .B(n5836), .Z(n7970) );
  XNOR2_X1 U7387 ( .A(n8437), .B(n5850), .ZN(n5835) );
  NOR2_X1 U7388 ( .A1(n5835), .A2(n8062), .ZN(n7986) );
  AOI21_X1 U7389 ( .B1(n5835), .B2(n8062), .A(n7986), .ZN(n7909) );
  INV_X1 U7390 ( .A(n5836), .ZN(n5837) );
  INV_X1 U7391 ( .A(n8297), .ZN(n8063) );
  NAND2_X1 U7392 ( .A1(n5837), .A2(n8063), .ZN(n7910) );
  NAND2_X1 U7393 ( .A1(n7969), .A2(n5838), .ZN(n7908) );
  INV_X1 U7394 ( .A(n7986), .ZN(n5839) );
  NAND2_X1 U7395 ( .A1(n7908), .A2(n5839), .ZN(n5841) );
  XNOR2_X1 U7396 ( .A(n5840), .B(n8231), .ZN(n7985) );
  OAI21_X2 U7397 ( .B1(n5842), .B2(n8231), .A(n7988), .ZN(n7927) );
  XNOR2_X1 U7398 ( .A(n8220), .B(n5850), .ZN(n5846) );
  NAND2_X1 U7399 ( .A1(n5846), .A2(n8232), .ZN(n7930) );
  INV_X1 U7400 ( .A(n7930), .ZN(n5844) );
  NOR2_X1 U7401 ( .A1(n7928), .A2(n8248), .ZN(n5843) );
  NAND2_X1 U7402 ( .A1(n7928), .A2(n8248), .ZN(n5845) );
  INV_X1 U7403 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U7404 ( .A1(n5847), .A2(n7938), .ZN(n7931) );
  XNOR2_X1 U7405 ( .A(n8206), .B(n5824), .ZN(n5849) );
  XNOR2_X1 U7406 ( .A(n5849), .B(n8215), .ZN(n7932) );
  XNOR2_X1 U7407 ( .A(n8195), .B(n5850), .ZN(n5851) );
  XNOR2_X2 U7408 ( .A(n5853), .B(n5851), .ZN(n8035) );
  NAND2_X1 U7409 ( .A1(n8035), .A2(n8036), .ZN(n5885) );
  INV_X1 U7410 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U7411 ( .A1(n5853), .A2(n5852), .ZN(n5882) );
  NAND2_X1 U7412 ( .A1(n5885), .A2(n5882), .ZN(n5854) );
  XNOR2_X1 U7413 ( .A(n8183), .B(n5824), .ZN(n7858) );
  XNOR2_X1 U7414 ( .A(n7858), .B(n7868), .ZN(n5881) );
  NAND2_X1 U7415 ( .A1(n5854), .A2(n5881), .ZN(n5887) );
  INV_X1 U7416 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U7417 ( .A1(n6718), .A2(n6710), .ZN(n5857) );
  INV_X1 U7418 ( .A(n5855), .ZN(n8567) );
  NAND2_X1 U7419 ( .A1(n8567), .A2(n7700), .ZN(n5856) );
  INV_X1 U7420 ( .A(n6708), .ZN(n5858) );
  NAND2_X1 U7421 ( .A1(n5858), .A2(n6586), .ZN(n7028) );
  NOR2_X1 U7422 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .ZN(
        n5862) );
  NOR4_X1 U7423 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5861) );
  NOR4_X1 U7424 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5860) );
  NOR4_X1 U7425 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5859) );
  AND4_X1 U7426 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n5868)
         );
  NOR4_X1 U7427 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5866) );
  NOR4_X1 U7428 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5865) );
  NOR4_X1 U7429 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5864) );
  NOR4_X1 U7430 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5863) );
  AND4_X1 U7431 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n5867)
         );
  NAND2_X1 U7432 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U7433 ( .A1(n6718), .A2(n5869), .ZN(n6582) );
  INV_X1 U7434 ( .A(n6582), .ZN(n5895) );
  OR2_X1 U7435 ( .A1(n7028), .A2(n5895), .ZN(n5902) );
  INV_X1 U7436 ( .A(n6554), .ZN(n5872) );
  INV_X1 U7437 ( .A(n5870), .ZN(n5871) );
  NAND2_X1 U7438 ( .A1(n5872), .A2(n5871), .ZN(n5876) );
  INV_X1 U7439 ( .A(n5876), .ZN(n6572) );
  NAND2_X1 U7440 ( .A1(n6570), .A2(n6572), .ZN(n5880) );
  INV_X1 U7441 ( .A(n6586), .ZN(n5873) );
  NAND2_X1 U7442 ( .A1(n6708), .A2(n5873), .ZN(n6591) );
  INV_X1 U7443 ( .A(n6591), .ZN(n5875) );
  NOR2_X1 U7444 ( .A1(n6581), .A2(n5895), .ZN(n5874) );
  NOR2_X1 U7445 ( .A1(n9914), .A2(n6561), .ZN(n5877) );
  NAND2_X1 U7446 ( .A1(n5877), .A2(n5876), .ZN(n5894) );
  INV_X1 U7447 ( .A(n5894), .ZN(n5878) );
  NAND2_X1 U7448 ( .A1(n6571), .A2(n5878), .ZN(n5879) );
  INV_X1 U7449 ( .A(n5881), .ZN(n5883) );
  AND2_X1 U7450 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  NAND2_X1 U7451 ( .A1(n5885), .A2(n5884), .ZN(n7861) );
  NAND3_X1 U7452 ( .A1(n5887), .A2(n5886), .A3(n7861), .ZN(n5912) );
  NAND2_X1 U7453 ( .A1(n6571), .A2(n9914), .ZN(n5889) );
  NAND2_X1 U7454 ( .A1(n9914), .A2(n7201), .ZN(n6590) );
  INV_X1 U7455 ( .A(n6590), .ZN(n5888) );
  OR2_X1 U7456 ( .A1(n5771), .A2(n7877), .ZN(n5890) );
  NAND2_X1 U7457 ( .A1(n6562), .A2(n5890), .ZN(n6563) );
  INV_X1 U7458 ( .A(n6559), .ZN(n7033) );
  AND2_X1 U7459 ( .A1(n6563), .A2(n7033), .ZN(n5891) );
  INV_X1 U7460 ( .A(n8182), .ZN(n5907) );
  NAND2_X1 U7461 ( .A1(n5902), .A2(n6572), .ZN(n5899) );
  INV_X1 U7462 ( .A(n5892), .ZN(n6557) );
  NOR2_X1 U7463 ( .A1(n6580), .A2(n5972), .ZN(n5898) );
  INV_X1 U7464 ( .A(n7201), .ZN(n5893) );
  NAND2_X1 U7465 ( .A1(n9914), .A2(n5893), .ZN(n7031) );
  NAND2_X1 U7466 ( .A1(n5894), .A2(n7031), .ZN(n6569) );
  NAND2_X1 U7467 ( .A1(n6569), .A2(n6591), .ZN(n5897) );
  NAND2_X1 U7468 ( .A1(n6569), .A2(n5895), .ZN(n5896) );
  NAND4_X1 U7469 ( .A1(n5899), .A2(n5898), .A3(n5897), .A4(n5896), .ZN(n5900)
         );
  NAND2_X1 U7470 ( .A1(n5900), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5904) );
  NOR2_X1 U7471 ( .A1(n6581), .A2(n6559), .ZN(n5901) );
  NAND2_X1 U7472 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  NOR2_X1 U7473 ( .A1(n6563), .A2(n6559), .ZN(n5905) );
  NAND2_X1 U7474 ( .A1(n6570), .A2(n5905), .ZN(n8049) );
  AOI22_X1 U7475 ( .A1(n8202), .A2(n8038), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n5906) );
  OAI21_X1 U7476 ( .B1(n5907), .B2(n8040), .A(n5906), .ZN(n5908) );
  AOI21_X1 U7477 ( .B1(n8043), .B2(n8179), .A(n5908), .ZN(n5909) );
  NAND2_X1 U7478 ( .A1(n5912), .A2(n5911), .ZN(P2_U3154) );
  OAI21_X1 U7479 ( .B1(n6561), .B2(n5972), .A(n5973), .ZN(n6022) );
  NAND2_X1 U7480 ( .A1(n6022), .A2(n6562), .ZN(n5913) );
  NAND2_X1 U7481 ( .A1(n5913), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7482 ( .A(n5972), .ZN(n5914) );
  INV_X1 U7483 ( .A(n8150), .ZN(n8159) );
  NAND2_X1 U7484 ( .A1(n8159), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5940) );
  OAI21_X1 U7485 ( .B1(n8159), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5940), .ZN(
        n8152) );
  INV_X1 U7486 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9821) );
  INV_X1 U7487 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5915) );
  OAI21_X1 U7488 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n5915), .A(n5992), .ZN(n5916) );
  NAND2_X1 U7489 ( .A1(n5004), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7490 ( .A1(n5916), .A2(n5917), .ZN(n6667) );
  INV_X1 U7491 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6668) );
  NOR2_X1 U7492 ( .A1(n6667), .A2(n6668), .ZN(n6666) );
  INV_X1 U7493 ( .A(n5917), .ZN(n5918) );
  INV_X1 U7494 ( .A(n5919), .ZN(n7181) );
  XNOR2_X1 U7495 ( .A(n7190), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7182) );
  INV_X1 U7496 ( .A(n6678), .ZN(n7348) );
  INV_X1 U7497 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7333) );
  INV_X1 U7498 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5920) );
  AOI22_X1 U7499 ( .A1(n5998), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n5920), .B2(
        n7402), .ZN(n7404) );
  NOR2_X1 U7500 ( .A1(n9821), .A2(n9820), .ZN(n9819) );
  NOR2_X1 U7501 ( .A1(n9825), .A2(n5922), .ZN(n5923) );
  INV_X1 U7502 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7476) );
  MUX2_X1 U7503 ( .A(n7476), .B(P2_REG2_REG_8__SCAN_IN), .S(n6701), .Z(n7606)
         );
  NAND2_X1 U7504 ( .A1(n6701), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5924) );
  INV_X1 U7505 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7726) );
  INV_X1 U7506 ( .A(n5986), .ZN(n7794) );
  INV_X1 U7507 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5927) );
  AOI22_X1 U7508 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n5986), .B1(n7794), .B2(
        n5927), .ZN(n7785) );
  NOR2_X1 U7509 ( .A1(n5986), .A2(n5927), .ZN(n5928) );
  INV_X1 U7510 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U7511 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6764), .ZN(n5931) );
  OAI21_X1 U7512 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6764), .A(n5931), .ZN(
        n7817) );
  AND2_X1 U7513 ( .A1(n6764), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5932) );
  INV_X1 U7514 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9843) );
  INV_X1 U7515 ( .A(n9836), .ZN(n6821) );
  XOR2_X1 U7516 ( .A(n6821), .B(n5933), .Z(n9842) );
  NAND2_X1 U7517 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8085), .ZN(n5934) );
  OAI21_X1 U7518 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8085), .A(n5934), .ZN(
        n8079) );
  NOR2_X1 U7519 ( .A1(n8100), .A2(n5935), .ZN(n5936) );
  INV_X1 U7520 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8352) );
  INV_X1 U7521 ( .A(n8100), .ZN(n6910) );
  INV_X1 U7522 ( .A(n5977), .ZN(n8120) );
  INV_X1 U7523 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8342) );
  OAI21_X1 U7524 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8120), .A(n4442), .ZN(
        n8113) );
  OAI21_X1 U7525 ( .B1(n5937), .B2(n8138), .A(n5938), .ZN(n8131) );
  INV_X1 U7526 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8130) );
  NOR2_X1 U7527 ( .A1(n8131), .A2(n8130), .ZN(n8129) );
  INV_X1 U7528 ( .A(n5938), .ZN(n5939) );
  INV_X1 U7529 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8301) );
  XNOR2_X1 U7530 ( .A(n6556), .B(n8301), .ZN(n6018) );
  NOR2_X1 U7531 ( .A1(n5771), .A2(P2_U3151), .ZN(n8561) );
  NAND2_X1 U7532 ( .A1(n8561), .A2(n6022), .ZN(n7053) );
  INV_X1 U7533 ( .A(n9844), .ZN(n6975) );
  NAND2_X1 U7534 ( .A1(n8159), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U7535 ( .B1(n8159), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5968), .ZN(
        n8156) );
  INV_X1 U7536 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7537 ( .A1(n5986), .A2(n5955), .ZN(n5956) );
  INV_X1 U7538 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9922) );
  MUX2_X1 U7539 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9922), .S(n9800), .Z(n9813)
         );
  INV_X1 U7540 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7057) );
  NAND2_X1 U7541 ( .A1(n7057), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7542 ( .A1(n5992), .A2(n5942), .ZN(n5943) );
  NAND2_X1 U7543 ( .A1(n5004), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7544 ( .A1(n5943), .A2(n5945), .ZN(n6663) );
  INV_X1 U7545 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7546 ( .A1(n6663), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U7547 ( .A1(n5946), .A2(n5945), .ZN(n9812) );
  NAND2_X1 U7548 ( .A1(n9800), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7549 ( .A1(n5948), .A2(n6979), .ZN(n7171) );
  INV_X1 U7550 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7551 ( .A(n7190), .B(n5950), .ZN(n7172) );
  NAND2_X1 U7552 ( .A1(n7190), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5951) );
  INV_X1 U7553 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7457) );
  AOI22_X1 U7554 ( .A1(n5998), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n7457), .B2(
        n7402), .ZN(n7407) );
  NOR2_X1 U7555 ( .A1(n7408), .A2(n7407), .ZN(n7406) );
  INV_X1 U7556 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9928) );
  INV_X1 U7557 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5990) );
  MUX2_X1 U7558 ( .A(n5990), .B(P2_REG1_REG_8__SCAN_IN), .S(n6701), .Z(n7615)
         );
  INV_X1 U7559 ( .A(n5953), .ZN(n5954) );
  INV_X1 U7560 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U7561 ( .A1(n7724), .A2(n9931), .ZN(n7723) );
  MUX2_X1 U7562 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n5955), .S(n5986), .Z(n7782)
         );
  NAND2_X1 U7563 ( .A1(n5957), .A2(n7807), .ZN(n5958) );
  OR2_X1 U7564 ( .A1(n6764), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7565 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6764), .ZN(n5959) );
  NAND2_X1 U7566 ( .A1(n5960), .A2(n5959), .ZN(n7822) );
  NOR2_X1 U7567 ( .A1(n9836), .A2(n4385), .ZN(n5961) );
  INV_X1 U7568 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U7569 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8085), .ZN(n5962) );
  OAI21_X1 U7570 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8085), .A(n5962), .ZN(
        n8087) );
  NOR2_X1 U7571 ( .A1(n8088), .A2(n8087), .ZN(n8086) );
  NOR2_X1 U7572 ( .A1(n8100), .A2(n5963), .ZN(n5964) );
  INV_X1 U7573 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8454) );
  INV_X1 U7574 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5965) );
  AOI22_X1 U7575 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n5977), .B1(n8120), .B2(
        n5965), .ZN(n8122) );
  INV_X1 U7576 ( .A(n5966), .ZN(n5967) );
  INV_X1 U7577 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8450) );
  NOR2_X1 U7578 ( .A1(n8156), .A2(n8157), .ZN(n8155) );
  INV_X1 U7579 ( .A(n5968), .ZN(n5969) );
  NOR2_X1 U7580 ( .A1(n8155), .A2(n5969), .ZN(n5970) );
  XNOR2_X1 U7581 ( .A(n5770), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6017) );
  INV_X1 U7582 ( .A(n9853), .ZN(n9815) );
  AND2_X1 U7583 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7584 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7902) );
  MUX2_X1 U7585 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n7877), .Z(n6013) );
  XNOR2_X1 U7586 ( .A(n6013), .B(n5976), .ZN(n8134) );
  MUX2_X1 U7587 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n7877), .Z(n5978) );
  OR2_X1 U7588 ( .A1(n5978), .A2(n8120), .ZN(n6012) );
  XNOR2_X1 U7589 ( .A(n5978), .B(n5977), .ZN(n8116) );
  MUX2_X1 U7590 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n7877), .Z(n5979) );
  OR2_X1 U7591 ( .A1(n5979), .A2(n6910), .ZN(n6011) );
  XNOR2_X1 U7592 ( .A(n5979), .B(n8100), .ZN(n8099) );
  MUX2_X1 U7593 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n7877), .Z(n5981) );
  OR2_X1 U7594 ( .A1(n5981), .A2(n8085), .ZN(n6010) );
  XNOR2_X1 U7595 ( .A(n5981), .B(n5980), .ZN(n8082) );
  MUX2_X1 U7596 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n7877), .Z(n5982) );
  OR2_X1 U7597 ( .A1(n5982), .A2(n6821), .ZN(n6009) );
  XNOR2_X1 U7598 ( .A(n5982), .B(n9836), .ZN(n9848) );
  MUX2_X1 U7599 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n7877), .Z(n5983) );
  OR2_X1 U7600 ( .A1(n5983), .A2(n6764), .ZN(n6008) );
  XNOR2_X1 U7601 ( .A(n5983), .B(n7823), .ZN(n7820) );
  MUX2_X1 U7602 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n7877), .Z(n5985) );
  OR2_X1 U7603 ( .A1(n5985), .A2(n7807), .ZN(n6007) );
  XNOR2_X1 U7604 ( .A(n5985), .B(n5984), .ZN(n7801) );
  MUX2_X1 U7605 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n7877), .Z(n5987) );
  OR2_X1 U7606 ( .A1(n5987), .A2(n7794), .ZN(n6006) );
  XNOR2_X1 U7607 ( .A(n5987), .B(n5986), .ZN(n7790) );
  MUX2_X1 U7608 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n7877), .Z(n5989) );
  OR2_X1 U7609 ( .A1(n5989), .A2(n7735), .ZN(n6005) );
  XNOR2_X1 U7610 ( .A(n5989), .B(n5988), .ZN(n7730) );
  MUX2_X1 U7611 ( .A(n7476), .B(n5990), .S(n7877), .Z(n6002) );
  XNOR2_X1 U7612 ( .A(n6002), .B(n6701), .ZN(n7609) );
  MUX2_X1 U7613 ( .A(n9821), .B(n9928), .S(n7877), .Z(n5991) );
  NAND2_X1 U7614 ( .A1(n5991), .A2(n9825), .ZN(n6001) );
  XNOR2_X1 U7615 ( .A(n5991), .B(n6697), .ZN(n9831) );
  MUX2_X1 U7616 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n7877), .Z(n5999) );
  OR2_X1 U7617 ( .A1(n5999), .A2(n7402), .ZN(n6000) );
  MUX2_X1 U7618 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n7877), .Z(n5997) );
  MUX2_X1 U7619 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n7877), .Z(n5996) );
  MUX2_X1 U7620 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n7877), .Z(n5995) );
  MUX2_X1 U7621 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n7877), .Z(n5994) );
  AOI21_X1 U7622 ( .B1(n5993), .B2(n4504), .A(n6661), .ZN(n9808) );
  XNOR2_X1 U7623 ( .A(n5994), .B(n9800), .ZN(n9809) );
  NOR2_X1 U7624 ( .A1(n9808), .A2(n9809), .ZN(n9806) );
  XOR2_X1 U7625 ( .A(n5995), .B(n6979), .Z(n6972) );
  XNOR2_X1 U7626 ( .A(n5996), .B(n7190), .ZN(n7169) );
  AOI21_X1 U7627 ( .B1(n5996), .B2(n7190), .A(n7167), .ZN(n7344) );
  XNOR2_X1 U7628 ( .A(n5997), .B(n6678), .ZN(n7345) );
  NOR2_X1 U7629 ( .A1(n7344), .A2(n7345), .ZN(n7343) );
  XNOR2_X1 U7630 ( .A(n5999), .B(n5998), .ZN(n7399) );
  NAND2_X1 U7631 ( .A1(n6001), .A2(n9829), .ZN(n7608) );
  NAND2_X1 U7632 ( .A1(n7609), .A2(n7608), .ZN(n6004) );
  INV_X1 U7633 ( .A(n6701), .ZN(n7610) );
  NAND2_X1 U7634 ( .A1(n6002), .A2(n7610), .ZN(n6003) );
  NAND2_X1 U7635 ( .A1(n6004), .A2(n6003), .ZN(n7731) );
  NAND2_X1 U7636 ( .A1(n7730), .A2(n7731), .ZN(n7729) );
  NAND2_X1 U7637 ( .A1(n6005), .A2(n7729), .ZN(n7789) );
  NAND2_X1 U7638 ( .A1(n7790), .A2(n7789), .ZN(n7788) );
  NAND2_X1 U7639 ( .A1(n6006), .A2(n7788), .ZN(n7800) );
  NAND2_X1 U7640 ( .A1(n7801), .A2(n7800), .ZN(n7799) );
  NAND2_X1 U7641 ( .A1(n6007), .A2(n7799), .ZN(n7819) );
  NAND2_X1 U7642 ( .A1(n7820), .A2(n7819), .ZN(n7818) );
  NAND2_X1 U7643 ( .A1(n6008), .A2(n7818), .ZN(n9847) );
  NAND2_X1 U7644 ( .A1(n9848), .A2(n9847), .ZN(n9846) );
  NAND2_X1 U7645 ( .A1(n6009), .A2(n9846), .ZN(n8081) );
  NAND2_X1 U7646 ( .A1(n8082), .A2(n8081), .ZN(n8080) );
  NAND2_X1 U7647 ( .A1(n6010), .A2(n8080), .ZN(n8098) );
  NAND2_X1 U7648 ( .A1(n8099), .A2(n8098), .ZN(n8097) );
  NAND2_X1 U7649 ( .A1(n6011), .A2(n8097), .ZN(n8115) );
  NAND2_X1 U7650 ( .A1(n8116), .A2(n8115), .ZN(n8114) );
  NAND2_X1 U7651 ( .A1(n6012), .A2(n8114), .ZN(n8133) );
  INV_X1 U7652 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10121) );
  INV_X1 U7653 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8444) );
  MUX2_X1 U7654 ( .A(n10121), .B(n8444), .S(n7877), .Z(n6014) );
  NOR2_X1 U7655 ( .A1(n6015), .A2(n6014), .ZN(n8149) );
  OAI21_X1 U7656 ( .B1(n8149), .B2(n8159), .A(n6016), .ZN(n6020) );
  MUX2_X1 U7657 ( .A(n6018), .B(n6017), .S(n7877), .Z(n6019) );
  XNOR2_X1 U7658 ( .A(n6020), .B(n6019), .ZN(n6021) );
  AND2_X1 U7659 ( .A1(n6022), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6023) );
  MUX2_X1 U7660 ( .A(P2_U3893), .B(n6023), .S(n5771), .Z(n6024) );
  NAND2_X1 U7661 ( .A1(n6024), .A2(n6562), .ZN(n8139) );
  NAND2_X1 U7662 ( .A1(n9837), .A2(n6556), .ZN(n6025) );
  NOR2_X1 U7663 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6034) );
  NOR2_X1 U7664 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6033) );
  NOR2_X1 U7665 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6032) );
  NOR2_X1 U7666 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6031) );
  NAND4_X1 U7667 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n6036)
         );
  NAND4_X1 U7668 ( .A1(n6269), .A2(n10117), .A3(n6415), .A4(n6465), .ZN(n6035)
         );
  NOR2_X1 U7669 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U7670 ( .A1(n6469), .A2(n6039), .ZN(n6063) );
  NAND2_X1 U7671 ( .A1(n6058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6042) );
  MUX2_X1 U7672 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6042), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n6044) );
  INV_X1 U7673 ( .A(n6043), .ZN(n9611) );
  INV_X1 U7674 ( .A(n6048), .ZN(n6045) );
  NOR2_X1 U7675 ( .A1(n6047), .A2(n6045), .ZN(n6077) );
  INV_X1 U7676 ( .A(n6077), .ZN(n6046) );
  NAND2_X1 U7677 ( .A1(n6116), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7678 ( .A1(n6076), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7679 ( .A1(n4346), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7680 ( .A1(n6075), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6049) );
  NAND4_X2 U7681 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .ZN(n6863)
         );
  NAND2_X1 U7682 ( .A1(n4325), .A2(SI_0_), .ZN(n6054) );
  INV_X1 U7683 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7684 ( .A1(n6054), .A2(n6053), .ZN(n6056) );
  AND2_X1 U7685 ( .A1(n6056), .A2(n6055), .ZN(n9628) );
  OR3_X1 U7686 ( .A1(n6057), .A2(n6040), .A3(n9610), .ZN(n6062) );
  NAND2_X2 U7687 ( .A1(n6062), .A2(n6061), .ZN(n6459) );
  NAND2_X1 U7688 ( .A1(n6863), .A2(n9473), .ZN(n6877) );
  NAND2_X1 U7689 ( .A1(n6394), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7690 ( .A1(n6075), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7691 ( .A1(n6077), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7692 ( .A1(n6076), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6066) );
  INV_X1 U7693 ( .A(n6856), .ZN(n9198) );
  INV_X1 U7694 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6692) );
  INV_X1 U7695 ( .A(n6071), .ZN(n6691) );
  INV_X1 U7696 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7697 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6072) );
  XNOR2_X1 U7698 ( .A(n6073), .B(n6072), .ZN(n6690) );
  NAND2_X1 U7699 ( .A1(n9198), .A2(n7078), .ZN(n9110) );
  NAND2_X1 U7700 ( .A1(n6877), .A2(n6419), .ZN(n6879) );
  NAND2_X1 U7701 ( .A1(n6856), .A2(n7078), .ZN(n6074) );
  NAND2_X1 U7702 ( .A1(n6879), .A2(n6074), .ZN(n6925) );
  NAND2_X1 U7703 ( .A1(n4346), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7704 ( .A1(n6075), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7705 ( .A1(n6076), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7706 ( .A1(n6077), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7707 ( .A1(n6082), .A2(n9610), .ZN(n6107) );
  INV_X1 U7708 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7709 ( .A1(n6091), .A2(n6686), .ZN(n6084) );
  OR2_X1 U7710 ( .A1(n6112), .A2(n6687), .ZN(n6083) );
  OAI211_X2 U7711 ( .C1(n6632), .C2(n6685), .A(n6084), .B(n6083), .ZN(n6932)
         );
  NAND2_X1 U7712 ( .A1(n6938), .A2(n6932), .ZN(n6421) );
  INV_X1 U7713 ( .A(n6938), .ZN(n9197) );
  NAND2_X1 U7714 ( .A1(n6925), .A2(n9033), .ZN(n6924) );
  NAND2_X1 U7715 ( .A1(n6938), .A2(n7087), .ZN(n6085) );
  NAND2_X1 U7716 ( .A1(n6924), .A2(n6085), .ZN(n6936) );
  INV_X1 U7717 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7718 ( .A1(n4345), .A2(n6086), .ZN(n6090) );
  NAND2_X1 U7719 ( .A1(n6075), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7720 ( .A1(n6608), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7721 ( .A1(n6116), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6087) );
  NAND4_X1 U7722 ( .A1(n6090), .A2(n6089), .A3(n6088), .A4(n6087), .ZN(n9196)
         );
  OR2_X1 U7723 ( .A1(n6091), .A2(n6694), .ZN(n6098) );
  INV_X1 U7724 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6693) );
  OR2_X1 U7725 ( .A1(n6112), .A2(n6693), .ZN(n6097) );
  NAND2_X1 U7726 ( .A1(n6107), .A2(n6092), .ZN(n6093) );
  NAND2_X1 U7727 ( .A1(n6093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6095) );
  INV_X1 U7728 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6094) );
  XNOR2_X1 U7729 ( .A(n6095), .B(n6094), .ZN(n6695) );
  OR2_X1 U7730 ( .A1(n6632), .A2(n6695), .ZN(n6096) );
  NAND2_X1 U7731 ( .A1(n6936), .A2(n9034), .ZN(n6935) );
  INV_X1 U7732 ( .A(n9196), .ZN(n6904) );
  NAND2_X1 U7733 ( .A1(n6904), .A2(n6961), .ZN(n6099) );
  NAND2_X1 U7734 ( .A1(n6608), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6103) );
  NOR2_X1 U7735 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6100) );
  NOR2_X1 U7736 ( .A1(n6117), .A2(n6100), .ZN(n8846) );
  NAND2_X1 U7737 ( .A1(n4346), .A2(n8846), .ZN(n6102) );
  NAND2_X1 U7738 ( .A1(n6116), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6101) );
  NAND3_X1 U7739 ( .A1(n6103), .A2(n6102), .A3(n6101), .ZN(n6104) );
  OR2_X1 U7740 ( .A1(n6105), .A2(n9610), .ZN(n6106) );
  AND2_X1 U7741 ( .A1(n6107), .A2(n6106), .ZN(n6109) );
  INV_X1 U7742 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7743 ( .A1(n6109), .A2(n6108), .ZN(n6123) );
  INV_X1 U7744 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7745 ( .A1(n6110), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7746 ( .A1(n6123), .A2(n6111), .ZN(n6742) );
  OR2_X1 U7747 ( .A1(n6091), .A2(n6676), .ZN(n6114) );
  INV_X1 U7748 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6675) );
  OR2_X1 U7749 ( .A1(n6112), .A2(n6675), .ZN(n6113) );
  OAI211_X1 U7750 ( .C1(n6632), .C2(n6742), .A(n6114), .B(n6113), .ZN(n8847)
         );
  NAND2_X1 U7751 ( .A1(n7279), .A2(n8847), .ZN(n6425) );
  INV_X1 U7752 ( .A(n7279), .ZN(n9195) );
  INV_X1 U7753 ( .A(n8847), .ZN(n7277) );
  NAND2_X1 U7754 ( .A1(n9195), .A2(n7277), .ZN(n9108) );
  NAND2_X1 U7755 ( .A1(n6425), .A2(n9108), .ZN(n7018) );
  NAND2_X1 U7756 ( .A1(n7015), .A2(n7018), .ZN(n7014) );
  NAND2_X1 U7757 ( .A1(n7279), .A2(n7277), .ZN(n6115) );
  NAND2_X1 U7758 ( .A1(n7014), .A2(n6115), .ZN(n7121) );
  NAND2_X1 U7759 ( .A1(n9013), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7760 ( .A1(n9012), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6121) );
  NOR2_X1 U7761 ( .A1(n6117), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6118) );
  NOR2_X1 U7762 ( .A1(n6129), .A2(n6118), .ZN(n9757) );
  NAND2_X1 U7763 ( .A1(n4346), .A2(n9757), .ZN(n6120) );
  NAND2_X1 U7764 ( .A1(n6608), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7765 ( .A1(n6123), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6125) );
  INV_X1 U7766 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6124) );
  XNOR2_X1 U7767 ( .A(n6125), .B(n6124), .ZN(n6745) );
  OR2_X1 U7768 ( .A1(n6091), .A2(n6689), .ZN(n6127) );
  OR2_X1 U7769 ( .A1(n6112), .A2(n6688), .ZN(n6126) );
  OAI211_X1 U7770 ( .C1(n6632), .C2(n6745), .A(n6127), .B(n6126), .ZN(n7290)
         );
  NAND2_X1 U7771 ( .A1(n7097), .A2(n7290), .ZN(n6427) );
  INV_X1 U7772 ( .A(n7097), .ZN(n9194) );
  INV_X1 U7773 ( .A(n7290), .ZN(n9761) );
  NAND2_X1 U7774 ( .A1(n9194), .A2(n9761), .ZN(n9115) );
  NAND2_X1 U7775 ( .A1(n6427), .A2(n9115), .ZN(n9039) );
  NAND2_X1 U7776 ( .A1(n7121), .A2(n9039), .ZN(n7120) );
  NAND2_X1 U7777 ( .A1(n7097), .A2(n9761), .ZN(n6128) );
  NAND2_X1 U7778 ( .A1(n7120), .A2(n6128), .ZN(n7093) );
  NAND2_X1 U7779 ( .A1(n6608), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6135) );
  NOR2_X1 U7780 ( .A1(n6129), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6130) );
  NOR2_X1 U7781 ( .A1(n6143), .A2(n6130), .ZN(n7359) );
  NAND2_X1 U7782 ( .A1(n4345), .A2(n7359), .ZN(n6134) );
  NAND2_X1 U7783 ( .A1(n9012), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6133) );
  INV_X1 U7784 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6131) );
  OR2_X1 U7785 ( .A1(n6395), .A2(n6131), .ZN(n6132) );
  NAND2_X1 U7786 ( .A1(n6136), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6137) );
  MUX2_X1 U7787 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6137), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6139) );
  NAND2_X1 U7788 ( .A1(n6139), .A2(n6138), .ZN(n6746) );
  OR2_X1 U7789 ( .A1(n6091), .A2(n6684), .ZN(n6141) );
  OR2_X1 U7790 ( .A1(n6112), .A2(n6683), .ZN(n6140) );
  OAI211_X1 U7791 ( .C1(n6632), .C2(n6746), .A(n6141), .B(n6140), .ZN(n7364)
         );
  NAND2_X1 U7792 ( .A1(n7355), .A2(n7364), .ZN(n6429) );
  INV_X1 U7793 ( .A(n7355), .ZN(n9193) );
  NAND2_X1 U7794 ( .A1(n9193), .A2(n7354), .ZN(n7238) );
  NAND2_X1 U7795 ( .A1(n6429), .A2(n7238), .ZN(n7096) );
  NAND2_X1 U7796 ( .A1(n7355), .A2(n7354), .ZN(n6142) );
  NAND2_X1 U7797 ( .A1(n9013), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7798 ( .A1(n9012), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7799 ( .A1(n6143), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6168) );
  OAI21_X1 U7800 ( .B1(n6143), .B2(P1_REG3_REG_7__SCAN_IN), .A(n6168), .ZN(
        n7450) );
  INV_X1 U7801 ( .A(n7450), .ZN(n7245) );
  NAND2_X1 U7802 ( .A1(n4345), .A2(n7245), .ZN(n6145) );
  NAND2_X1 U7803 ( .A1(n6608), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7804 ( .A1(n6138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6149) );
  INV_X1 U7805 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6148) );
  XNOR2_X1 U7806 ( .A(n6149), .B(n6148), .ZN(n6747) );
  NAND2_X1 U7807 ( .A1(n7501), .A2(n7452), .ZN(n7502) );
  INV_X1 U7808 ( .A(n7501), .ZN(n9192) );
  NAND2_X1 U7809 ( .A1(n9192), .A2(n7247), .ZN(n7372) );
  NAND2_X1 U7810 ( .A1(n9013), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7811 ( .A1(n6608), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6152) );
  XNOR2_X1 U7812 ( .A(n6168), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U7813 ( .A1(n4345), .A2(n9744), .ZN(n6151) );
  NAND2_X1 U7814 ( .A1(n9012), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6150) );
  OR2_X1 U7815 ( .A1(n6702), .A2(n6091), .ZN(n6160) );
  OR2_X1 U7816 ( .A1(n6154), .A2(n9610), .ZN(n6157) );
  INV_X1 U7817 ( .A(n6157), .ZN(n6155) );
  NAND2_X1 U7818 ( .A1(n6155), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6158) );
  INV_X1 U7819 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7820 ( .A1(n6157), .A2(n6156), .ZN(n6162) );
  AND2_X1 U7821 ( .A1(n6158), .A2(n6162), .ZN(n6813) );
  AOI22_X1 U7822 ( .A1(n6300), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6299), .B2(
        n6813), .ZN(n6159) );
  NAND2_X1 U7823 ( .A1(n7570), .A2(n9746), .ZN(n7374) );
  INV_X1 U7824 ( .A(n9746), .ZN(n7510) );
  INV_X1 U7825 ( .A(n7570), .ZN(n9191) );
  NAND2_X1 U7826 ( .A1(n4574), .A2(n9191), .ZN(n7373) );
  NAND2_X1 U7827 ( .A1(n7374), .A2(n7373), .ZN(n7504) );
  NAND2_X1 U7828 ( .A1(n7500), .A2(n7504), .ZN(n7499) );
  NAND2_X1 U7829 ( .A1(n7570), .A2(n7510), .ZN(n6161) );
  NAND2_X1 U7830 ( .A1(n6704), .A2(n6602), .ZN(n6165) );
  NAND2_X1 U7831 ( .A1(n6162), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6163) );
  XNOR2_X1 U7832 ( .A(n6163), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6995) );
  AOI22_X1 U7833 ( .A1(n6300), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6299), .B2(
        n6995), .ZN(n6164) );
  NAND2_X1 U7834 ( .A1(n6165), .A2(n6164), .ZN(n7687) );
  NAND2_X1 U7835 ( .A1(n9013), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7836 ( .A1(n9012), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6172) );
  INV_X1 U7837 ( .A(n6168), .ZN(n6166) );
  AOI21_X1 U7838 ( .B1(n6166), .B2(P1_REG3_REG_8__SCAN_IN), .A(
        P1_REG3_REG_9__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7839 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n6167) );
  NOR2_X1 U7840 ( .A1(n6168), .A2(n6167), .ZN(n6182) );
  OR2_X1 U7841 ( .A1(n6169), .A2(n6182), .ZN(n7685) );
  INV_X1 U7842 ( .A(n7685), .ZN(n7383) );
  NAND2_X1 U7843 ( .A1(n4346), .A2(n7383), .ZN(n6171) );
  NAND2_X1 U7844 ( .A1(n6608), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6170) );
  OR2_X1 U7845 ( .A1(n7687), .A2(n7676), .ZN(n8941) );
  NAND2_X1 U7846 ( .A1(n7687), .A2(n7676), .ZN(n8938) );
  NAND2_X1 U7847 ( .A1(n8941), .A2(n8938), .ZN(n7379) );
  INV_X1 U7848 ( .A(n7676), .ZN(n9190) );
  OR2_X1 U7849 ( .A1(n7687), .A2(n9190), .ZN(n6174) );
  NAND2_X1 U7850 ( .A1(n6711), .A2(n6602), .ZN(n6181) );
  NOR2_X1 U7851 ( .A1(n6255), .A2(n9610), .ZN(n6175) );
  MUX2_X1 U7852 ( .A(n9610), .B(n6175), .S(P1_IR_REG_10__SCAN_IN), .Z(n6176)
         );
  INV_X1 U7853 ( .A(n6176), .ZN(n6179) );
  INV_X1 U7854 ( .A(n6177), .ZN(n6178) );
  AOI22_X1 U7855 ( .A1(n6300), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6299), .B2(
        n9637), .ZN(n6180) );
  NAND2_X1 U7856 ( .A1(n6181), .A2(n6180), .ZN(n9651) );
  NAND2_X1 U7857 ( .A1(n9013), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7858 ( .A1(n9012), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7859 ( .A1(n6182), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6196) );
  OR2_X1 U7860 ( .A1(n6182), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7861 ( .A1(n6196), .A2(n6183), .ZN(n9654) );
  INV_X1 U7862 ( .A(n9654), .ZN(n6184) );
  NAND2_X1 U7863 ( .A1(n4346), .A2(n6184), .ZN(n6187) );
  INV_X1 U7864 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7312) );
  OR2_X1 U7865 ( .A1(n6185), .A2(n7312), .ZN(n6186) );
  OR2_X1 U7866 ( .A1(n9651), .A2(n8585), .ZN(n9117) );
  NAND2_X1 U7867 ( .A1(n9651), .A2(n8585), .ZN(n8943) );
  NAND2_X1 U7868 ( .A1(n9117), .A2(n8943), .ZN(n9032) );
  NAND2_X1 U7869 ( .A1(n6721), .A2(n6602), .ZN(n6195) );
  NOR2_X1 U7870 ( .A1(n6177), .A2(n9610), .ZN(n6190) );
  MUX2_X1 U7871 ( .A(n9610), .B(n6190), .S(P1_IR_REG_11__SCAN_IN), .Z(n6191)
         );
  INV_X1 U7872 ( .A(n6191), .ZN(n6193) );
  AND2_X1 U7873 ( .A1(n6193), .A2(n6192), .ZN(n9655) );
  AOI22_X1 U7874 ( .A1(n6300), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6299), .B2(
        n9655), .ZN(n6194) );
  NAND2_X1 U7875 ( .A1(n6196), .A2(n8884), .ZN(n6197) );
  AND2_X1 U7876 ( .A1(n6210), .A2(n6197), .ZN(n8887) );
  NAND2_X1 U7877 ( .A1(n4345), .A2(n8887), .ZN(n6201) );
  NAND2_X1 U7878 ( .A1(n9013), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7879 ( .A1(n6608), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7880 ( .A1(n9012), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6198) );
  NAND4_X1 U7881 ( .A1(n6201), .A2(n6200), .A3(n6199), .A4(n6198), .ZN(n9188)
         );
  NAND2_X1 U7882 ( .A1(n8592), .A2(n9188), .ZN(n6202) );
  NAND2_X1 U7883 ( .A1(n7486), .A2(n6202), .ZN(n6204) );
  OR2_X1 U7884 ( .A1(n8592), .A2(n9188), .ZN(n6203) );
  NAND2_X1 U7885 ( .A1(n6763), .A2(n6602), .ZN(n6208) );
  NAND2_X1 U7886 ( .A1(n6192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6205) );
  MUX2_X1 U7887 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6205), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6206) );
  OR2_X1 U7888 ( .A1(n6192), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6228) );
  AOI22_X1 U7889 ( .A1(n6300), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6299), .B2(
        n7710), .ZN(n6207) );
  NAND2_X1 U7890 ( .A1(n9012), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6216) );
  AND2_X1 U7891 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  NOR2_X1 U7892 ( .A1(n6221), .A2(n6211), .ZN(n9731) );
  NAND2_X1 U7893 ( .A1(n4346), .A2(n9731), .ZN(n6215) );
  NAND2_X1 U7894 ( .A1(n6608), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6214) );
  INV_X1 U7895 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6212) );
  OR2_X1 U7896 ( .A1(n6395), .A2(n6212), .ZN(n6213) );
  OR2_X1 U7897 ( .A1(n9785), .A2(n7527), .ZN(n8949) );
  NAND2_X1 U7898 ( .A1(n9785), .A2(n7527), .ZN(n9125) );
  NAND2_X1 U7899 ( .A1(n9785), .A2(n9187), .ZN(n6217) );
  NAND2_X1 U7900 ( .A1(n6805), .A2(n6602), .ZN(n6220) );
  NAND2_X1 U7901 ( .A1(n6228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6218) );
  XNOR2_X1 U7902 ( .A(n6218), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9681) );
  AOI22_X1 U7903 ( .A1(n6300), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6299), .B2(
        n9681), .ZN(n6219) );
  NAND2_X2 U7904 ( .A1(n6220), .A2(n6219), .ZN(n8867) );
  NAND2_X1 U7905 ( .A1(n9012), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7906 ( .A1(n9013), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6225) );
  NOR2_X1 U7907 ( .A1(n6221), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6222) );
  OR2_X1 U7908 ( .A1(n6233), .A2(n6222), .ZN(n8865) );
  INV_X1 U7909 ( .A(n8865), .ZN(n7532) );
  NAND2_X1 U7910 ( .A1(n4345), .A2(n7532), .ZN(n6224) );
  NAND2_X1 U7911 ( .A1(n6608), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6223) );
  OR2_X1 U7912 ( .A1(n8867), .A2(n8790), .ZN(n8956) );
  NAND2_X1 U7913 ( .A1(n8867), .A2(n8790), .ZN(n9124) );
  NAND2_X1 U7914 ( .A1(n8956), .A2(n9124), .ZN(n9047) );
  INV_X1 U7915 ( .A(n8790), .ZN(n9186) );
  NAND2_X1 U7916 ( .A1(n8867), .A2(n9186), .ZN(n6227) );
  NAND2_X1 U7917 ( .A1(n6850), .A2(n6602), .ZN(n6232) );
  OAI21_X1 U7918 ( .B1(n6228), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7919 ( .A1(n6229), .A2(n10117), .ZN(n6241) );
  OR2_X1 U7920 ( .A1(n6229), .A2(n10117), .ZN(n6230) );
  AOI22_X1 U7921 ( .A1(n6300), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6299), .B2(
        n9693), .ZN(n6231) );
  NAND2_X2 U7922 ( .A1(n6232), .A2(n6231), .ZN(n8738) );
  NAND2_X1 U7923 ( .A1(n9013), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7924 ( .A1(n9012), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7925 ( .A1(n6233), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6246) );
  OR2_X1 U7926 ( .A1(n6233), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6234) );
  AND2_X1 U7927 ( .A1(n6246), .A2(n6234), .ZN(n8733) );
  NAND2_X1 U7928 ( .A1(n4345), .A2(n8733), .ZN(n6236) );
  NAND2_X1 U7929 ( .A1(n6608), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6235) );
  NAND4_X1 U7930 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n9185)
         );
  AND2_X1 U7931 ( .A1(n8738), .A2(n9185), .ZN(n6240) );
  OR2_X1 U7932 ( .A1(n8738), .A2(n9185), .ZN(n6239) );
  NAND2_X1 U7933 ( .A1(n6908), .A2(n6602), .ZN(n6245) );
  NAND2_X1 U7934 ( .A1(n6241), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6243) );
  INV_X1 U7935 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6242) );
  XNOR2_X1 U7936 ( .A(n6243), .B(n6242), .ZN(n7713) );
  INV_X1 U7937 ( .A(n7713), .ZN(n9706) );
  AOI22_X1 U7938 ( .A1(n6300), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6299), .B2(
        n9706), .ZN(n6244) );
  NAND2_X2 U7939 ( .A1(n6245), .A2(n6244), .ZN(n8609) );
  NAND2_X1 U7940 ( .A1(n9012), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7941 ( .A1(n9013), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7942 ( .A1(n6246), .A2(n8922), .ZN(n6247) );
  AND2_X1 U7943 ( .A1(n6261), .A2(n6247), .ZN(n8928) );
  NAND2_X1 U7944 ( .A1(n4346), .A2(n8928), .ZN(n6249) );
  NAND2_X1 U7945 ( .A1(n6608), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6248) );
  NAND4_X1 U7946 ( .A1(n6251), .A2(n6250), .A3(n6249), .A4(n6248), .ZN(n9184)
         );
  NAND2_X1 U7947 ( .A1(n7002), .A2(n6602), .ZN(n6259) );
  NOR2_X1 U7948 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6254) );
  NOR2_X1 U7949 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6253) );
  INV_X1 U7950 ( .A(n6270), .ZN(n6256) );
  NAND2_X1 U7951 ( .A1(n6256), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6257) );
  XNOR2_X1 U7952 ( .A(n6257), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7749) );
  AOI22_X1 U7953 ( .A1(n6300), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6299), .B2(
        n7749), .ZN(n6258) );
  NAND2_X1 U7954 ( .A1(n9012), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7955 ( .A1(n9013), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6265) );
  INV_X1 U7956 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7957 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  AND2_X1 U7958 ( .A1(n6274), .A2(n6262), .ZN(n9461) );
  NAND2_X1 U7959 ( .A1(n4346), .A2(n9461), .ZN(n6264) );
  NAND2_X1 U7960 ( .A1(n6608), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7961 ( .A1(n9603), .A2(n8821), .ZN(n8965) );
  NAND2_X1 U7962 ( .A1(n8966), .A2(n8965), .ZN(n9452) );
  NAND2_X1 U7963 ( .A1(n9451), .A2(n9452), .ZN(n6268) );
  INV_X1 U7964 ( .A(n8821), .ZN(n9183) );
  NAND2_X1 U7965 ( .A1(n9603), .A2(n9183), .ZN(n6267) );
  NAND2_X1 U7966 ( .A1(n7060), .A2(n6602), .ZN(n6272) );
  XNOR2_X1 U7967 ( .A(n6282), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9243) );
  AOI22_X1 U7968 ( .A1(n6300), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6299), .B2(
        n9243), .ZN(n6271) );
  NAND2_X1 U7969 ( .A1(n9013), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7970 ( .A1(n6608), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6278) );
  INV_X1 U7971 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6273) );
  AND2_X1 U7972 ( .A1(n6274), .A2(n6273), .ZN(n6275) );
  NOR2_X1 U7973 ( .A1(n6289), .A2(n6275), .ZN(n9445) );
  NAND2_X1 U7974 ( .A1(n4345), .A2(n9445), .ZN(n6277) );
  NAND2_X1 U7975 ( .A1(n9012), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6276) );
  NAND4_X1 U7976 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n9182)
         );
  OR2_X1 U7977 ( .A1(n9545), .A2(n9182), .ZN(n6280) );
  NAND2_X1 U7978 ( .A1(n7064), .A2(n6602), .ZN(n6288) );
  INV_X1 U7979 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7980 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  OR2_X1 U7981 ( .A1(n6285), .A2(n6284), .ZN(n6286) );
  AND2_X1 U7982 ( .A1(n6297), .A2(n6286), .ZN(n9713) );
  AOI22_X1 U7983 ( .A1(n6300), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6299), .B2(
        n9713), .ZN(n6287) );
  NAND2_X1 U7984 ( .A1(n9013), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7985 ( .A1(n9012), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6293) );
  OR2_X1 U7986 ( .A1(n6289), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7987 ( .A1(n6289), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6303) );
  AND2_X1 U7988 ( .A1(n6290), .A2(n6303), .ZN(n9431) );
  NAND2_X1 U7989 ( .A1(n4346), .A2(n9431), .ZN(n6292) );
  NAND2_X1 U7990 ( .A1(n6608), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6291) );
  NAND4_X1 U7991 ( .A1(n6294), .A2(n6293), .A3(n6292), .A4(n6291), .ZN(n8822)
         );
  NAND2_X1 U7992 ( .A1(n9594), .A2(n8822), .ZN(n6295) );
  NAND2_X1 U7993 ( .A1(n6296), .A2(n6295), .ZN(n9406) );
  INV_X1 U7994 ( .A(n9406), .ZN(n6309) );
  NAND2_X1 U7995 ( .A1(n7252), .A2(n6602), .ZN(n6302) );
  AOI22_X1 U7996 ( .A1(n6300), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9430), .B2(
        n6299), .ZN(n6301) );
  NAND2_X1 U7997 ( .A1(n9013), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7998 ( .A1(n9012), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6307) );
  INV_X1 U7999 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U8000 ( .A1(n6303), .A2(n8752), .ZN(n6304) );
  AND2_X1 U8001 ( .A1(n6315), .A2(n6304), .ZN(n9414) );
  NAND2_X1 U8002 ( .A1(n4346), .A2(n9414), .ZN(n6306) );
  NAND2_X1 U8003 ( .A1(n6608), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6305) );
  NAND4_X1 U8004 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n8854)
         );
  NAND2_X1 U8005 ( .A1(n6309), .A2(n4427), .ZN(n6311) );
  OR2_X1 U8006 ( .A1(n8648), .A2(n8854), .ZN(n6310) );
  NAND2_X1 U8007 ( .A1(n6311), .A2(n6310), .ZN(n9389) );
  NAND2_X1 U8008 ( .A1(n7367), .A2(n6602), .ZN(n6314) );
  OR2_X1 U8009 ( .A1(n6112), .A2(n6312), .ZN(n6313) );
  INV_X1 U8010 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8856) );
  AND2_X1 U8011 ( .A1(n6315), .A2(n8856), .ZN(n6316) );
  OR2_X1 U8012 ( .A1(n6316), .A2(n6325), .ZN(n9402) );
  NAND2_X1 U8013 ( .A1(n9013), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8014 ( .A1(n9012), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6317) );
  AND2_X1 U8015 ( .A1(n6318), .A2(n6317), .ZN(n6320) );
  NAND2_X1 U8016 ( .A1(n6608), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6319) );
  OAI211_X1 U8017 ( .C1(n9402), .C2(n6367), .A(n6320), .B(n6319), .ZN(n9181)
         );
  NOR2_X1 U8018 ( .A1(n9530), .A2(n9181), .ZN(n6321) );
  NAND2_X1 U8019 ( .A1(n9530), .A2(n9181), .ZN(n6322) );
  NAND2_X1 U8020 ( .A1(n7483), .A2(n6602), .ZN(n6324) );
  OR2_X1 U8021 ( .A1(n6112), .A2(n7832), .ZN(n6323) );
  NOR2_X1 U8022 ( .A1(n6325), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6326) );
  OR2_X1 U8023 ( .A1(n6333), .A2(n6326), .ZN(n9383) );
  AOI22_X1 U8024 ( .A1(n9012), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n9013), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U8025 ( .A1(n6608), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6327) );
  OAI211_X1 U8026 ( .C1(n9383), .C2(n6367), .A(n6328), .B(n6327), .ZN(n9180)
         );
  OR2_X1 U8027 ( .A1(n9382), .A2(n9180), .ZN(n6329) );
  NAND2_X1 U8028 ( .A1(n7520), .A2(n6602), .ZN(n6332) );
  OR2_X1 U8029 ( .A1(n6112), .A2(n10146), .ZN(n6331) );
  OR2_X1 U8030 ( .A1(n6333), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U8031 ( .A1(n6343), .A2(n6334), .ZN(n8875) );
  AOI22_X1 U8032 ( .A1(n9012), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n9013), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8033 ( .A1(n6608), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6335) );
  OAI211_X1 U8034 ( .C1(n8875), .C2(n6367), .A(n6336), .B(n6335), .ZN(n9179)
         );
  NOR2_X1 U8035 ( .A1(n9516), .A2(n9179), .ZN(n6337) );
  NAND2_X1 U8036 ( .A1(n9516), .A2(n9179), .ZN(n6338) );
  NAND2_X1 U8037 ( .A1(n6339), .A2(n6602), .ZN(n6341) );
  OR2_X1 U8038 ( .A1(n6112), .A2(n7559), .ZN(n6340) );
  INV_X1 U8039 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U8040 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  AND2_X1 U8041 ( .A1(n6353), .A2(n6344), .ZN(n9351) );
  NAND2_X1 U8042 ( .A1(n9351), .A2(n4345), .ZN(n6349) );
  INV_X1 U8043 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U8044 ( .A1(n9013), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U8045 ( .A1(n6608), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6345) );
  OAI211_X1 U8046 ( .C1(n6046), .C2(n9514), .A(n6346), .B(n6345), .ZN(n6347)
         );
  INV_X1 U8047 ( .A(n6347), .ZN(n6348) );
  NAND2_X1 U8048 ( .A1(n6349), .A2(n6348), .ZN(n9178) );
  AND2_X1 U8049 ( .A1(n9513), .A2(n9178), .ZN(n6350) );
  NAND2_X1 U8050 ( .A1(n7643), .A2(n6602), .ZN(n6352) );
  OR2_X1 U8051 ( .A1(n6112), .A2(n7646), .ZN(n6351) );
  INV_X1 U8052 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8836) );
  AND2_X1 U8053 ( .A1(n6353), .A2(n8836), .ZN(n6354) );
  OR2_X1 U8054 ( .A1(n6354), .A2(n6365), .ZN(n9340) );
  INV_X1 U8055 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U8056 ( .A1(n9013), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8057 ( .A1(n6608), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6355) );
  OAI211_X1 U8058 ( .C1(n6046), .C2(n6357), .A(n6356), .B(n6355), .ZN(n6358)
         );
  INV_X1 U8059 ( .A(n6358), .ZN(n6359) );
  NOR2_X1 U8060 ( .A1(n9504), .A2(n9177), .ZN(n6360) );
  NAND2_X1 U8061 ( .A1(n9504), .A2(n9177), .ZN(n6361) );
  NAND2_X1 U8062 ( .A1(n7699), .A2(n6602), .ZN(n6364) );
  OR2_X1 U8063 ( .A1(n6112), .A2(n7701), .ZN(n6363) );
  NAND2_X1 U8064 ( .A1(n6365), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6377) );
  OR2_X1 U8065 ( .A1(n6365), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U8066 ( .A1(n6377), .A2(n6366), .ZN(n9318) );
  INV_X1 U8067 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U8068 ( .A1(n6608), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U8069 ( .A1(n9013), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6368) );
  OAI211_X1 U8070 ( .C1(n6046), .C2(n10013), .A(n6369), .B(n6368), .ZN(n6370)
         );
  INV_X1 U8071 ( .A(n6370), .ZN(n6371) );
  AND2_X1 U8072 ( .A1(n9499), .A2(n9176), .ZN(n6373) );
  NAND2_X1 U8073 ( .A1(n8564), .A2(n6602), .ZN(n6375) );
  OR2_X1 U8074 ( .A1(n6112), .A2(n9624), .ZN(n6374) );
  NAND2_X1 U8075 ( .A1(n9013), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U8076 ( .A1(n9012), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U8077 ( .A1(n6608), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6379) );
  INV_X1 U8078 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6376) );
  AOI21_X1 U8079 ( .B1(n6377), .B2(n6376), .A(n6385), .ZN(n9310) );
  NAND2_X1 U8080 ( .A1(n4346), .A2(n9310), .ZN(n6378) );
  NAND4_X1 U8081 ( .A1(n6381), .A2(n6380), .A3(n6379), .A4(n6378), .ZN(n9175)
         );
  NOR2_X1 U8082 ( .A1(n8913), .A2(n9175), .ZN(n6382) );
  OR2_X1 U8083 ( .A1(n6112), .A2(n9621), .ZN(n6383) );
  NAND2_X1 U8084 ( .A1(n9013), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U8085 ( .A1(n9012), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6389) );
  INV_X1 U8086 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8725) );
  INV_X1 U8087 ( .A(n6385), .ZN(n6384) );
  NAND2_X1 U8088 ( .A1(n8725), .A2(n6384), .ZN(n6386) );
  NAND2_X1 U8089 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n6385), .ZN(n6454) );
  NAND2_X1 U8090 ( .A1(n4345), .A2(n9297), .ZN(n6388) );
  NAND2_X1 U8091 ( .A1(n6608), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8092 ( .A1(n9296), .A2(n8908), .ZN(n9007) );
  INV_X1 U8093 ( .A(n8908), .ZN(n9174) );
  NAND2_X1 U8094 ( .A1(n6391), .A2(n6602), .ZN(n6393) );
  OR2_X1 U8095 ( .A1(n6112), .A2(n9618), .ZN(n6392) );
  NAND2_X1 U8096 ( .A1(n9012), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6399) );
  XNOR2_X1 U8097 ( .A(n6454), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U8098 ( .A1(n4346), .A2(n8768), .ZN(n6398) );
  NAND2_X1 U8099 ( .A1(n6608), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6397) );
  OR2_X1 U8100 ( .A1(n6395), .A2(n6498), .ZN(n6396) );
  OR2_X1 U8101 ( .A1(n8773), .A2(n9277), .ZN(n9064) );
  NAND2_X1 U8102 ( .A1(n8773), .A2(n9277), .ZN(n9269) );
  NAND2_X1 U8103 ( .A1(n6400), .A2(n9267), .ZN(n6401) );
  NAND2_X1 U8104 ( .A1(n9265), .A2(n6401), .ZN(n7835) );
  INV_X1 U8105 ( .A(n6402), .ZN(n6403) );
  AND2_X1 U8106 ( .A1(n6415), .A2(n6408), .ZN(n6404) );
  NAND2_X1 U8107 ( .A1(n6416), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U8108 ( .A1(n6416), .A2(n6415), .ZN(n6407) );
  NAND2_X1 U8109 ( .A1(n6407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U8110 ( .A1(n6622), .A2(n9156), .ZN(n6417) );
  INV_X1 U8111 ( .A(n6836), .ZN(n9468) );
  AND2_X1 U8112 ( .A1(n6417), .A2(n9468), .ZN(n6418) );
  NAND2_X1 U8113 ( .A1(n6831), .A2(n9166), .ZN(n9467) );
  NAND2_X1 U8114 ( .A1(n6418), .A2(n9467), .ZN(n7491) );
  NAND2_X1 U8115 ( .A1(n9029), .A2(n9430), .ZN(n9161) );
  INV_X1 U8116 ( .A(n6863), .ZN(n6628) );
  NAND2_X1 U8117 ( .A1(n6628), .A2(n9473), .ZN(n6881) );
  INV_X1 U8118 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U8119 ( .A1(n6904), .A2(n7191), .ZN(n6423) );
  NAND2_X1 U8120 ( .A1(n9196), .A2(n6961), .ZN(n9107) );
  NAND2_X1 U8121 ( .A1(n6424), .A2(n9107), .ZN(n7019) );
  NAND2_X1 U8122 ( .A1(n7019), .A2(n6425), .ZN(n6426) );
  NAND2_X1 U8123 ( .A1(n8941), .A2(n7373), .ZN(n6431) );
  AND2_X1 U8124 ( .A1(n7502), .A2(n7374), .ZN(n6428) );
  OAI21_X1 U8125 ( .B1(n6431), .B2(n6428), .A(n8938), .ZN(n6432) );
  INV_X1 U8126 ( .A(n6429), .ZN(n7236) );
  NAND2_X1 U8127 ( .A1(n7372), .A2(n7238), .ZN(n6430) );
  NOR2_X1 U8128 ( .A1(n6431), .A2(n6430), .ZN(n9041) );
  OR2_X1 U8129 ( .A1(n6432), .A2(n9041), .ZN(n9118) );
  NAND2_X1 U8130 ( .A1(n7305), .A2(n8943), .ZN(n7488) );
  INV_X1 U8131 ( .A(n9188), .ZN(n6433) );
  OR2_X1 U8132 ( .A1(n8592), .A2(n6433), .ZN(n8944) );
  NAND2_X1 U8133 ( .A1(n8592), .A2(n6433), .ZN(n8947) );
  NAND2_X1 U8134 ( .A1(n8944), .A2(n8947), .ZN(n7487) );
  OAI21_X1 U8135 ( .B1(n7488), .B2(n7487), .A(n8944), .ZN(n9726) );
  INV_X1 U8136 ( .A(n9732), .ZN(n9725) );
  INV_X1 U8137 ( .A(n9124), .ZN(n6435) );
  INV_X1 U8138 ( .A(n9185), .ZN(n6436) );
  OR2_X1 U8139 ( .A1(n8738), .A2(n6436), .ZN(n9129) );
  NAND2_X1 U8140 ( .A1(n8738), .A2(n6436), .ZN(n8958) );
  NAND2_X1 U8141 ( .A1(n9129), .A2(n8958), .ZN(n9048) );
  INV_X1 U8142 ( .A(n9184), .ZN(n8613) );
  OR2_X1 U8143 ( .A1(n8609), .A2(n8613), .ZN(n8960) );
  NAND2_X1 U8144 ( .A1(n8609), .A2(n8613), .ZN(n8963) );
  INV_X1 U8145 ( .A(n8958), .ZN(n6437) );
  NOR2_X1 U8146 ( .A1(n9051), .A2(n6437), .ZN(n6438) );
  INV_X1 U8147 ( .A(n9452), .ZN(n9454) );
  NAND2_X1 U8148 ( .A1(n9455), .A2(n9454), .ZN(n9453) );
  NAND2_X1 U8149 ( .A1(n9453), .A2(n8966), .ZN(n9441) );
  XNOR2_X1 U8150 ( .A(n9545), .B(n9182), .ZN(n9440) );
  NAND2_X1 U8151 ( .A1(n9441), .A2(n9440), .ZN(n9439) );
  INV_X1 U8152 ( .A(n9182), .ZN(n8972) );
  OR2_X1 U8153 ( .A1(n9545), .A2(n8972), .ZN(n9422) );
  NAND2_X1 U8154 ( .A1(n9439), .A2(n9422), .ZN(n6440) );
  INV_X1 U8155 ( .A(n8822), .ZN(n6439) );
  NAND2_X1 U8156 ( .A1(n9594), .A2(n6439), .ZN(n8974) );
  NAND2_X1 U8157 ( .A1(n6440), .A2(n9424), .ZN(n9429) );
  INV_X1 U8158 ( .A(n8854), .ZN(n8894) );
  OR2_X1 U8159 ( .A1(n8648), .A2(n8894), .ZN(n8979) );
  NAND2_X1 U8160 ( .A1(n8648), .A2(n8894), .ZN(n9105) );
  NAND2_X1 U8161 ( .A1(n8979), .A2(n9105), .ZN(n9409) );
  INV_X1 U8162 ( .A(n9408), .ZN(n6441) );
  NOR2_X1 U8163 ( .A1(n9409), .A2(n6441), .ZN(n6442) );
  NAND2_X1 U8164 ( .A1(n9429), .A2(n6442), .ZN(n6443) );
  INV_X1 U8165 ( .A(n9181), .ZN(n6444) );
  OR2_X1 U8166 ( .A1(n9530), .A2(n6444), .ZN(n8980) );
  NAND2_X1 U8167 ( .A1(n9530), .A2(n6444), .ZN(n8988) );
  XNOR2_X1 U8168 ( .A(n9382), .B(n9180), .ZN(n9373) );
  INV_X1 U8169 ( .A(n9180), .ZN(n8932) );
  NAND2_X1 U8170 ( .A1(n9382), .A2(n8932), .ZN(n8991) );
  INV_X1 U8171 ( .A(n9179), .ZN(n6445) );
  OR2_X1 U8172 ( .A1(n9516), .A2(n6445), .ZN(n8982) );
  NAND2_X1 U8173 ( .A1(n9516), .A2(n6445), .ZN(n9078) );
  NAND2_X1 U8174 ( .A1(n9359), .A2(n9360), .ZN(n9358) );
  NAND2_X1 U8175 ( .A1(n9358), .A2(n9078), .ZN(n9345) );
  INV_X1 U8176 ( .A(n9178), .ZN(n8678) );
  OR2_X1 U8177 ( .A1(n9513), .A2(n8678), .ZN(n8984) );
  NAND2_X1 U8178 ( .A1(n9513), .A2(n8678), .ZN(n9077) );
  NAND2_X1 U8179 ( .A1(n9345), .A2(n9346), .ZN(n6446) );
  NAND2_X1 U8180 ( .A1(n6446), .A2(n9077), .ZN(n9337) );
  INV_X1 U8181 ( .A(n9177), .ZN(n6447) );
  NAND2_X1 U8182 ( .A1(n9504), .A2(n6447), .ZN(n9076) );
  NAND2_X1 U8183 ( .A1(n9068), .A2(n9076), .ZN(n9057) );
  NAND2_X1 U8184 ( .A1(n6448), .A2(n9068), .ZN(n9322) );
  INV_X1 U8185 ( .A(n9176), .ZN(n6449) );
  NAND2_X1 U8186 ( .A1(n9499), .A2(n6449), .ZN(n9083) );
  INV_X1 U8187 ( .A(n9175), .ZN(n6450) );
  XNOR2_X1 U8188 ( .A(n8913), .B(n6450), .ZN(n9304) );
  NAND2_X1 U8189 ( .A1(n8913), .A2(n6450), .ZN(n9146) );
  NAND2_X1 U8190 ( .A1(n9291), .A2(n9290), .ZN(n6451) );
  NAND2_X1 U8191 ( .A1(n6451), .A2(n9007), .ZN(n9268) );
  XNOR2_X1 U8192 ( .A(n9268), .B(n9267), .ZN(n6462) );
  OR2_X1 U8193 ( .A1(n9029), .A2(n9101), .ZN(n6452) );
  NAND2_X1 U8194 ( .A1(n9109), .A2(n6835), .ZN(n9158) );
  NAND2_X1 U8195 ( .A1(n9013), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8196 ( .A1(n9012), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6457) );
  INV_X1 U8197 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6453) );
  NOR2_X1 U8198 ( .A1(n6454), .A2(n6453), .ZN(n9284) );
  NAND2_X1 U8199 ( .A1(n4345), .A2(n9284), .ZN(n6456) );
  NAND2_X1 U8200 ( .A1(n6608), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6455) );
  NAND4_X1 U8201 ( .A1(n6458), .A2(n6457), .A3(n6456), .A4(n6455), .ZN(n9172)
         );
  NAND2_X1 U8202 ( .A1(n9172), .A2(n8874), .ZN(n6461) );
  INV_X1 U8203 ( .A(n6459), .ZN(n6648) );
  NAND2_X1 U8204 ( .A1(n9174), .A2(n9167), .ZN(n6460) );
  NAND2_X1 U8205 ( .A1(n6461), .A2(n6460), .ZN(n8769) );
  AOI21_X1 U8206 ( .B1(n6462), .B2(n9729), .A(n8769), .ZN(n7836) );
  NAND2_X1 U8207 ( .A1(n6940), .A2(n6961), .ZN(n7017) );
  OR2_X1 U8208 ( .A1(n7017), .A2(n8847), .ZN(n7123) );
  INV_X1 U8209 ( .A(n9651), .ZN(n9780) );
  INV_X1 U8210 ( .A(n9594), .ZN(n9433) );
  NAND2_X1 U8211 ( .A1(n9420), .A2(n9535), .ZN(n9407) );
  INV_X1 U8212 ( .A(n9516), .ZN(n9369) );
  INV_X1 U8213 ( .A(n9513), .ZN(n9354) );
  NAND2_X1 U8214 ( .A1(n9566), .A2(n9317), .ZN(n9309) );
  AOI21_X1 U8215 ( .B1(n8773), .B2(n9295), .A(n9736), .ZN(n6463) );
  NAND2_X1 U8216 ( .A1(n6463), .A2(n9281), .ZN(n7837) );
  NAND2_X1 U8217 ( .A1(n6473), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6475) );
  OAI211_X1 U8218 ( .C1(n9166), .C2(n9099), .A(n7557), .B(n6827), .ZN(n6477)
         );
  INV_X1 U8219 ( .A(n6477), .ZN(n6825) );
  NOR4_X1 U8220 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6481) );
  NOR4_X1 U8221 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6480) );
  NOR4_X1 U8222 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6479) );
  NOR4_X1 U8223 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6478) );
  NAND4_X1 U8224 ( .A1(n6481), .A2(n6480), .A3(n6479), .A4(n6478), .ZN(n6490)
         );
  NOR2_X1 U8225 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n6485) );
  NOR4_X1 U8226 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6484) );
  NOR4_X1 U8227 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6483) );
  NOR4_X1 U8228 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6482) );
  NAND4_X1 U8229 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n6489)
         );
  NAND2_X1 U8230 ( .A1(n7703), .A2(P1_B_REG_SCAN_IN), .ZN(n6487) );
  INV_X1 U8231 ( .A(n7648), .ZN(n6486) );
  MUX2_X1 U8232 ( .A(n6487), .B(P1_B_REG_SCAN_IN), .S(n6486), .Z(n6488) );
  OAI21_X1 U8233 ( .B1(n6490), .B2(n6489), .A(n6494), .ZN(n6824) );
  INV_X1 U8234 ( .A(n6491), .ZN(n9627) );
  NAND2_X1 U8235 ( .A1(n9627), .A2(n7703), .ZN(n6492) );
  NAND2_X1 U8236 ( .A1(n9505), .A2(n9430), .ZN(n6837) );
  INV_X1 U8237 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8238 ( .A1(n6494), .A2(n6493), .ZN(n6496) );
  NAND2_X1 U8239 ( .A1(n9627), .A2(n7648), .ZN(n6495) );
  INV_X1 U8240 ( .A(n9608), .ZN(n6497) );
  NAND2_X1 U8241 ( .A1(n6614), .A2(n6498), .ZN(n6499) );
  INV_X1 U8242 ( .A(n8773), .ZN(n6500) );
  INV_X1 U8243 ( .A(n9604), .ZN(n6501) );
  NAND2_X1 U8244 ( .A1(n6503), .A2(n6502), .ZN(P1_U3518) );
  INV_X1 U8245 ( .A(n9553), .ZN(n6505) );
  NAND2_X1 U8246 ( .A1(n8773), .A2(n9553), .ZN(n6506) );
  INV_X1 U8247 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6575) );
  INV_X1 U8248 ( .A(n8175), .ZN(n6568) );
  AND2_X1 U8249 ( .A1(n7521), .A2(n7201), .ZN(n9880) );
  INV_X1 U8250 ( .A(n8220), .ZN(n8495) );
  INV_X1 U8251 ( .A(n8533), .ZN(n7947) );
  OR2_X1 U8252 ( .A1(n4366), .A2(n7041), .ZN(n7008) );
  NAND2_X1 U8253 ( .A1(n6508), .A2(n7008), .ZN(n6511) );
  NAND2_X1 U8254 ( .A1(n6509), .A2(n7011), .ZN(n6510) );
  NAND2_X1 U8255 ( .A1(n5789), .A2(n6953), .ZN(n6512) );
  AND2_X1 U8256 ( .A1(n7210), .A2(n6513), .ZN(n6514) );
  OR2_X1 U8257 ( .A1(n7210), .A2(n6513), .ZN(n6516) );
  NAND2_X1 U8258 ( .A1(n4367), .A2(n7261), .ZN(n6520) );
  OR2_X1 U8259 ( .A1(n7225), .A2(n6515), .ZN(n6518) );
  NAND2_X1 U8260 ( .A1(n6520), .A2(n6519), .ZN(n7321) );
  INV_X1 U8261 ( .A(n6521), .ZN(n6523) );
  INV_X1 U8262 ( .A(n7461), .ZN(n8029) );
  AND2_X1 U8263 ( .A1(n8071), .A2(n8029), .ZN(n6526) );
  INV_X1 U8264 ( .A(n8071), .ZN(n6524) );
  NAND2_X1 U8265 ( .A1(n6524), .A2(n7461), .ZN(n6525) );
  NAND2_X1 U8266 ( .A1(n8069), .A2(n7478), .ZN(n6527) );
  AND2_X1 U8267 ( .A1(n7465), .A2(n6527), .ZN(n6529) );
  INV_X1 U8268 ( .A(n6527), .ZN(n6528) );
  NAND2_X1 U8269 ( .A1(n8026), .A2(n9882), .ZN(n7467) );
  AND2_X1 U8270 ( .A1(n7479), .A2(n7467), .ZN(n7470) );
  NOR2_X1 U8271 ( .A1(n7599), .A2(n9894), .ZN(n6530) );
  NAND2_X1 U8272 ( .A1(n6532), .A2(n5815), .ZN(n7665) );
  INV_X1 U8273 ( .A(n8388), .ZN(n8066) );
  NAND2_X1 U8274 ( .A1(n9908), .A2(n8066), .ZN(n6533) );
  OR2_X1 U8275 ( .A1(n9913), .A2(n8378), .ZN(n6534) );
  NAND2_X1 U8276 ( .A1(n9913), .A2(n8378), .ZN(n6535) );
  INV_X1 U8277 ( .A(n8374), .ZN(n8372) );
  OR2_X1 U8278 ( .A1(n8549), .A2(n8065), .ZN(n8357) );
  AND2_X1 U8279 ( .A1(n6536), .A2(n8357), .ZN(n6537) );
  NAND2_X1 U8280 ( .A1(n8368), .A2(n8376), .ZN(n8347) );
  INV_X1 U8281 ( .A(n8332), .ZN(n8336) );
  NAND2_X1 U8282 ( .A1(n8059), .A2(n8362), .ZN(n8334) );
  NAND2_X1 U8283 ( .A1(n8333), .A2(n6540), .ZN(n8335) );
  OAI21_X1 U8284 ( .B1(n8326), .B2(n7947), .A(n8335), .ZN(n8322) );
  INV_X1 U8285 ( .A(n8522), .ZN(n8017) );
  NAND2_X1 U8286 ( .A1(n8017), .A2(n8325), .ZN(n8294) );
  INV_X1 U8287 ( .A(n8278), .ZN(n8311) );
  NAND2_X1 U8288 ( .A1(n8518), .A2(n8311), .ZN(n8274) );
  INV_X1 U8289 ( .A(n8513), .ZN(n7976) );
  NAND2_X1 U8290 ( .A1(n7976), .A2(n8297), .ZN(n8259) );
  NAND2_X1 U8291 ( .A1(n8258), .A2(n8259), .ZN(n8241) );
  NOR2_X1 U8292 ( .A1(n8243), .A2(n8260), .ZN(n6543) );
  OR2_X1 U8293 ( .A1(n8437), .A2(n8062), .ZN(n8244) );
  OAI22_X1 U8294 ( .A1(n8243), .A2(n8244), .B1(n8231), .B2(n8252), .ZN(n6542)
         );
  INV_X1 U8295 ( .A(n6544), .ZN(n6545) );
  AOI21_X1 U8296 ( .B1(n8201), .B2(n6546), .A(n6545), .ZN(n8190) );
  OAI21_X1 U8297 ( .B1(n8202), .B2(n8195), .A(n8190), .ZN(n6547) );
  INV_X2 U8298 ( .A(n7868), .ZN(n8191) );
  NOR2_X1 U8299 ( .A1(n7872), .A2(n8179), .ZN(n6550) );
  INV_X1 U8300 ( .A(n6553), .ZN(n6555) );
  OR2_X1 U8301 ( .A1(n7521), .A2(n6556), .ZN(n6585) );
  NAND2_X1 U8302 ( .A1(n6585), .A2(n6557), .ZN(n6558) );
  NAND3_X1 U8303 ( .A1(n6559), .A2(n9893), .A3(n6558), .ZN(n9901) );
  INV_X1 U8304 ( .A(n6560), .ZN(n8060) );
  AOI21_X1 U8305 ( .B1(P2_B_REG_SCAN_IN), .B2(n6562), .A(n8389), .ZN(n8161) );
  AOI22_X1 U8306 ( .A1(n8060), .A2(n8161), .B1(n8377), .B2(n8179), .ZN(n6564)
         );
  OAI21_X1 U8307 ( .B1(n8175), .B2(n9901), .A(n6564), .ZN(n6565) );
  INV_X1 U8308 ( .A(n6565), .ZN(n6566) );
  NAND2_X1 U8309 ( .A1(n6567), .A2(n6566), .ZN(n8168) );
  AOI21_X1 U8310 ( .B1(n6568), .B2(n9880), .A(n8168), .ZN(n6592) );
  NAND2_X1 U8311 ( .A1(n6570), .A2(n6569), .ZN(n6574) );
  OAI21_X1 U8312 ( .B1(n7033), .B2(n6572), .A(n6571), .ZN(n6573) );
  MUX2_X1 U8313 ( .A(n6575), .B(n6592), .S(n9919), .Z(n6579) );
  NAND2_X1 U8314 ( .A1(n6576), .A2(n6577), .ZN(n6578) );
  NAND2_X1 U8315 ( .A1(n6579), .A2(n6578), .ZN(P2_U3456) );
  INV_X1 U8316 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6593) );
  NOR2_X1 U8317 ( .A1(n6581), .A2(n6580), .ZN(n6583) );
  OAI21_X1 U8318 ( .B1(n7390), .B2(n6585), .A(n6584), .ZN(n6587) );
  OR2_X1 U8319 ( .A1(n6587), .A2(n6586), .ZN(n6589) );
  NAND2_X1 U8320 ( .A1(n6587), .A2(n6708), .ZN(n6588) );
  MUX2_X1 U8321 ( .A(n6593), .B(n6592), .S(n9938), .Z(n6596) );
  NAND2_X1 U8322 ( .A1(n6576), .A2(n6594), .ZN(n6595) );
  NAND2_X1 U8323 ( .A1(n6596), .A2(n6595), .ZN(P2_U3488) );
  NAND2_X1 U8324 ( .A1(n9609), .A2(n6602), .ZN(n6599) );
  INV_X1 U8325 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6597) );
  OR2_X1 U8326 ( .A1(n6112), .A2(n6597), .ZN(n6598) );
  NAND2_X1 U8327 ( .A1(n7844), .A2(n6602), .ZN(n6601) );
  OR2_X1 U8328 ( .A1(n6112), .A2(n7845), .ZN(n6600) );
  NAND2_X1 U8329 ( .A1(n7882), .A2(n6602), .ZN(n6604) );
  INV_X1 U8330 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9616) );
  OR2_X1 U8331 ( .A1(n6112), .A2(n9616), .ZN(n6603) );
  XNOR2_X1 U8332 ( .A(n9481), .B(n9259), .ZN(n6607) );
  NOR2_X2 U8333 ( .A1(n6607), .A2(n9736), .ZN(n9257) );
  NAND2_X1 U8334 ( .A1(n9012), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8335 ( .A1(n6608), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U8336 ( .A1(n9013), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6609) );
  AND3_X1 U8337 ( .A1(n6611), .A2(n6610), .A3(n6609), .ZN(n9060) );
  INV_X1 U8338 ( .A(n6612), .ZN(n9165) );
  NAND2_X1 U8339 ( .A1(n9165), .A2(P1_B_REG_SCAN_IN), .ZN(n6613) );
  NAND2_X1 U8340 ( .A1(n8874), .A2(n6613), .ZN(n9274) );
  NOR2_X1 U8341 ( .A1(n9060), .A2(n9274), .ZN(n9482) );
  NOR2_X1 U8342 ( .A1(n9257), .A2(n9482), .ZN(n9478) );
  OR2_X1 U8343 ( .A1(n9478), .A2(n6614), .ZN(n6618) );
  INV_X1 U8344 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6615) );
  INV_X1 U8345 ( .A(n6616), .ZN(n6617) );
  NAND2_X1 U8346 ( .A1(n6618), .A2(n6617), .ZN(P1_U3521) );
  NOR2_X1 U8347 ( .A1(n6827), .A2(P1_U3086), .ZN(n6619) );
  NAND2_X1 U8348 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6636) );
  INV_X1 U8349 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6625) );
  INV_X1 U8350 ( .A(n6621), .ZN(n6620) );
  NAND2_X1 U8351 ( .A1(n6827), .A2(n6620), .ZN(n6626) );
  NAND2_X1 U8352 ( .A1(n6863), .A2(n6895), .ZN(n6624) );
  NAND2_X1 U8353 ( .A1(n9473), .A2(n7289), .ZN(n6623) );
  AND2_X1 U8354 ( .A1(n6624), .A2(n6623), .ZN(n6853) );
  OAI21_X1 U8355 ( .B1(n6827), .B2(n6625), .A(n6853), .ZN(n6854) );
  INV_X1 U8356 ( .A(n9473), .ZN(n6872) );
  INV_X1 U8357 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6735) );
  OAI222_X1 U8358 ( .A1(n8764), .A2(n6872), .B1(n8677), .B2(n6628), .C1(n6827), 
        .C2(n6735), .ZN(n6855) );
  XOR2_X1 U8359 ( .A(n6854), .B(n6855), .Z(n6833) );
  MUX2_X1 U8360 ( .A(n6636), .B(n6833), .S(n6612), .Z(n6630) );
  OAI21_X1 U8361 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n6612), .A(n6648), .ZN(
        n6733) );
  NAND2_X1 U8362 ( .A1(n6733), .A2(n6735), .ZN(n6629) );
  OAI211_X1 U8363 ( .C1(n6630), .C2(n6459), .A(P1_U3973), .B(n6629), .ZN(n9224) );
  INV_X1 U8364 ( .A(n9224), .ZN(n6660) );
  INV_X1 U8365 ( .A(n6827), .ZN(n6631) );
  AOI21_X1 U8366 ( .B1(n6631), .B2(n7557), .A(P1_U3086), .ZN(n6642) );
  NAND2_X1 U8367 ( .A1(n7557), .A2(n6831), .ZN(n6633) );
  NAND2_X1 U8368 ( .A1(n6633), .A2(n6632), .ZN(n6640) );
  INV_X1 U8369 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6647) );
  XNOR2_X1 U8370 ( .A(n6742), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6645) );
  INV_X1 U8371 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6634) );
  MUX2_X1 U8372 ( .A(n6634), .B(P1_REG2_REG_2__SCAN_IN), .S(n6685), .Z(n9217)
         );
  INV_X1 U8373 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6635) );
  MUX2_X1 U8374 ( .A(n6635), .B(P1_REG2_REG_1__SCAN_IN), .S(n6690), .Z(n9204)
         );
  INV_X1 U8375 ( .A(n6636), .ZN(n9203) );
  NAND2_X1 U8376 ( .A1(n9204), .A2(n9203), .ZN(n9202) );
  INV_X1 U8377 ( .A(n6690), .ZN(n9206) );
  NAND2_X1 U8378 ( .A1(n9206), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U8379 ( .A1(n9202), .A2(n6637), .ZN(n9216) );
  NAND2_X1 U8380 ( .A1(n9217), .A2(n9216), .ZN(n9215) );
  INV_X1 U8381 ( .A(n6685), .ZN(n9214) );
  NAND2_X1 U8382 ( .A1(n9214), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U8383 ( .A1(n9215), .A2(n6638), .ZN(n9230) );
  XNOR2_X1 U8384 ( .A(n6695), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U8385 ( .A1(n9230), .A2(n9231), .ZN(n9229) );
  INV_X1 U8386 ( .A(n6695), .ZN(n9228) );
  NAND2_X1 U8387 ( .A1(n9228), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U8388 ( .A1(n9229), .A2(n6639), .ZN(n6644) );
  INV_X1 U8389 ( .A(n6640), .ZN(n6641) );
  NAND2_X1 U8390 ( .A1(n6642), .A2(n6641), .ZN(n6649) );
  INV_X1 U8391 ( .A(n6649), .ZN(n6739) );
  NOR2_X1 U8392 ( .A1(n6459), .A2(n6612), .ZN(n6643) );
  NAND2_X1 U8393 ( .A1(n6644), .A2(n6645), .ZN(n6755) );
  OAI211_X1 U8394 ( .C1(n6645), .C2(n6644), .A(n9716), .B(n6755), .ZN(n6646)
         );
  NAND2_X1 U8395 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n8850) );
  OAI211_X1 U8396 ( .C1(n9724), .C2(n6647), .A(n6646), .B(n8850), .ZN(n6659)
         );
  XNOR2_X1 U8397 ( .A(n6742), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6656) );
  INV_X1 U8398 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6650) );
  MUX2_X1 U8399 ( .A(n6650), .B(P1_REG1_REG_2__SCAN_IN), .S(n6685), .Z(n9220)
         );
  INV_X1 U8400 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6651) );
  MUX2_X1 U8401 ( .A(n6651), .B(P1_REG1_REG_1__SCAN_IN), .S(n6690), .Z(n9201)
         );
  AND2_X1 U8402 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9200) );
  NAND2_X1 U8403 ( .A1(n9206), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U8404 ( .A1(n9199), .A2(n6652), .ZN(n9219) );
  NAND2_X1 U8405 ( .A1(n9220), .A2(n9219), .ZN(n9218) );
  NAND2_X1 U8406 ( .A1(n9214), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U8407 ( .A1(n9218), .A2(n6653), .ZN(n9233) );
  XNOR2_X1 U8408 ( .A(n6695), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U8409 ( .A1(n9233), .A2(n9234), .ZN(n9232) );
  NAND2_X1 U8410 ( .A1(n9228), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U8411 ( .A1(n9232), .A2(n6654), .ZN(n6655) );
  NAND2_X1 U8412 ( .A1(n6655), .A2(n6656), .ZN(n6743) );
  OAI21_X1 U8413 ( .B1(n6656), .B2(n6655), .A(n6743), .ZN(n6657) );
  OAI22_X1 U8414 ( .A1(n6742), .A2(n9668), .B1(n9709), .B2(n6657), .ZN(n6658)
         );
  OR3_X1 U8415 ( .A1(n6660), .A2(n6659), .A3(n6658), .ZN(P1_U3247) );
  AOI211_X1 U8416 ( .C1(n6662), .C2(n7050), .A(n9807), .B(n6661), .ZN(n6674)
         );
  NOR2_X1 U8417 ( .A1(n8139), .A2(n4504), .ZN(n6673) );
  XNOR2_X1 U8418 ( .A(n6663), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6665) );
  INV_X1 U8419 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6664) );
  OAI22_X1 U8420 ( .A1(n9853), .A2(n6665), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6664), .ZN(n6672) );
  INV_X1 U8421 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6670) );
  AOI21_X1 U8422 ( .B1(n6668), .B2(n6667), .A(n6666), .ZN(n6669) );
  OAI22_X1 U8423 ( .A1(n9805), .A2(n6670), .B1(n9844), .B2(n6669), .ZN(n6671)
         );
  OR4_X1 U8424 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(P2_U3183)
         );
  NAND2_X1 U8425 ( .A1(n4325), .A2(P2_U3151), .ZN(n8565) );
  NOR2_X1 U8426 ( .A1(n4325), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8559) );
  OAI222_X1 U8427 ( .A1(n8565), .A2(n4732), .B1(n8568), .B2(n6691), .C1(
        P2_U3151), .C2(n4504), .ZN(P2_U3294) );
  INV_X1 U8428 ( .A(n9613), .ZN(n9623) );
  OAI222_X1 U8429 ( .A1(n6742), .A2(P1_U3086), .B1(n9626), .B2(n6676), .C1(
        n6675), .C2(n9623), .ZN(P1_U3351) );
  INV_X1 U8430 ( .A(n8565), .ZN(n8562) );
  INV_X1 U8431 ( .A(n8562), .ZN(n8555) );
  OAI222_X1 U8432 ( .A1(n8555), .A2(n6677), .B1(n8568), .B2(n6676), .C1(
        P2_U3151), .C2(n7190), .ZN(P2_U3291) );
  OAI222_X1 U8433 ( .A1(n8555), .A2(n6679), .B1(n8568), .B2(n6689), .C1(
        P2_U3151), .C2(n6678), .ZN(P2_U3290) );
  OAI222_X1 U8434 ( .A1(n8555), .A2(n6680), .B1(n8568), .B2(n6686), .C1(
        P2_U3151), .C2(n9800), .ZN(P2_U3293) );
  OAI222_X1 U8435 ( .A1(n8555), .A2(n6681), .B1(n8568), .B2(n6694), .C1(
        P2_U3151), .C2(n6979), .ZN(P2_U3292) );
  OAI222_X1 U8436 ( .A1(n8555), .A2(n6682), .B1(n8568), .B2(n6684), .C1(
        P2_U3151), .C2(n7402), .ZN(P2_U3289) );
  OAI222_X1 U8437 ( .A1(n6746), .A2(P1_U3086), .B1(n9626), .B2(n6684), .C1(
        n6683), .C2(n9623), .ZN(P1_U3349) );
  INV_X1 U8438 ( .A(n9626), .ZN(n7556) );
  INV_X1 U8439 ( .A(n7556), .ZN(n9620) );
  OAI222_X1 U8440 ( .A1(n9623), .A2(n6687), .B1(n9620), .B2(n6686), .C1(n6685), 
        .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U8441 ( .A1(n6745), .A2(P1_U3086), .B1(n9620), .B2(n6689), .C1(
        n6688), .C2(n9623), .ZN(P1_U3350) );
  OAI222_X1 U8442 ( .A1(n9623), .A2(n6692), .B1(n9620), .B2(n6691), .C1(n6690), 
        .C2(P1_U3086), .ZN(P1_U3354) );
  OAI222_X1 U8443 ( .A1(n6695), .A2(P1_U3086), .B1(n9620), .B2(n6694), .C1(
        n6693), .C2(n9623), .ZN(P1_U3352) );
  OAI222_X1 U8444 ( .A1(n6747), .A2(P1_U3086), .B1(n9620), .B2(n6698), .C1(
        n6696), .C2(n9623), .ZN(P1_U3348) );
  OAI222_X1 U8445 ( .A1(n8555), .A2(n6699), .B1(n8568), .B2(n6698), .C1(
        P2_U3151), .C2(n6697), .ZN(P2_U3288) );
  AOI22_X1 U8446 ( .A1(n6813), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9613), .ZN(n6700) );
  OAI21_X1 U8447 ( .B1(n6702), .B2(n9620), .A(n6700), .ZN(P1_U3347) );
  OAI222_X1 U8448 ( .A1(n8555), .A2(n6703), .B1(n8568), .B2(n6702), .C1(
        P2_U3151), .C2(n6701), .ZN(P2_U3287) );
  INV_X1 U8449 ( .A(n6704), .ZN(n6707) );
  AOI22_X1 U8450 ( .A1(n6995), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9613), .ZN(n6705) );
  OAI21_X1 U8451 ( .B1(n6707), .B2(n9626), .A(n6705), .ZN(P1_U3346) );
  OAI222_X1 U8452 ( .A1(n8568), .A2(n6707), .B1(n7735), .B2(P2_U3151), .C1(
        n6706), .C2(n8555), .ZN(P2_U3286) );
  INV_X1 U8453 ( .A(n9724), .ZN(n9205) );
  NOR2_X1 U8454 ( .A1(n9205), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8455 ( .A1(n6720), .A2(n6708), .ZN(n6709) );
  OAI21_X1 U8456 ( .B1(n6720), .B2(n6710), .A(n6709), .ZN(P2_U3377) );
  INV_X1 U8457 ( .A(n6711), .ZN(n6713) );
  OAI222_X1 U8458 ( .A1(n8568), .A2(n6713), .B1(n7794), .B2(P2_U3151), .C1(
        n6712), .C2(n8555), .ZN(P2_U3285) );
  INV_X1 U8459 ( .A(n9637), .ZN(n6714) );
  OAI222_X1 U8460 ( .A1(P1_U3086), .A2(n6714), .B1(n9620), .B2(n6713), .C1(
        n10120), .C2(n9623), .ZN(P1_U3345) );
  INV_X1 U8461 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U8462 ( .A1(n8822), .A2(P1_U3973), .ZN(n6715) );
  OAI21_X1 U8463 ( .B1(n10087), .B2(P1_U3973), .A(n6715), .ZN(P1_U3572) );
  INV_X1 U8464 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7253) );
  NAND2_X1 U8465 ( .A1(n8854), .A2(P1_U3973), .ZN(n6716) );
  OAI21_X1 U8466 ( .B1(n7253), .B2(P1_U3973), .A(n6716), .ZN(P1_U3573) );
  INV_X1 U8467 ( .A(n9060), .ZN(n9094) );
  NAND2_X1 U8468 ( .A1(n9094), .A2(P1_U3973), .ZN(n6717) );
  OAI21_X1 U8469 ( .B1(P1_U3973), .B2(n8556), .A(n6717), .ZN(P1_U3585) );
  INV_X1 U8470 ( .A(n6718), .ZN(n6719) );
  AND2_X1 U8471 ( .A1(n6729), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8472 ( .A1(n6729), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8473 ( .A1(n6729), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8474 ( .A1(n6729), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8475 ( .A1(n6729), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8476 ( .A1(n6729), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8477 ( .A1(n6729), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8478 ( .A1(n6729), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8479 ( .A1(n6729), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8480 ( .A1(n6729), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8481 ( .A1(n6729), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8482 ( .A1(n6729), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8483 ( .A1(n6729), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8484 ( .A1(n6729), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8485 ( .A1(n6729), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8486 ( .A1(n6729), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8487 ( .A1(n6729), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8488 ( .A1(n6729), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8489 ( .A1(n6729), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8490 ( .A1(n6729), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8491 ( .A1(n6729), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8492 ( .A1(n6729), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8493 ( .A1(n6729), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8494 ( .A1(n6729), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8495 ( .A1(n6729), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  INV_X1 U8496 ( .A(n6721), .ZN(n6727) );
  AOI22_X1 U8497 ( .A1(n9655), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9613), .ZN(n6722) );
  OAI21_X1 U8498 ( .B1(n6727), .B2(n9626), .A(n6722), .ZN(P1_U3344) );
  INV_X1 U8499 ( .A(n6723), .ZN(n6843) );
  INV_X1 U8500 ( .A(n6724), .ZN(n6725) );
  AOI22_X1 U8501 ( .A1(n6729), .A2(n6726), .B1(n6843), .B2(n6725), .ZN(
        P2_U3376) );
  OAI222_X1 U8502 ( .A1(n8555), .A2(n6728), .B1(n8568), .B2(n6727), .C1(
        P2_U3151), .C2(n7807), .ZN(P2_U3284) );
  INV_X1 U8503 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U8504 ( .A1(n6731), .A2(n10130), .ZN(P2_U3262) );
  INV_X1 U8505 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9988) );
  NOR2_X1 U8506 ( .A1(n6731), .A2(n9988), .ZN(P2_U3258) );
  INV_X1 U8507 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10102) );
  NOR2_X1 U8508 ( .A1(n6731), .A2(n10102), .ZN(P2_U3263) );
  INV_X1 U8509 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6730) );
  NOR2_X1 U8510 ( .A1(n6731), .A2(n6730), .ZN(P2_U3261) );
  INV_X1 U8511 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10147) );
  NOR2_X1 U8512 ( .A1(n6731), .A2(n10147), .ZN(P2_U3243) );
  AOI21_X1 U8513 ( .B1(n6625), .B2(n6612), .A(n6733), .ZN(n6732) );
  MUX2_X1 U8514 ( .A(n6733), .B(n6732), .S(n6735), .Z(n6738) );
  INV_X1 U8515 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6734) );
  INV_X1 U8516 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6842) );
  OAI22_X1 U8517 ( .A1(n9724), .A2(n6734), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6842), .ZN(n6737) );
  NOR3_X1 U8518 ( .A1(n9709), .A2(n6735), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6736) );
  AOI211_X1 U8519 ( .C1(n6739), .C2(n6738), .A(n6737), .B(n6736), .ZN(n6740)
         );
  INV_X1 U8520 ( .A(n6740), .ZN(P1_U3243) );
  NOR2_X1 U8521 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6995), .ZN(n6741) );
  AOI21_X1 U8522 ( .B1(n6995), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6741), .ZN(
        n6749) );
  INV_X1 U8523 ( .A(n6747), .ZN(n6784) );
  INV_X1 U8524 ( .A(n6746), .ZN(n6771) );
  INV_X1 U8525 ( .A(n6745), .ZN(n6797) );
  INV_X1 U8526 ( .A(n6742), .ZN(n6757) );
  INV_X1 U8527 ( .A(n6743), .ZN(n6744) );
  XOR2_X1 U8528 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6745), .Z(n6795) );
  NOR2_X1 U8529 ( .A1(n6796), .A2(n6795), .ZN(n6794) );
  AOI21_X1 U8530 ( .B1(n6797), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6794), .ZN(
        n6770) );
  XOR2_X1 U8531 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6746), .Z(n6769) );
  NOR2_X1 U8532 ( .A1(n6770), .A2(n6769), .ZN(n6768) );
  XOR2_X1 U8533 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6747), .Z(n6782) );
  NOR2_X1 U8534 ( .A1(n6783), .A2(n6782), .ZN(n6781) );
  AOI21_X1 U8535 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6784), .A(n6781), .ZN(
        n6809) );
  XNOR2_X1 U8536 ( .A(n6813), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6808) );
  NOR2_X1 U8537 ( .A1(n6809), .A2(n6808), .ZN(n6807) );
  NAND2_X1 U8538 ( .A1(n6748), .A2(n6749), .ZN(n6984) );
  OAI21_X1 U8539 ( .B1(n6749), .B2(n6748), .A(n6984), .ZN(n6753) );
  INV_X1 U8540 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6751) );
  INV_X1 U8541 ( .A(n9668), .ZN(n9712) );
  NAND2_X1 U8542 ( .A1(n9712), .A2(n6995), .ZN(n6750) );
  NAND2_X1 U8543 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7683) );
  OAI211_X1 U8544 ( .C1(n9724), .C2(n6751), .A(n6750), .B(n7683), .ZN(n6752)
         );
  AOI21_X1 U8545 ( .B1(n6753), .B2(n9660), .A(n6752), .ZN(n6762) );
  NOR2_X1 U8546 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6995), .ZN(n6754) );
  AOI21_X1 U8547 ( .B1(n6995), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6754), .ZN(
        n6759) );
  INV_X1 U8548 ( .A(n6755), .ZN(n6756) );
  XNOR2_X1 U8549 ( .A(n6797), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6792) );
  NOR2_X1 U8550 ( .A1(n6793), .A2(n6792), .ZN(n6791) );
  AOI21_X1 U8551 ( .B1(n6797), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6791), .ZN(
        n6767) );
  XNOR2_X1 U8552 ( .A(n6771), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6766) );
  NOR2_X1 U8553 ( .A1(n6767), .A2(n6766), .ZN(n6765) );
  XNOR2_X1 U8554 ( .A(n6784), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6779) );
  NOR2_X1 U8555 ( .A1(n6780), .A2(n6779), .ZN(n6778) );
  AOI21_X1 U8556 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6784), .A(n6778), .ZN(
        n6812) );
  XNOR2_X1 U8557 ( .A(n6813), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6811) );
  NOR2_X1 U8558 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  NAND2_X1 U8559 ( .A1(n6758), .A2(n6759), .ZN(n6994) );
  OAI21_X1 U8560 ( .B1(n6759), .B2(n6758), .A(n6994), .ZN(n6760) );
  NAND2_X1 U8561 ( .A1(n6760), .A2(n9716), .ZN(n6761) );
  NAND2_X1 U8562 ( .A1(n6762), .A2(n6761), .ZN(P1_U3252) );
  INV_X1 U8563 ( .A(n6763), .ZN(n6804) );
  OAI222_X1 U8564 ( .A1(n8568), .A2(n6804), .B1(n6764), .B2(P2_U3151), .C1(
        n10105), .C2(n8555), .ZN(P2_U3283) );
  AOI211_X1 U8565 ( .C1(n6767), .C2(n6766), .A(n6765), .B(n9700), .ZN(n6777)
         );
  AOI211_X1 U8566 ( .C1(n6770), .C2(n6769), .A(n6768), .B(n9709), .ZN(n6776)
         );
  INV_X1 U8567 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U8568 ( .A1(n9712), .A2(n6771), .ZN(n6773) );
  NAND2_X1 U8569 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6772) );
  OAI211_X1 U8570 ( .C1(n6774), .C2(n9724), .A(n6773), .B(n6772), .ZN(n6775)
         );
  OR3_X1 U8571 ( .A1(n6777), .A2(n6776), .A3(n6775), .ZN(P1_U3249) );
  AOI211_X1 U8572 ( .C1(n6780), .C2(n6779), .A(n9700), .B(n6778), .ZN(n6790)
         );
  AOI211_X1 U8573 ( .C1(n6783), .C2(n6782), .A(n9709), .B(n6781), .ZN(n6789)
         );
  INV_X1 U8574 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U8575 ( .A1(n9712), .A2(n6784), .ZN(n6786) );
  NAND2_X1 U8576 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6785) );
  OAI211_X1 U8577 ( .C1(n6787), .C2(n9724), .A(n6786), .B(n6785), .ZN(n6788)
         );
  OR3_X1 U8578 ( .A1(n6790), .A2(n6789), .A3(n6788), .ZN(P1_U3250) );
  AOI211_X1 U8579 ( .C1(n6793), .C2(n6792), .A(n6791), .B(n9700), .ZN(n6802)
         );
  AOI211_X1 U8580 ( .C1(n6796), .C2(n6795), .A(n6794), .B(n9709), .ZN(n6801)
         );
  INV_X1 U8581 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8582 ( .A1(n9712), .A2(n6797), .ZN(n6798) );
  NAND2_X1 U8583 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7296) );
  OAI211_X1 U8584 ( .C1(n6799), .C2(n9724), .A(n6798), .B(n7296), .ZN(n6800)
         );
  OR3_X1 U8585 ( .A1(n6802), .A2(n6801), .A3(n6800), .ZN(P1_U3248) );
  INV_X1 U8586 ( .A(n7710), .ZN(n6989) );
  OAI222_X1 U8587 ( .A1(P1_U3086), .A2(n6989), .B1(n9620), .B2(n6804), .C1(
        n6803), .C2(n9623), .ZN(P1_U3343) );
  INV_X1 U8588 ( .A(n6805), .ZN(n6822) );
  AOI22_X1 U8589 ( .A1(n9681), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9613), .ZN(n6806) );
  OAI21_X1 U8590 ( .B1(n6822), .B2(n9626), .A(n6806), .ZN(P1_U3342) );
  AOI211_X1 U8591 ( .C1(n6809), .C2(n6808), .A(n9709), .B(n6807), .ZN(n6819)
         );
  AOI211_X1 U8592 ( .C1(n6812), .C2(n6811), .A(n9700), .B(n6810), .ZN(n6818)
         );
  INV_X1 U8593 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U8594 ( .A1(n9712), .A2(n6813), .ZN(n6815) );
  NAND2_X1 U8595 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n6814) );
  OAI211_X1 U8596 ( .C1(n6816), .C2(n9724), .A(n6815), .B(n6814), .ZN(n6817)
         );
  OR3_X1 U8597 ( .A1(n6819), .A2(n6818), .A3(n6817), .ZN(P1_U3251) );
  NAND2_X1 U8598 ( .A1(n8073), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n6820) );
  OAI21_X1 U8599 ( .B1(n8362), .B2(n8073), .A(n6820), .ZN(P2_U3506) );
  INV_X1 U8600 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6823) );
  OAI222_X1 U8601 ( .A1(n8555), .A2(n6823), .B1(n8568), .B2(n6822), .C1(
        P2_U3151), .C2(n6821), .ZN(P2_U3282) );
  NAND2_X1 U8602 ( .A1(n9608), .A2(n6824), .ZN(n6830) );
  NOR2_X1 U8603 ( .A1(n9103), .A2(P1_U3086), .ZN(n7368) );
  OAI22_X1 U8604 ( .A1(n6830), .A2(n7066), .B1(n7368), .B2(n9787), .ZN(n6826)
         );
  NAND2_X1 U8605 ( .A1(n6826), .A2(n6825), .ZN(n6966) );
  NOR2_X1 U8606 ( .A1(n6966), .A2(P1_U3086), .ZN(n6907) );
  INV_X1 U8607 ( .A(n7066), .ZN(n6829) );
  AND2_X1 U8608 ( .A1(n6827), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6828) );
  NAND2_X1 U8609 ( .A1(n6829), .A2(n9771), .ZN(n9769) );
  OR2_X1 U8610 ( .A1(n6830), .A2(n9769), .ZN(n6839) );
  OR2_X1 U8611 ( .A1(n9546), .A2(n6831), .ZN(n6832) );
  NAND2_X1 U8612 ( .A1(n6833), .A2(n8905), .ZN(n6841) );
  NOR2_X1 U8613 ( .A1(n6856), .A2(n8907), .ZN(n9471) );
  INV_X1 U8614 ( .A(n6839), .ZN(n6834) );
  NAND2_X1 U8615 ( .A1(n6836), .A2(n6835), .ZN(n7072) );
  INV_X1 U8616 ( .A(n6837), .ZN(n6838) );
  AOI22_X1 U8617 ( .A1(n9471), .A2(n8895), .B1(n9473), .B2(n9650), .ZN(n6840)
         );
  OAI211_X1 U8618 ( .C1(n6907), .C2(n6842), .A(n6841), .B(n6840), .ZN(P1_U3232) );
  NAND2_X1 U8619 ( .A1(n6844), .A2(n6843), .ZN(n6911) );
  NAND2_X1 U8620 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n6911), .ZN(n6847) );
  NAND2_X1 U8621 ( .A1(n8030), .A2(n6845), .ZN(n6846) );
  OAI211_X1 U8622 ( .C1(n6509), .C2(n8052), .A(n6847), .B(n6846), .ZN(n6848)
         );
  AOI21_X1 U8623 ( .B1(n7032), .B2(n5886), .A(n6848), .ZN(n6849) );
  INV_X1 U8624 ( .A(n6849), .ZN(P2_U3172) );
  INV_X1 U8625 ( .A(n6850), .ZN(n6868) );
  AOI22_X1 U8626 ( .A1(n9693), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9613), .ZN(n6851) );
  OAI21_X1 U8627 ( .B1(n6868), .B2(n9626), .A(n6851), .ZN(P1_U3341) );
  INV_X1 U8628 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U8629 ( .A1(n6890), .A2(n6895), .ZN(n6858) );
  OAI21_X1 U8630 ( .B1(n6861), .B2(n6860), .A(n6902), .ZN(n6862) );
  NAND2_X1 U8631 ( .A1(n6862), .A2(n8905), .ZN(n6867) );
  OR2_X1 U8632 ( .A1(n6938), .A2(n8907), .ZN(n6865) );
  NAND2_X1 U8633 ( .A1(n6863), .A2(n9167), .ZN(n6864) );
  NAND2_X1 U8634 ( .A1(n6865), .A2(n6864), .ZN(n6885) );
  AOI22_X1 U8635 ( .A1(n6885), .A2(n8895), .B1(n9650), .B2(n6890), .ZN(n6866)
         );
  OAI211_X1 U8636 ( .C1(n6907), .C2(n7073), .A(n6867), .B(n6866), .ZN(P1_U3222) );
  INV_X1 U8637 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6869) );
  OAI222_X1 U8638 ( .A1(n8565), .A2(n6869), .B1(n8568), .B2(n6868), .C1(
        P2_U3151), .C2(n8085), .ZN(P2_U3281) );
  INV_X1 U8639 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6874) );
  INV_X1 U8640 ( .A(n9471), .ZN(n6871) );
  NAND2_X1 U8641 ( .A1(n6863), .A2(n6872), .ZN(n9106) );
  NAND2_X1 U8642 ( .A1(n6881), .A2(n9106), .ZN(n9469) );
  OAI21_X1 U8643 ( .B1(n9729), .B2(n9791), .A(n9469), .ZN(n6870) );
  OAI211_X1 U8644 ( .C1(n9468), .C2(n6872), .A(n6871), .B(n6870), .ZN(n6875)
         );
  NAND2_X1 U8645 ( .A1(n6875), .A2(n9793), .ZN(n6873) );
  OAI21_X1 U8646 ( .B1(n9793), .B2(n6874), .A(n6873), .ZN(P1_U3453) );
  NAND2_X1 U8647 ( .A1(n6875), .A2(n9799), .ZN(n6876) );
  OAI21_X1 U8648 ( .B1(n9799), .B2(n6625), .A(n6876), .ZN(P1_U3522) );
  INV_X1 U8649 ( .A(n7511), .ZN(n7551) );
  OR2_X1 U8650 ( .A1(n6419), .A2(n6877), .ZN(n6878) );
  NAND2_X1 U8651 ( .A1(n6879), .A2(n6878), .ZN(n7080) );
  NAND2_X1 U8652 ( .A1(n6890), .A2(n9473), .ZN(n6880) );
  AND3_X1 U8653 ( .A1(n6926), .A2(n9505), .A3(n6880), .ZN(n7075) );
  INV_X1 U8654 ( .A(n7491), .ZN(n7508) );
  NAND2_X1 U8655 ( .A1(n7080), .A2(n7508), .ZN(n6888) );
  NAND2_X1 U8656 ( .A1(n6419), .A2(n6881), .ZN(n6882) );
  NAND2_X1 U8657 ( .A1(n6883), .A2(n6882), .ZN(n6884) );
  NAND2_X1 U8658 ( .A1(n6884), .A2(n9729), .ZN(n6887) );
  INV_X1 U8659 ( .A(n6885), .ZN(n6886) );
  NAND3_X1 U8660 ( .A1(n6888), .A2(n6887), .A3(n6886), .ZN(n7069) );
  AOI211_X1 U8661 ( .C1(n7551), .C2(n7080), .A(n7075), .B(n7069), .ZN(n6892)
         );
  AOI22_X1 U8662 ( .A1(n9604), .A2(n6890), .B1(n6614), .B2(
        P1_REG0_REG_1__SCAN_IN), .ZN(n6889) );
  OAI21_X1 U8663 ( .B1(n6892), .B2(n6614), .A(n6889), .ZN(P1_U3456) );
  AOI22_X1 U8664 ( .A1(n9553), .A2(n6890), .B1(n4846), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6891) );
  OAI21_X1 U8665 ( .B1(n6892), .B2(n4846), .A(n6891), .ZN(P1_U3523) );
  INV_X1 U8666 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9211) );
  INV_X1 U8667 ( .A(n6893), .ZN(n6901) );
  XNOR2_X1 U8668 ( .A(n6894), .B(n8761), .ZN(n6899) );
  OR2_X1 U8669 ( .A1(n6938), .A2(n8677), .ZN(n6897) );
  NAND2_X1 U8670 ( .A1(n6932), .A2(n6895), .ZN(n6896) );
  AND2_X1 U8671 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8672 ( .A1(n6899), .A2(n6898), .ZN(n6959) );
  AND3_X1 U8673 ( .A1(n6902), .A2(n6901), .A3(n6900), .ZN(n6903) );
  OAI21_X1 U8674 ( .B1(n6960), .B2(n6903), .A(n8905), .ZN(n6906) );
  OAI22_X1 U8675 ( .A1(n6904), .A2(n8907), .B1(n6856), .B2(n9276), .ZN(n6928)
         );
  AOI22_X1 U8676 ( .A1(n6928), .A2(n8895), .B1(n6932), .B2(n9650), .ZN(n6905)
         );
  OAI211_X1 U8677 ( .C1(n6907), .C2(n9211), .A(n6906), .B(n6905), .ZN(P1_U3237) );
  INV_X1 U8678 ( .A(n6908), .ZN(n6923) );
  OAI222_X1 U8679 ( .A1(n8568), .A2(n6923), .B1(n6910), .B2(P2_U3151), .C1(
        n6909), .C2(n8555), .ZN(P2_U3280) );
  INV_X1 U8680 ( .A(n6911), .ZN(n6958) );
  OAI21_X1 U8681 ( .B1(n6914), .B2(n6913), .A(n6912), .ZN(n6915) );
  NAND2_X1 U8682 ( .A1(n6915), .A2(n5886), .ZN(n6918) );
  OAI22_X1 U8683 ( .A1(n5789), .A2(n8052), .B1(n8058), .B2(n7011), .ZN(n6916)
         );
  AOI21_X1 U8684 ( .B1(n8038), .B2(n8078), .A(n6916), .ZN(n6917) );
  OAI211_X1 U8685 ( .C1(n6958), .C2(n6664), .A(n6918), .B(n6917), .ZN(P2_U3162) );
  INV_X1 U8686 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6921) );
  INV_X1 U8687 ( .A(n9880), .ZN(n9902) );
  OAI21_X1 U8688 ( .B1(n8392), .B2(n9915), .A(n7032), .ZN(n6919) );
  NAND2_X1 U8689 ( .A1(n8077), .A2(n8375), .ZN(n7035) );
  OAI211_X1 U8690 ( .C1(n9893), .C2(n7041), .A(n6919), .B(n7035), .ZN(n8463)
         );
  NAND2_X1 U8691 ( .A1(n8463), .A2(n9919), .ZN(n6920) );
  OAI21_X1 U8692 ( .B1(n6921), .B2(n9919), .A(n6920), .ZN(P2_U3390) );
  OAI222_X1 U8693 ( .A1(P1_U3086), .A2(n7713), .B1(n9620), .B2(n6923), .C1(
        n6922), .C2(n9623), .ZN(P1_U3340) );
  OAI21_X1 U8694 ( .B1(n6925), .B2(n9033), .A(n6924), .ZN(n7084) );
  AOI211_X1 U8695 ( .C1(n6932), .C2(n6926), .A(n9736), .B(n6940), .ZN(n7089)
         );
  XNOR2_X1 U8696 ( .A(n6927), .B(n9033), .ZN(n6930) );
  INV_X1 U8697 ( .A(n6928), .ZN(n6929) );
  OAI21_X1 U8698 ( .B1(n6930), .B2(n9425), .A(n6929), .ZN(n7085) );
  AOI211_X1 U8699 ( .C1(n9791), .C2(n7084), .A(n7089), .B(n7085), .ZN(n6934)
         );
  AOI22_X1 U8700 ( .A1(n9604), .A2(n6932), .B1(n6614), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n6931) );
  OAI21_X1 U8701 ( .B1(n6934), .B2(n6614), .A(n6931), .ZN(P1_U3459) );
  AOI22_X1 U8702 ( .A1(n9553), .A2(n6932), .B1(n4846), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6933) );
  OAI21_X1 U8703 ( .B1(n6934), .B2(n4846), .A(n6933), .ZN(P1_U3524) );
  INV_X1 U8704 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6944) );
  OAI21_X1 U8705 ( .B1(n6936), .B2(n9034), .A(n6935), .ZN(n7196) );
  INV_X1 U8706 ( .A(n7196), .ZN(n6941) );
  XNOR2_X1 U8707 ( .A(n6937), .B(n9034), .ZN(n6939) );
  OAI22_X1 U8708 ( .A1(n7279), .A2(n8907), .B1(n6938), .B2(n9276), .ZN(n6967)
         );
  AOI21_X1 U8709 ( .B1(n6939), .B2(n9729), .A(n6967), .ZN(n7198) );
  OAI211_X1 U8710 ( .C1(n6940), .C2(n6961), .A(n7017), .B(n9505), .ZN(n7194)
         );
  OAI211_X1 U8711 ( .C1(n9509), .C2(n6941), .A(n7198), .B(n7194), .ZN(n6945)
         );
  NAND2_X1 U8712 ( .A1(n6945), .A2(n9793), .ZN(n6943) );
  NAND2_X1 U8713 ( .A1(n9604), .A2(n7191), .ZN(n6942) );
  OAI211_X1 U8714 ( .C1(n9793), .C2(n6944), .A(n6943), .B(n6942), .ZN(P1_U3462) );
  INV_X1 U8715 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U8716 ( .A1(n6945), .A2(n9799), .ZN(n6947) );
  NAND2_X1 U8717 ( .A1(n9553), .A2(n7191), .ZN(n6946) );
  OAI211_X1 U8718 ( .C1(n9799), .C2(n6948), .A(n6947), .B(n6946), .ZN(P1_U3525) );
  INV_X1 U8719 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6957) );
  OAI21_X1 U8720 ( .B1(n6951), .B2(n6950), .A(n6949), .ZN(n6952) );
  NAND2_X1 U8721 ( .A1(n6952), .A2(n5886), .ZN(n6956) );
  OAI22_X1 U8722 ( .A1(n7210), .A2(n8052), .B1(n8058), .B2(n6953), .ZN(n6954)
         );
  AOI21_X1 U8723 ( .B1(n8038), .B2(n8077), .A(n6954), .ZN(n6955) );
  OAI211_X1 U8724 ( .C1(n6958), .C2(n6957), .A(n6956), .B(n6955), .ZN(P2_U3177) );
  NAND2_X1 U8725 ( .A1(n9196), .A2(n8758), .ZN(n6963) );
  OR2_X1 U8726 ( .A1(n6961), .A2(n8764), .ZN(n6962) );
  NAND2_X1 U8727 ( .A1(n6963), .A2(n6962), .ZN(n7275) );
  AOI22_X1 U8728 ( .A1(n6895), .A2(n9196), .B1(n7191), .B2(n8709), .ZN(n6964)
         );
  XNOR2_X1 U8729 ( .A(n6964), .B(n8695), .ZN(n7274) );
  XOR2_X1 U8730 ( .A(n7275), .B(n7274), .Z(n6965) );
  AOI22_X1 U8731 ( .A1(n9650), .A2(n7191), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n6969) );
  AOI22_X1 U8732 ( .A1(n6967), .A2(n8895), .B1(n8929), .B2(n6086), .ZN(n6968)
         );
  OAI211_X1 U8733 ( .C1(n6970), .C2(n9646), .A(n6969), .B(n6968), .ZN(P1_U3218) );
  OAI21_X1 U8734 ( .B1(n6973), .B2(n6972), .A(n6971), .ZN(n6981) );
  AOI22_X1 U8735 ( .A1(n9835), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n6975), .B2(
        n6974), .ZN(n6978) );
  OAI21_X1 U8736 ( .B1(n4441), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7176), .ZN(
        n6976) );
  AND2_X1 U8737 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7047) );
  AOI21_X1 U8738 ( .B1(n9815), .B2(n6976), .A(n7047), .ZN(n6977) );
  OAI211_X1 U8739 ( .C1(n6979), .C2(n8139), .A(n6978), .B(n6977), .ZN(n6980)
         );
  AOI21_X1 U8740 ( .B1(n6981), .B2(n9849), .A(n6980), .ZN(n6982) );
  INV_X1 U8741 ( .A(n6982), .ZN(P2_U3185) );
  INV_X1 U8742 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6983) );
  MUX2_X1 U8743 ( .A(n6983), .B(P1_REG1_REG_10__SCAN_IN), .S(n9637), .Z(n9633)
         );
  NOR2_X1 U8744 ( .A1(n9633), .A2(n9634), .ZN(n9632) );
  INV_X1 U8745 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6985) );
  MUX2_X1 U8746 ( .A(n6985), .B(P1_REG1_REG_11__SCAN_IN), .S(n9655), .Z(n9658)
         );
  NOR2_X1 U8747 ( .A1(n9657), .A2(n9658), .ZN(n9656) );
  AOI21_X1 U8748 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9655), .A(n9656), .ZN(
        n6987) );
  INV_X1 U8749 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U8750 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7710), .B1(n6989), .B2(
        n9797), .ZN(n6986) );
  NAND2_X1 U8751 ( .A1(n6987), .A2(n6986), .ZN(n7704) );
  OAI21_X1 U8752 ( .B1(n6987), .B2(n6986), .A(n7704), .ZN(n6991) );
  NAND2_X1 U8753 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U8754 ( .A1(n9205), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6988) );
  OAI211_X1 U8755 ( .C1(n9668), .C2(n6989), .A(n8794), .B(n6988), .ZN(n6990)
         );
  AOI21_X1 U8756 ( .B1(n6991), .B2(n9660), .A(n6990), .ZN(n7001) );
  NOR2_X1 U8757 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7710), .ZN(n6992) );
  AOI21_X1 U8758 ( .B1(n7710), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6992), .ZN(
        n6998) );
  NAND2_X1 U8759 ( .A1(n9637), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6993) );
  OAI21_X1 U8760 ( .B1(n9637), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6993), .ZN(
        n9630) );
  NOR2_X1 U8761 ( .A1(n9630), .A2(n9631), .ZN(n9629) );
  NAND2_X1 U8762 ( .A1(n9655), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6996) );
  OAI21_X1 U8763 ( .B1(n9655), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6996), .ZN(
        n9663) );
  NOR2_X1 U8764 ( .A1(n9662), .A2(n9663), .ZN(n9661) );
  AOI21_X1 U8765 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9655), .A(n9661), .ZN(
        n6997) );
  NAND2_X1 U8766 ( .A1(n6998), .A2(n6997), .ZN(n7709) );
  OAI21_X1 U8767 ( .B1(n6998), .B2(n6997), .A(n7709), .ZN(n6999) );
  NAND2_X1 U8768 ( .A1(n6999), .A2(n9716), .ZN(n7000) );
  NAND2_X1 U8769 ( .A1(n7001), .A2(n7000), .ZN(P1_U3255) );
  INV_X1 U8770 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7003) );
  INV_X1 U8771 ( .A(n7002), .ZN(n7004) );
  OAI222_X1 U8772 ( .A1(n8565), .A2(n7003), .B1(n8568), .B2(n7004), .C1(
        P2_U3151), .C2(n8120), .ZN(P2_U3279) );
  INV_X1 U8773 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7005) );
  INV_X1 U8774 ( .A(n7749), .ZN(n7707) );
  OAI222_X1 U8775 ( .A1(n9623), .A2(n7005), .B1(n9620), .B2(n7004), .C1(n7707), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  OAI21_X1 U8776 ( .B1(n4999), .B2(n4998), .A(n7007), .ZN(n7217) );
  XNOR2_X1 U8777 ( .A(n4999), .B(n7008), .ZN(n7009) );
  OAI222_X1 U8778 ( .A1(n8389), .A2(n5789), .B1(n8387), .B2(n4366), .C1(n8323), 
        .C2(n7009), .ZN(n7218) );
  AOI21_X1 U8779 ( .B1(n9915), .B2(n7217), .A(n7218), .ZN(n7059) );
  INV_X1 U8780 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7010) );
  OAI22_X1 U8781 ( .A1(n7011), .A2(n8543), .B1(n9919), .B2(n7010), .ZN(n7012)
         );
  INV_X1 U8782 ( .A(n7012), .ZN(n7013) );
  OAI21_X1 U8783 ( .B1(n7059), .B2(n9921), .A(n7013), .ZN(P2_U3393) );
  OAI21_X1 U8784 ( .B1(n7015), .B2(n7018), .A(n7014), .ZN(n7154) );
  INV_X1 U8785 ( .A(n7123), .ZN(n7016) );
  AOI211_X1 U8786 ( .C1(n8847), .C2(n7017), .A(n9736), .B(n7016), .ZN(n7150)
         );
  INV_X1 U8787 ( .A(n7018), .ZN(n9037) );
  XNOR2_X1 U8788 ( .A(n7019), .B(n9037), .ZN(n7023) );
  OR2_X1 U8789 ( .A1(n7097), .A2(n8907), .ZN(n7021) );
  NAND2_X1 U8790 ( .A1(n9196), .A2(n9167), .ZN(n7020) );
  NAND2_X1 U8791 ( .A1(n7021), .A2(n7020), .ZN(n8845) );
  INV_X1 U8792 ( .A(n8845), .ZN(n7022) );
  OAI21_X1 U8793 ( .B1(n7023), .B2(n9425), .A(n7022), .ZN(n7149) );
  AOI211_X1 U8794 ( .C1(n9791), .C2(n7154), .A(n7150), .B(n7149), .ZN(n7026)
         );
  AOI22_X1 U8795 ( .A1(n9604), .A2(n8847), .B1(n6614), .B2(
        P1_REG0_REG_4__SCAN_IN), .ZN(n7024) );
  OAI21_X1 U8796 ( .B1(n7026), .B2(n6614), .A(n7024), .ZN(P1_U3465) );
  AOI22_X1 U8797 ( .A1(n9553), .A2(n8847), .B1(n4846), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7025) );
  OAI21_X1 U8798 ( .B1(n7026), .B2(n4846), .A(n7025), .ZN(P1_U3526) );
  INV_X1 U8799 ( .A(n7027), .ZN(n7030) );
  NAND3_X1 U8800 ( .A1(n7030), .A2(n7029), .A3(n7028), .ZN(n7036) );
  INV_X1 U8801 ( .A(n7036), .ZN(n7203) );
  INV_X1 U8802 ( .A(n7031), .ZN(n8219) );
  INV_X1 U8803 ( .A(n7032), .ZN(n7034) );
  NOR3_X1 U8804 ( .A1(n7034), .A2(n7033), .A3(n9914), .ZN(n7038) );
  INV_X1 U8805 ( .A(n7035), .ZN(n7037) );
  OAI21_X1 U8806 ( .B1(n7038), .B2(n7037), .A(n8401), .ZN(n7040) );
  AOI22_X1 U8807 ( .A1(n8408), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n8396), .ZN(n7039) );
  OAI211_X1 U8808 ( .C1(n8403), .C2(n7041), .A(n7040), .B(n7039), .ZN(P2_U3233) );
  AOI21_X1 U8809 ( .B1(n7043), .B2(n7042), .A(n7983), .ZN(n7045) );
  NAND2_X1 U8810 ( .A1(n7045), .A2(n7044), .ZN(n7049) );
  OAI22_X1 U8811 ( .A1(n7261), .A2(n8052), .B1(n5789), .B2(n8049), .ZN(n7046)
         );
  AOI211_X1 U8812 ( .C1(n9865), .C2(n8030), .A(n7047), .B(n7046), .ZN(n7048)
         );
  OAI211_X1 U8813 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8040), .A(n7049), .B(
        n7048), .ZN(P2_U3158) );
  AOI21_X1 U8814 ( .B1(n7057), .B2(n7051), .A(n7050), .ZN(n7052) );
  AOI21_X1 U8815 ( .B1(n7053), .B2(n9807), .A(n7052), .ZN(n7054) );
  AOI21_X1 U8816 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n7054), .ZN(
        n7056) );
  NAND2_X1 U8817 ( .A1(n9835), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n7055) );
  OAI211_X1 U8818 ( .C1(n8139), .C2(n7057), .A(n7056), .B(n7055), .ZN(P2_U3182) );
  AOI22_X1 U8819 ( .A1(n6594), .A2(n5783), .B1(n9935), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7058) );
  OAI21_X1 U8820 ( .B1(n7059), .B2(n9935), .A(n7058), .ZN(P2_U3460) );
  INV_X1 U8821 ( .A(n7060), .ZN(n7063) );
  AOI22_X1 U8822 ( .A1(n9243), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9613), .ZN(n7061) );
  OAI21_X1 U8823 ( .B1(n7063), .B2(n9626), .A(n7061), .ZN(P1_U3338) );
  INV_X1 U8824 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7062) );
  OAI222_X1 U8825 ( .A1(n8568), .A2(n7063), .B1(n8138), .B2(P2_U3151), .C1(
        n7062), .C2(n8555), .ZN(P2_U3278) );
  INV_X1 U8826 ( .A(n7064), .ZN(n7119) );
  AOI22_X1 U8827 ( .A1(n9713), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9613), .ZN(n7065) );
  OAI21_X1 U8828 ( .B1(n7119), .B2(n9626), .A(n7065), .ZN(P1_U3337) );
  NOR2_X1 U8829 ( .A1(n9608), .A2(n7066), .ZN(n7067) );
  NAND2_X1 U8830 ( .A1(n7068), .A2(n7067), .ZN(n7074) );
  MUX2_X1 U8831 ( .A(n7069), .B(P1_REG2_REG_1__SCAN_IN), .S(n9767), .Z(n7070)
         );
  INV_X1 U8832 ( .A(n7070), .ZN(n7082) );
  INV_X1 U8833 ( .A(n7498), .ZN(n9749) );
  OR2_X1 U8834 ( .A1(n9401), .A2(n7073), .ZN(n7077) );
  NAND2_X1 U8835 ( .A1(n9754), .A2(n7075), .ZN(n7076) );
  OAI211_X1 U8836 ( .C1(n9760), .C2(n7078), .A(n7077), .B(n7076), .ZN(n7079)
         );
  AOI21_X1 U8837 ( .B1(n7080), .B2(n9749), .A(n7079), .ZN(n7081) );
  NAND2_X1 U8838 ( .A1(n7082), .A2(n7081), .ZN(P1_U3292) );
  OR2_X1 U8839 ( .A1(n9767), .A2(n7491), .ZN(n7083) );
  INV_X1 U8840 ( .A(n7084), .ZN(n7092) );
  INV_X1 U8841 ( .A(n7085), .ZN(n7086) );
  MUX2_X1 U8842 ( .A(n6634), .B(n7086), .S(n9470), .Z(n7091) );
  OAI22_X1 U8843 ( .A1(n9760), .A2(n7087), .B1(n9211), .B2(n9401), .ZN(n7088)
         );
  AOI21_X1 U8844 ( .B1(n7089), .B2(n9754), .A(n7088), .ZN(n7090) );
  OAI211_X1 U8845 ( .C1(n9466), .C2(n7092), .A(n7091), .B(n7090), .ZN(P1_U3291) );
  OR2_X1 U8846 ( .A1(n7093), .A2(n7096), .ZN(n7094) );
  NAND2_X1 U8847 ( .A1(n7095), .A2(n7094), .ZN(n7116) );
  INV_X1 U8848 ( .A(n7116), .ZN(n7107) );
  XNOR2_X1 U8849 ( .A(n7237), .B(n7096), .ZN(n7101) );
  OR2_X1 U8850 ( .A1(n7097), .A2(n9276), .ZN(n7099) );
  OR2_X1 U8851 ( .A1(n7501), .A2(n8907), .ZN(n7098) );
  NAND2_X1 U8852 ( .A1(n7099), .A2(n7098), .ZN(n7360) );
  INV_X1 U8853 ( .A(n7360), .ZN(n7100) );
  OAI21_X1 U8854 ( .B1(n7101), .B2(n9425), .A(n7100), .ZN(n7109) );
  NAND2_X1 U8855 ( .A1(n7109), .A2(n9470), .ZN(n7106) );
  INV_X1 U8856 ( .A(n7122), .ZN(n7102) );
  AOI211_X1 U8857 ( .C1(n7364), .C2(n7102), .A(n9736), .B(n7243), .ZN(n7108)
         );
  INV_X2 U8858 ( .A(n9401), .ZN(n9756) );
  AOI22_X1 U8859 ( .A1(n9767), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7359), .B2(
        n9756), .ZN(n7103) );
  OAI21_X1 U8860 ( .B1(n9760), .B2(n7354), .A(n7103), .ZN(n7104) );
  AOI21_X1 U8861 ( .B1(n7108), .B2(n9754), .A(n7104), .ZN(n7105) );
  OAI211_X1 U8862 ( .C1(n9466), .C2(n7107), .A(n7106), .B(n7105), .ZN(P1_U3287) );
  NOR2_X1 U8863 ( .A1(n7109), .A2(n7108), .ZN(n7118) );
  INV_X1 U8864 ( .A(n9555), .ZN(n7112) );
  INV_X1 U8865 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7110) );
  OAI22_X1 U8866 ( .A1(n6505), .A2(n7354), .B1(n9799), .B2(n7110), .ZN(n7111)
         );
  AOI21_X1 U8867 ( .B1(n7116), .B2(n7112), .A(n7111), .ZN(n7113) );
  OAI21_X1 U8868 ( .B1(n7118), .B2(n4846), .A(n7113), .ZN(P1_U3528) );
  INV_X1 U8869 ( .A(n9606), .ZN(n7115) );
  OAI22_X1 U8870 ( .A1(n6501), .A2(n7354), .B1(n9793), .B2(n6131), .ZN(n7114)
         );
  AOI21_X1 U8871 ( .B1(n7116), .B2(n7115), .A(n7114), .ZN(n7117) );
  OAI21_X1 U8872 ( .B1(n7118), .B2(n6614), .A(n7117), .ZN(P1_U3471) );
  OAI222_X1 U8873 ( .A1(n8568), .A2(n7119), .B1(n8555), .B2(n10087), .C1(
        P2_U3151), .C2(n8159), .ZN(P2_U3277) );
  OAI21_X1 U8874 ( .B1(n7121), .B2(n9039), .A(n7120), .ZN(n9763) );
  AOI211_X1 U8875 ( .C1(n7290), .C2(n7123), .A(n9736), .B(n7122), .ZN(n9755)
         );
  XNOR2_X1 U8876 ( .A(n7124), .B(n9039), .ZN(n7126) );
  OR2_X1 U8877 ( .A1(n7279), .A2(n9276), .ZN(n7125) );
  OAI21_X1 U8878 ( .B1(n7355), .B2(n8907), .A(n7125), .ZN(n7295) );
  AOI21_X1 U8879 ( .B1(n7126), .B2(n9729), .A(n7295), .ZN(n9766) );
  INV_X1 U8880 ( .A(n9766), .ZN(n7127) );
  AOI211_X1 U8881 ( .C1(n9791), .C2(n9763), .A(n9755), .B(n7127), .ZN(n7130)
         );
  AOI22_X1 U8882 ( .A1(n9553), .A2(n7290), .B1(n4846), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7128) );
  OAI21_X1 U8883 ( .B1(n7130), .B2(n4846), .A(n7128), .ZN(P1_U3527) );
  AOI22_X1 U8884 ( .A1(n9604), .A2(n7290), .B1(n6614), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n7129) );
  OAI21_X1 U8885 ( .B1(n7130), .B2(n6614), .A(n7129), .ZN(P1_U3468) );
  INV_X1 U8886 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9944) );
  INV_X1 U8887 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9977) );
  INV_X1 U8888 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8135) );
  AOI22_X1 U8889 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9977), .B2(n8135), .ZN(n9950) );
  NOR2_X1 U8890 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7131) );
  AOI21_X1 U8891 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7131), .ZN(n9953) );
  INV_X1 U8892 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10001) );
  INV_X1 U8893 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8103) );
  AOI22_X1 U8894 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .B1(n10001), .B2(n8103), .ZN(n9956) );
  NOR2_X1 U8895 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7132) );
  AOI21_X1 U8896 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7132), .ZN(n9959) );
  NOR2_X1 U8897 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7133) );
  AOI21_X1 U8898 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7133), .ZN(n9962) );
  NOR2_X1 U8899 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7134) );
  AOI21_X1 U8900 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7134), .ZN(n9965) );
  NOR2_X1 U8901 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7135) );
  AOI21_X1 U8902 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7135), .ZN(n9968) );
  NOR2_X1 U8903 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7136) );
  AOI21_X1 U8904 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7136), .ZN(n9971) );
  NOR2_X1 U8905 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7137) );
  AOI21_X1 U8906 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7137), .ZN(n10170) );
  NOR2_X1 U8907 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7138) );
  AOI21_X1 U8908 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7138), .ZN(n10176) );
  NOR2_X1 U8909 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7139) );
  AOI21_X1 U8910 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7139), .ZN(n10173) );
  NOR2_X1 U8911 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n7140) );
  AOI21_X1 U8912 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n7140), .ZN(n10179) );
  NOR2_X1 U8913 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7141) );
  AOI21_X1 U8914 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7141), .ZN(n10167) );
  AND2_X1 U8915 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7142) );
  NOR2_X1 U8916 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7142), .ZN(n9940) );
  INV_X1 U8917 ( .A(n9940), .ZN(n9941) );
  NAND3_X1 U8918 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U8919 ( .A1(n6670), .A2(n9942), .ZN(n9939) );
  NAND2_X1 U8920 ( .A1(n9941), .A2(n9939), .ZN(n10182) );
  NAND2_X1 U8921 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7143) );
  OAI21_X1 U8922 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7143), .ZN(n10181) );
  NOR2_X1 U8923 ( .A1(n10182), .A2(n10181), .ZN(n10180) );
  AOI21_X1 U8924 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10180), .ZN(n10185) );
  NAND2_X1 U8925 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7144) );
  OAI21_X1 U8926 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7144), .ZN(n10184) );
  NOR2_X1 U8927 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  AOI21_X1 U8928 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10183), .ZN(n10188) );
  NOR2_X1 U8929 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7145) );
  AOI21_X1 U8930 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7145), .ZN(n10187) );
  NAND2_X1 U8931 ( .A1(n10188), .A2(n10187), .ZN(n10186) );
  OAI21_X1 U8932 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10186), .ZN(n10166) );
  NAND2_X1 U8933 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  OAI21_X1 U8934 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10165), .ZN(n10178) );
  NAND2_X1 U8935 ( .A1(n10179), .A2(n10178), .ZN(n10177) );
  OAI21_X1 U8936 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10177), .ZN(n10172) );
  NAND2_X1 U8937 ( .A1(n10173), .A2(n10172), .ZN(n10171) );
  OAI21_X1 U8938 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10171), .ZN(n10175) );
  NAND2_X1 U8939 ( .A1(n10176), .A2(n10175), .ZN(n10174) );
  OAI21_X1 U8940 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10174), .ZN(n10169) );
  NAND2_X1 U8941 ( .A1(n10170), .A2(n10169), .ZN(n10168) );
  OAI21_X1 U8942 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10168), .ZN(n9970) );
  NAND2_X1 U8943 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  OAI21_X1 U8944 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9969), .ZN(n9967) );
  NAND2_X1 U8945 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  OAI21_X1 U8946 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9966), .ZN(n9964) );
  NAND2_X1 U8947 ( .A1(n9965), .A2(n9964), .ZN(n9963) );
  OAI21_X1 U8948 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9963), .ZN(n9961) );
  NAND2_X1 U8949 ( .A1(n9962), .A2(n9961), .ZN(n9960) );
  OAI21_X1 U8950 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9960), .ZN(n9958) );
  NAND2_X1 U8951 ( .A1(n9959), .A2(n9958), .ZN(n9957) );
  OAI21_X1 U8952 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9957), .ZN(n9955) );
  NAND2_X1 U8953 ( .A1(n9956), .A2(n9955), .ZN(n9954) );
  OAI21_X1 U8954 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9954), .ZN(n9952) );
  NAND2_X1 U8955 ( .A1(n9953), .A2(n9952), .ZN(n9951) );
  OAI21_X1 U8956 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9951), .ZN(n9949) );
  NAND2_X1 U8957 ( .A1(n9950), .A2(n9949), .ZN(n9948) );
  OAI21_X1 U8958 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9948), .ZN(n9945) );
  NOR2_X1 U8959 ( .A1(n9944), .A2(n9945), .ZN(n7146) );
  NAND2_X1 U8960 ( .A1(n9944), .A2(n9945), .ZN(n9943) );
  OAI21_X1 U8961 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7146), .A(n9943), .ZN(
        n7148) );
  XNOR2_X1 U8962 ( .A(n4569), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7147) );
  XNOR2_X1 U8963 ( .A(n7148), .B(n7147), .ZN(ADD_1068_U4) );
  INV_X1 U8964 ( .A(n7149), .ZN(n7156) );
  NAND2_X1 U8965 ( .A1(n7150), .A2(n9754), .ZN(n7152) );
  AOI22_X1 U8966 ( .A1(n9767), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n8846), .B2(
        n9756), .ZN(n7151) );
  OAI211_X1 U8967 ( .C1(n7277), .C2(n9760), .A(n7152), .B(n7151), .ZN(n7153)
         );
  AOI21_X1 U8968 ( .B1(n9764), .B2(n7154), .A(n7153), .ZN(n7155) );
  OAI21_X1 U8969 ( .B1(n7156), .B2(n9767), .A(n7155), .ZN(P1_U3289) );
  INV_X1 U8970 ( .A(n7270), .ZN(n7166) );
  OAI21_X1 U8971 ( .B1(n7159), .B2(n7158), .A(n7157), .ZN(n7160) );
  NAND2_X1 U8972 ( .A1(n7160), .A2(n5886), .ZN(n7165) );
  NAND2_X1 U8973 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7178) );
  INV_X1 U8974 ( .A(n7178), .ZN(n7163) );
  OAI22_X1 U8975 ( .A1(n7161), .A2(n8052), .B1(n7210), .B2(n8049), .ZN(n7162)
         );
  AOI211_X1 U8976 ( .C1(n7271), .C2(n8030), .A(n7163), .B(n7162), .ZN(n7164)
         );
  OAI211_X1 U8977 ( .C1(n7166), .C2(n8040), .A(n7165), .B(n7164), .ZN(P2_U3170) );
  AOI211_X1 U8978 ( .C1(n7169), .C2(n7168), .A(n9807), .B(n7167), .ZN(n7170)
         );
  INV_X1 U8979 ( .A(n7170), .ZN(n7189) );
  INV_X1 U8980 ( .A(n7171), .ZN(n7173) );
  NOR2_X1 U8981 ( .A1(n7173), .A2(n7172), .ZN(n7177) );
  INV_X1 U8982 ( .A(n7174), .ZN(n7175) );
  AOI21_X1 U8983 ( .B1(n7177), .B2(n7176), .A(n7175), .ZN(n7179) );
  OAI21_X1 U8984 ( .B1(n9853), .B2(n7179), .A(n7178), .ZN(n7187) );
  INV_X1 U8985 ( .A(n7180), .ZN(n7185) );
  NAND3_X1 U8986 ( .A1(n7183), .A2(n7182), .A3(n7181), .ZN(n7184) );
  AOI21_X1 U8987 ( .B1(n7185), .B2(n7184), .A(n9844), .ZN(n7186) );
  AOI211_X1 U8988 ( .C1(n9835), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7187), .B(
        n7186), .ZN(n7188) );
  OAI211_X1 U8989 ( .C1(n8139), .C2(n7190), .A(n7189), .B(n7188), .ZN(P2_U3186) );
  AOI22_X1 U8990 ( .A1(n9767), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9756), .B2(
        n6086), .ZN(n7193) );
  NAND2_X1 U8991 ( .A1(n9745), .A2(n7191), .ZN(n7192) );
  OAI211_X1 U8992 ( .C1(n7194), .C2(n9740), .A(n7193), .B(n7192), .ZN(n7195)
         );
  AOI21_X1 U8993 ( .B1(n7196), .B2(n9764), .A(n7195), .ZN(n7197) );
  OAI21_X1 U8994 ( .B1(n7198), .B2(n9767), .A(n7197), .ZN(P1_U3290) );
  NAND2_X1 U8995 ( .A1(n8073), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7199) );
  OAI21_X1 U8996 ( .B1(n8163), .B2(n8073), .A(n7199), .ZN(P2_U3522) );
  AND2_X1 U8997 ( .A1(n7201), .A2(n7200), .ZN(n7202) );
  NAND2_X1 U8998 ( .A1(n7203), .A2(n7202), .ZN(n8174) );
  NAND2_X1 U8999 ( .A1(n8174), .A2(n9901), .ZN(n7204) );
  OAI21_X1 U9000 ( .B1(n7207), .B2(n7206), .A(n7205), .ZN(n9860) );
  INV_X1 U9001 ( .A(n9860), .ZN(n7216) );
  XNOR2_X1 U9002 ( .A(n7209), .B(n7208), .ZN(n7212) );
  OAI22_X1 U9003 ( .A1(n6509), .A2(n8387), .B1(n7210), .B2(n8389), .ZN(n7211)
         );
  AOI21_X1 U9004 ( .B1(n7212), .B2(n8392), .A(n7211), .ZN(n9861) );
  AOI22_X1 U9005 ( .A1(n8219), .A2(n9858), .B1(n8396), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7213) );
  AND2_X1 U9006 ( .A1(n9861), .A2(n7213), .ZN(n7214) );
  MUX2_X1 U9007 ( .A(n7214), .B(n4799), .S(n8408), .Z(n7215) );
  OAI21_X1 U9008 ( .B1(n8384), .B2(n7216), .A(n7215), .ZN(P2_U3231) );
  INV_X1 U9009 ( .A(n7217), .ZN(n7222) );
  INV_X1 U9010 ( .A(n7218), .ZN(n7219) );
  MUX2_X1 U9011 ( .A(n6668), .B(n7219), .S(n8401), .Z(n7221) );
  AOI22_X1 U9012 ( .A1(n8381), .A2(n5783), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8396), .ZN(n7220) );
  OAI211_X1 U9013 ( .C1(n8384), .C2(n7222), .A(n7221), .B(n7220), .ZN(P2_U3232) );
  OAI21_X1 U9014 ( .B1(n7224), .B2(n7226), .A(n7223), .ZN(n9866) );
  INV_X1 U9015 ( .A(n9866), .ZN(n7232) );
  INV_X1 U9016 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7228) );
  XOR2_X1 U9017 ( .A(n7226), .B(n7225), .Z(n7227) );
  AOI222_X1 U9018 ( .A1(n8392), .A2(n7227), .B1(n8074), .B2(n8375), .C1(n8076), 
        .C2(n8377), .ZN(n9868) );
  MUX2_X1 U9019 ( .A(n7228), .B(n9868), .S(n8401), .Z(n7231) );
  AOI22_X1 U9020 ( .A1(n8381), .A2(n9865), .B1(n8396), .B2(n7229), .ZN(n7230)
         );
  OAI211_X1 U9021 ( .C1(n7232), .C2(n8384), .A(n7231), .B(n7230), .ZN(P2_U3230) );
  OAI21_X1 U9022 ( .B1(n7234), .B2(n7235), .A(n7233), .ZN(n7394) );
  INV_X1 U9023 ( .A(n7394), .ZN(n7251) );
  INV_X1 U9024 ( .A(n7235), .ZN(n7370) );
  NAND2_X1 U9025 ( .A1(n7239), .A2(n7370), .ZN(n7503) );
  OAI21_X1 U9026 ( .B1(n7370), .B2(n7239), .A(n7503), .ZN(n7241) );
  OR2_X1 U9027 ( .A1(n7570), .A2(n8907), .ZN(n7240) );
  OAI21_X1 U9028 ( .B1(n7355), .B2(n9276), .A(n7240), .ZN(n7448) );
  AOI21_X1 U9029 ( .B1(n7241), .B2(n9729), .A(n7448), .ZN(n7242) );
  OAI21_X1 U9030 ( .B1(n7251), .B2(n7491), .A(n7242), .ZN(n7392) );
  NAND2_X1 U9031 ( .A1(n7392), .A2(n9470), .ZN(n7250) );
  INV_X1 U9032 ( .A(n7243), .ZN(n7244) );
  AOI211_X1 U9033 ( .C1(n7452), .C2(n7244), .A(n9736), .B(n4437), .ZN(n7393)
         );
  AOI22_X1 U9034 ( .A1(n9767), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7245), .B2(
        n9756), .ZN(n7246) );
  OAI21_X1 U9035 ( .B1(n9760), .B2(n7247), .A(n7246), .ZN(n7248) );
  AOI21_X1 U9036 ( .B1(n7393), .B2(n9754), .A(n7248), .ZN(n7249) );
  OAI211_X1 U9037 ( .C1(n7251), .C2(n7498), .A(n7250), .B(n7249), .ZN(P1_U3286) );
  INV_X1 U9038 ( .A(n7252), .ZN(n7843) );
  OAI222_X1 U9039 ( .A1(n5770), .A2(P2_U3151), .B1(n8568), .B2(n7843), .C1(
        n8565), .C2(n7253), .ZN(P2_U3276) );
  INV_X1 U9040 ( .A(n7254), .ZN(n7325) );
  INV_X1 U9041 ( .A(n7157), .ZN(n7258) );
  INV_X1 U9042 ( .A(n7255), .ZN(n7257) );
  NOR3_X1 U9043 ( .A1(n7258), .A2(n7257), .A3(n7256), .ZN(n7260) );
  INV_X1 U9044 ( .A(n7259), .ZN(n8020) );
  OAI21_X1 U9045 ( .B1(n7260), .B2(n8020), .A(n5886), .ZN(n7265) );
  NAND2_X1 U9046 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7334) );
  INV_X1 U9047 ( .A(n7334), .ZN(n7263) );
  OAI22_X1 U9048 ( .A1(n7261), .A2(n8049), .B1(n8058), .B2(n9876), .ZN(n7262)
         );
  AOI211_X1 U9049 ( .C1(n8043), .C2(n8071), .A(n7263), .B(n7262), .ZN(n7264)
         );
  OAI211_X1 U9050 ( .C1(n7325), .C2(n8040), .A(n7265), .B(n7264), .ZN(P2_U3167) );
  XNOR2_X1 U9051 ( .A(n7266), .B(n7267), .ZN(n9870) );
  INV_X1 U9052 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7269) );
  XNOR2_X1 U9053 ( .A(n4367), .B(n7267), .ZN(n7268) );
  AOI222_X1 U9054 ( .A1(n8392), .A2(n7268), .B1(n8072), .B2(n8375), .C1(n8075), 
        .C2(n8377), .ZN(n9871) );
  MUX2_X1 U9055 ( .A(n7269), .B(n9871), .S(n8401), .Z(n7273) );
  AOI22_X1 U9056 ( .A1(n8381), .A2(n7271), .B1(n8396), .B2(n7270), .ZN(n7272)
         );
  OAI211_X1 U9057 ( .C1(n8384), .C2(n9870), .A(n7273), .B(n7272), .ZN(P2_U3229) );
  AOI22_X1 U9058 ( .A1(n9194), .A2(n8758), .B1(n6895), .B2(n7290), .ZN(n7294)
         );
  INV_X1 U9059 ( .A(n7274), .ZN(n7276) );
  NOR2_X1 U9060 ( .A1(n7276), .A2(n7275), .ZN(n8842) );
  OAI22_X1 U9061 ( .A1(n7279), .A2(n8764), .B1(n7277), .B2(n7352), .ZN(n7278)
         );
  XNOR2_X1 U9062 ( .A(n7278), .B(n8695), .ZN(n7287) );
  OR2_X1 U9063 ( .A1(n7279), .A2(n8677), .ZN(n7281) );
  NAND2_X1 U9064 ( .A1(n8847), .A2(n6895), .ZN(n7280) );
  NAND2_X1 U9065 ( .A1(n7281), .A2(n7280), .ZN(n7286) );
  XNOR2_X1 U9066 ( .A(n7287), .B(n7286), .ZN(n8841) );
  NAND2_X1 U9067 ( .A1(n7283), .A2(n7282), .ZN(n7284) );
  NAND2_X1 U9068 ( .A1(n7287), .A2(n7286), .ZN(n7288) );
  AOI22_X1 U9069 ( .A1(n9194), .A2(n6895), .B1(n7290), .B2(n8709), .ZN(n7291)
         );
  XNOR2_X1 U9070 ( .A(n7291), .B(n8695), .ZN(n7293) );
  INV_X1 U9071 ( .A(n7293), .ZN(n7292) );
  NOR2_X1 U9072 ( .A1(n8924), .A2(n9761), .ZN(n7300) );
  INV_X1 U9073 ( .A(n9757), .ZN(n7298) );
  NAND2_X1 U9074 ( .A1(n7295), .A2(n8895), .ZN(n7297) );
  OAI211_X1 U9075 ( .C1(n9653), .C2(n7298), .A(n7297), .B(n7296), .ZN(n7299)
         );
  AOI211_X1 U9076 ( .C1(n7301), .C2(n8905), .A(n7300), .B(n7299), .ZN(n7302)
         );
  INV_X1 U9077 ( .A(n7302), .ZN(P1_U3227) );
  NAND2_X1 U9078 ( .A1(n7303), .A2(n9032), .ZN(n7304) );
  NAND2_X1 U9079 ( .A1(n7305), .A2(n7304), .ZN(n7309) );
  OR2_X1 U9080 ( .A1(n7676), .A2(n9276), .ZN(n7307) );
  NAND2_X1 U9081 ( .A1(n9188), .A2(n8874), .ZN(n7306) );
  AND2_X1 U9082 ( .A1(n7307), .A2(n7306), .ZN(n9642) );
  INV_X1 U9083 ( .A(n9642), .ZN(n7308) );
  AOI21_X1 U9084 ( .B1(n7309), .B2(n9729), .A(n7308), .ZN(n9779) );
  OAI21_X1 U9085 ( .B1(n7311), .B2(n9032), .A(n7310), .ZN(n9782) );
  NAND2_X1 U9086 ( .A1(n9782), .A2(n9764), .ZN(n7318) );
  OAI22_X1 U9087 ( .A1(n9470), .A2(n7312), .B1(n9654), .B2(n9401), .ZN(n7316)
         );
  INV_X1 U9088 ( .A(n7313), .ZN(n7493) );
  OAI211_X1 U9089 ( .C1(n9780), .C2(n7314), .A(n7493), .B(n9505), .ZN(n9778)
         );
  NOR2_X1 U9090 ( .A1(n9778), .A2(n9740), .ZN(n7315) );
  AOI211_X1 U9091 ( .C1(n9745), .C2(n9651), .A(n7316), .B(n7315), .ZN(n7317)
         );
  OAI211_X1 U9092 ( .C1(n9767), .C2(n9779), .A(n7318), .B(n7317), .ZN(P1_U3283) );
  XNOR2_X1 U9093 ( .A(n7319), .B(n7320), .ZN(n9879) );
  INV_X1 U9094 ( .A(n9879), .ZN(n7330) );
  XNOR2_X1 U9095 ( .A(n7321), .B(n7320), .ZN(n7324) );
  INV_X1 U9096 ( .A(n9901), .ZN(n9899) );
  NAND2_X1 U9097 ( .A1(n9879), .A2(n9899), .ZN(n7323) );
  AOI22_X1 U9098 ( .A1(n8377), .A2(n8074), .B1(n8071), .B2(n8375), .ZN(n7322)
         );
  OAI211_X1 U9099 ( .C1(n8323), .C2(n7324), .A(n7323), .B(n7322), .ZN(n9877)
         );
  NAND2_X1 U9100 ( .A1(n9877), .A2(n8401), .ZN(n7329) );
  OAI22_X1 U9101 ( .A1(n8401), .A2(n7333), .B1(n7325), .B2(n8227), .ZN(n7326)
         );
  AOI21_X1 U9102 ( .B1(n8381), .B2(n7327), .A(n7326), .ZN(n7328) );
  OAI211_X1 U9103 ( .C1(n7330), .C2(n8174), .A(n7329), .B(n7328), .ZN(P2_U3228) );
  AOI21_X1 U9104 ( .B1(n7333), .B2(n7332), .A(n7331), .ZN(n7342) );
  INV_X1 U9105 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U9106 ( .B1(n9805), .B2(n7335), .A(n7334), .ZN(n7336) );
  INV_X1 U9107 ( .A(n7336), .ZN(n7341) );
  NOR2_X1 U9108 ( .A1(n7337), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7338) );
  OAI21_X1 U9109 ( .B1(n7339), .B2(n7338), .A(n9815), .ZN(n7340) );
  OAI211_X1 U9110 ( .C1(n7342), .C2(n9844), .A(n7341), .B(n7340), .ZN(n7347)
         );
  AOI211_X1 U9111 ( .C1(n7345), .C2(n7344), .A(n9807), .B(n7343), .ZN(n7346)
         );
  AOI211_X1 U9112 ( .C1(n9837), .C2(n7348), .A(n7347), .B(n7346), .ZN(n7349)
         );
  INV_X1 U9113 ( .A(n7349), .ZN(P2_U3187) );
  OAI22_X1 U9114 ( .A1(n7355), .A2(n8764), .B1(n7354), .B2(n7352), .ZN(n7353)
         );
  XNOR2_X1 U9115 ( .A(n7353), .B(n8695), .ZN(n7357) );
  OAI22_X1 U9116 ( .A1(n7355), .A2(n8677), .B1(n7354), .B2(n8764), .ZN(n7356)
         );
  NAND2_X1 U9117 ( .A1(n7357), .A2(n7356), .ZN(n7443) );
  NAND2_X1 U9118 ( .A1(n4748), .A2(n7443), .ZN(n7358) );
  XNOR2_X1 U9119 ( .A(n7444), .B(n7358), .ZN(n7366) );
  INV_X1 U9120 ( .A(n7359), .ZN(n7362) );
  AOI22_X1 U9121 ( .A1(n7360), .A2(n8895), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7361) );
  OAI21_X1 U9122 ( .B1(n7362), .B2(n9653), .A(n7361), .ZN(n7363) );
  AOI21_X1 U9123 ( .B1(n7364), .B2(n9650), .A(n7363), .ZN(n7365) );
  OAI21_X1 U9124 ( .B1(n7366), .B2(n9646), .A(n7365), .ZN(P1_U3239) );
  INV_X1 U9125 ( .A(n7367), .ZN(n7391) );
  AOI21_X1 U9126 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(n9613), .A(n7368), .ZN(
        n7369) );
  OAI21_X1 U9127 ( .B1(n7391), .B2(n9626), .A(n7369), .ZN(P1_U3335) );
  AND2_X1 U9128 ( .A1(n7373), .A2(n7372), .ZN(n7376) );
  INV_X1 U9129 ( .A(n7374), .ZN(n7375) );
  XOR2_X1 U9130 ( .A(n8935), .B(n7379), .Z(n7377) );
  OR2_X1 U9131 ( .A1(n7570), .A2(n9276), .ZN(n7680) );
  OAI21_X1 U9132 ( .B1(n7377), .B2(n9425), .A(n7680), .ZN(n9774) );
  INV_X1 U9133 ( .A(n9774), .ZN(n7388) );
  OAI21_X1 U9134 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n9776) );
  INV_X1 U9135 ( .A(n7687), .ZN(n9773) );
  XNOR2_X1 U9136 ( .A(n7509), .B(n9773), .ZN(n7382) );
  NAND2_X1 U9137 ( .A1(n9189), .A2(n8874), .ZN(n7681) );
  INV_X1 U9138 ( .A(n7681), .ZN(n7381) );
  AOI21_X1 U9139 ( .B1(n7382), .B2(n9505), .A(n7381), .ZN(n9772) );
  AOI22_X1 U9140 ( .A1(n9767), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7383), .B2(
        n9756), .ZN(n7385) );
  NAND2_X1 U9141 ( .A1(n9745), .A2(n7687), .ZN(n7384) );
  OAI211_X1 U9142 ( .C1(n9772), .C2(n9740), .A(n7385), .B(n7384), .ZN(n7386)
         );
  AOI21_X1 U9143 ( .B1(n9776), .B2(n9764), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9144 ( .B1(n7388), .B2(n9767), .A(n7387), .ZN(P1_U3284) );
  OAI222_X1 U9145 ( .A1(n8568), .A2(n7391), .B1(n7390), .B2(P2_U3151), .C1(
        n7389), .C2(n8555), .ZN(P2_U3275) );
  AOI211_X1 U9146 ( .C1(n7551), .C2(n7394), .A(n7393), .B(n7392), .ZN(n7397)
         );
  AOI22_X1 U9147 ( .A1(n9553), .A2(n7452), .B1(n4846), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7395) );
  OAI21_X1 U9148 ( .B1(n7397), .B2(n4846), .A(n7395), .ZN(P1_U3529) );
  AOI22_X1 U9149 ( .A1(n9604), .A2(n7452), .B1(n6614), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n7396) );
  OAI21_X1 U9150 ( .B1(n7397), .B2(n6614), .A(n7396), .ZN(P1_U3474) );
  OAI21_X1 U9151 ( .B1(n7400), .B2(n7399), .A(n7398), .ZN(n7413) );
  NAND2_X1 U9152 ( .A1(n9835), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U9153 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8024) );
  OAI211_X1 U9154 ( .C1(n8139), .C2(n7402), .A(n7401), .B(n8024), .ZN(n7412)
         );
  AOI21_X1 U9155 ( .B1(n7405), .B2(n7404), .A(n7403), .ZN(n7410) );
  AOI21_X1 U9156 ( .B1(n7408), .B2(n7407), .A(n7406), .ZN(n7409) );
  OAI22_X1 U9157 ( .A1(n7410), .A2(n9844), .B1(n7409), .B2(n9853), .ZN(n7411)
         );
  AOI211_X1 U9158 ( .C1(n7413), .C2(n9849), .A(n7412), .B(n7411), .ZN(n7414)
         );
  INV_X1 U9159 ( .A(n7414), .ZN(P2_U3188) );
  OR2_X1 U9160 ( .A1(n7416), .A2(n7415), .ZN(n7417) );
  NAND2_X1 U9161 ( .A1(n7418), .A2(n7417), .ZN(n9883) );
  XNOR2_X1 U9162 ( .A(n7466), .B(n7465), .ZN(n7419) );
  NAND2_X1 U9163 ( .A1(n7419), .A2(n8392), .ZN(n7421) );
  AOI22_X1 U9164 ( .A1(n8377), .A2(n8071), .B1(n8069), .B2(n8375), .ZN(n7420)
         );
  NAND2_X1 U9165 ( .A1(n7421), .A2(n7420), .ZN(n9886) );
  NAND2_X1 U9166 ( .A1(n9886), .A2(n8401), .ZN(n7425) );
  INV_X1 U9167 ( .A(n7422), .ZN(n7432) );
  OAI22_X1 U9168 ( .A1(n8401), .A2(n9821), .B1(n7432), .B2(n8227), .ZN(n7423)
         );
  AOI21_X1 U9169 ( .B1(n8381), .B2(n7434), .A(n7423), .ZN(n7424) );
  OAI211_X1 U9170 ( .C1(n8384), .C2(n9883), .A(n7425), .B(n7424), .ZN(P2_U3226) );
  INV_X1 U9171 ( .A(n7426), .ZN(n7427) );
  AOI21_X1 U9172 ( .B1(n7429), .B2(n7428), .A(n7427), .ZN(n7436) );
  AND2_X1 U9173 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9824) );
  AOI21_X1 U9174 ( .B1(n8043), .B2(n8069), .A(n9824), .ZN(n7431) );
  NAND2_X1 U9175 ( .A1(n8038), .A2(n8071), .ZN(n7430) );
  OAI211_X1 U9176 ( .C1(n8040), .C2(n7432), .A(n7431), .B(n7430), .ZN(n7433)
         );
  AOI21_X1 U9177 ( .B1(n7434), .B2(n8030), .A(n7433), .ZN(n7435) );
  OAI21_X1 U9178 ( .B1(n7436), .B2(n7983), .A(n7435), .ZN(P2_U3153) );
  XNOR2_X1 U9179 ( .A(n7437), .B(n7438), .ZN(n7456) );
  XOR2_X1 U9180 ( .A(n7439), .B(n7438), .Z(n7440) );
  AOI222_X1 U9181 ( .A1(n8392), .A2(n7440), .B1(n8070), .B2(n8375), .C1(n8072), 
        .C2(n8377), .ZN(n7455) );
  MUX2_X1 U9182 ( .A(n5920), .B(n7455), .S(n8401), .Z(n7442) );
  AOI22_X1 U9183 ( .A1(n8381), .A2(n8029), .B1(n8396), .B2(n8028), .ZN(n7441)
         );
  OAI211_X1 U9184 ( .C1(n8384), .C2(n7456), .A(n7442), .B(n7441), .ZN(P2_U3227) );
  OR2_X1 U9185 ( .A1(n7501), .A2(n8677), .ZN(n7446) );
  NAND2_X1 U9186 ( .A1(n7452), .A2(n6895), .ZN(n7445) );
  NAND2_X1 U9187 ( .A1(n7446), .A2(n7445), .ZN(n7564) );
  AOI22_X1 U9188 ( .A1(n9192), .A2(n6895), .B1(n7452), .B2(n8709), .ZN(n7447)
         );
  XNOR2_X1 U9189 ( .A(n7447), .B(n8695), .ZN(n7563) );
  XOR2_X1 U9190 ( .A(n7564), .B(n7563), .Z(n7566) );
  XOR2_X1 U9191 ( .A(n7567), .B(n7566), .Z(n7454) );
  AOI22_X1 U9192 ( .A1(n7448), .A2(n8895), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7449) );
  OAI21_X1 U9193 ( .B1(n7450), .B2(n9653), .A(n7449), .ZN(n7451) );
  AOI21_X1 U9194 ( .B1(n7452), .B2(n8912), .A(n7451), .ZN(n7453) );
  OAI21_X1 U9195 ( .B1(n7454), .B2(n9646), .A(n7453), .ZN(P1_U3213) );
  INV_X1 U9196 ( .A(n9915), .ZN(n8473) );
  OAI21_X1 U9197 ( .B1(n8473), .B2(n7456), .A(n7455), .ZN(n7463) );
  OAI22_X1 U9198 ( .A1(n8457), .A2(n7461), .B1(n9938), .B2(n7457), .ZN(n7458)
         );
  AOI21_X1 U9199 ( .B1(n7463), .B2(n9938), .A(n7458), .ZN(n7459) );
  INV_X1 U9200 ( .A(n7459), .ZN(P2_U3465) );
  INV_X1 U9201 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7460) );
  OAI22_X1 U9202 ( .A1(n7461), .A2(n8543), .B1(n9919), .B2(n7460), .ZN(n7462)
         );
  AOI21_X1 U9203 ( .B1(n7463), .B2(n9919), .A(n7462), .ZN(n7464) );
  INV_X1 U9204 ( .A(n7464), .ZN(P2_U3408) );
  NAND2_X1 U9205 ( .A1(n7466), .A2(n7465), .ZN(n7471) );
  NAND2_X1 U9206 ( .A1(n7471), .A2(n7467), .ZN(n7469) );
  INV_X1 U9207 ( .A(n7479), .ZN(n7468) );
  AOI21_X1 U9208 ( .B1(n7469), .B2(n7468), .A(n8323), .ZN(n7474) );
  NAND2_X1 U9209 ( .A1(n7471), .A2(n7470), .ZN(n7473) );
  OAI22_X1 U9210 ( .A1(n8026), .A2(n8387), .B1(n7599), .B2(n8389), .ZN(n7472)
         );
  AOI21_X1 U9211 ( .B1(n7474), .B2(n7473), .A(n7472), .ZN(n9888) );
  INV_X1 U9212 ( .A(n7544), .ZN(n7475) );
  OAI22_X1 U9213 ( .A1(n8401), .A2(n7476), .B1(n7475), .B2(n8227), .ZN(n7477)
         );
  AOI21_X1 U9214 ( .B1(n8381), .B2(n7478), .A(n7477), .ZN(n7482) );
  XNOR2_X1 U9215 ( .A(n7480), .B(n7479), .ZN(n9891) );
  NAND2_X1 U9216 ( .A1(n9891), .A2(n8406), .ZN(n7481) );
  OAI211_X1 U9217 ( .C1(n9888), .C2(n8408), .A(n7482), .B(n7481), .ZN(P2_U3225) );
  INV_X1 U9218 ( .A(n7483), .ZN(n7833) );
  OAI222_X1 U9219 ( .A1(n8568), .A2(n7833), .B1(n7485), .B2(P2_U3151), .C1(
        n7484), .C2(n8555), .ZN(P2_U3274) );
  INV_X1 U9220 ( .A(n7487), .ZN(n9046) );
  XNOR2_X1 U9221 ( .A(n7486), .B(n9046), .ZN(n7547) );
  AOI22_X1 U9222 ( .A1(n9167), .A2(n9189), .B1(n9187), .B2(n8874), .ZN(n8885)
         );
  XNOR2_X1 U9223 ( .A(n7488), .B(n9046), .ZN(n7489) );
  NAND2_X1 U9224 ( .A1(n7489), .A2(n9729), .ZN(n7490) );
  OAI211_X1 U9225 ( .C1(n7547), .C2(n7491), .A(n8885), .B(n7490), .ZN(n7548)
         );
  NAND2_X1 U9226 ( .A1(n7548), .A2(n9470), .ZN(n7497) );
  INV_X1 U9227 ( .A(n9737), .ZN(n7492) );
  AOI211_X1 U9228 ( .C1(n8592), .C2(n7493), .A(n9736), .B(n7492), .ZN(n7549)
         );
  AOI22_X1 U9229 ( .A1(n9767), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8887), .B2(
        n9756), .ZN(n7494) );
  OAI21_X1 U9230 ( .B1(n8890), .B2(n9760), .A(n7494), .ZN(n7495) );
  AOI21_X1 U9231 ( .B1(n7549), .B2(n9754), .A(n7495), .ZN(n7496) );
  OAI211_X1 U9232 ( .C1(n7547), .C2(n7498), .A(n7497), .B(n7496), .ZN(P1_U3282) );
  INV_X1 U9233 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7515) );
  OAI21_X1 U9234 ( .B1(n7500), .B2(n7504), .A(n7499), .ZN(n9750) );
  INV_X1 U9235 ( .A(n9750), .ZN(n7512) );
  OAI22_X1 U9236 ( .A1(n7676), .A2(n8907), .B1(n7501), .B2(n9276), .ZN(n7575)
         );
  NAND2_X1 U9237 ( .A1(n7503), .A2(n7502), .ZN(n7505) );
  XNOR2_X1 U9238 ( .A(n7505), .B(n7504), .ZN(n7506) );
  NOR2_X1 U9239 ( .A1(n7506), .A2(n9425), .ZN(n7507) );
  AOI211_X1 U9240 ( .C1(n7508), .C2(n9750), .A(n7575), .B(n7507), .ZN(n9753)
         );
  OAI211_X1 U9241 ( .C1(n4437), .C2(n7510), .A(n9505), .B(n7509), .ZN(n9747)
         );
  OAI211_X1 U9242 ( .C1(n7512), .C2(n7511), .A(n9753), .B(n9747), .ZN(n7516)
         );
  NAND2_X1 U9243 ( .A1(n7516), .A2(n9793), .ZN(n7514) );
  NAND2_X1 U9244 ( .A1(n9604), .A2(n9746), .ZN(n7513) );
  OAI211_X1 U9245 ( .C1(n9793), .C2(n7515), .A(n7514), .B(n7513), .ZN(P1_U3477) );
  INV_X1 U9246 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U9247 ( .A1(n7516), .A2(n9799), .ZN(n7518) );
  NAND2_X1 U9248 ( .A1(n9553), .A2(n9746), .ZN(n7517) );
  OAI211_X1 U9249 ( .C1(n9799), .C2(n7519), .A(n7518), .B(n7517), .ZN(P1_U3530) );
  INV_X1 U9250 ( .A(n7520), .ZN(n7881) );
  OAI222_X1 U9251 ( .A1(n8565), .A2(n7522), .B1(n8568), .B2(n7881), .C1(
        P2_U3151), .C2(n7521), .ZN(P2_U3273) );
  OAI21_X1 U9252 ( .B1(n7524), .B2(n9047), .A(n7523), .ZN(n7642) );
  XNOR2_X1 U9253 ( .A(n7525), .B(n9047), .ZN(n7529) );
  NAND2_X1 U9254 ( .A1(n9185), .A2(n8874), .ZN(n7526) );
  OAI21_X1 U9255 ( .B1(n7527), .B2(n9276), .A(n7526), .ZN(n8863) );
  INV_X1 U9256 ( .A(n8863), .ZN(n7528) );
  OAI21_X1 U9257 ( .B1(n7529), .B2(n9425), .A(n7528), .ZN(n7635) );
  INV_X1 U9258 ( .A(n8867), .ZN(n7535) );
  INV_X1 U9259 ( .A(n7589), .ZN(n7531) );
  AOI211_X1 U9260 ( .C1(n8867), .C2(n9738), .A(n9736), .B(n7531), .ZN(n7636)
         );
  NAND2_X1 U9261 ( .A1(n7636), .A2(n9754), .ZN(n7534) );
  AOI22_X1 U9262 ( .A1(n9767), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7532), .B2(
        n9756), .ZN(n7533) );
  OAI211_X1 U9263 ( .C1(n7535), .C2(n9760), .A(n7534), .B(n7533), .ZN(n7536)
         );
  AOI21_X1 U9264 ( .B1(n7635), .B2(n9470), .A(n7536), .ZN(n7537) );
  OAI21_X1 U9265 ( .B1(n7642), .B2(n9466), .A(n7537), .ZN(P1_U3280) );
  OAI21_X1 U9266 ( .B1(n7629), .B2(n7539), .A(n7538), .ZN(n7540) );
  NAND2_X1 U9267 ( .A1(n7540), .A2(n5886), .ZN(n7546) );
  OR2_X1 U9268 ( .A1(n8026), .A2(n8049), .ZN(n7542) );
  INV_X1 U9269 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7541) );
  OR2_X1 U9270 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7541), .ZN(n7611) );
  OAI211_X1 U9271 ( .C1(n7599), .C2(n8052), .A(n7542), .B(n7611), .ZN(n7543)
         );
  AOI21_X1 U9272 ( .B1(n8055), .B2(n7544), .A(n7543), .ZN(n7545) );
  OAI211_X1 U9273 ( .C1(n9889), .C2(n8058), .A(n7546), .B(n7545), .ZN(P2_U3161) );
  INV_X1 U9274 ( .A(n7547), .ZN(n7550) );
  AOI211_X1 U9275 ( .C1(n7551), .C2(n7550), .A(n7549), .B(n7548), .ZN(n7553)
         );
  MUX2_X1 U9276 ( .A(n6985), .B(n7553), .S(n9799), .Z(n7552) );
  OAI21_X1 U9277 ( .B1(n8890), .B2(n6505), .A(n7552), .ZN(P1_U3533) );
  INV_X1 U9278 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7554) );
  MUX2_X1 U9279 ( .A(n7554), .B(n7553), .S(n9793), .Z(n7555) );
  OAI21_X1 U9280 ( .B1(n8890), .B2(n6501), .A(n7555), .ZN(P1_U3486) );
  NAND2_X1 U9281 ( .A1(n6339), .A2(n7556), .ZN(n7558) );
  OR2_X1 U9282 ( .A1(n7557), .A2(P1_U3086), .ZN(n9170) );
  OAI211_X1 U9283 ( .C1(n7559), .C2(n9623), .A(n7558), .B(n9170), .ZN(P1_U3332) );
  NAND2_X1 U9284 ( .A1(n6339), .A2(n8559), .ZN(n7561) );
  OAI211_X1 U9285 ( .C1(n7562), .C2(n8555), .A(n7561), .B(n7560), .ZN(P2_U3272) );
  INV_X1 U9286 ( .A(n7563), .ZN(n7565) );
  NAND2_X1 U9287 ( .A1(n9746), .A2(n8709), .ZN(n7568) );
  OAI21_X1 U9288 ( .B1(n7570), .B2(n8764), .A(n7568), .ZN(n7569) );
  XNOR2_X1 U9289 ( .A(n7569), .B(n8761), .ZN(n8577) );
  XNOR2_X1 U9290 ( .A(n8580), .B(n8577), .ZN(n7574) );
  OR2_X1 U9291 ( .A1(n7570), .A2(n8677), .ZN(n7572) );
  NAND2_X1 U9292 ( .A1(n9746), .A2(n6895), .ZN(n7571) );
  INV_X1 U9293 ( .A(n8575), .ZN(n7573) );
  NOR2_X1 U9294 ( .A1(n7574), .A2(n7573), .ZN(n7677) );
  AOI21_X1 U9295 ( .B1(n7574), .B2(n7573), .A(n7677), .ZN(n7580) );
  INV_X1 U9296 ( .A(n9744), .ZN(n7577) );
  AOI22_X1 U9297 ( .A1(n7575), .A2(n8895), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7576) );
  OAI21_X1 U9298 ( .B1(n7577), .B2(n9653), .A(n7576), .ZN(n7578) );
  AOI21_X1 U9299 ( .B1(n9746), .B2(n8912), .A(n7578), .ZN(n7579) );
  OAI21_X1 U9300 ( .B1(n7580), .B2(n9646), .A(n7579), .ZN(P1_U3221) );
  XOR2_X1 U9301 ( .A(n9048), .B(n7581), .Z(n7692) );
  INV_X1 U9302 ( .A(n7692), .ZN(n7594) );
  NAND2_X1 U9303 ( .A1(n7582), .A2(n9048), .ZN(n7583) );
  NAND2_X1 U9304 ( .A1(n7652), .A2(n7583), .ZN(n7584) );
  NAND2_X1 U9305 ( .A1(n7584), .A2(n9729), .ZN(n7588) );
  OR2_X1 U9306 ( .A1(n8790), .A2(n9276), .ZN(n7586) );
  NAND2_X1 U9307 ( .A1(n9184), .A2(n8874), .ZN(n7585) );
  NAND2_X1 U9308 ( .A1(n7586), .A2(n7585), .ZN(n8734) );
  INV_X1 U9309 ( .A(n8734), .ZN(n7587) );
  NAND2_X1 U9310 ( .A1(n7588), .A2(n7587), .ZN(n7690) );
  INV_X1 U9311 ( .A(n8738), .ZN(n7698) );
  AOI211_X1 U9312 ( .C1(n8738), .C2(n7589), .A(n9736), .B(n4421), .ZN(n7691)
         );
  NAND2_X1 U9313 ( .A1(n7691), .A2(n9754), .ZN(n7591) );
  AOI22_X1 U9314 ( .A1(n9767), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8733), .B2(
        n9756), .ZN(n7590) );
  OAI211_X1 U9315 ( .C1(n7698), .C2(n9760), .A(n7591), .B(n7590), .ZN(n7592)
         );
  AOI21_X1 U9316 ( .B1(n7690), .B2(n9470), .A(n7592), .ZN(n7593) );
  OAI21_X1 U9317 ( .B1(n7594), .B2(n9466), .A(n7593), .ZN(P1_U3279) );
  XNOR2_X1 U9318 ( .A(n7595), .B(n7596), .ZN(n9900) );
  XNOR2_X1 U9319 ( .A(n7597), .B(n7596), .ZN(n7598) );
  OAI222_X1 U9320 ( .A1(n8389), .A2(n8388), .B1(n8387), .B2(n7599), .C1(n7598), 
        .C2(n8323), .ZN(n9903) );
  NAND2_X1 U9321 ( .A1(n9903), .A2(n8401), .ZN(n7603) );
  INV_X1 U9322 ( .A(n7774), .ZN(n7600) );
  OAI22_X1 U9323 ( .A1(n8401), .A2(n5927), .B1(n7600), .B2(n8227), .ZN(n7601)
         );
  AOI21_X1 U9324 ( .B1(n8381), .B2(n9905), .A(n7601), .ZN(n7602) );
  OAI211_X1 U9325 ( .C1(n8384), .C2(n9900), .A(n7603), .B(n7602), .ZN(P2_U3223) );
  INV_X1 U9326 ( .A(n7604), .ZN(n7605) );
  AOI21_X1 U9327 ( .B1(n7607), .B2(n7606), .A(n7605), .ZN(n7622) );
  XNOR2_X1 U9328 ( .A(n7609), .B(n7608), .ZN(n7620) );
  INV_X1 U9329 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9330 ( .A1(n9837), .A2(n7610), .ZN(n7612) );
  OAI211_X1 U9331 ( .C1(n7613), .C2(n9805), .A(n7612), .B(n7611), .ZN(n7619)
         );
  AOI21_X1 U9332 ( .B1(n7616), .B2(n7615), .A(n7614), .ZN(n7617) );
  NOR2_X1 U9333 ( .A1(n7617), .A2(n9853), .ZN(n7618) );
  AOI211_X1 U9334 ( .C1(n9849), .C2(n7620), .A(n7619), .B(n7618), .ZN(n7621)
         );
  OAI21_X1 U9335 ( .B1(n7622), .B2(n9844), .A(n7621), .ZN(P2_U3190) );
  INV_X1 U9336 ( .A(n7623), .ZN(n7624) );
  AOI21_X1 U9337 ( .B1(n7625), .B2(n7626), .A(n7624), .ZN(n9898) );
  INV_X1 U9338 ( .A(n9898), .ZN(n9895) );
  XNOR2_X1 U9339 ( .A(n7627), .B(n7626), .ZN(n7628) );
  OAI222_X1 U9340 ( .A1(n8389), .A2(n7630), .B1(n8387), .B2(n7629), .C1(n7628), 
        .C2(n8323), .ZN(n9896) );
  NAND2_X1 U9341 ( .A1(n9896), .A2(n8401), .ZN(n7634) );
  INV_X1 U9342 ( .A(n7631), .ZN(n7755) );
  OAI22_X1 U9343 ( .A1(n8401), .A2(n7726), .B1(n7755), .B2(n8227), .ZN(n7632)
         );
  AOI21_X1 U9344 ( .B1(n8381), .B2(n7762), .A(n7632), .ZN(n7633) );
  OAI211_X1 U9345 ( .C1(n9895), .C2(n8384), .A(n7634), .B(n7633), .ZN(P2_U3224) );
  INV_X1 U9346 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7637) );
  AOI211_X1 U9347 ( .C1(n9546), .C2(n8867), .A(n7636), .B(n7635), .ZN(n7639)
         );
  MUX2_X1 U9348 ( .A(n7637), .B(n7639), .S(n9799), .Z(n7638) );
  OAI21_X1 U9349 ( .B1(n9555), .B2(n7642), .A(n7638), .ZN(P1_U3535) );
  INV_X1 U9350 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7640) );
  MUX2_X1 U9351 ( .A(n7640), .B(n7639), .S(n9793), .Z(n7641) );
  OAI21_X1 U9352 ( .B1(n7642), .B2(n9606), .A(n7641), .ZN(P1_U3492) );
  INV_X1 U9353 ( .A(n7643), .ZN(n7647) );
  OAI222_X1 U9354 ( .A1(n8568), .A2(n7647), .B1(P2_U3151), .B2(n7645), .C1(
        n7644), .C2(n8555), .ZN(P2_U3271) );
  OAI222_X1 U9355 ( .A1(P1_U3086), .A2(n7648), .B1(n9620), .B2(n7647), .C1(
        n7646), .C2(n9623), .ZN(P1_U3331) );
  XOR2_X1 U9356 ( .A(n7649), .B(n9051), .Z(n7771) );
  NAND2_X1 U9357 ( .A1(n7650), .A2(n9729), .ZN(n7656) );
  INV_X1 U9358 ( .A(n9051), .ZN(n7651) );
  AOI21_X1 U9359 ( .B1(n7652), .B2(n8958), .A(n7651), .ZN(n7655) );
  OR2_X1 U9360 ( .A1(n8821), .A2(n8907), .ZN(n7654) );
  NAND2_X1 U9361 ( .A1(n9185), .A2(n9167), .ZN(n7653) );
  AND2_X1 U9362 ( .A1(n7654), .A2(n7653), .ZN(n8923) );
  OAI21_X1 U9363 ( .B1(n7656), .B2(n7655), .A(n8923), .ZN(n7765) );
  OAI211_X1 U9364 ( .C1(n4421), .C2(n8925), .A(n9458), .B(n9505), .ZN(n7764)
         );
  AOI22_X1 U9365 ( .A1(n9767), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8928), .B2(
        n9756), .ZN(n7658) );
  NAND2_X1 U9366 ( .A1(n8609), .A2(n9745), .ZN(n7657) );
  OAI211_X1 U9367 ( .C1(n7764), .C2(n9740), .A(n7658), .B(n7657), .ZN(n7659)
         );
  AOI21_X1 U9368 ( .B1(n7765), .B2(n9470), .A(n7659), .ZN(n7660) );
  OAI21_X1 U9369 ( .B1(n7771), .B2(n9466), .A(n7660), .ZN(P1_U3278) );
  XNOR2_X1 U9370 ( .A(n7661), .B(n7662), .ZN(n9907) );
  INV_X1 U9371 ( .A(n9907), .ZN(n7672) );
  INV_X1 U9372 ( .A(n8005), .ZN(n7668) );
  NAND2_X1 U9373 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  NAND3_X1 U9374 ( .A1(n7665), .A2(n8392), .A3(n7664), .ZN(n7667) );
  AOI22_X1 U9375 ( .A1(n8378), .A2(n8375), .B1(n8377), .B2(n8067), .ZN(n7666)
         );
  AND2_X1 U9376 ( .A1(n7667), .A2(n7666), .ZN(n9911) );
  OAI21_X1 U9377 ( .B1(n7668), .B2(n8227), .A(n9911), .ZN(n7670) );
  INV_X1 U9378 ( .A(n9908), .ZN(n8008) );
  OAI22_X1 U9379 ( .A1(n8008), .A2(n8403), .B1(n7809), .B2(n8401), .ZN(n7669)
         );
  AOI21_X1 U9380 ( .B1(n7670), .B2(n8401), .A(n7669), .ZN(n7671) );
  OAI21_X1 U9381 ( .B1(n8384), .B2(n7672), .A(n7671), .ZN(P2_U3222) );
  NAND2_X1 U9382 ( .A1(n7687), .A2(n8709), .ZN(n7674) );
  OR2_X1 U9383 ( .A1(n7676), .A2(n8764), .ZN(n7673) );
  NAND2_X1 U9384 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  XNOR2_X1 U9385 ( .A(n7675), .B(n8695), .ZN(n8573) );
  OAI22_X1 U9386 ( .A1(n9773), .A2(n8764), .B1(n7676), .B2(n8677), .ZN(n8572)
         );
  NAND2_X1 U9387 ( .A1(n8573), .A2(n8572), .ZN(n8570) );
  OAI21_X1 U9388 ( .B1(n8573), .B2(n8572), .A(n8570), .ZN(n7679) );
  AOI21_X1 U9389 ( .B1(n8577), .B2(n8580), .A(n7677), .ZN(n7678) );
  XOR2_X1 U9390 ( .A(n7679), .B(n7678), .Z(n7689) );
  NAND2_X1 U9391 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  NAND2_X1 U9392 ( .A1(n7682), .A2(n8895), .ZN(n7684) );
  OAI211_X1 U9393 ( .C1(n9653), .C2(n7685), .A(n7684), .B(n7683), .ZN(n7686)
         );
  AOI21_X1 U9394 ( .B1(n7687), .B2(n9650), .A(n7686), .ZN(n7688) );
  OAI21_X1 U9395 ( .B1(n7689), .B2(n9646), .A(n7688), .ZN(P1_U3231) );
  INV_X1 U9396 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7693) );
  AOI211_X1 U9397 ( .C1(n7692), .C2(n9791), .A(n7691), .B(n7690), .ZN(n7695)
         );
  MUX2_X1 U9398 ( .A(n7693), .B(n7695), .S(n9793), .Z(n7694) );
  OAI21_X1 U9399 ( .B1(n7698), .B2(n6501), .A(n7694), .ZN(P1_U3495) );
  INV_X1 U9400 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7696) );
  MUX2_X1 U9401 ( .A(n7696), .B(n7695), .S(n9799), .Z(n7697) );
  OAI21_X1 U9402 ( .B1(n7698), .B2(n6505), .A(n7697), .ZN(P1_U3536) );
  INV_X1 U9403 ( .A(n7699), .ZN(n7702) );
  OAI222_X1 U9404 ( .A1(n8568), .A2(n7702), .B1(P2_U3151), .B2(n7700), .C1(
        n10114), .C2(n8555), .ZN(P2_U3270) );
  OAI222_X1 U9405 ( .A1(P1_U3086), .A2(n7703), .B1(n9626), .B2(n7702), .C1(
        n7701), .C2(n9623), .ZN(P1_U3330) );
  XNOR2_X1 U9406 ( .A(n9243), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9244) );
  OAI21_X1 U9407 ( .B1(n7710), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7704), .ZN(
        n9674) );
  XNOR2_X1 U9408 ( .A(n9681), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9675) );
  NOR2_X1 U9409 ( .A1(n9674), .A2(n9675), .ZN(n9673) );
  XNOR2_X1 U9410 ( .A(n9693), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9689) );
  NOR2_X1 U9411 ( .A1(n9690), .A2(n9689), .ZN(n9688) );
  NOR2_X1 U9412 ( .A1(n7705), .A2(n7713), .ZN(n7706) );
  INV_X1 U9413 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9698) );
  XNOR2_X1 U9414 ( .A(n7713), .B(n7705), .ZN(n9699) );
  NOR2_X1 U9415 ( .A1(n9698), .A2(n9699), .ZN(n9697) );
  NOR2_X1 U9416 ( .A1(n7706), .A2(n9697), .ZN(n7740) );
  XOR2_X1 U9417 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n7749), .Z(n7741) );
  INV_X1 U9418 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7708) );
  AOI22_X1 U9419 ( .A1(n7740), .A2(n7741), .B1(n7708), .B2(n7707), .ZN(n9245)
         );
  XOR2_X1 U9420 ( .A(n9244), .B(n9245), .Z(n7722) );
  XNOR2_X1 U9421 ( .A(n9243), .B(n10142), .ZN(n7717) );
  XNOR2_X1 U9422 ( .A(n9681), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n9677) );
  NOR2_X1 U9423 ( .A1(n9678), .A2(n9677), .ZN(n9676) );
  NAND2_X1 U9424 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9693), .ZN(n7711) );
  OAI21_X1 U9425 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9693), .A(n7711), .ZN(
        n9686) );
  NOR2_X1 U9426 ( .A1(n9687), .A2(n9686), .ZN(n9685) );
  NOR2_X1 U9427 ( .A1(n7712), .A2(n7713), .ZN(n7714) );
  INV_X1 U9428 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9702) );
  XNOR2_X1 U9429 ( .A(n7713), .B(n7712), .ZN(n9703) );
  NOR2_X1 U9430 ( .A1(n9702), .A2(n9703), .ZN(n9701) );
  NOR2_X1 U9431 ( .A1(n7714), .A2(n9701), .ZN(n7746) );
  XNOR2_X1 U9432 ( .A(n7749), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U9433 ( .A1(n7749), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U9434 ( .A1(n7716), .A2(n7717), .ZN(n9239) );
  OAI21_X1 U9435 ( .B1(n7717), .B2(n7716), .A(n9239), .ZN(n7720) );
  NAND2_X1 U9436 ( .A1(n9712), .A2(n9243), .ZN(n7718) );
  NAND2_X1 U9437 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8826) );
  OAI211_X1 U9438 ( .C1(n9724), .C2(n9977), .A(n7718), .B(n8826), .ZN(n7719)
         );
  AOI21_X1 U9439 ( .B1(n7720), .B2(n9716), .A(n7719), .ZN(n7721) );
  OAI21_X1 U9440 ( .B1(n7722), .B2(n9709), .A(n7721), .ZN(P1_U3260) );
  AOI21_X1 U9441 ( .B1(n9931), .B2(n7724), .A(n7723), .ZN(n7739) );
  AOI21_X1 U9442 ( .B1(n7727), .B2(n7726), .A(n7725), .ZN(n7728) );
  NOR2_X1 U9443 ( .A1(n7728), .A2(n9844), .ZN(n7737) );
  OAI21_X1 U9444 ( .B1(n7731), .B2(n7730), .A(n7729), .ZN(n7732) );
  NAND2_X1 U9445 ( .A1(n7732), .A2(n9849), .ZN(n7734) );
  AND2_X1 U9446 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7752) );
  AOI21_X1 U9447 ( .B1(n9835), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7752), .ZN(
        n7733) );
  OAI211_X1 U9448 ( .C1(n8139), .C2(n7735), .A(n7734), .B(n7733), .ZN(n7736)
         );
  NOR2_X1 U9449 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  OAI21_X1 U9450 ( .B1(n7739), .B2(n9853), .A(n7738), .ZN(P2_U3191) );
  XOR2_X1 U9451 ( .A(n7741), .B(n7740), .Z(n7751) );
  INV_X1 U9452 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U9453 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8811) );
  OAI21_X1 U9454 ( .B1(n9724), .B2(n7742), .A(n8811), .ZN(n7748) );
  INV_X1 U9455 ( .A(n7743), .ZN(n7744) );
  AOI211_X1 U9456 ( .C1(n7746), .C2(n7745), .A(n9700), .B(n7744), .ZN(n7747)
         );
  AOI211_X1 U9457 ( .C1(n9712), .C2(n7749), .A(n7748), .B(n7747), .ZN(n7750)
         );
  OAI21_X1 U9458 ( .B1(n7751), .B2(n9709), .A(n7750), .ZN(P1_U3259) );
  AOI21_X1 U9459 ( .B1(n8038), .B2(n8069), .A(n7752), .ZN(n7754) );
  NAND2_X1 U9460 ( .A1(n8043), .A2(n8067), .ZN(n7753) );
  OAI211_X1 U9461 ( .C1(n8040), .C2(n7755), .A(n7754), .B(n7753), .ZN(n7761)
         );
  INV_X1 U9462 ( .A(n7756), .ZN(n7757) );
  AOI211_X1 U9463 ( .C1(n7759), .C2(n7758), .A(n7983), .B(n7757), .ZN(n7760)
         );
  AOI211_X1 U9464 ( .C1(n7762), .C2(n8030), .A(n7761), .B(n7760), .ZN(n7763)
         );
  INV_X1 U9465 ( .A(n7763), .ZN(P2_U3171) );
  INV_X1 U9466 ( .A(n7764), .ZN(n7766) );
  AOI211_X1 U9467 ( .C1(n9546), .C2(n8609), .A(n7766), .B(n7765), .ZN(n7768)
         );
  MUX2_X1 U9468 ( .A(n9698), .B(n7768), .S(n9799), .Z(n7767) );
  OAI21_X1 U9469 ( .B1(n7771), .B2(n9555), .A(n7767), .ZN(P1_U3537) );
  INV_X1 U9470 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7769) );
  MUX2_X1 U9471 ( .A(n7769), .B(n7768), .S(n9793), .Z(n7770) );
  OAI21_X1 U9472 ( .B1(n7771), .B2(n9606), .A(n7770), .ZN(P1_U3498) );
  XNOR2_X1 U9473 ( .A(n7916), .B(n8067), .ZN(n7772) );
  NOR2_X1 U9474 ( .A1(n7772), .A2(n7773), .ZN(n7998) );
  AOI21_X1 U9475 ( .B1(n7773), .B2(n7772), .A(n7998), .ZN(n7780) );
  NAND2_X1 U9476 ( .A1(n8055), .A2(n7774), .ZN(n7777) );
  INV_X1 U9477 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7775) );
  NOR2_X1 U9478 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7775), .ZN(n7787) );
  AOI21_X1 U9479 ( .B1(n8068), .B2(n8038), .A(n7787), .ZN(n7776) );
  OAI211_X1 U9480 ( .C1(n8388), .C2(n8052), .A(n7777), .B(n7776), .ZN(n7778)
         );
  AOI21_X1 U9481 ( .B1(n9905), .B2(n8030), .A(n7778), .ZN(n7779) );
  OAI21_X1 U9482 ( .B1(n7780), .B2(n7983), .A(n7779), .ZN(P2_U3157) );
  AOI21_X1 U9483 ( .B1(n7783), .B2(n7782), .A(n7781), .ZN(n7798) );
  AOI21_X1 U9484 ( .B1(n4363), .B2(n7785), .A(n7784), .ZN(n7786) );
  NOR2_X1 U9485 ( .A1(n7786), .A2(n9844), .ZN(n7796) );
  AOI21_X1 U9486 ( .B1(n9835), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7787), .ZN(
        n7793) );
  OAI21_X1 U9487 ( .B1(n7790), .B2(n7789), .A(n7788), .ZN(n7791) );
  NAND2_X1 U9488 ( .A1(n7791), .A2(n9849), .ZN(n7792) );
  OAI211_X1 U9489 ( .C1(n8139), .C2(n7794), .A(n7793), .B(n7792), .ZN(n7795)
         );
  NOR2_X1 U9490 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  OAI21_X1 U9491 ( .B1(n7798), .B2(n9853), .A(n7797), .ZN(P2_U3192) );
  OAI21_X1 U9492 ( .B1(n7801), .B2(n7800), .A(n7799), .ZN(n7814) );
  AND2_X1 U9493 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8001) );
  AOI21_X1 U9494 ( .B1(n9835), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8001), .ZN(
        n7806) );
  OAI21_X1 U9495 ( .B1(n7803), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7802), .ZN(
        n7804) );
  NAND2_X1 U9496 ( .A1(n9815), .A2(n7804), .ZN(n7805) );
  OAI211_X1 U9497 ( .C1(n8139), .C2(n7807), .A(n7806), .B(n7805), .ZN(n7813)
         );
  AOI21_X1 U9498 ( .B1(n7810), .B2(n7809), .A(n7808), .ZN(n7811) );
  NOR2_X1 U9499 ( .A1(n7811), .A2(n9844), .ZN(n7812) );
  AOI211_X1 U9500 ( .C1(n9849), .C2(n7814), .A(n7813), .B(n7812), .ZN(n7815)
         );
  INV_X1 U9501 ( .A(n7815), .ZN(P2_U3193) );
  AOI21_X1 U9502 ( .B1(n4438), .B2(n7817), .A(n7816), .ZN(n7831) );
  OAI21_X1 U9503 ( .B1(n7820), .B2(n7819), .A(n7818), .ZN(n7829) );
  AOI21_X1 U9504 ( .B1(n4433), .B2(n7822), .A(n7821), .ZN(n7827) );
  NAND2_X1 U9505 ( .A1(n9837), .A2(n7823), .ZN(n7826) );
  NOR2_X1 U9506 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7824), .ZN(n7921) );
  AOI21_X1 U9507 ( .B1(n9835), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7921), .ZN(
        n7825) );
  OAI211_X1 U9508 ( .C1(n7827), .C2(n9853), .A(n7826), .B(n7825), .ZN(n7828)
         );
  AOI21_X1 U9509 ( .B1(n9849), .B2(n7829), .A(n7828), .ZN(n7830) );
  OAI21_X1 U9510 ( .B1(n7831), .B2(n9844), .A(n7830), .ZN(P2_U3194) );
  OAI222_X1 U9511 ( .A1(P1_U3086), .A2(n7834), .B1(n9620), .B2(n7833), .C1(
        n7832), .C2(n9623), .ZN(P1_U3334) );
  INV_X1 U9512 ( .A(n7836), .ZN(n7841) );
  NOR2_X1 U9513 ( .A1(n7837), .A2(n9740), .ZN(n7840) );
  AOI22_X1 U9514 ( .A1(n9767), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8768), .B2(
        n9756), .ZN(n7838) );
  OAI21_X1 U9515 ( .B1(n6500), .B2(n9760), .A(n7838), .ZN(n7839) );
  AOI211_X1 U9516 ( .C1(n7841), .C2(n9470), .A(n7840), .B(n7839), .ZN(n7842)
         );
  OAI21_X1 U9517 ( .B1(n7835), .B2(n9466), .A(n7842), .ZN(P1_U3265) );
  INV_X1 U9518 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9987) );
  OAI222_X1 U9519 ( .A1(n9101), .A2(P1_U3086), .B1(n9620), .B2(n7843), .C1(
        n9987), .C2(n9623), .ZN(P1_U3336) );
  INV_X1 U9520 ( .A(n7844), .ZN(n7879) );
  OAI222_X1 U9521 ( .A1(n7846), .A2(P1_U3086), .B1(n9626), .B2(n7879), .C1(
        n7845), .C2(n9623), .ZN(P1_U3325) );
  INV_X1 U9522 ( .A(n7869), .ZN(n8061) );
  NAND2_X1 U9523 ( .A1(n8061), .A2(n8375), .ZN(n7850) );
  NAND2_X1 U9524 ( .A1(n8191), .A2(n8377), .ZN(n7849) );
  OAI21_X1 U9525 ( .B1(n7854), .B2(n7862), .A(n7853), .ZN(n8415) );
  AOI22_X1 U9526 ( .A1(n7865), .A2(n8396), .B1(n8408), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n7855) );
  OAI21_X1 U9527 ( .B1(n8418), .B2(n8403), .A(n7855), .ZN(n7856) );
  AOI21_X1 U9528 ( .B1(n8415), .B2(n8406), .A(n7856), .ZN(n7857) );
  OAI21_X1 U9529 ( .B1(n8417), .B2(n8408), .A(n7857), .ZN(P2_U3205) );
  INV_X1 U9530 ( .A(n7858), .ZN(n7859) );
  NAND2_X1 U9531 ( .A1(n7859), .A2(n8191), .ZN(n7860) );
  NAND2_X1 U9532 ( .A1(n7861), .A2(n7860), .ZN(n7864) );
  XNOR2_X1 U9533 ( .A(n7862), .B(n5824), .ZN(n7863) );
  XNOR2_X1 U9534 ( .A(n7864), .B(n7863), .ZN(n7874) );
  INV_X1 U9535 ( .A(n7865), .ZN(n7867) );
  INV_X1 U9536 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7866) );
  OAI22_X1 U9537 ( .A1(n7867), .A2(n8040), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7866), .ZN(n7871) );
  OAI22_X1 U9538 ( .A1(n7869), .A2(n8052), .B1(n7868), .B2(n8049), .ZN(n7870)
         );
  AOI211_X1 U9539 ( .C1(n7872), .C2(n8030), .A(n7871), .B(n7870), .ZN(n7873)
         );
  OAI21_X1 U9540 ( .B1(n7874), .B2(n7983), .A(n7873), .ZN(P2_U3160) );
  INV_X1 U9541 ( .A(n7875), .ZN(n9622) );
  OAI222_X1 U9542 ( .A1(n8568), .A2(n9622), .B1(n7877), .B2(P2_U3151), .C1(
        n7876), .C2(n8565), .ZN(P2_U3268) );
  OAI222_X1 U9543 ( .A1(n8555), .A2(n7880), .B1(n8568), .B2(n7879), .C1(
        P2_U3151), .C2(n7878), .ZN(P2_U3265) );
  OAI222_X1 U9544 ( .A1(n9029), .A2(P1_U3086), .B1(n9620), .B2(n7881), .C1(
        n10146), .C2(n9623), .ZN(P1_U3333) );
  INV_X1 U9545 ( .A(n7882), .ZN(n9617) );
  OAI222_X1 U9546 ( .A1(n8568), .A2(n9617), .B1(n7884), .B2(P2_U3151), .C1(
        n7883), .C2(n8565), .ZN(P2_U3266) );
  XOR2_X1 U9547 ( .A(n7885), .B(n7886), .Z(n7891) );
  NAND2_X1 U9548 ( .A1(n8065), .A2(n8038), .ZN(n7887) );
  NAND2_X1 U9549 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8083) );
  OAI211_X1 U9550 ( .C1(n8362), .C2(n8052), .A(n7887), .B(n8083), .ZN(n7889)
         );
  INV_X1 U9551 ( .A(n8368), .ZN(n8544) );
  NOR2_X1 U9552 ( .A1(n8544), .A2(n8058), .ZN(n7888) );
  AOI211_X1 U9553 ( .C1(n8367), .C2(n8055), .A(n7889), .B(n7888), .ZN(n7890)
         );
  OAI21_X1 U9554 ( .B1(n7891), .B2(n7983), .A(n7890), .ZN(P2_U3155) );
  XNOR2_X1 U9555 ( .A(n7927), .B(n7928), .ZN(n7929) );
  XNOR2_X1 U9556 ( .A(n7929), .B(n8248), .ZN(n7897) );
  AOI22_X1 U9557 ( .A1(n8232), .A2(n8043), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7893) );
  NAND2_X1 U9558 ( .A1(n8055), .A2(n8226), .ZN(n7892) );
  OAI211_X1 U9559 ( .C1(n8264), .C2(n8049), .A(n7893), .B(n7892), .ZN(n7894)
         );
  AOI21_X1 U9560 ( .B1(n7895), .B2(n8030), .A(n7894), .ZN(n7896) );
  OAI21_X1 U9561 ( .B1(n7897), .B2(n7983), .A(n7896), .ZN(P2_U3156) );
  INV_X1 U9562 ( .A(n8518), .ZN(n7907) );
  AND3_X1 U9563 ( .A1(n8009), .A2(n7899), .A3(n7898), .ZN(n7900) );
  OAI21_X1 U9564 ( .B1(n7901), .B2(n7900), .A(n5886), .ZN(n7906) );
  NOR2_X1 U9565 ( .A1(n8325), .A2(n8049), .ZN(n7904) );
  OAI21_X1 U9566 ( .B1(n8297), .B2(n8052), .A(n7902), .ZN(n7903) );
  AOI211_X1 U9567 ( .C1(n8302), .C2(n8055), .A(n7904), .B(n7903), .ZN(n7905)
         );
  OAI211_X1 U9568 ( .C1(n7907), .C2(n8058), .A(n7906), .B(n7905), .ZN(P2_U3159) );
  INV_X1 U9569 ( .A(n8437), .ZN(n8267) );
  INV_X1 U9570 ( .A(n7908), .ZN(n7987) );
  AOI21_X1 U9571 ( .B1(n7969), .B2(n7910), .A(n7909), .ZN(n7911) );
  OAI21_X1 U9572 ( .B1(n7987), .B2(n7911), .A(n5886), .ZN(n7915) );
  AOI22_X1 U9573 ( .A1(n8231), .A2(n8043), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7912) );
  OAI21_X1 U9574 ( .B1(n8297), .B2(n8049), .A(n7912), .ZN(n7913) );
  AOI21_X1 U9575 ( .B1(n8265), .B2(n8055), .A(n7913), .ZN(n7914) );
  OAI211_X1 U9576 ( .C1(n8267), .C2(n8058), .A(n7915), .B(n7914), .ZN(P2_U3163) );
  NOR2_X1 U9577 ( .A1(n7916), .A2(n8067), .ZN(n7997) );
  NOR3_X1 U9578 ( .A1(n7998), .A2(n7997), .A3(n7996), .ZN(n7995) );
  AOI21_X1 U9579 ( .B1(n8066), .B2(n7996), .A(n7995), .ZN(n7920) );
  NAND2_X1 U9580 ( .A1(n7918), .A2(n7917), .ZN(n7919) );
  XNOR2_X1 U9581 ( .A(n7920), .B(n7919), .ZN(n7926) );
  NAND2_X1 U9582 ( .A1(n8055), .A2(n8395), .ZN(n7923) );
  AOI21_X1 U9583 ( .B1(n8066), .B2(n8038), .A(n7921), .ZN(n7922) );
  OAI211_X1 U9584 ( .C1(n8390), .C2(n8052), .A(n7923), .B(n7922), .ZN(n7924)
         );
  AOI21_X1 U9585 ( .B1(n9913), .B2(n8030), .A(n7924), .ZN(n7925) );
  OAI21_X1 U9586 ( .B1(n7926), .B2(n7983), .A(n7925), .ZN(P2_U3164) );
  INV_X1 U9587 ( .A(n8206), .ZN(n8489) );
  OAI22_X1 U9588 ( .A1(n7929), .A2(n8248), .B1(n7928), .B2(n7927), .ZN(n7961)
         );
  NAND2_X1 U9589 ( .A1(n7930), .A2(n7931), .ZN(n7962) );
  NOR2_X1 U9590 ( .A1(n7961), .A2(n7962), .ZN(n7960) );
  INV_X1 U9591 ( .A(n7931), .ZN(n7933) );
  NOR3_X1 U9592 ( .A1(n7960), .A2(n7933), .A3(n7932), .ZN(n7936) );
  INV_X1 U9593 ( .A(n7934), .ZN(n7935) );
  OAI21_X1 U9594 ( .B1(n7936), .B2(n7935), .A(n5886), .ZN(n7942) );
  OAI22_X1 U9595 ( .A1(n7938), .A2(n8049), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7937), .ZN(n7940) );
  NOR2_X1 U9596 ( .A1(n8036), .A2(n8052), .ZN(n7939) );
  AOI211_X1 U9597 ( .C1(n8205), .C2(n8055), .A(n7940), .B(n7939), .ZN(n7941)
         );
  OAI211_X1 U9598 ( .C1(n8489), .C2(n8058), .A(n7942), .B(n7941), .ZN(P2_U3165) );
  AOI21_X1 U9599 ( .B1(n7945), .B2(n7944), .A(n7943), .ZN(n7951) );
  NAND2_X1 U9600 ( .A1(n8312), .A2(n8043), .ZN(n7946) );
  NAND2_X1 U9601 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8119) );
  OAI211_X1 U9602 ( .C1(n8362), .C2(n8049), .A(n7946), .B(n8119), .ZN(n7949)
         );
  NOR2_X1 U9603 ( .A1(n7947), .A2(n8058), .ZN(n7948) );
  AOI211_X1 U9604 ( .C1(n8343), .C2(n8055), .A(n7949), .B(n7948), .ZN(n7950)
         );
  OAI21_X1 U9605 ( .B1(n7951), .B2(n7983), .A(n7950), .ZN(P2_U3166) );
  XNOR2_X1 U9606 ( .A(n7952), .B(n8312), .ZN(n7953) );
  XNOR2_X1 U9607 ( .A(n4430), .B(n7953), .ZN(n7959) );
  NAND2_X1 U9608 ( .A1(n8064), .A2(n8043), .ZN(n7954) );
  NAND2_X1 U9609 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8137) );
  OAI211_X1 U9610 ( .C1(n8326), .C2(n8049), .A(n7954), .B(n8137), .ZN(n7957)
         );
  INV_X1 U9611 ( .A(n7955), .ZN(n8530) );
  NOR2_X1 U9612 ( .A1(n8530), .A2(n8058), .ZN(n7956) );
  AOI211_X1 U9613 ( .C1(n8327), .C2(n8055), .A(n7957), .B(n7956), .ZN(n7958)
         );
  OAI21_X1 U9614 ( .B1(n7959), .B2(n7983), .A(n7958), .ZN(P2_U3168) );
  AOI21_X1 U9615 ( .B1(n7962), .B2(n7961), .A(n7960), .ZN(n7968) );
  AOI22_X1 U9616 ( .A1(n8216), .A2(n8038), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7964) );
  NAND2_X1 U9617 ( .A1(n8055), .A2(n8218), .ZN(n7963) );
  OAI211_X1 U9618 ( .C1(n7965), .C2(n8052), .A(n7964), .B(n7963), .ZN(n7966)
         );
  AOI21_X1 U9619 ( .B1(n8220), .B2(n8030), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9620 ( .B1(n7968), .B2(n7983), .A(n7967), .ZN(P2_U3169) );
  OAI211_X1 U9621 ( .C1(n7971), .C2(n7970), .A(n7969), .B(n5886), .ZN(n7975)
         );
  AOI22_X1 U9622 ( .A1(n8062), .A2(n8043), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7972) );
  OAI21_X1 U9623 ( .B1(n8278), .B2(n8049), .A(n7972), .ZN(n7973) );
  AOI21_X1 U9624 ( .B1(n8282), .B2(n8055), .A(n7973), .ZN(n7974) );
  OAI211_X1 U9625 ( .C1(n7976), .C2(n8058), .A(n7975), .B(n7974), .ZN(P2_U3173) );
  XOR2_X1 U9626 ( .A(n7977), .B(n7978), .Z(n7984) );
  NAND2_X1 U9627 ( .A1(n8055), .A2(n8380), .ZN(n7980) );
  AOI22_X1 U9628 ( .A1(n8378), .A2(n8038), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n7979) );
  OAI211_X1 U9629 ( .C1(n8050), .C2(n8052), .A(n7980), .B(n7979), .ZN(n7981)
         );
  AOI21_X1 U9630 ( .B1(n8549), .B2(n8030), .A(n7981), .ZN(n7982) );
  OAI21_X1 U9631 ( .B1(n7984), .B2(n7983), .A(n7982), .ZN(P2_U3174) );
  INV_X1 U9632 ( .A(n8252), .ZN(n8503) );
  NOR3_X1 U9633 ( .A1(n7987), .A2(n7986), .A3(n7985), .ZN(n7990) );
  INV_X1 U9634 ( .A(n7988), .ZN(n7989) );
  OAI21_X1 U9635 ( .B1(n7990), .B2(n7989), .A(n5886), .ZN(n7994) );
  AOI22_X1 U9636 ( .A1(n8062), .A2(n8038), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7991) );
  OAI21_X1 U9637 ( .B1(n8248), .B2(n8052), .A(n7991), .ZN(n7992) );
  AOI21_X1 U9638 ( .B1(n8251), .B2(n8055), .A(n7992), .ZN(n7993) );
  OAI211_X1 U9639 ( .C1(n8503), .C2(n8058), .A(n7994), .B(n7993), .ZN(P2_U3175) );
  INV_X1 U9640 ( .A(n7995), .ZN(n8000) );
  OAI21_X1 U9641 ( .B1(n7998), .B2(n7997), .A(n7996), .ZN(n7999) );
  NAND3_X1 U9642 ( .A1(n8000), .A2(n5886), .A3(n7999), .ZN(n8007) );
  AOI21_X1 U9643 ( .B1(n8038), .B2(n8067), .A(n8001), .ZN(n8002) );
  OAI21_X1 U9644 ( .B1(n8003), .B2(n8052), .A(n8002), .ZN(n8004) );
  AOI21_X1 U9645 ( .B1(n8005), .B2(n8055), .A(n8004), .ZN(n8006) );
  OAI211_X1 U9646 ( .C1(n8008), .C2(n8058), .A(n8007), .B(n8006), .ZN(P2_U3176) );
  OAI21_X1 U9647 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8012) );
  NAND2_X1 U9648 ( .A1(n8012), .A2(n5886), .ZN(n8016) );
  NAND2_X1 U9649 ( .A1(n8311), .A2(n8043), .ZN(n8013) );
  NAND2_X1 U9650 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8154) );
  OAI211_X1 U9651 ( .C1(n8340), .C2(n8049), .A(n8013), .B(n8154), .ZN(n8014)
         );
  AOI21_X1 U9652 ( .B1(n8314), .B2(n8055), .A(n8014), .ZN(n8015) );
  OAI211_X1 U9653 ( .C1(n8017), .C2(n8058), .A(n8016), .B(n8015), .ZN(P2_U3178) );
  INV_X1 U9654 ( .A(n8018), .ZN(n8019) );
  NOR2_X1 U9655 ( .A1(n8020), .A2(n8019), .ZN(n8023) );
  OAI211_X1 U9656 ( .C1(n8023), .C2(n8022), .A(n8021), .B(n5886), .ZN(n8034)
         );
  NAND2_X1 U9657 ( .A1(n8038), .A2(n8072), .ZN(n8025) );
  OAI211_X1 U9658 ( .C1(n8026), .C2(n8052), .A(n8025), .B(n8024), .ZN(n8027)
         );
  INV_X1 U9659 ( .A(n8027), .ZN(n8033) );
  NAND2_X1 U9660 ( .A1(n8055), .A2(n8028), .ZN(n8032) );
  NAND2_X1 U9661 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NAND4_X1 U9662 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(
        P2_U3179) );
  OAI21_X1 U9663 ( .B1(n8036), .B2(n8035), .A(n5885), .ZN(n8037) );
  NAND2_X1 U9664 ( .A1(n8037), .A2(n5886), .ZN(n8045) );
  INV_X1 U9665 ( .A(n8194), .ZN(n8041) );
  AOI22_X1 U9666 ( .A1(n8215), .A2(n8038), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8039) );
  OAI21_X1 U9667 ( .B1(n8041), .B2(n8040), .A(n8039), .ZN(n8042) );
  AOI21_X1 U9668 ( .B1(n8043), .B2(n8191), .A(n8042), .ZN(n8044) );
  OAI211_X1 U9669 ( .C1(n8483), .C2(n8058), .A(n8045), .B(n8044), .ZN(P2_U3180) );
  OAI211_X1 U9670 ( .C1(n8048), .C2(n8047), .A(n8046), .B(n5886), .ZN(n8057)
         );
  NOR2_X1 U9671 ( .A1(n8050), .A2(n8049), .ZN(n8054) );
  NAND2_X1 U9672 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8101) );
  OAI21_X1 U9673 ( .B1(n8326), .B2(n8052), .A(n8101), .ZN(n8053) );
  AOI211_X1 U9674 ( .C1(n8353), .C2(n8055), .A(n8054), .B(n8053), .ZN(n8056)
         );
  OAI211_X1 U9675 ( .C1(n8059), .C2(n8058), .A(n8057), .B(n8056), .ZN(P2_U3181) );
  MUX2_X1 U9676 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8060), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9677 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8061), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9678 ( .A(n8179), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8073), .Z(
        P2_U3519) );
  MUX2_X1 U9679 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8191), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9680 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8202), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9681 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8215), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9682 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8232), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9683 ( .A(n8216), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8073), .Z(
        P2_U3514) );
  MUX2_X1 U9684 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8231), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9685 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8062), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9686 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8063), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9687 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8311), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9688 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8064), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9689 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8312), .S(P2_U3893), .Z(
        P2_U3508) );
  INV_X1 U9690 ( .A(n8326), .ZN(n8350) );
  MUX2_X1 U9691 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8350), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9692 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8376), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9693 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8065), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9694 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8378), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9695 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8066), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9696 ( .A(n8067), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8073), .Z(
        P2_U3501) );
  MUX2_X1 U9697 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8068), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9698 ( .A(n8069), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8073), .Z(
        P2_U3499) );
  MUX2_X1 U9699 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8070), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9700 ( .A(n8071), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8073), .Z(
        P2_U3497) );
  MUX2_X1 U9701 ( .A(n8072), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8073), .Z(
        P2_U3496) );
  MUX2_X1 U9702 ( .A(n8074), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8073), .Z(
        P2_U3495) );
  MUX2_X1 U9703 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8075), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9704 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8076), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9705 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8077), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9706 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8078), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U9707 ( .B1(n4432), .B2(n8079), .A(n4360), .ZN(n8094) );
  OAI21_X1 U9708 ( .B1(n8082), .B2(n8081), .A(n8080), .ZN(n8092) );
  NAND2_X1 U9709 ( .A1(n9835), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8084) );
  OAI211_X1 U9710 ( .C1(n8139), .C2(n8085), .A(n8084), .B(n8083), .ZN(n8091)
         );
  AOI21_X1 U9711 ( .B1(n8088), .B2(n8087), .A(n8086), .ZN(n8089) );
  NOR2_X1 U9712 ( .A1(n8089), .A2(n9853), .ZN(n8090) );
  AOI211_X1 U9713 ( .C1(n9849), .C2(n8092), .A(n8091), .B(n8090), .ZN(n8093)
         );
  OAI21_X1 U9714 ( .B1(n8094), .B2(n9844), .A(n8093), .ZN(P2_U3196) );
  AOI21_X1 U9715 ( .B1(n8096), .B2(n8454), .A(n8095), .ZN(n8111) );
  OAI21_X1 U9716 ( .B1(n8099), .B2(n8098), .A(n8097), .ZN(n8109) );
  NAND2_X1 U9717 ( .A1(n9837), .A2(n8100), .ZN(n8102) );
  OAI211_X1 U9718 ( .C1(n8103), .C2(n9805), .A(n8102), .B(n8101), .ZN(n8108)
         );
  AOI21_X1 U9719 ( .B1(n8352), .B2(n8105), .A(n8104), .ZN(n8106) );
  NOR2_X1 U9720 ( .A1(n8106), .A2(n9844), .ZN(n8107) );
  AOI211_X1 U9721 ( .C1(n9849), .C2(n8109), .A(n8108), .B(n8107), .ZN(n8110)
         );
  OAI21_X1 U9722 ( .B1(n8111), .B2(n9853), .A(n8110), .ZN(P2_U3197) );
  AOI21_X1 U9723 ( .B1(n4424), .B2(n8113), .A(n8112), .ZN(n8128) );
  OAI21_X1 U9724 ( .B1(n8116), .B2(n8115), .A(n8114), .ZN(n8126) );
  INV_X1 U9725 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8117) );
  OR2_X1 U9726 ( .A1(n9805), .A2(n8117), .ZN(n8118) );
  OAI211_X1 U9727 ( .C1(n8139), .C2(n8120), .A(n8119), .B(n8118), .ZN(n8125)
         );
  AOI21_X1 U9728 ( .B1(n4388), .B2(n8122), .A(n8121), .ZN(n8123) );
  NOR2_X1 U9729 ( .A1(n8123), .A2(n9853), .ZN(n8124) );
  AOI211_X1 U9730 ( .C1(n9849), .C2(n8126), .A(n8125), .B(n8124), .ZN(n8127)
         );
  OAI21_X1 U9731 ( .B1(n8128), .B2(n9844), .A(n8127), .ZN(P2_U3198) );
  AOI21_X1 U9732 ( .B1(n8131), .B2(n8130), .A(n8129), .ZN(n8147) );
  OAI21_X1 U9733 ( .B1(n8134), .B2(n8133), .A(n8132), .ZN(n8145) );
  OR2_X1 U9734 ( .A1(n9805), .A2(n8135), .ZN(n8136) );
  OAI211_X1 U9735 ( .C1(n8139), .C2(n8138), .A(n8137), .B(n8136), .ZN(n8144)
         );
  AOI21_X1 U9736 ( .B1(n8450), .B2(n8141), .A(n8140), .ZN(n8142) );
  NOR2_X1 U9737 ( .A1(n8142), .A2(n9853), .ZN(n8143) );
  AOI211_X1 U9738 ( .C1(n9849), .C2(n8145), .A(n8144), .B(n8143), .ZN(n8146)
         );
  OAI21_X1 U9739 ( .B1(n8147), .B2(n9844), .A(n8146), .ZN(P2_U3199) );
  NOR2_X1 U9740 ( .A1(n8149), .A2(n8148), .ZN(n8151) );
  AOI21_X1 U9741 ( .B1(n8151), .B2(P2_U3893), .A(n9837), .ZN(n8160) );
  NOR3_X1 U9742 ( .A1(n8151), .A2(n8150), .A3(n9807), .ZN(n8158) );
  INV_X1 U9743 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9946) );
  INV_X1 U9744 ( .A(n8161), .ZN(n8162) );
  NOR2_X1 U9745 ( .A1(n8163), .A2(n8162), .ZN(n8464) );
  NOR2_X1 U9746 ( .A1(n8164), .A2(n8227), .ZN(n8171) );
  AOI21_X1 U9747 ( .B1(n8464), .B2(n8401), .A(n8171), .ZN(n8167) );
  NAND2_X1 U9748 ( .A1(n8408), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8165) );
  OAI211_X1 U9749 ( .C1(n8466), .C2(n8403), .A(n8167), .B(n8165), .ZN(P2_U3202) );
  NAND2_X1 U9750 ( .A1(n8408), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8166) );
  OAI211_X1 U9751 ( .C1(n8469), .C2(n8403), .A(n8167), .B(n8166), .ZN(P2_U3203) );
  NAND2_X1 U9752 ( .A1(n8168), .A2(n8401), .ZN(n8173) );
  NOR2_X1 U9753 ( .A1(n8169), .A2(n8403), .ZN(n8170) );
  AOI211_X1 U9754 ( .C1(n8408), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8171), .B(
        n8170), .ZN(n8172) );
  OAI211_X1 U9755 ( .C1(n8175), .C2(n8174), .A(n8173), .B(n8172), .ZN(P2_U3204) );
  XOR2_X1 U9756 ( .A(n8177), .B(n8176), .Z(n8474) );
  INV_X1 U9757 ( .A(n8474), .ZN(n8186) );
  INV_X1 U9758 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8181) );
  XNOR2_X1 U9759 ( .A(n8178), .B(n8177), .ZN(n8180) );
  AOI222_X1 U9760 ( .A1(n8392), .A2(n8180), .B1(n8179), .B2(n8375), .C1(n8202), 
        .C2(n8377), .ZN(n8471) );
  MUX2_X1 U9761 ( .A(n8181), .B(n8471), .S(n8401), .Z(n8185) );
  AOI22_X1 U9762 ( .A1(n8183), .A2(n8381), .B1(n8396), .B2(n8182), .ZN(n8184)
         );
  OAI211_X1 U9763 ( .C1(n8186), .C2(n8384), .A(n8185), .B(n8184), .ZN(P2_U3206) );
  XNOR2_X1 U9764 ( .A(n8187), .B(n8188), .ZN(n8480) );
  INV_X1 U9765 ( .A(n8480), .ZN(n8198) );
  INV_X1 U9766 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8193) );
  XNOR2_X1 U9767 ( .A(n8190), .B(n8189), .ZN(n8192) );
  AOI222_X1 U9768 ( .A1(n8392), .A2(n8192), .B1(n8215), .B2(n8377), .C1(n8191), 
        .C2(n8375), .ZN(n8478) );
  MUX2_X1 U9769 ( .A(n8193), .B(n8478), .S(n8401), .Z(n8197) );
  AOI22_X1 U9770 ( .A1(n8195), .A2(n8381), .B1(n8396), .B2(n8194), .ZN(n8196)
         );
  OAI211_X1 U9771 ( .C1(n8198), .C2(n8384), .A(n8197), .B(n8196), .ZN(P2_U3207) );
  XNOR2_X1 U9772 ( .A(n8199), .B(n8200), .ZN(n8486) );
  INV_X1 U9773 ( .A(n8486), .ZN(n8209) );
  INV_X1 U9774 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8204) );
  XNOR2_X1 U9775 ( .A(n8201), .B(n8200), .ZN(n8203) );
  AOI222_X1 U9776 ( .A1(n8392), .A2(n8203), .B1(n8202), .B2(n8375), .C1(n8232), 
        .C2(n8377), .ZN(n8484) );
  MUX2_X1 U9777 ( .A(n8204), .B(n8484), .S(n8401), .Z(n8208) );
  AOI22_X1 U9778 ( .A1(n8206), .A2(n8381), .B1(n8396), .B2(n8205), .ZN(n8207)
         );
  OAI211_X1 U9779 ( .C1(n8209), .C2(n8384), .A(n8208), .B(n8207), .ZN(P2_U3208) );
  NAND2_X1 U9780 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  XOR2_X1 U9781 ( .A(n8213), .B(n8212), .Z(n8492) );
  INV_X1 U9782 ( .A(n8492), .ZN(n8224) );
  XNOR2_X1 U9783 ( .A(n8214), .B(n8213), .ZN(n8217) );
  AOI222_X1 U9784 ( .A1(n8392), .A2(n8217), .B1(n8216), .B2(n8377), .C1(n8215), 
        .C2(n8375), .ZN(n8490) );
  AOI22_X1 U9785 ( .A1(n8220), .A2(n8219), .B1(n8396), .B2(n8218), .ZN(n8221)
         );
  AOI21_X1 U9786 ( .B1(n8490), .B2(n8221), .A(n8408), .ZN(n8222) );
  AOI21_X1 U9787 ( .B1(n8408), .B2(P2_REG2_REG_24__SCAN_IN), .A(n8222), .ZN(
        n8223) );
  OAI21_X1 U9788 ( .B1(n8384), .B2(n8224), .A(n8223), .ZN(P2_U3209) );
  XOR2_X1 U9789 ( .A(n8225), .B(n8229), .Z(n8498) );
  INV_X1 U9790 ( .A(n8226), .ZN(n8228) );
  OAI22_X1 U9791 ( .A1(n8501), .A2(n8403), .B1(n8228), .B2(n8227), .ZN(n8236)
         );
  XNOR2_X1 U9792 ( .A(n8230), .B(n8229), .ZN(n8233) );
  AOI222_X1 U9793 ( .A1(n8392), .A2(n8233), .B1(n8232), .B2(n8375), .C1(n8231), 
        .C2(n8377), .ZN(n8496) );
  INV_X1 U9794 ( .A(n8496), .ZN(n8234) );
  MUX2_X1 U9795 ( .A(P2_REG2_REG_23__SCAN_IN), .B(n8234), .S(n8401), .Z(n8235)
         );
  AOI211_X1 U9796 ( .C1(n8406), .C2(n8498), .A(n8236), .B(n8235), .ZN(n8237)
         );
  INV_X1 U9797 ( .A(n8237), .ZN(P2_U3210) );
  XNOR2_X1 U9798 ( .A(n8238), .B(n8243), .ZN(n8504) );
  INV_X1 U9799 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8250) );
  INV_X1 U9800 ( .A(n8243), .ZN(n8240) );
  INV_X1 U9801 ( .A(n8244), .ZN(n8239) );
  NOR2_X1 U9802 ( .A1(n8240), .A2(n8239), .ZN(n8246) );
  INV_X1 U9803 ( .A(n8260), .ZN(n8242) );
  NAND2_X1 U9804 ( .A1(n8241), .A2(n8242), .ZN(n8262) );
  AOI21_X1 U9805 ( .B1(n8262), .B2(n8244), .A(n8243), .ZN(n8245) );
  AOI21_X1 U9806 ( .B1(n8246), .B2(n8262), .A(n8245), .ZN(n8247) );
  INV_X1 U9807 ( .A(n8502), .ZN(n8249) );
  MUX2_X1 U9808 ( .A(n8250), .B(n8249), .S(n8401), .Z(n8254) );
  AOI22_X1 U9809 ( .A1(n8252), .A2(n8381), .B1(n8396), .B2(n8251), .ZN(n8253)
         );
  OAI211_X1 U9810 ( .C1(n8504), .C2(n8384), .A(n8254), .B(n8253), .ZN(P2_U3211) );
  NAND2_X1 U9811 ( .A1(n8256), .A2(n8255), .ZN(n8257) );
  XOR2_X1 U9812 ( .A(n8260), .B(n8257), .Z(n8510) );
  NAND3_X1 U9813 ( .A1(n8258), .A2(n8260), .A3(n8259), .ZN(n8261) );
  AND2_X1 U9814 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  OAI222_X1 U9815 ( .A1(n8387), .A2(n8297), .B1(n8389), .B2(n8264), .C1(n8323), 
        .C2(n8263), .ZN(n8436) );
  AOI22_X1 U9816 ( .A1(n8408), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8396), .B2(
        n8265), .ZN(n8266) );
  OAI21_X1 U9817 ( .B1(n8267), .B2(n8403), .A(n8266), .ZN(n8268) );
  AOI21_X1 U9818 ( .B1(n8436), .B2(n8401), .A(n8268), .ZN(n8269) );
  OAI21_X1 U9819 ( .B1(n8384), .B2(n8510), .A(n8269), .ZN(P2_U3212) );
  AND2_X1 U9820 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  XNOR2_X1 U9821 ( .A(n8272), .B(n8273), .ZN(n8515) );
  INV_X1 U9822 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8281) );
  INV_X1 U9823 ( .A(n8258), .ZN(n8276) );
  AOI21_X1 U9824 ( .B1(n8292), .B2(n8274), .A(n8273), .ZN(n8275) );
  NOR2_X1 U9825 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  OAI222_X1 U9826 ( .A1(n8389), .A2(n8279), .B1(n8387), .B2(n8278), .C1(n8323), 
        .C2(n8277), .ZN(n8511) );
  INV_X1 U9827 ( .A(n8511), .ZN(n8280) );
  MUX2_X1 U9828 ( .A(n8281), .B(n8280), .S(n8401), .Z(n8284) );
  AOI22_X1 U9829 ( .A1(n8513), .A2(n8381), .B1(n8396), .B2(n8282), .ZN(n8283)
         );
  OAI211_X1 U9830 ( .C1(n8515), .C2(n8384), .A(n8284), .B(n8283), .ZN(P2_U3213) );
  NAND2_X1 U9831 ( .A1(n8285), .A2(n8286), .ZN(n8319) );
  NAND2_X1 U9832 ( .A1(n8319), .A2(n8287), .ZN(n8306) );
  NAND2_X1 U9833 ( .A1(n8306), .A2(n8288), .ZN(n8290) );
  NAND2_X1 U9834 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  XOR2_X1 U9835 ( .A(n8293), .B(n8291), .Z(n8520) );
  INV_X1 U9836 ( .A(n8292), .ZN(n8296) );
  AOI21_X1 U9837 ( .B1(n8308), .B2(n8294), .A(n8293), .ZN(n8295) );
  NOR3_X1 U9838 ( .A1(n8296), .A2(n8295), .A3(n8323), .ZN(n8299) );
  OAI22_X1 U9839 ( .A1(n8325), .A2(n8387), .B1(n8297), .B2(n8389), .ZN(n8298)
         );
  OR2_X1 U9840 ( .A1(n8299), .A2(n8298), .ZN(n8516) );
  INV_X1 U9841 ( .A(n8516), .ZN(n8300) );
  MUX2_X1 U9842 ( .A(n8301), .B(n8300), .S(n8401), .Z(n8304) );
  AOI22_X1 U9843 ( .A1(n8518), .A2(n8381), .B1(n8396), .B2(n8302), .ZN(n8303)
         );
  OAI211_X1 U9844 ( .C1(n8520), .C2(n8384), .A(n8304), .B(n8303), .ZN(P2_U3214) );
  NAND2_X1 U9845 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  XOR2_X1 U9846 ( .A(n8309), .B(n8307), .Z(n8524) );
  INV_X1 U9847 ( .A(n8524), .ZN(n8317) );
  OAI21_X1 U9848 ( .B1(n8310), .B2(n8309), .A(n8308), .ZN(n8313) );
  AOI222_X1 U9849 ( .A1(n8392), .A2(n8313), .B1(n8312), .B2(n8377), .C1(n8311), 
        .C2(n8375), .ZN(n8521) );
  MUX2_X1 U9850 ( .A(n10121), .B(n8521), .S(n8401), .Z(n8316) );
  AOI22_X1 U9851 ( .A1(n8522), .A2(n8381), .B1(n8396), .B2(n8314), .ZN(n8315)
         );
  OAI211_X1 U9852 ( .C1(n8317), .C2(n8384), .A(n8316), .B(n8315), .ZN(P2_U3215) );
  NAND2_X1 U9853 ( .A1(n8319), .A2(n8318), .ZN(n8320) );
  XNOR2_X1 U9854 ( .A(n8320), .B(n8321), .ZN(n8449) );
  INV_X1 U9855 ( .A(n8449), .ZN(n8331) );
  XNOR2_X1 U9856 ( .A(n8322), .B(n8321), .ZN(n8324) );
  OAI222_X1 U9857 ( .A1(n8387), .A2(n8326), .B1(n8389), .B2(n8325), .C1(n8324), 
        .C2(n8323), .ZN(n8448) );
  AOI22_X1 U9858 ( .A1(n8408), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8327), .B2(
        n8396), .ZN(n8328) );
  OAI21_X1 U9859 ( .B1(n8530), .B2(n8403), .A(n8328), .ZN(n8329) );
  AOI21_X1 U9860 ( .B1(n8448), .B2(n8401), .A(n8329), .ZN(n8330) );
  OAI21_X1 U9861 ( .B1(n8331), .B2(n8384), .A(n8330), .ZN(P2_U3216) );
  XNOR2_X1 U9862 ( .A(n8285), .B(n8332), .ZN(n8535) );
  AND2_X1 U9863 ( .A1(n8333), .A2(n8334), .ZN(n8337) );
  OAI211_X1 U9864 ( .C1(n8337), .C2(n8336), .A(n8335), .B(n8392), .ZN(n8339)
         );
  OR2_X1 U9865 ( .A1(n8362), .A2(n8387), .ZN(n8338) );
  OAI211_X1 U9866 ( .C1(n8340), .C2(n8389), .A(n8339), .B(n8338), .ZN(n8531)
         );
  INV_X1 U9867 ( .A(n8531), .ZN(n8341) );
  MUX2_X1 U9868 ( .A(n8342), .B(n8341), .S(n8401), .Z(n8345) );
  AOI22_X1 U9869 ( .A1(n8533), .A2(n8381), .B1(n8396), .B2(n8343), .ZN(n8344)
         );
  OAI211_X1 U9870 ( .C1(n8535), .C2(n8384), .A(n8345), .B(n8344), .ZN(P2_U3217) );
  XNOR2_X1 U9871 ( .A(n8346), .B(n8348), .ZN(n8541) );
  AND2_X1 U9872 ( .A1(n8360), .A2(n8347), .ZN(n8349) );
  OAI21_X1 U9873 ( .B1(n8349), .B2(n8348), .A(n8333), .ZN(n8351) );
  AOI222_X1 U9874 ( .A1(n8392), .A2(n8351), .B1(n8350), .B2(n8375), .C1(n8376), 
        .C2(n8377), .ZN(n8536) );
  MUX2_X1 U9875 ( .A(n8352), .B(n8536), .S(n8401), .Z(n8355) );
  AOI22_X1 U9876 ( .A1(n8538), .A2(n8381), .B1(n8396), .B2(n8353), .ZN(n8354)
         );
  OAI211_X1 U9877 ( .C1(n8541), .C2(n8384), .A(n8355), .B(n8354), .ZN(P2_U3218) );
  XNOR2_X1 U9878 ( .A(n8356), .B(n8358), .ZN(n8545) );
  NAND2_X1 U9879 ( .A1(n8373), .A2(n8357), .ZN(n8359) );
  NAND2_X1 U9880 ( .A1(n8359), .A2(n8358), .ZN(n8361) );
  NAND3_X1 U9881 ( .A1(n8361), .A2(n8392), .A3(n8360), .ZN(n8365) );
  OAI22_X1 U9882 ( .A1(n8362), .A2(n8389), .B1(n8390), .B2(n8387), .ZN(n8363)
         );
  INV_X1 U9883 ( .A(n8363), .ZN(n8364) );
  NAND2_X1 U9884 ( .A1(n8365), .A2(n8364), .ZN(n8542) );
  MUX2_X1 U9885 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n8542), .S(n8401), .Z(n8366)
         );
  INV_X1 U9886 ( .A(n8366), .ZN(n8370) );
  AOI22_X1 U9887 ( .A1(n8368), .A2(n8381), .B1(n8396), .B2(n8367), .ZN(n8369)
         );
  OAI211_X1 U9888 ( .C1(n8545), .C2(n8384), .A(n8370), .B(n8369), .ZN(P2_U3219) );
  XNOR2_X1 U9889 ( .A(n8371), .B(n8372), .ZN(n8553) );
  OAI21_X1 U9890 ( .B1(n4425), .B2(n8374), .A(n8373), .ZN(n8379) );
  AOI222_X1 U9891 ( .A1(n8392), .A2(n8379), .B1(n8378), .B2(n8377), .C1(n8376), 
        .C2(n8375), .ZN(n8548) );
  MUX2_X1 U9892 ( .A(n9843), .B(n8548), .S(n8401), .Z(n8383) );
  AOI22_X1 U9893 ( .A1(n8549), .A2(n8381), .B1(n8396), .B2(n8380), .ZN(n8382)
         );
  OAI211_X1 U9894 ( .C1(n8553), .C2(n8384), .A(n8383), .B(n8382), .ZN(P2_U3220) );
  XNOR2_X1 U9895 ( .A(n8386), .B(n8385), .ZN(n8393) );
  OAI22_X1 U9896 ( .A1(n8390), .A2(n8389), .B1(n8388), .B2(n8387), .ZN(n8391)
         );
  AOI21_X1 U9897 ( .B1(n8393), .B2(n8392), .A(n8391), .ZN(n9917) );
  INV_X1 U9898 ( .A(n9917), .ZN(n8394) );
  AOI21_X1 U9899 ( .B1(n8396), .B2(n8395), .A(n8394), .ZN(n8409) );
  INV_X1 U9900 ( .A(n8397), .ZN(n8398) );
  AOI21_X1 U9901 ( .B1(n8400), .B2(n8399), .A(n8398), .ZN(n9916) );
  INV_X1 U9902 ( .A(n9913), .ZN(n8404) );
  INV_X1 U9903 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8402) );
  OAI22_X1 U9904 ( .A1(n8404), .A2(n8403), .B1(n8402), .B2(n8401), .ZN(n8405)
         );
  AOI21_X1 U9905 ( .B1(n9916), .B2(n8406), .A(n8405), .ZN(n8407) );
  OAI21_X1 U9906 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(P2_U3221) );
  NAND2_X1 U9907 ( .A1(n8410), .A2(n6594), .ZN(n8411) );
  NAND2_X1 U9908 ( .A1(n8464), .A2(n9938), .ZN(n8413) );
  OAI211_X1 U9909 ( .C1(n9938), .C2(n5542), .A(n8411), .B(n8413), .ZN(P2_U3490) );
  NAND2_X1 U9910 ( .A1(n8412), .A2(n6594), .ZN(n8414) );
  OAI211_X1 U9911 ( .C1(n9938), .C2(n5554), .A(n8414), .B(n8413), .ZN(P2_U3489) );
  NAND2_X1 U9912 ( .A1(n8415), .A2(n9915), .ZN(n8416) );
  OAI211_X1 U9913 ( .C1(n8418), .C2(n9893), .A(n8417), .B(n8416), .ZN(n8470)
         );
  MUX2_X1 U9914 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8470), .S(n9938), .Z(
        P2_U3487) );
  MUX2_X1 U9915 ( .A(n8419), .B(n8471), .S(n9938), .Z(n8421) );
  NAND2_X1 U9916 ( .A1(n8474), .A2(n8445), .ZN(n8420) );
  OAI211_X1 U9917 ( .C1(n8477), .C2(n8457), .A(n8421), .B(n8420), .ZN(P2_U3486) );
  INV_X1 U9918 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8422) );
  MUX2_X1 U9919 ( .A(n8422), .B(n8478), .S(n9938), .Z(n8424) );
  NAND2_X1 U9920 ( .A1(n8480), .A2(n8445), .ZN(n8423) );
  OAI211_X1 U9921 ( .C1(n8483), .C2(n8457), .A(n8424), .B(n8423), .ZN(P2_U3485) );
  MUX2_X1 U9922 ( .A(n8425), .B(n8484), .S(n9938), .Z(n8427) );
  NAND2_X1 U9923 ( .A1(n8486), .A2(n8445), .ZN(n8426) );
  OAI211_X1 U9924 ( .C1(n8489), .C2(n8457), .A(n8427), .B(n8426), .ZN(P2_U3484) );
  MUX2_X1 U9925 ( .A(n8428), .B(n8490), .S(n9938), .Z(n8430) );
  NAND2_X1 U9926 ( .A1(n8492), .A2(n8445), .ZN(n8429) );
  OAI211_X1 U9927 ( .C1(n8495), .C2(n8457), .A(n8430), .B(n8429), .ZN(P2_U3483) );
  MUX2_X1 U9928 ( .A(n8431), .B(n8496), .S(n9938), .Z(n8433) );
  NAND2_X1 U9929 ( .A1(n8498), .A2(n8445), .ZN(n8432) );
  OAI211_X1 U9930 ( .C1(n8501), .C2(n8457), .A(n8433), .B(n8432), .ZN(P2_U3482) );
  MUX2_X1 U9931 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8502), .S(n9938), .Z(n8435)
         );
  INV_X1 U9932 ( .A(n8445), .ZN(n8462) );
  OAI22_X1 U9933 ( .A1(n8504), .A2(n8462), .B1(n8503), .B2(n8457), .ZN(n8434)
         );
  OR2_X1 U9934 ( .A1(n8435), .A2(n8434), .ZN(P2_U3481) );
  INV_X1 U9935 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8438) );
  AOI21_X1 U9936 ( .B1(n9914), .B2(n8437), .A(n8436), .ZN(n8507) );
  MUX2_X1 U9937 ( .A(n8438), .B(n8507), .S(n9938), .Z(n8439) );
  OAI21_X1 U9938 ( .B1(n8462), .B2(n8510), .A(n8439), .ZN(P2_U3480) );
  MUX2_X1 U9939 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8511), .S(n9938), .Z(n8440)
         );
  AOI21_X1 U9940 ( .B1(n6594), .B2(n8513), .A(n8440), .ZN(n8441) );
  OAI21_X1 U9941 ( .B1(n8462), .B2(n8515), .A(n8441), .ZN(P2_U3479) );
  MUX2_X1 U9942 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8516), .S(n9938), .Z(n8442)
         );
  AOI21_X1 U9943 ( .B1(n6594), .B2(n8518), .A(n8442), .ZN(n8443) );
  OAI21_X1 U9944 ( .B1(n8520), .B2(n8462), .A(n8443), .ZN(P2_U3478) );
  MUX2_X1 U9945 ( .A(n8444), .B(n8521), .S(n9938), .Z(n8447) );
  AOI22_X1 U9946 ( .A1(n8524), .A2(n8445), .B1(n6594), .B2(n8522), .ZN(n8446)
         );
  NAND2_X1 U9947 ( .A1(n8447), .A2(n8446), .ZN(P2_U3477) );
  AOI21_X1 U9948 ( .B1(n9915), .B2(n8449), .A(n8448), .ZN(n8527) );
  MUX2_X1 U9949 ( .A(n8450), .B(n8527), .S(n9938), .Z(n8451) );
  OAI21_X1 U9950 ( .B1(n8530), .B2(n8457), .A(n8451), .ZN(P2_U3476) );
  MUX2_X1 U9951 ( .A(n8531), .B(P2_REG1_REG_16__SCAN_IN), .S(n9935), .Z(n8452)
         );
  AOI21_X1 U9952 ( .B1(n6594), .B2(n8533), .A(n8452), .ZN(n8453) );
  OAI21_X1 U9953 ( .B1(n8535), .B2(n8462), .A(n8453), .ZN(P2_U3475) );
  MUX2_X1 U9954 ( .A(n8454), .B(n8536), .S(n9938), .Z(n8456) );
  NAND2_X1 U9955 ( .A1(n8538), .A2(n6594), .ZN(n8455) );
  OAI211_X1 U9956 ( .C1(n8462), .C2(n8541), .A(n8456), .B(n8455), .ZN(P2_U3474) );
  MUX2_X1 U9957 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8542), .S(n9938), .Z(n8459)
         );
  OAI22_X1 U9958 ( .A1(n8545), .A2(n8462), .B1(n8544), .B2(n8457), .ZN(n8458)
         );
  OR2_X1 U9959 ( .A1(n8459), .A2(n8458), .ZN(P2_U3473) );
  MUX2_X1 U9960 ( .A(n9840), .B(n8548), .S(n9938), .Z(n8461) );
  NAND2_X1 U9961 ( .A1(n8549), .A2(n6594), .ZN(n8460) );
  OAI211_X1 U9962 ( .C1(n8553), .C2(n8462), .A(n8461), .B(n8460), .ZN(P2_U3472) );
  MUX2_X1 U9963 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8463), .S(n9938), .Z(
        P2_U3459) );
  NAND2_X1 U9964 ( .A1(n8464), .A2(n9919), .ZN(n8467) );
  NAND2_X1 U9965 ( .A1(n9921), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8465) );
  OAI211_X1 U9966 ( .C1(n8466), .C2(n8543), .A(n8467), .B(n8465), .ZN(P2_U3458) );
  NAND2_X1 U9967 ( .A1(n9921), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8468) );
  OAI211_X1 U9968 ( .C1(n8469), .C2(n8543), .A(n8468), .B(n8467), .ZN(P2_U3457) );
  MUX2_X1 U9969 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8470), .S(n9919), .Z(
        P2_U3455) );
  INV_X1 U9970 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8472) );
  MUX2_X1 U9971 ( .A(n8472), .B(n8471), .S(n9919), .Z(n8476) );
  NAND2_X1 U9972 ( .A1(n8474), .A2(n8523), .ZN(n8475) );
  OAI211_X1 U9973 ( .C1(n8477), .C2(n8543), .A(n8476), .B(n8475), .ZN(P2_U3454) );
  MUX2_X1 U9974 ( .A(n8479), .B(n8478), .S(n9919), .Z(n8482) );
  NAND2_X1 U9975 ( .A1(n8480), .A2(n8523), .ZN(n8481) );
  OAI211_X1 U9976 ( .C1(n8483), .C2(n8543), .A(n8482), .B(n8481), .ZN(P2_U3453) );
  INV_X1 U9977 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8485) );
  MUX2_X1 U9978 ( .A(n8485), .B(n8484), .S(n9919), .Z(n8488) );
  NAND2_X1 U9979 ( .A1(n8486), .A2(n8523), .ZN(n8487) );
  OAI211_X1 U9980 ( .C1(n8489), .C2(n8543), .A(n8488), .B(n8487), .ZN(P2_U3452) );
  INV_X1 U9981 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8491) );
  MUX2_X1 U9982 ( .A(n8491), .B(n8490), .S(n9919), .Z(n8494) );
  NAND2_X1 U9983 ( .A1(n8492), .A2(n8523), .ZN(n8493) );
  OAI211_X1 U9984 ( .C1(n8495), .C2(n8543), .A(n8494), .B(n8493), .ZN(P2_U3451) );
  INV_X1 U9985 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8497) );
  MUX2_X1 U9986 ( .A(n8497), .B(n8496), .S(n9919), .Z(n8500) );
  NAND2_X1 U9987 ( .A1(n8498), .A2(n8523), .ZN(n8499) );
  OAI211_X1 U9988 ( .C1(n8501), .C2(n8543), .A(n8500), .B(n8499), .ZN(P2_U3450) );
  MUX2_X1 U9989 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8502), .S(n9919), .Z(n8506)
         );
  OAI22_X1 U9990 ( .A1(n8504), .A2(n8552), .B1(n8503), .B2(n8543), .ZN(n8505)
         );
  OR2_X1 U9991 ( .A1(n8506), .A2(n8505), .ZN(P2_U3449) );
  INV_X1 U9992 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8508) );
  MUX2_X1 U9993 ( .A(n8508), .B(n8507), .S(n9919), .Z(n8509) );
  OAI21_X1 U9994 ( .B1(n8510), .B2(n8552), .A(n8509), .ZN(P2_U3448) );
  MUX2_X1 U9995 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8511), .S(n9919), .Z(n8512)
         );
  AOI21_X1 U9996 ( .B1(n6577), .B2(n8513), .A(n8512), .ZN(n8514) );
  OAI21_X1 U9997 ( .B1(n8552), .B2(n8515), .A(n8514), .ZN(P2_U3447) );
  MUX2_X1 U9998 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8516), .S(n9919), .Z(n8517)
         );
  AOI21_X1 U9999 ( .B1(n6577), .B2(n8518), .A(n8517), .ZN(n8519) );
  OAI21_X1 U10000 ( .B1(n8520), .B2(n8552), .A(n8519), .ZN(P2_U3446) );
  INV_X1 U10001 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10115) );
  MUX2_X1 U10002 ( .A(n10115), .B(n8521), .S(n9919), .Z(n8526) );
  AOI22_X1 U10003 ( .A1(n8524), .A2(n8523), .B1(n6577), .B2(n8522), .ZN(n8525)
         );
  NAND2_X1 U10004 ( .A1(n8526), .A2(n8525), .ZN(P2_U3444) );
  INV_X1 U10005 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8528) );
  MUX2_X1 U10006 ( .A(n8528), .B(n8527), .S(n9919), .Z(n8529) );
  OAI21_X1 U10007 ( .B1(n8530), .B2(n8543), .A(n8529), .ZN(P2_U3441) );
  MUX2_X1 U10008 ( .A(n8531), .B(P2_REG0_REG_16__SCAN_IN), .S(n9921), .Z(n8532) );
  AOI21_X1 U10009 ( .B1(n6577), .B2(n8533), .A(n8532), .ZN(n8534) );
  OAI21_X1 U10010 ( .B1(n8535), .B2(n8552), .A(n8534), .ZN(P2_U3438) );
  INV_X1 U10011 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8537) );
  MUX2_X1 U10012 ( .A(n8537), .B(n8536), .S(n9919), .Z(n8540) );
  NAND2_X1 U10013 ( .A1(n8538), .A2(n6577), .ZN(n8539) );
  OAI211_X1 U10014 ( .C1(n8541), .C2(n8552), .A(n8540), .B(n8539), .ZN(
        P2_U3435) );
  MUX2_X1 U10015 ( .A(n8542), .B(P2_REG0_REG_14__SCAN_IN), .S(n9921), .Z(n8547) );
  OAI22_X1 U10016 ( .A1(n8545), .A2(n8552), .B1(n8544), .B2(n8543), .ZN(n8546)
         );
  OR2_X1 U10017 ( .A1(n8547), .A2(n8546), .ZN(P2_U3432) );
  INV_X1 U10018 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9999) );
  MUX2_X1 U10019 ( .A(n9999), .B(n8548), .S(n9919), .Z(n8551) );
  NAND2_X1 U10020 ( .A1(n8549), .A2(n6577), .ZN(n8550) );
  OAI211_X1 U10021 ( .C1(n8553), .C2(n8552), .A(n8551), .B(n8550), .ZN(
        P2_U3429) );
  INV_X1 U10022 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8554) );
  NAND3_X1 U10023 ( .A1(n8554), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8557) );
  OAI22_X1 U10024 ( .A1(n4968), .A2(n8557), .B1(n8556), .B2(n8555), .ZN(n8558)
         );
  AOI21_X1 U10025 ( .B1(n9609), .B2(n8559), .A(n8558), .ZN(n8560) );
  INV_X1 U10026 ( .A(n8560), .ZN(P2_U3264) );
  INV_X1 U10027 ( .A(n6391), .ZN(n9619) );
  AOI21_X1 U10028 ( .B1(n8562), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8561), .ZN(
        n8563) );
  OAI21_X1 U10029 ( .B1(n9619), .B2(n8568), .A(n8563), .ZN(P2_U3267) );
  INV_X1 U10030 ( .A(n8564), .ZN(n9625) );
  OAI222_X1 U10031 ( .A1(n8568), .A2(n9625), .B1(P2_U3151), .B2(n8567), .C1(
        n8566), .C2(n8565), .ZN(P2_U3269) );
  MUX2_X1 U10032 ( .A(n8569), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10033 ( .B1(n8575), .B2(n8577), .A(n8570), .ZN(n8571) );
  INV_X1 U10034 ( .A(n8572), .ZN(n8576) );
  AOI21_X1 U10035 ( .B1(n8577), .B2(n8575), .A(n8576), .ZN(n8574) );
  NAND3_X1 U10036 ( .A1(n8577), .A2(n8576), .A3(n8575), .ZN(n8578) );
  AOI22_X1 U10037 ( .A1(n9651), .A2(n8709), .B1(n6895), .B2(n9189), .ZN(n8581)
         );
  XNOR2_X1 U10038 ( .A(n8581), .B(n8695), .ZN(n8582) );
  NAND2_X1 U10039 ( .A1(n8583), .A2(n8582), .ZN(n8586) );
  OAI22_X1 U10040 ( .A1(n9780), .A2(n8764), .B1(n8585), .B2(n8677), .ZN(n9645)
         );
  INV_X1 U10041 ( .A(n8586), .ZN(n8587) );
  NAND2_X1 U10042 ( .A1(n8592), .A2(n8709), .ZN(n8589) );
  NAND2_X1 U10043 ( .A1(n9188), .A2(n6895), .ZN(n8588) );
  NAND2_X1 U10044 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  XNOR2_X1 U10045 ( .A(n8590), .B(n8761), .ZN(n8594) );
  AND2_X1 U10046 ( .A1(n9188), .A2(n8758), .ZN(n8591) );
  AOI21_X1 U10047 ( .B1(n8592), .B2(n6895), .A(n8591), .ZN(n8593) );
  NOR2_X1 U10048 ( .A1(n8594), .A2(n8593), .ZN(n8880) );
  AND2_X1 U10049 ( .A1(n8594), .A2(n8593), .ZN(n8882) );
  AOI22_X1 U10050 ( .A1(n9785), .A2(n6895), .B1(n8758), .B2(n9187), .ZN(n8598)
         );
  NAND2_X1 U10051 ( .A1(n9785), .A2(n8709), .ZN(n8596) );
  NAND2_X1 U10052 ( .A1(n9187), .A2(n6895), .ZN(n8595) );
  NAND2_X1 U10053 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  XNOR2_X1 U10054 ( .A(n8597), .B(n8695), .ZN(n8600) );
  XOR2_X1 U10055 ( .A(n8598), .B(n8600), .Z(n8789) );
  INV_X1 U10056 ( .A(n8598), .ZN(n8599) );
  NAND2_X1 U10057 ( .A1(n8867), .A2(n8709), .ZN(n8602) );
  OR2_X1 U10058 ( .A1(n8790), .A2(n8764), .ZN(n8601) );
  NAND2_X1 U10059 ( .A1(n8602), .A2(n8601), .ZN(n8603) );
  XNOR2_X1 U10060 ( .A(n8603), .B(n8695), .ZN(n8604) );
  AOI22_X1 U10061 ( .A1(n8867), .A2(n6895), .B1(n8758), .B2(n9186), .ZN(n8605)
         );
  XNOR2_X1 U10062 ( .A(n8604), .B(n8605), .ZN(n8861) );
  NAND2_X1 U10063 ( .A1(n8862), .A2(n8861), .ZN(n8608) );
  INV_X1 U10064 ( .A(n8604), .ZN(n8606) );
  NAND2_X1 U10065 ( .A1(n8606), .A2(n8605), .ZN(n8607) );
  NAND2_X1 U10066 ( .A1(n8608), .A2(n8607), .ZN(n8730) );
  NAND2_X1 U10067 ( .A1(n8609), .A2(n8709), .ZN(n8611) );
  NAND2_X1 U10068 ( .A1(n9184), .A2(n6895), .ZN(n8610) );
  NAND2_X1 U10069 ( .A1(n8611), .A2(n8610), .ZN(n8612) );
  XNOR2_X1 U10070 ( .A(n8612), .B(n8695), .ZN(n8918) );
  OAI22_X1 U10071 ( .A1(n8925), .A2(n8764), .B1(n8613), .B2(n8677), .ZN(n8621)
         );
  NAND2_X1 U10072 ( .A1(n8738), .A2(n6895), .ZN(n8615) );
  NAND2_X1 U10073 ( .A1(n9185), .A2(n8758), .ZN(n8614) );
  NAND2_X1 U10074 ( .A1(n8615), .A2(n8614), .ZN(n8731) );
  NAND2_X1 U10075 ( .A1(n8738), .A2(n8709), .ZN(n8617) );
  NAND2_X1 U10076 ( .A1(n9185), .A2(n6895), .ZN(n8616) );
  NAND2_X1 U10077 ( .A1(n8617), .A2(n8616), .ZN(n8618) );
  XNOR2_X1 U10078 ( .A(n8618), .B(n8695), .ZN(n8620) );
  AOI22_X1 U10079 ( .A1(n8918), .A2(n8621), .B1(n8731), .B2(n8620), .ZN(n8619)
         );
  NAND2_X1 U10080 ( .A1(n8730), .A2(n8619), .ZN(n8627) );
  INV_X1 U10081 ( .A(n8731), .ZN(n8623) );
  INV_X1 U10082 ( .A(n8621), .ZN(n8919) );
  AOI21_X1 U10083 ( .B1(n8917), .B2(n8623), .A(n8919), .ZN(n8622) );
  NAND3_X1 U10084 ( .A1(n8919), .A2(n8623), .A3(n8917), .ZN(n8624) );
  NAND2_X1 U10085 ( .A1(n8627), .A2(n8626), .ZN(n8808) );
  NOR2_X1 U10086 ( .A1(n8821), .A2(n8677), .ZN(n8628) );
  AOI21_X1 U10087 ( .B1(n9603), .B2(n6895), .A(n8628), .ZN(n8639) );
  AOI22_X1 U10088 ( .A1(n9603), .A2(n8709), .B1(n6895), .B2(n9183), .ZN(n8629)
         );
  XNOR2_X1 U10089 ( .A(n8629), .B(n8695), .ZN(n8640) );
  XOR2_X1 U10090 ( .A(n8639), .B(n8640), .Z(n8816) );
  NAND2_X1 U10091 ( .A1(n9545), .A2(n8709), .ZN(n8631) );
  NAND2_X1 U10092 ( .A1(n9182), .A2(n6895), .ZN(n8630) );
  NAND2_X1 U10093 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  XNOR2_X1 U10094 ( .A(n8632), .B(n8695), .ZN(n8635) );
  INV_X1 U10095 ( .A(n8635), .ZN(n8633) );
  AOI22_X1 U10096 ( .A1(n9545), .A2(n6895), .B1(n8758), .B2(n9182), .ZN(n8634)
         );
  NAND2_X1 U10097 ( .A1(n8633), .A2(n8634), .ZN(n8641) );
  INV_X1 U10098 ( .A(n8641), .ZN(n8636) );
  XNOR2_X1 U10099 ( .A(n8635), .B(n8634), .ZN(n8820) );
  OR2_X1 U10100 ( .A1(n8636), .A2(n8820), .ZN(n8638) );
  AND2_X1 U10101 ( .A1(n8816), .A2(n8638), .ZN(n8637) );
  NAND2_X1 U10102 ( .A1(n8808), .A2(n8637), .ZN(n8645) );
  INV_X1 U10103 ( .A(n8638), .ZN(n8643) );
  NAND2_X1 U10104 ( .A1(n8640), .A2(n8639), .ZN(n8817) );
  AND2_X1 U10105 ( .A1(n8817), .A2(n8641), .ZN(n8642) );
  OR2_X1 U10106 ( .A1(n8643), .A2(n8642), .ZN(n8644) );
  AOI22_X1 U10107 ( .A1(n9594), .A2(n8709), .B1(n6895), .B2(n8822), .ZN(n8646)
         );
  XNOR2_X1 U10108 ( .A(n8646), .B(n8695), .ZN(n8892) );
  AOI22_X1 U10109 ( .A1(n9594), .A2(n6895), .B1(n8758), .B2(n8822), .ZN(n8891)
         );
  OAI22_X1 U10110 ( .A1(n9535), .A2(n8764), .B1(n8894), .B2(n8677), .ZN(n8653)
         );
  NAND2_X1 U10111 ( .A1(n8648), .A2(n8709), .ZN(n8650) );
  NAND2_X1 U10112 ( .A1(n8854), .A2(n6895), .ZN(n8649) );
  NAND2_X1 U10113 ( .A1(n8650), .A2(n8649), .ZN(n8651) );
  XNOR2_X1 U10114 ( .A(n8651), .B(n8695), .ZN(n8652) );
  XOR2_X1 U10115 ( .A(n8653), .B(n8652), .Z(n8750) );
  INV_X1 U10116 ( .A(n8652), .ZN(n8655) );
  INV_X1 U10117 ( .A(n8653), .ZN(n8654) );
  NAND2_X1 U10118 ( .A1(n9530), .A2(n8709), .ZN(n8657) );
  NAND2_X1 U10119 ( .A1(n9181), .A2(n6895), .ZN(n8656) );
  NAND2_X1 U10120 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  XNOR2_X1 U10121 ( .A(n8658), .B(n8695), .ZN(n8659) );
  AOI22_X1 U10122 ( .A1(n9530), .A2(n6895), .B1(n8758), .B2(n9181), .ZN(n8660)
         );
  XNOR2_X1 U10123 ( .A(n8659), .B(n8660), .ZN(n8852) );
  INV_X1 U10124 ( .A(n8659), .ZN(n8661) );
  NAND2_X1 U10125 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  NAND2_X1 U10126 ( .A1(n9382), .A2(n8709), .ZN(n8665) );
  NAND2_X1 U10127 ( .A1(n9180), .A2(n6895), .ZN(n8664) );
  NAND2_X1 U10128 ( .A1(n8665), .A2(n8664), .ZN(n8666) );
  XNOR2_X1 U10129 ( .A(n8666), .B(n8695), .ZN(n8670) );
  NAND2_X1 U10130 ( .A1(n9382), .A2(n6895), .ZN(n8668) );
  NAND2_X1 U10131 ( .A1(n9180), .A2(n8758), .ZN(n8667) );
  NAND2_X1 U10132 ( .A1(n8668), .A2(n8667), .ZN(n8669) );
  NAND2_X1 U10133 ( .A1(n8670), .A2(n8669), .ZN(n8672) );
  OAI21_X1 U10134 ( .B1(n8670), .B2(n8669), .A(n8672), .ZN(n8785) );
  INV_X1 U10135 ( .A(n8785), .ZN(n8671) );
  AOI22_X1 U10136 ( .A1(n9516), .A2(n8709), .B1(n6895), .B2(n9179), .ZN(n8673)
         );
  XOR2_X1 U10137 ( .A(n8695), .B(n8673), .Z(n8674) );
  AOI22_X1 U10138 ( .A1(n9516), .A2(n6895), .B1(n8758), .B2(n9179), .ZN(n8872)
         );
  AOI22_X1 U10139 ( .A1(n9513), .A2(n8709), .B1(n6895), .B2(n9178), .ZN(n8676)
         );
  XOR2_X1 U10140 ( .A(n8695), .B(n8676), .Z(n8679) );
  OAI22_X1 U10141 ( .A1(n9354), .A2(n8764), .B1(n8678), .B2(n8677), .ZN(n8680)
         );
  NAND2_X1 U10142 ( .A1(n8679), .A2(n8680), .ZN(n8743) );
  INV_X1 U10143 ( .A(n8679), .ZN(n8682) );
  INV_X1 U10144 ( .A(n8680), .ZN(n8681) );
  NAND2_X1 U10145 ( .A1(n8682), .A2(n8681), .ZN(n8742) );
  NAND2_X1 U10146 ( .A1(n8683), .A2(n8742), .ZN(n8831) );
  NAND2_X1 U10147 ( .A1(n9504), .A2(n8709), .ZN(n8685) );
  NAND2_X1 U10148 ( .A1(n9177), .A2(n6895), .ZN(n8684) );
  NAND2_X1 U10149 ( .A1(n8685), .A2(n8684), .ZN(n8686) );
  XNOR2_X1 U10150 ( .A(n8686), .B(n8695), .ZN(n8690) );
  NAND2_X1 U10151 ( .A1(n9504), .A2(n6895), .ZN(n8688) );
  NAND2_X1 U10152 ( .A1(n9177), .A2(n8758), .ZN(n8687) );
  NAND2_X1 U10153 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  NOR2_X1 U10154 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  AOI21_X1 U10155 ( .B1(n8690), .B2(n8689), .A(n8691), .ZN(n8832) );
  NAND2_X1 U10156 ( .A1(n8831), .A2(n8832), .ZN(n8830) );
  INV_X1 U10157 ( .A(n8691), .ZN(n8692) );
  NAND2_X1 U10158 ( .A1(n9499), .A2(n8709), .ZN(n8694) );
  NAND2_X1 U10159 ( .A1(n9176), .A2(n6895), .ZN(n8693) );
  NAND2_X1 U10160 ( .A1(n8694), .A2(n8693), .ZN(n8696) );
  XNOR2_X1 U10161 ( .A(n8696), .B(n8695), .ZN(n8703) );
  AOI22_X1 U10162 ( .A1(n9499), .A2(n6895), .B1(n8758), .B2(n9176), .ZN(n8701)
         );
  XNOR2_X1 U10163 ( .A(n8703), .B(n8701), .ZN(n8800) );
  NAND2_X1 U10164 ( .A1(n8913), .A2(n8709), .ZN(n8698) );
  NAND2_X1 U10165 ( .A1(n9175), .A2(n6895), .ZN(n8697) );
  NAND2_X1 U10166 ( .A1(n8698), .A2(n8697), .ZN(n8699) );
  XNOR2_X1 U10167 ( .A(n8699), .B(n8761), .ZN(n8705) );
  AND2_X1 U10168 ( .A1(n9175), .A2(n8758), .ZN(n8700) );
  AOI21_X1 U10169 ( .B1(n8913), .B2(n6895), .A(n8700), .ZN(n8706) );
  XNOR2_X1 U10170 ( .A(n8705), .B(n8706), .ZN(n8901) );
  INV_X1 U10171 ( .A(n8701), .ZN(n8702) );
  NOR2_X1 U10172 ( .A1(n8703), .A2(n8702), .ZN(n8902) );
  NOR2_X1 U10173 ( .A1(n8901), .A2(n8902), .ZN(n8704) );
  INV_X1 U10174 ( .A(n8705), .ZN(n8708) );
  INV_X1 U10175 ( .A(n8706), .ZN(n8707) );
  NAND2_X1 U10176 ( .A1(n8708), .A2(n8707), .ZN(n8719) );
  NAND2_X1 U10177 ( .A1(n9296), .A2(n8709), .ZN(n8711) );
  OR2_X1 U10178 ( .A1(n8908), .A2(n8764), .ZN(n8710) );
  NAND2_X1 U10179 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  XNOR2_X1 U10180 ( .A(n8712), .B(n8761), .ZN(n8715) );
  INV_X1 U10181 ( .A(n8715), .ZN(n8717) );
  NOR2_X1 U10182 ( .A1(n8908), .A2(n8677), .ZN(n8713) );
  AOI21_X1 U10183 ( .B1(n9296), .B2(n6895), .A(n8713), .ZN(n8714) );
  INV_X1 U10184 ( .A(n8714), .ZN(n8716) );
  AOI21_X1 U10185 ( .B1(n8717), .B2(n8716), .A(n8774), .ZN(n8718) );
  INV_X1 U10186 ( .A(n8718), .ZN(n8721) );
  INV_X1 U10187 ( .A(n8719), .ZN(n8720) );
  NOR2_X1 U10188 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  INV_X1 U10189 ( .A(n9277), .ZN(n9173) );
  AND2_X1 U10190 ( .A1(n9175), .A2(n9167), .ZN(n8724) );
  AOI21_X1 U10191 ( .B1(n9173), .B2(n8874), .A(n8724), .ZN(n9293) );
  OAI22_X1 U10192 ( .A1(n9293), .A2(n9641), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8725), .ZN(n8726) );
  AOI21_X1 U10193 ( .B1(n9297), .B2(n8929), .A(n8726), .ZN(n8728) );
  NAND2_X1 U10194 ( .A1(n9296), .A2(n8912), .ZN(n8727) );
  NAND3_X1 U10195 ( .A1(n8729), .A2(n8728), .A3(n8727), .ZN(P1_U3214) );
  XNOR2_X1 U10196 ( .A(n8730), .B(n8917), .ZN(n8732) );
  NOR2_X1 U10197 ( .A1(n8732), .A2(n8731), .ZN(n8916) );
  AOI21_X1 U10198 ( .B1(n8732), .B2(n8731), .A(n8916), .ZN(n8740) );
  INV_X1 U10199 ( .A(n8733), .ZN(n8736) );
  AOI22_X1 U10200 ( .A1(n8734), .A2(n8895), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8735) );
  OAI21_X1 U10201 ( .B1(n8736), .B2(n9653), .A(n8735), .ZN(n8737) );
  AOI21_X1 U10202 ( .B1(n8738), .B2(n8912), .A(n8737), .ZN(n8739) );
  OAI21_X1 U10203 ( .B1(n8740), .B2(n9646), .A(n8739), .ZN(P1_U3215) );
  NAND2_X1 U10204 ( .A1(n8743), .A2(n8742), .ZN(n8744) );
  XNOR2_X1 U10205 ( .A(n8741), .B(n8744), .ZN(n8749) );
  AND2_X1 U10206 ( .A1(n9179), .A2(n9167), .ZN(n8745) );
  AOI21_X1 U10207 ( .B1(n9177), .B2(n8874), .A(n8745), .ZN(n9347) );
  AOI22_X1 U10208 ( .A1(n8929), .A2(n9351), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8746) );
  OAI21_X1 U10209 ( .B1(n9347), .B2(n9641), .A(n8746), .ZN(n8747) );
  AOI21_X1 U10210 ( .B1(n9513), .B2(n8912), .A(n8747), .ZN(n8748) );
  OAI21_X1 U10211 ( .B1(n8749), .B2(n9646), .A(n8748), .ZN(P1_U3216) );
  XOR2_X1 U10212 ( .A(n8751), .B(n8750), .Z(n8756) );
  AOI22_X1 U10213 ( .A1(n9181), .A2(n8874), .B1(n9167), .B2(n8822), .ZN(n9411)
         );
  OAI22_X1 U10214 ( .A1(n9411), .A2(n9641), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8752), .ZN(n8754) );
  NOR2_X1 U10215 ( .A1(n9535), .A2(n8924), .ZN(n8753) );
  AOI211_X1 U10216 ( .C1(n8929), .C2(n9414), .A(n8754), .B(n8753), .ZN(n8755)
         );
  OAI21_X1 U10217 ( .B1(n8756), .B2(n9646), .A(n8755), .ZN(P1_U3219) );
  NAND2_X1 U10218 ( .A1(n8773), .A2(n6895), .ZN(n8760) );
  NAND2_X1 U10219 ( .A1(n9173), .A2(n8758), .ZN(n8759) );
  NAND2_X1 U10220 ( .A1(n8760), .A2(n8759), .ZN(n8762) );
  XNOR2_X1 U10221 ( .A(n8762), .B(n8761), .ZN(n8766) );
  NAND2_X1 U10222 ( .A1(n8773), .A2(n8709), .ZN(n8763) );
  OAI21_X1 U10223 ( .B1(n9277), .B2(n8764), .A(n8763), .ZN(n8765) );
  XNOR2_X1 U10224 ( .A(n8766), .B(n8765), .ZN(n8775) );
  NAND3_X1 U10225 ( .A1(n8767), .A2(n8905), .A3(n8775), .ZN(n8778) );
  INV_X1 U10226 ( .A(n8768), .ZN(n8771) );
  AOI22_X1 U10227 ( .A1(n8895), .A2(n8769), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8770) );
  OAI21_X1 U10228 ( .B1(n8771), .B2(n9653), .A(n8770), .ZN(n8772) );
  AOI21_X1 U10229 ( .B1(n8773), .B2(n8912), .A(n8772), .ZN(n8777) );
  NAND3_X1 U10230 ( .A1(n8775), .A2(n8905), .A3(n8774), .ZN(n8776) );
  NAND2_X1 U10231 ( .A1(n9179), .A2(n8874), .ZN(n8780) );
  NAND2_X1 U10232 ( .A1(n9181), .A2(n9167), .ZN(n8779) );
  NAND2_X1 U10233 ( .A1(n8780), .A2(n8779), .ZN(n9376) );
  AOI22_X1 U10234 ( .A1(n9376), .A2(n8895), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8781) );
  OAI21_X1 U10235 ( .B1(n9383), .B2(n9653), .A(n8781), .ZN(n8787) );
  INV_X1 U10236 ( .A(n8782), .ZN(n8783) );
  AOI211_X1 U10237 ( .C1(n8785), .C2(n8784), .A(n9646), .B(n8783), .ZN(n8786)
         );
  AOI211_X1 U10238 ( .C1(n9382), .C2(n9650), .A(n8787), .B(n8786), .ZN(n8788)
         );
  INV_X1 U10239 ( .A(n8788), .ZN(P1_U3223) );
  OR2_X1 U10240 ( .A1(n8790), .A2(n8907), .ZN(n8792) );
  NAND2_X1 U10241 ( .A1(n9188), .A2(n9167), .ZN(n8791) );
  AND2_X1 U10242 ( .A1(n8792), .A2(n8791), .ZN(n9727) );
  NAND2_X1 U10243 ( .A1(n8929), .A2(n9731), .ZN(n8793) );
  OAI211_X1 U10244 ( .C1(n9727), .C2(n9641), .A(n8794), .B(n8793), .ZN(n8795)
         );
  AOI21_X1 U10245 ( .B1(n9785), .B2(n8912), .A(n8795), .ZN(n8796) );
  OAI21_X1 U10246 ( .B1(n8797), .B2(n9646), .A(n8796), .ZN(P1_U3224) );
  INV_X1 U10247 ( .A(n9499), .ZN(n9321) );
  OAI21_X1 U10248 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8801) );
  NAND2_X1 U10249 ( .A1(n8801), .A2(n8905), .ZN(n8807) );
  NAND2_X1 U10250 ( .A1(n9177), .A2(n9167), .ZN(n8803) );
  NAND2_X1 U10251 ( .A1(n9175), .A2(n8874), .ZN(n8802) );
  NAND2_X1 U10252 ( .A1(n8803), .A2(n8802), .ZN(n9326) );
  INV_X1 U10253 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8804) );
  OAI22_X1 U10254 ( .A1(n9318), .A2(n9653), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8804), .ZN(n8805) );
  AOI21_X1 U10255 ( .B1(n9326), .B2(n8895), .A(n8805), .ZN(n8806) );
  OAI211_X1 U10256 ( .C1(n9321), .C2(n8924), .A(n8807), .B(n8806), .ZN(
        P1_U3225) );
  XOR2_X1 U10257 ( .A(n8808), .B(n8816), .Z(n8815) );
  NAND2_X1 U10258 ( .A1(n9184), .A2(n9167), .ZN(n8810) );
  NAND2_X1 U10259 ( .A1(n9182), .A2(n8874), .ZN(n8809) );
  AND2_X1 U10260 ( .A1(n8810), .A2(n8809), .ZN(n9456) );
  NAND2_X1 U10261 ( .A1(n8929), .A2(n9461), .ZN(n8812) );
  OAI211_X1 U10262 ( .C1(n9456), .C2(n9641), .A(n8812), .B(n8811), .ZN(n8813)
         );
  AOI21_X1 U10263 ( .B1(n9603), .B2(n8912), .A(n8813), .ZN(n8814) );
  OAI21_X1 U10264 ( .B1(n8815), .B2(n9646), .A(n8814), .ZN(P1_U3226) );
  NAND2_X1 U10265 ( .A1(n8808), .A2(n8816), .ZN(n8818) );
  NAND2_X1 U10266 ( .A1(n8818), .A2(n8817), .ZN(n8819) );
  XOR2_X1 U10267 ( .A(n8820), .B(n8819), .Z(n8829) );
  OR2_X1 U10268 ( .A1(n8821), .A2(n9276), .ZN(n8824) );
  NAND2_X1 U10269 ( .A1(n8822), .A2(n8874), .ZN(n8823) );
  AND2_X1 U10270 ( .A1(n8824), .A2(n8823), .ZN(n9442) );
  NAND2_X1 U10271 ( .A1(n8929), .A2(n9445), .ZN(n8825) );
  OAI211_X1 U10272 ( .C1(n9442), .C2(n9641), .A(n8826), .B(n8825), .ZN(n8827)
         );
  AOI21_X1 U10273 ( .B1(n9545), .B2(n9650), .A(n8827), .ZN(n8828) );
  OAI21_X1 U10274 ( .B1(n8829), .B2(n9646), .A(n8828), .ZN(P1_U3228) );
  INV_X1 U10275 ( .A(n9504), .ZN(n9334) );
  OAI21_X1 U10276 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n8833) );
  NAND2_X1 U10277 ( .A1(n8833), .A2(n8905), .ZN(n8839) );
  NAND2_X1 U10278 ( .A1(n9176), .A2(n8874), .ZN(n8835) );
  NAND2_X1 U10279 ( .A1(n9178), .A2(n9167), .ZN(n8834) );
  NAND2_X1 U10280 ( .A1(n8835), .A2(n8834), .ZN(n9338) );
  OAI22_X1 U10281 ( .A1(n9340), .A2(n9653), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8836), .ZN(n8837) );
  AOI21_X1 U10282 ( .B1(n9338), .B2(n8895), .A(n8837), .ZN(n8838) );
  OAI211_X1 U10283 ( .C1(n9334), .C2(n8924), .A(n8839), .B(n8838), .ZN(
        P1_U3229) );
  OAI21_X1 U10284 ( .B1(n8843), .B2(n8842), .A(n8841), .ZN(n8844) );
  NAND3_X1 U10285 ( .A1(n8840), .A2(n8905), .A3(n8844), .ZN(n8851) );
  AOI22_X1 U10286 ( .A1(n8846), .A2(n8929), .B1(n8845), .B2(n8895), .ZN(n8849)
         );
  NAND2_X1 U10287 ( .A1(n8912), .A2(n8847), .ZN(n8848) );
  NAND4_X1 U10288 ( .A1(n8851), .A2(n8850), .A3(n8849), .A4(n8848), .ZN(
        P1_U3230) );
  XOR2_X1 U10289 ( .A(n8853), .B(n8852), .Z(n8860) );
  NOR2_X1 U10290 ( .A1(n9653), .A2(n9402), .ZN(n8858) );
  AND2_X1 U10291 ( .A1(n8854), .A2(n9167), .ZN(n8855) );
  AOI21_X1 U10292 ( .B1(n9180), .B2(n8874), .A(n8855), .ZN(n9399) );
  OAI22_X1 U10293 ( .A1(n9399), .A2(n9641), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8856), .ZN(n8857) );
  AOI211_X1 U10294 ( .C1(n9530), .C2(n8912), .A(n8858), .B(n8857), .ZN(n8859)
         );
  OAI21_X1 U10295 ( .B1(n8860), .B2(n9646), .A(n8859), .ZN(P1_U3233) );
  XOR2_X1 U10296 ( .A(n8862), .B(n8861), .Z(n8869) );
  AOI22_X1 U10297 ( .A1(n8863), .A2(n8895), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n8864) );
  OAI21_X1 U10298 ( .B1(n8865), .B2(n9653), .A(n8864), .ZN(n8866) );
  AOI21_X1 U10299 ( .B1(n8867), .B2(n8912), .A(n8866), .ZN(n8868) );
  OAI21_X1 U10300 ( .B1(n8869), .B2(n9646), .A(n8868), .ZN(P1_U3234) );
  NAND2_X1 U10301 ( .A1(n8871), .A2(n8870), .ZN(n8873) );
  XNOR2_X1 U10302 ( .A(n8873), .B(n8872), .ZN(n8879) );
  AOI22_X1 U10303 ( .A1(n9178), .A2(n8874), .B1(n9167), .B2(n9180), .ZN(n9362)
         );
  INV_X1 U10304 ( .A(n8875), .ZN(n9366) );
  AOI22_X1 U10305 ( .A1(n8929), .A2(n9366), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8876) );
  OAI21_X1 U10306 ( .B1(n9362), .B2(n9641), .A(n8876), .ZN(n8877) );
  AOI21_X1 U10307 ( .B1(n9516), .B2(n8912), .A(n8877), .ZN(n8878) );
  OAI21_X1 U10308 ( .B1(n8879), .B2(n9646), .A(n8878), .ZN(P1_U3235) );
  OAI21_X1 U10309 ( .B1(n8880), .B2(n8882), .A(n4435), .ZN(n8881) );
  OAI21_X1 U10310 ( .B1(n4429), .B2(n8882), .A(n8881), .ZN(n8883) );
  NAND2_X1 U10311 ( .A1(n8883), .A2(n8905), .ZN(n8889) );
  OAI22_X1 U10312 ( .A1(n8885), .A2(n9641), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8884), .ZN(n8886) );
  AOI21_X1 U10313 ( .B1(n8887), .B2(n8929), .A(n8886), .ZN(n8888) );
  OAI211_X1 U10314 ( .C1(n8890), .C2(n8924), .A(n8889), .B(n8888), .ZN(
        P1_U3236) );
  XNOR2_X1 U10315 ( .A(n8892), .B(n8891), .ZN(n8893) );
  XNOR2_X1 U10316 ( .A(n8647), .B(n8893), .ZN(n8900) );
  INV_X1 U10317 ( .A(n9431), .ZN(n8897) );
  OAI22_X1 U10318 ( .A1(n8972), .A2(n9276), .B1(n8894), .B2(n8907), .ZN(n9427)
         );
  AOI22_X1 U10319 ( .A1(n9427), .A2(n8895), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8896) );
  OAI21_X1 U10320 ( .B1(n8897), .B2(n9653), .A(n8896), .ZN(n8898) );
  AOI21_X1 U10321 ( .B1(n9594), .B2(n8912), .A(n8898), .ZN(n8899) );
  OAI21_X1 U10322 ( .B1(n8900), .B2(n9646), .A(n8899), .ZN(P1_U3238) );
  INV_X1 U10323 ( .A(n8798), .ZN(n8903) );
  OAI21_X1 U10324 ( .B1(n8903), .B2(n8902), .A(n8901), .ZN(n8906) );
  NAND3_X1 U10325 ( .A1(n8906), .A2(n8905), .A3(n8904), .ZN(n8915) );
  NOR2_X1 U10326 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  AOI21_X1 U10327 ( .B1(n9176), .B2(n9167), .A(n8909), .ZN(n9306) );
  AOI22_X1 U10328 ( .A1(n8929), .A2(n9310), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8910) );
  OAI21_X1 U10329 ( .B1(n9306), .B2(n9641), .A(n8910), .ZN(n8911) );
  AOI21_X1 U10330 ( .B1(n8913), .B2(n8912), .A(n8911), .ZN(n8914) );
  NAND2_X1 U10331 ( .A1(n8915), .A2(n8914), .ZN(P1_U3240) );
  AOI21_X1 U10332 ( .B1(n8917), .B2(n8730), .A(n8916), .ZN(n8921) );
  XNOR2_X1 U10333 ( .A(n8919), .B(n8918), .ZN(n8920) );
  XNOR2_X1 U10334 ( .A(n8921), .B(n8920), .ZN(n8931) );
  OAI22_X1 U10335 ( .A1(n8923), .A2(n9641), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8922), .ZN(n8927) );
  NOR2_X1 U10336 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  AOI211_X1 U10337 ( .C1(n8929), .C2(n8928), .A(n8927), .B(n8926), .ZN(n8930)
         );
  OAI21_X1 U10338 ( .B1(n8931), .B2(n9646), .A(n8930), .ZN(P1_U3241) );
  INV_X1 U10339 ( .A(n9161), .ZN(n9023) );
  NOR2_X1 U10340 ( .A1(n9382), .A2(n8932), .ZN(n8987) );
  INV_X1 U10341 ( .A(n8980), .ZN(n8933) );
  INV_X1 U10342 ( .A(n8941), .ZN(n8934) );
  NOR2_X1 U10343 ( .A1(n8935), .A2(n8934), .ZN(n8937) );
  OAI21_X1 U10344 ( .B1(n8935), .B2(n9161), .A(n8938), .ZN(n8936) );
  NAND2_X1 U10345 ( .A1(n8942), .A2(n8938), .ZN(n8939) );
  NAND2_X1 U10346 ( .A1(n8947), .A2(n8943), .ZN(n9122) );
  AOI21_X1 U10347 ( .B1(n8939), .B2(n9117), .A(n9122), .ZN(n8940) );
  NAND2_X1 U10348 ( .A1(n8949), .A2(n8944), .ZN(n9126) );
  OAI21_X1 U10349 ( .B1(n8940), .B2(n9126), .A(n9125), .ZN(n8952) );
  NAND2_X1 U10350 ( .A1(n8946), .A2(n8945), .ZN(n8948) );
  NAND3_X1 U10351 ( .A1(n8948), .A2(n8947), .A3(n9125), .ZN(n8950) );
  NAND2_X1 U10352 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  AOI21_X1 U10353 ( .B1(n8957), .B2(n9124), .A(n9048), .ZN(n8954) );
  NAND2_X1 U10354 ( .A1(n8963), .A2(n8958), .ZN(n9128) );
  OR2_X1 U10355 ( .A1(n9128), .A2(n8956), .ZN(n8953) );
  AND2_X1 U10356 ( .A1(n8953), .A2(n8960), .ZN(n9131) );
  OAI21_X1 U10357 ( .B1(n8954), .B2(n9128), .A(n9131), .ZN(n8955) );
  INV_X1 U10358 ( .A(n8966), .ZN(n9133) );
  AOI21_X1 U10359 ( .B1(n8955), .B2(n8965), .A(n9133), .ZN(n8968) );
  NAND2_X1 U10360 ( .A1(n8957), .A2(n8956), .ZN(n8959) );
  NAND3_X1 U10361 ( .A1(n8959), .A2(n8958), .A3(n9124), .ZN(n8962) );
  NAND2_X1 U10362 ( .A1(n8962), .A2(n8961), .ZN(n8964) );
  NAND2_X1 U10363 ( .A1(n8964), .A2(n8963), .ZN(n8967) );
  INV_X1 U10364 ( .A(n8965), .ZN(n9135) );
  INV_X1 U10365 ( .A(n9440), .ZN(n9438) );
  INV_X1 U10366 ( .A(n8975), .ZN(n8971) );
  NAND2_X1 U10367 ( .A1(n9545), .A2(n8972), .ZN(n8973) );
  NAND2_X1 U10368 ( .A1(n8974), .A2(n8973), .ZN(n9137) );
  NAND2_X1 U10369 ( .A1(n8979), .A2(n9408), .ZN(n9138) );
  OAI211_X1 U10370 ( .C1(n8976), .C2(n9138), .A(n9105), .B(n8988), .ZN(n8977)
         );
  AOI21_X1 U10371 ( .B1(n8980), .B2(n8979), .A(n9161), .ZN(n8981) );
  INV_X1 U10372 ( .A(n9360), .ZN(n8993) );
  NAND2_X1 U10373 ( .A1(n9077), .A2(n9078), .ZN(n8983) );
  NAND2_X1 U10374 ( .A1(n8984), .A2(n8982), .ZN(n9066) );
  MUX2_X1 U10375 ( .A(n8983), .B(n9066), .S(n9023), .Z(n8995) );
  NAND2_X1 U10376 ( .A1(n9566), .A2(n9175), .ZN(n9073) );
  NAND2_X1 U10377 ( .A1(n9073), .A2(n9071), .ZN(n9001) );
  AOI211_X1 U10378 ( .C1(n8986), .C2(n9076), .A(n9023), .B(n9001), .ZN(n9006)
         );
  INV_X1 U10379 ( .A(n8987), .ZN(n8990) );
  INV_X1 U10380 ( .A(n8988), .ZN(n8989) );
  NAND2_X1 U10381 ( .A1(n8990), .A2(n8989), .ZN(n8992) );
  NAND2_X1 U10382 ( .A1(n8992), .A2(n8991), .ZN(n9079) );
  OAI211_X1 U10383 ( .C1(n8996), .C2(n8995), .A(n9336), .B(n9077), .ZN(n8998)
         );
  NAND3_X1 U10384 ( .A1(n9146), .A2(n9023), .A3(n9083), .ZN(n8997) );
  AOI21_X1 U10385 ( .B1(n8998), .B2(n9068), .A(n8997), .ZN(n9005) );
  INV_X1 U10386 ( .A(n9001), .ZN(n9000) );
  INV_X1 U10387 ( .A(n9083), .ZN(n8999) );
  NAND3_X1 U10388 ( .A1(n9000), .A2(n8999), .A3(n9161), .ZN(n9003) );
  NAND3_X1 U10389 ( .A1(n9001), .A2(n9023), .A3(n9146), .ZN(n9002) );
  OAI211_X1 U10390 ( .C1(n9023), .C2(n9146), .A(n9003), .B(n9002), .ZN(n9004)
         );
  NAND2_X1 U10391 ( .A1(n9269), .A2(n9007), .ZN(n9086) );
  INV_X1 U10392 ( .A(n9008), .ZN(n9075) );
  INV_X1 U10393 ( .A(n9172), .ZN(n9010) );
  NAND2_X1 U10394 ( .A1(n9011), .A2(n9010), .ZN(n9090) );
  NAND2_X1 U10395 ( .A1(n9012), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U10396 ( .A1(n6608), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U10397 ( .A1(n9013), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9014) );
  NOR3_X1 U10398 ( .A1(n9260), .A2(n9060), .A3(n9275), .ZN(n9019) );
  AND2_X1 U10399 ( .A1(n9260), .A2(n9275), .ZN(n9030) );
  NOR2_X1 U10400 ( .A1(n9065), .A2(n9161), .ZN(n9018) );
  NOR2_X1 U10401 ( .A1(n9090), .A2(n9023), .ZN(n9017) );
  NOR4_X1 U10402 ( .A1(n9019), .A2(n9030), .A3(n9018), .A4(n9017), .ZN(n9021)
         );
  OAI21_X1 U10403 ( .B1(n9094), .B2(n9260), .A(n9481), .ZN(n9020) );
  INV_X1 U10404 ( .A(n9275), .ZN(n9171) );
  NAND2_X1 U10405 ( .A1(n9171), .A2(n9161), .ZN(n9025) );
  NAND3_X1 U10406 ( .A1(n9260), .A2(n9023), .A3(n9275), .ZN(n9024) );
  OAI211_X1 U10407 ( .C1(n9260), .C2(n9025), .A(n9024), .B(n9094), .ZN(n9026)
         );
  INV_X1 U10408 ( .A(n9481), .ZN(n9061) );
  NAND2_X1 U10409 ( .A1(n9026), .A2(n9061), .ZN(n9027) );
  NAND2_X1 U10410 ( .A1(n9260), .A2(n9060), .ZN(n9095) );
  NOR2_X1 U10411 ( .A1(n9260), .A2(n9275), .ZN(n9151) );
  INV_X1 U10412 ( .A(n9151), .ZN(n9031) );
  NOR2_X1 U10413 ( .A1(n6419), .A2(n9033), .ZN(n9038) );
  NOR2_X1 U10414 ( .A1(n9469), .A2(n9109), .ZN(n9036) );
  INV_X1 U10415 ( .A(n9034), .ZN(n9035) );
  NAND4_X1 U10416 ( .A1(n9038), .A2(n9037), .A3(n9036), .A4(n9035), .ZN(n9040)
         );
  NOR2_X1 U10417 ( .A1(n9040), .A2(n9039), .ZN(n9042) );
  NAND3_X1 U10418 ( .A1(n4724), .A2(n9042), .A3(n9041), .ZN(n9044) );
  NOR2_X1 U10419 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NAND3_X1 U10420 ( .A1(n9732), .A2(n9046), .A3(n9045), .ZN(n9049) );
  OR3_X1 U10421 ( .A1(n9049), .A2(n9048), .A3(n9047), .ZN(n9050) );
  NOR2_X1 U10422 ( .A1(n9051), .A2(n9050), .ZN(n9052) );
  NAND4_X1 U10423 ( .A1(n9424), .A2(n9454), .A3(n9052), .A4(n9440), .ZN(n9053)
         );
  NOR2_X1 U10424 ( .A1(n9409), .A2(n9053), .ZN(n9054) );
  AND2_X1 U10425 ( .A1(n9397), .A2(n9054), .ZN(n9055) );
  NAND4_X1 U10426 ( .A1(n9346), .A2(n9360), .A3(n9055), .A4(n9373), .ZN(n9056)
         );
  NOR2_X1 U10427 ( .A1(n9057), .A2(n9056), .ZN(n9058) );
  INV_X1 U10428 ( .A(n9159), .ZN(n9059) );
  INV_X1 U10429 ( .A(n9098), .ZN(n9062) );
  NAND2_X1 U10430 ( .A1(n9061), .A2(n9060), .ZN(n9162) );
  AOI21_X1 U10431 ( .B1(n9062), .B2(n9162), .A(n9101), .ZN(n9063) );
  AND2_X1 U10432 ( .A1(n9065), .A2(n9064), .ZN(n9148) );
  NAND2_X1 U10433 ( .A1(n9066), .A2(n9077), .ZN(n9067) );
  NAND2_X1 U10434 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  NAND2_X1 U10435 ( .A1(n9069), .A2(n9076), .ZN(n9070) );
  NAND2_X1 U10436 ( .A1(n9071), .A2(n9070), .ZN(n9084) );
  NOR2_X1 U10437 ( .A1(n9084), .A2(n4422), .ZN(n9141) );
  INV_X1 U10438 ( .A(n9146), .ZN(n9072) );
  AOI21_X1 U10439 ( .B1(n9141), .B2(n9396), .A(n9072), .ZN(n9089) );
  INV_X1 U10440 ( .A(n9073), .ZN(n9074) );
  NOR2_X1 U10441 ( .A1(n9075), .A2(n9074), .ZN(n9088) );
  INV_X1 U10442 ( .A(n9088), .ZN(n9144) );
  INV_X1 U10443 ( .A(n9076), .ZN(n9082) );
  INV_X1 U10444 ( .A(n9077), .ZN(n9081) );
  INV_X1 U10445 ( .A(n9078), .ZN(n9080) );
  NOR4_X1 U10446 ( .A1(n9082), .A2(n9081), .A3(n9080), .A4(n9079), .ZN(n9085)
         );
  OAI21_X1 U10447 ( .B1(n9085), .B2(n9084), .A(n9083), .ZN(n9087) );
  AOI21_X1 U10448 ( .B1(n9088), .B2(n9087), .A(n9086), .ZN(n9147) );
  OAI21_X1 U10449 ( .B1(n9089), .B2(n9144), .A(n9147), .ZN(n9092) );
  NAND2_X1 U10450 ( .A1(n9091), .A2(n9090), .ZN(n9104) );
  AOI21_X1 U10451 ( .B1(n9148), .B2(n9092), .A(n9104), .ZN(n9093) );
  AOI21_X1 U10452 ( .B1(n9151), .B2(n9094), .A(n9093), .ZN(n9097) );
  INV_X1 U10453 ( .A(n9095), .ZN(n9096) );
  NOR3_X1 U10454 ( .A1(n9097), .A2(n9096), .A3(n9159), .ZN(n9100) );
  OAI21_X1 U10455 ( .B1(n9100), .B2(n9099), .A(n9098), .ZN(n9102) );
  NAND2_X1 U10456 ( .A1(n9430), .A2(n9103), .ZN(n9157) );
  INV_X1 U10457 ( .A(n9104), .ZN(n9153) );
  INV_X1 U10458 ( .A(n9105), .ZN(n9143) );
  NAND3_X1 U10459 ( .A1(n9108), .A2(n9107), .A3(n9106), .ZN(n9113) );
  NAND3_X1 U10460 ( .A1(n9111), .A2(n9110), .A3(n9109), .ZN(n9112) );
  NOR2_X1 U10461 ( .A1(n9113), .A2(n9112), .ZN(n9116) );
  AOI21_X1 U10462 ( .B1(n9116), .B2(n9115), .A(n9114), .ZN(n9121) );
  INV_X1 U10463 ( .A(n9117), .ZN(n9120) );
  INV_X1 U10464 ( .A(n9118), .ZN(n9119) );
  NOR3_X1 U10465 ( .A1(n9121), .A2(n9120), .A3(n9119), .ZN(n9123) );
  NOR2_X1 U10466 ( .A1(n9123), .A2(n9122), .ZN(n9127) );
  OAI211_X1 U10467 ( .C1(n9127), .C2(n9126), .A(n9125), .B(n9124), .ZN(n9130)
         );
  AOI21_X1 U10468 ( .B1(n9130), .B2(n9129), .A(n9128), .ZN(n9134) );
  INV_X1 U10469 ( .A(n9131), .ZN(n9132) );
  NOR3_X1 U10470 ( .A1(n9134), .A2(n9133), .A3(n9132), .ZN(n9136) );
  OAI21_X1 U10471 ( .B1(n9136), .B2(n9135), .A(n9422), .ZN(n9140) );
  INV_X1 U10472 ( .A(n9137), .ZN(n9139) );
  AOI21_X1 U10473 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9142) );
  OAI21_X1 U10474 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9145) );
  AOI21_X1 U10475 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9150) );
  INV_X1 U10476 ( .A(n9147), .ZN(n9149) );
  OAI21_X1 U10477 ( .B1(n9150), .B2(n9149), .A(n9148), .ZN(n9152) );
  AOI21_X1 U10478 ( .B1(n9153), .B2(n9152), .A(n9151), .ZN(n9154) );
  OAI21_X1 U10479 ( .B1(n9154), .B2(n9159), .A(n9162), .ZN(n9155) );
  MUX2_X1 U10480 ( .A(n9157), .B(n9156), .S(n9155), .Z(n9164) );
  AOI211_X1 U10481 ( .C1(n9159), .C2(n9430), .A(n6411), .B(n9158), .ZN(n9163)
         );
  NAND4_X1 U10482 ( .A1(n9771), .A2(n9167), .A3(n9166), .A4(n9165), .ZN(n9168)
         );
  OAI211_X1 U10483 ( .C1(n6411), .C2(n9170), .A(n9168), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9169) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9171), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10485 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9172), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9173), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9174), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9175), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10489 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9176), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10490 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9177), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10491 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9178), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9179), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9180), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9181), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10495 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9182), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9183), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9184), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9185), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9186), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10500 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9187), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9188), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9189), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9190), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9191), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9192), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10506 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9193), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9194), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9195), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10510 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9197), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9198), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10512 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6863), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10513 ( .C1(n9201), .C2(n9200), .A(n9660), .B(n9199), .ZN(n9210)
         );
  OAI211_X1 U10514 ( .C1(n9204), .C2(n9203), .A(n9716), .B(n9202), .ZN(n9209)
         );
  AOI22_X1 U10515 ( .A1(n9205), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9208) );
  NAND2_X1 U10516 ( .A1(n9712), .A2(n9206), .ZN(n9207) );
  NAND4_X1 U10517 ( .A1(n9210), .A2(n9209), .A3(n9208), .A4(n9207), .ZN(
        P1_U3244) );
  INV_X1 U10518 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9212) );
  OAI22_X1 U10519 ( .A1(n9724), .A2(n9212), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9211), .ZN(n9213) );
  AOI21_X1 U10520 ( .B1(n9712), .B2(n9214), .A(n9213), .ZN(n9223) );
  OAI211_X1 U10521 ( .C1(n9217), .C2(n9216), .A(n9716), .B(n9215), .ZN(n9222)
         );
  OAI211_X1 U10522 ( .C1(n9220), .C2(n9219), .A(n9660), .B(n9218), .ZN(n9221)
         );
  NAND4_X1 U10523 ( .A1(n9224), .A2(n9223), .A3(n9222), .A4(n9221), .ZN(
        P1_U3245) );
  INV_X1 U10524 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U10525 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9225) );
  OAI21_X1 U10526 ( .B1(n9724), .B2(n9226), .A(n9225), .ZN(n9227) );
  AOI21_X1 U10527 ( .B1(n9712), .B2(n9228), .A(n9227), .ZN(n9237) );
  OAI211_X1 U10528 ( .C1(n9231), .C2(n9230), .A(n9716), .B(n9229), .ZN(n9236)
         );
  OAI211_X1 U10529 ( .C1(n9234), .C2(n9233), .A(n9660), .B(n9232), .ZN(n9235)
         );
  NAND3_X1 U10530 ( .A1(n9237), .A2(n9236), .A3(n9235), .ZN(P1_U3246) );
  OR2_X1 U10531 ( .A1(n9243), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U10532 ( .A1(n9713), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9241) );
  OR2_X1 U10533 ( .A1(n9713), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9240) );
  AND2_X1 U10534 ( .A1(n9241), .A2(n9240), .ZN(n9718) );
  NAND2_X1 U10535 ( .A1(n9719), .A2(n9718), .ZN(n9717) );
  NAND2_X1 U10536 ( .A1(n9717), .A2(n9241), .ZN(n9242) );
  XNOR2_X1 U10537 ( .A(n9242), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9251) );
  INV_X1 U10538 ( .A(n9251), .ZN(n9248) );
  OAI22_X1 U10539 ( .A1(n9245), .A2(n9244), .B1(n9243), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U10540 ( .A1(n9713), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9246) );
  OAI21_X1 U10541 ( .B1(n9713), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9246), .ZN(
        n9710) );
  NAND2_X1 U10542 ( .A1(n9714), .A2(n9246), .ZN(n9247) );
  INV_X1 U10543 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9537) );
  XNOR2_X1 U10544 ( .A(n9247), .B(n9537), .ZN(n9249) );
  AOI22_X1 U10545 ( .A1(n9716), .A2(n9248), .B1(n9249), .B2(n9660), .ZN(n9253)
         );
  OAI21_X1 U10546 ( .B1(n9249), .B2(n9709), .A(n9668), .ZN(n9250) );
  AOI21_X1 U10547 ( .B1(n9716), .B2(n9251), .A(n9250), .ZN(n9252) );
  NAND2_X1 U10548 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9254) );
  NAND2_X1 U10549 ( .A1(n9767), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U10550 ( .A1(n9470), .A2(n9482), .ZN(n9261) );
  OAI211_X1 U10551 ( .C1(n9481), .C2(n9760), .A(n9255), .B(n9261), .ZN(n9256)
         );
  AOI21_X1 U10552 ( .B1(n9257), .B2(n9754), .A(n9256), .ZN(n9258) );
  INV_X1 U10553 ( .A(n9258), .ZN(P1_U3263) );
  AOI211_X1 U10554 ( .C1(n9260), .C2(n9282), .A(n9736), .B(n9259), .ZN(n9483)
         );
  NAND2_X1 U10555 ( .A1(n9483), .A2(n9754), .ZN(n9264) );
  INV_X1 U10556 ( .A(n9261), .ZN(n9262) );
  AOI21_X1 U10557 ( .B1(n9767), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9262), .ZN(
        n9263) );
  OAI211_X1 U10558 ( .C1(n9559), .C2(n9760), .A(n9264), .B(n9263), .ZN(
        P1_U3264) );
  OAI21_X1 U10559 ( .B1(n6500), .B2(n9277), .A(n9265), .ZN(n9266) );
  XNOR2_X1 U10560 ( .A(n9266), .B(n9271), .ZN(n9562) );
  NAND2_X1 U10561 ( .A1(n9268), .A2(n9267), .ZN(n9270) );
  NAND2_X1 U10562 ( .A1(n9270), .A2(n9269), .ZN(n9272) );
  XNOR2_X1 U10563 ( .A(n9272), .B(n4675), .ZN(n9273) );
  NAND2_X1 U10564 ( .A1(n9273), .A2(n9729), .ZN(n9280) );
  OAI22_X1 U10565 ( .A1(n9277), .A2(n9276), .B1(n9275), .B2(n9274), .ZN(n9278)
         );
  INV_X1 U10566 ( .A(n9278), .ZN(n9279) );
  NAND2_X1 U10567 ( .A1(n9280), .A2(n9279), .ZN(n9488) );
  AOI21_X1 U10568 ( .B1(n9011), .B2(n9281), .A(n9736), .ZN(n9283) );
  NAND2_X1 U10569 ( .A1(n9283), .A2(n9282), .ZN(n9486) );
  NOR2_X1 U10570 ( .A1(n9486), .A2(n9740), .ZN(n9287) );
  AOI22_X1 U10571 ( .A1(n9767), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9284), .B2(
        n9756), .ZN(n9285) );
  OAI21_X1 U10572 ( .B1(n6605), .B2(n9760), .A(n9285), .ZN(n9286) );
  OAI21_X1 U10573 ( .B1(n9562), .B2(n9466), .A(n9288), .ZN(P1_U3356) );
  XNOR2_X1 U10574 ( .A(n9289), .B(n9290), .ZN(n9492) );
  INV_X1 U10575 ( .A(n9492), .ZN(n9302) );
  XNOR2_X1 U10576 ( .A(n9291), .B(n9290), .ZN(n9292) );
  NAND2_X1 U10577 ( .A1(n9292), .A2(n9729), .ZN(n9294) );
  NAND2_X1 U10578 ( .A1(n9294), .A2(n9293), .ZN(n9490) );
  AOI211_X1 U10579 ( .C1(n9296), .C2(n9309), .A(n9736), .B(n4573), .ZN(n9491)
         );
  NAND2_X1 U10580 ( .A1(n9491), .A2(n9754), .ZN(n9299) );
  AOI22_X1 U10581 ( .A1(n9767), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9297), .B2(
        n9756), .ZN(n9298) );
  OAI211_X1 U10582 ( .C1(n4489), .C2(n9760), .A(n9299), .B(n9298), .ZN(n9300)
         );
  AOI21_X1 U10583 ( .B1(n9490), .B2(n9470), .A(n9300), .ZN(n9301) );
  OAI21_X1 U10584 ( .B1(n9302), .B2(n9466), .A(n9301), .ZN(P1_U3266) );
  XOR2_X1 U10585 ( .A(n9304), .B(n9303), .Z(n9567) );
  XNOR2_X1 U10586 ( .A(n9305), .B(n9304), .ZN(n9308) );
  INV_X1 U10587 ( .A(n9306), .ZN(n9307) );
  AOI21_X1 U10588 ( .B1(n9308), .B2(n9729), .A(n9307), .ZN(n9496) );
  INV_X1 U10589 ( .A(n9496), .ZN(n9314) );
  OAI211_X1 U10590 ( .C1(n9566), .C2(n9317), .A(n9505), .B(n9309), .ZN(n9495)
         );
  NOR2_X1 U10591 ( .A1(n9495), .A2(n9740), .ZN(n9313) );
  AOI22_X1 U10592 ( .A1(n9767), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9310), .B2(
        n9756), .ZN(n9311) );
  OAI21_X1 U10593 ( .B1(n9566), .B2(n9760), .A(n9311), .ZN(n9312) );
  AOI211_X1 U10594 ( .C1(n9314), .C2(n9470), .A(n9313), .B(n9312), .ZN(n9315)
         );
  OAI21_X1 U10595 ( .B1(n9567), .B2(n9466), .A(n9315), .ZN(P1_U3267) );
  XOR2_X1 U10596 ( .A(n9316), .B(n9323), .Z(n9503) );
  AOI21_X1 U10597 ( .B1(n9499), .B2(n4949), .A(n9317), .ZN(n9500) );
  NOR2_X1 U10598 ( .A1(n9740), .A2(n9736), .ZN(n9474) );
  INV_X1 U10599 ( .A(n9318), .ZN(n9319) );
  AOI22_X1 U10600 ( .A1(n9319), .A2(n9756), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9767), .ZN(n9320) );
  OAI21_X1 U10601 ( .B1(n9321), .B2(n9760), .A(n9320), .ZN(n9330) );
  INV_X1 U10602 ( .A(n9322), .ZN(n9325) );
  INV_X1 U10603 ( .A(n9323), .ZN(n9324) );
  AOI21_X1 U10604 ( .B1(n9325), .B2(n9324), .A(n9425), .ZN(n9328) );
  AOI21_X1 U10605 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(n9502) );
  NOR2_X1 U10606 ( .A1(n9502), .A2(n9767), .ZN(n9329) );
  AOI211_X1 U10607 ( .C1(n9500), .C2(n9474), .A(n9330), .B(n9329), .ZN(n9331)
         );
  OAI21_X1 U10608 ( .B1(n9503), .B2(n9466), .A(n9331), .ZN(P1_U3268) );
  XNOR2_X1 U10609 ( .A(n9332), .B(n9336), .ZN(n9510) );
  AOI21_X1 U10610 ( .B1(n9504), .B2(n9349), .A(n4582), .ZN(n9506) );
  INV_X1 U10611 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9333) );
  OAI22_X1 U10612 ( .A1(n9334), .A2(n9760), .B1(n9333), .B2(n9470), .ZN(n9335)
         );
  AOI21_X1 U10613 ( .B1(n9506), .B2(n9474), .A(n9335), .ZN(n9343) );
  XNOR2_X1 U10614 ( .A(n9337), .B(n9336), .ZN(n9339) );
  AOI21_X1 U10615 ( .B1(n9339), .B2(n9729), .A(n9338), .ZN(n9508) );
  OAI21_X1 U10616 ( .B1(n9340), .B2(n9401), .A(n9508), .ZN(n9341) );
  NAND2_X1 U10617 ( .A1(n9341), .A2(n9470), .ZN(n9342) );
  OAI211_X1 U10618 ( .C1(n9510), .C2(n9466), .A(n9343), .B(n9342), .ZN(
        P1_U3269) );
  XOR2_X1 U10619 ( .A(n9346), .B(n9344), .Z(n9576) );
  XOR2_X1 U10620 ( .A(n9345), .B(n9346), .Z(n9348) );
  OAI21_X1 U10621 ( .B1(n9348), .B2(n9425), .A(n9347), .ZN(n9511) );
  INV_X1 U10622 ( .A(n9364), .ZN(n9350) );
  AOI211_X1 U10623 ( .C1(n9513), .C2(n9350), .A(n9736), .B(n4583), .ZN(n9512)
         );
  NAND2_X1 U10624 ( .A1(n9512), .A2(n9754), .ZN(n9353) );
  AOI22_X1 U10625 ( .A1(n9351), .A2(n9756), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9767), .ZN(n9352) );
  OAI211_X1 U10626 ( .C1(n9354), .C2(n9760), .A(n9353), .B(n9352), .ZN(n9355)
         );
  AOI21_X1 U10627 ( .B1(n9511), .B2(n9470), .A(n9355), .ZN(n9356) );
  OAI21_X1 U10628 ( .B1(n9576), .B2(n9466), .A(n9356), .ZN(P1_U3270) );
  XNOR2_X1 U10629 ( .A(n9357), .B(n9360), .ZN(n9580) );
  OAI21_X1 U10630 ( .B1(n9360), .B2(n9359), .A(n9358), .ZN(n9361) );
  NAND2_X1 U10631 ( .A1(n9361), .A2(n9729), .ZN(n9363) );
  NAND2_X1 U10632 ( .A1(n9363), .A2(n9362), .ZN(n9519) );
  OAI21_X1 U10633 ( .B1(n9380), .B2(n9369), .A(n9505), .ZN(n9365) );
  NOR2_X1 U10634 ( .A1(n9365), .A2(n9364), .ZN(n9518) );
  NAND2_X1 U10635 ( .A1(n9518), .A2(n9754), .ZN(n9368) );
  AOI22_X1 U10636 ( .A1(n9366), .A2(n9756), .B1(n9767), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9367) );
  OAI211_X1 U10637 ( .C1(n9369), .C2(n9760), .A(n9368), .B(n9367), .ZN(n9370)
         );
  AOI21_X1 U10638 ( .B1(n9519), .B2(n9470), .A(n9370), .ZN(n9371) );
  OAI21_X1 U10639 ( .B1(n9580), .B2(n9466), .A(n9371), .ZN(P1_U3271) );
  XOR2_X1 U10640 ( .A(n9372), .B(n9373), .Z(n9583) );
  XNOR2_X1 U10641 ( .A(n9374), .B(n9373), .ZN(n9375) );
  NAND2_X1 U10642 ( .A1(n9375), .A2(n9729), .ZN(n9378) );
  INV_X1 U10643 ( .A(n9376), .ZN(n9377) );
  NAND2_X1 U10644 ( .A1(n9378), .A2(n9377), .ZN(n9525) );
  NAND2_X1 U10645 ( .A1(n9390), .A2(n9382), .ZN(n9379) );
  NAND2_X1 U10646 ( .A1(n9379), .A2(n9505), .ZN(n9381) );
  OR2_X1 U10647 ( .A1(n9381), .A2(n9380), .ZN(n9522) );
  NOR2_X1 U10648 ( .A1(n9522), .A2(n9740), .ZN(n9387) );
  INV_X1 U10649 ( .A(n9382), .ZN(n9523) );
  INV_X1 U10650 ( .A(n9383), .ZN(n9384) );
  AOI22_X1 U10651 ( .A1(n9767), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9384), .B2(
        n9756), .ZN(n9385) );
  OAI21_X1 U10652 ( .B1(n9523), .B2(n9760), .A(n9385), .ZN(n9386) );
  AOI211_X1 U10653 ( .C1(n9525), .C2(n9470), .A(n9387), .B(n9386), .ZN(n9388)
         );
  OAI21_X1 U10654 ( .B1(n9583), .B2(n9466), .A(n9388), .ZN(P1_U3272) );
  XNOR2_X1 U10655 ( .A(n9389), .B(n9397), .ZN(n9587) );
  INV_X1 U10656 ( .A(n9390), .ZN(n9391) );
  AOI211_X1 U10657 ( .C1(n9530), .C2(n9407), .A(n9736), .B(n9391), .ZN(n9529)
         );
  INV_X1 U10658 ( .A(n9530), .ZN(n9393) );
  INV_X1 U10659 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9392) );
  OAI22_X1 U10660 ( .A1(n9393), .A2(n9760), .B1(n9470), .B2(n9392), .ZN(n9394)
         );
  AOI21_X1 U10661 ( .B1(n9529), .B2(n9754), .A(n9394), .ZN(n9405) );
  OAI21_X1 U10662 ( .B1(n9397), .B2(n9396), .A(n9395), .ZN(n9398) );
  NAND2_X1 U10663 ( .A1(n9398), .A2(n9729), .ZN(n9400) );
  NAND2_X1 U10664 ( .A1(n9400), .A2(n9399), .ZN(n9528) );
  NOR2_X1 U10665 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  OAI21_X1 U10666 ( .B1(n9528), .B2(n9403), .A(n9470), .ZN(n9404) );
  OAI211_X1 U10667 ( .C1(n9587), .C2(n9466), .A(n9405), .B(n9404), .ZN(
        P1_U3273) );
  XNOR2_X1 U10668 ( .A(n9406), .B(n9409), .ZN(n9591) );
  OAI211_X1 U10669 ( .C1(n9420), .C2(n9535), .A(n9505), .B(n9407), .ZN(n9533)
         );
  NAND2_X1 U10670 ( .A1(n9429), .A2(n9408), .ZN(n9410) );
  XNOR2_X1 U10671 ( .A(n9410), .B(n9409), .ZN(n9413) );
  INV_X1 U10672 ( .A(n9411), .ZN(n9412) );
  AOI21_X1 U10673 ( .B1(n9413), .B2(n9729), .A(n9412), .ZN(n9534) );
  OAI21_X1 U10674 ( .B1(n9430), .B2(n9533), .A(n9534), .ZN(n9417) );
  AOI22_X1 U10675 ( .A1(n9767), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9414), .B2(
        n9756), .ZN(n9415) );
  OAI21_X1 U10676 ( .B1(n9535), .B2(n9760), .A(n9415), .ZN(n9416) );
  AOI21_X1 U10677 ( .B1(n9417), .B2(n9470), .A(n9416), .ZN(n9418) );
  OAI21_X1 U10678 ( .B1(n9591), .B2(n9466), .A(n9418), .ZN(P1_U3274) );
  XNOR2_X1 U10679 ( .A(n9419), .B(n9424), .ZN(n9596) );
  INV_X1 U10680 ( .A(n9420), .ZN(n9421) );
  OAI211_X1 U10681 ( .C1(n9433), .C2(n9444), .A(n9421), .B(n9505), .ZN(n9539)
         );
  INV_X1 U10682 ( .A(n9422), .ZN(n9423) );
  NOR2_X1 U10683 ( .A1(n9424), .A2(n9423), .ZN(n9426) );
  AOI21_X1 U10684 ( .B1(n9439), .B2(n9426), .A(n9425), .ZN(n9428) );
  AOI21_X1 U10685 ( .B1(n9429), .B2(n9428), .A(n9427), .ZN(n9540) );
  OAI21_X1 U10686 ( .B1(n9430), .B2(n9539), .A(n9540), .ZN(n9435) );
  AOI22_X1 U10687 ( .A1(n9767), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9431), .B2(
        n9756), .ZN(n9432) );
  OAI21_X1 U10688 ( .B1(n9433), .B2(n9760), .A(n9432), .ZN(n9434) );
  AOI21_X1 U10689 ( .B1(n9435), .B2(n9470), .A(n9434), .ZN(n9436) );
  OAI21_X1 U10690 ( .B1(n9596), .B2(n9466), .A(n9436), .ZN(P1_U3275) );
  XNOR2_X1 U10691 ( .A(n9437), .B(n9438), .ZN(n9600) );
  OAI211_X1 U10692 ( .C1(n9441), .C2(n9440), .A(n9439), .B(n9729), .ZN(n9443)
         );
  NAND2_X1 U10693 ( .A1(n9443), .A2(n9442), .ZN(n9543) );
  INV_X1 U10694 ( .A(n9545), .ZN(n9448) );
  AOI211_X1 U10695 ( .C1(n9545), .C2(n9459), .A(n9736), .B(n9444), .ZN(n9544)
         );
  NAND2_X1 U10696 ( .A1(n9544), .A2(n9754), .ZN(n9447) );
  AOI22_X1 U10697 ( .A1(n9767), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9445), .B2(
        n9756), .ZN(n9446) );
  OAI211_X1 U10698 ( .C1(n9448), .C2(n9760), .A(n9447), .B(n9446), .ZN(n9449)
         );
  AOI21_X1 U10699 ( .B1(n9543), .B2(n9470), .A(n9449), .ZN(n9450) );
  OAI21_X1 U10700 ( .B1(n9600), .B2(n9466), .A(n9450), .ZN(P1_U3276) );
  XNOR2_X1 U10701 ( .A(n9451), .B(n9452), .ZN(n9607) );
  OAI211_X1 U10702 ( .C1(n9455), .C2(n9454), .A(n9453), .B(n9729), .ZN(n9457)
         );
  NAND2_X1 U10703 ( .A1(n9457), .A2(n9456), .ZN(n9549) );
  INV_X1 U10704 ( .A(n9458), .ZN(n9460) );
  OAI211_X1 U10705 ( .C1(n4576), .C2(n9460), .A(n9459), .B(n9505), .ZN(n9550)
         );
  AOI22_X1 U10706 ( .A1(n9767), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9461), .B2(
        n9756), .ZN(n9463) );
  NAND2_X1 U10707 ( .A1(n9603), .A2(n9745), .ZN(n9462) );
  OAI211_X1 U10708 ( .C1(n9550), .C2(n9740), .A(n9463), .B(n9462), .ZN(n9464)
         );
  AOI21_X1 U10709 ( .B1(n9549), .B2(n9470), .A(n9464), .ZN(n9465) );
  OAI21_X1 U10710 ( .B1(n9607), .B2(n9466), .A(n9465), .ZN(P1_U3277) );
  AND3_X1 U10711 ( .A1(n9469), .A2(n9468), .A3(n9467), .ZN(n9472) );
  OAI21_X1 U10712 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n9477) );
  AOI22_X1 U10713 ( .A1(n9767), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9756), .ZN(n9476) );
  OAI21_X1 U10714 ( .B1(n9745), .B2(n9474), .A(n9473), .ZN(n9475) );
  NAND3_X1 U10715 ( .A1(n9477), .A2(n9476), .A3(n9475), .ZN(P1_U3293) );
  INV_X1 U10716 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9479) );
  MUX2_X1 U10717 ( .A(n9479), .B(n9478), .S(n9799), .Z(n9480) );
  OAI21_X1 U10718 ( .B1(n9481), .B2(n6505), .A(n9480), .ZN(P1_U3553) );
  INV_X1 U10719 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9484) );
  NOR2_X1 U10720 ( .A1(n9483), .A2(n9482), .ZN(n9556) );
  MUX2_X1 U10721 ( .A(n9484), .B(n9556), .S(n9799), .Z(n9485) );
  OAI21_X1 U10722 ( .B1(n9559), .B2(n6505), .A(n9485), .ZN(P1_U3552) );
  INV_X1 U10723 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9489) );
  OAI21_X1 U10724 ( .B1(n6605), .B2(n9787), .A(n9486), .ZN(n9487) );
  NOR2_X1 U10725 ( .A1(n9488), .A2(n9487), .ZN(n9560) );
  INV_X1 U10726 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U10727 ( .A(n9493), .B(n9563), .S(n9799), .Z(n9494) );
  OAI21_X1 U10728 ( .B1(n4489), .B2(n6505), .A(n9494), .ZN(P1_U3549) );
  OAI22_X1 U10729 ( .A1(n9567), .A2(n9555), .B1(n9566), .B2(n6505), .ZN(n9498)
         );
  NAND2_X1 U10730 ( .A1(n9496), .A2(n9495), .ZN(n9568) );
  MUX2_X1 U10731 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9568), .S(n9799), .Z(n9497) );
  OR2_X1 U10732 ( .A1(n9498), .A2(n9497), .ZN(P1_U3548) );
  AOI22_X1 U10733 ( .A1(n9500), .A2(n9505), .B1(n9546), .B2(n9499), .ZN(n9501)
         );
  OAI211_X1 U10734 ( .C1(n9503), .C2(n9509), .A(n9502), .B(n9501), .ZN(n9571)
         );
  MUX2_X1 U10735 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9571), .S(n9799), .Z(
        P1_U3547) );
  AOI22_X1 U10736 ( .A1(n9506), .A2(n9505), .B1(n9546), .B2(n9504), .ZN(n9507)
         );
  OAI211_X1 U10737 ( .C1(n9510), .C2(n9509), .A(n9508), .B(n9507), .ZN(n9572)
         );
  MUX2_X1 U10738 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9572), .S(n9799), .Z(
        P1_U3546) );
  AOI211_X1 U10739 ( .C1(n9546), .C2(n9513), .A(n9512), .B(n9511), .ZN(n9573)
         );
  MUX2_X1 U10740 ( .A(n9514), .B(n9573), .S(n9799), .Z(n9515) );
  OAI21_X1 U10741 ( .B1(n9576), .B2(n9555), .A(n9515), .ZN(P1_U3545) );
  AND2_X1 U10742 ( .A1(n9516), .A2(n9546), .ZN(n9517) );
  MUX2_X1 U10743 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9577), .S(n9799), .Z(n9520) );
  INV_X1 U10744 ( .A(n9520), .ZN(n9521) );
  OAI21_X1 U10745 ( .B1(n9580), .B2(n9555), .A(n9521), .ZN(P1_U3544) );
  INV_X1 U10746 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9526) );
  OAI21_X1 U10747 ( .B1(n9523), .B2(n9787), .A(n9522), .ZN(n9524) );
  NOR2_X1 U10748 ( .A1(n9525), .A2(n9524), .ZN(n9581) );
  MUX2_X1 U10749 ( .A(n9526), .B(n9581), .S(n9799), .Z(n9527) );
  OAI21_X1 U10750 ( .B1(n9583), .B2(n9555), .A(n9527), .ZN(P1_U3543) );
  INV_X1 U10751 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9531) );
  AOI211_X1 U10752 ( .C1(n9546), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9584)
         );
  MUX2_X1 U10753 ( .A(n9531), .B(n9584), .S(n9799), .Z(n9532) );
  OAI21_X1 U10754 ( .B1(n9587), .B2(n9555), .A(n9532), .ZN(P1_U3542) );
  OAI211_X1 U10755 ( .C1(n9535), .C2(n9787), .A(n9534), .B(n9533), .ZN(n9536)
         );
  INV_X1 U10756 ( .A(n9536), .ZN(n9588) );
  MUX2_X1 U10757 ( .A(n9537), .B(n9588), .S(n9799), .Z(n9538) );
  OAI21_X1 U10758 ( .B1(n9591), .B2(n9555), .A(n9538), .ZN(P1_U3541) );
  NAND2_X1 U10759 ( .A1(n9540), .A2(n9539), .ZN(n9592) );
  MUX2_X1 U10760 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9592), .S(n9799), .Z(n9541) );
  AOI21_X1 U10761 ( .B1(n9553), .B2(n9594), .A(n9541), .ZN(n9542) );
  OAI21_X1 U10762 ( .B1(n9596), .B2(n9555), .A(n9542), .ZN(P1_U3540) );
  INV_X1 U10763 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9547) );
  AOI211_X1 U10764 ( .C1(n9546), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9597)
         );
  MUX2_X1 U10765 ( .A(n9547), .B(n9597), .S(n9799), .Z(n9548) );
  OAI21_X1 U10766 ( .B1(n9600), .B2(n9555), .A(n9548), .ZN(P1_U3539) );
  INV_X1 U10767 ( .A(n9549), .ZN(n9551) );
  NAND2_X1 U10768 ( .A1(n9551), .A2(n9550), .ZN(n9601) );
  MUX2_X1 U10769 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9601), .S(n9799), .Z(n9552) );
  AOI21_X1 U10770 ( .B1(n9553), .B2(n9603), .A(n9552), .ZN(n9554) );
  OAI21_X1 U10771 ( .B1(n9607), .B2(n9555), .A(n9554), .ZN(P1_U3538) );
  INV_X1 U10772 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9557) );
  MUX2_X1 U10773 ( .A(n9557), .B(n9556), .S(n9793), .Z(n9558) );
  OAI21_X1 U10774 ( .B1(n9559), .B2(n6501), .A(n9558), .ZN(P1_U3520) );
  INV_X1 U10775 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9561) );
  INV_X1 U10776 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9564) );
  MUX2_X1 U10777 ( .A(n9564), .B(n9563), .S(n9793), .Z(n9565) );
  OAI21_X1 U10778 ( .B1(n4489), .B2(n6501), .A(n9565), .ZN(P1_U3517) );
  OAI22_X1 U10779 ( .A1(n9567), .A2(n9606), .B1(n9566), .B2(n6501), .ZN(n9570)
         );
  MUX2_X1 U10780 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9568), .S(n9793), .Z(n9569) );
  OR2_X1 U10781 ( .A1(n9570), .A2(n9569), .ZN(P1_U3516) );
  MUX2_X1 U10782 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9571), .S(n9793), .Z(
        P1_U3515) );
  MUX2_X1 U10783 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9572), .S(n9793), .Z(
        P1_U3514) );
  INV_X1 U10784 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9574) );
  MUX2_X1 U10785 ( .A(n9574), .B(n9573), .S(n9793), .Z(n9575) );
  OAI21_X1 U10786 ( .B1(n9576), .B2(n9606), .A(n9575), .ZN(P1_U3513) );
  MUX2_X1 U10787 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9577), .S(n9793), .Z(n9578) );
  INV_X1 U10788 ( .A(n9578), .ZN(n9579) );
  OAI21_X1 U10789 ( .B1(n9580), .B2(n9606), .A(n9579), .ZN(P1_U3512) );
  INV_X1 U10790 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10143) );
  MUX2_X1 U10791 ( .A(n10143), .B(n9581), .S(n9793), .Z(n9582) );
  OAI21_X1 U10792 ( .B1(n9583), .B2(n9606), .A(n9582), .ZN(P1_U3511) );
  INV_X1 U10793 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9585) );
  MUX2_X1 U10794 ( .A(n9585), .B(n9584), .S(n9793), .Z(n9586) );
  OAI21_X1 U10795 ( .B1(n9587), .B2(n9606), .A(n9586), .ZN(P1_U3510) );
  INV_X1 U10796 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9589) );
  MUX2_X1 U10797 ( .A(n9589), .B(n9588), .S(n9793), .Z(n9590) );
  OAI21_X1 U10798 ( .B1(n9591), .B2(n9606), .A(n9590), .ZN(P1_U3509) );
  MUX2_X1 U10799 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9592), .S(n9793), .Z(n9593) );
  AOI21_X1 U10800 ( .B1(n9604), .B2(n9594), .A(n9593), .ZN(n9595) );
  OAI21_X1 U10801 ( .B1(n9596), .B2(n9606), .A(n9595), .ZN(P1_U3507) );
  INV_X1 U10802 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9598) );
  MUX2_X1 U10803 ( .A(n9598), .B(n9597), .S(n9793), .Z(n9599) );
  OAI21_X1 U10804 ( .B1(n9600), .B2(n9606), .A(n9599), .ZN(P1_U3504) );
  MUX2_X1 U10805 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9601), .S(n9793), .Z(n9602) );
  AOI21_X1 U10806 ( .B1(n9604), .B2(n9603), .A(n9602), .ZN(n9605) );
  OAI21_X1 U10807 ( .B1(n9607), .B2(n9606), .A(n9605), .ZN(P1_U3501) );
  MUX2_X1 U10808 ( .A(P1_D_REG_0__SCAN_IN), .B(n9608), .S(n9771), .Z(P1_U3439)
         );
  INV_X1 U10809 ( .A(n9609), .ZN(n9615) );
  NOR4_X1 U10810 ( .A1(n9611), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9610), .ZN(n9612) );
  AOI21_X1 U10811 ( .B1(n9613), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9612), .ZN(
        n9614) );
  OAI21_X1 U10812 ( .B1(n9615), .B2(n9626), .A(n9614), .ZN(P1_U3324) );
  OAI222_X1 U10813 ( .A1(P1_U3086), .A2(n6045), .B1(n9626), .B2(n9617), .C1(
        n9616), .C2(n9623), .ZN(P1_U3326) );
  OAI222_X1 U10814 ( .A1(P1_U3086), .A2(n6459), .B1(n9620), .B2(n9619), .C1(
        n9618), .C2(n9623), .ZN(P1_U3327) );
  OAI222_X1 U10815 ( .A1(P1_U3086), .A2(n6612), .B1(n9626), .B2(n9622), .C1(
        n9621), .C2(n9623), .ZN(P1_U3328) );
  OAI222_X1 U10816 ( .A1(P1_U3086), .A2(n9627), .B1(n9626), .B2(n9625), .C1(
        n9624), .C2(n9623), .ZN(P1_U3329) );
  MUX2_X1 U10817 ( .A(n9628), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10818 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9639) );
  AOI211_X1 U10819 ( .C1(n9631), .C2(n9630), .A(n9629), .B(n9700), .ZN(n9636)
         );
  AOI211_X1 U10820 ( .C1(n9634), .C2(n9633), .A(n9632), .B(n9709), .ZN(n9635)
         );
  AOI211_X1 U10821 ( .C1(n9712), .C2(n9637), .A(n9636), .B(n9635), .ZN(n9638)
         );
  NAND2_X1 U10822 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9640) );
  OAI211_X1 U10823 ( .C1(n9724), .C2(n9639), .A(n9638), .B(n9640), .ZN(
        P1_U3253) );
  OAI21_X1 U10824 ( .B1(n9642), .B2(n9641), .A(n9640), .ZN(n9649) );
  AOI21_X1 U10825 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9647) );
  NOR2_X1 U10826 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  AOI211_X1 U10827 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(n9652)
         );
  OAI21_X1 U10828 ( .B1(n9654), .B2(n9653), .A(n9652), .ZN(P1_U3217) );
  XNOR2_X1 U10829 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10830 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10831 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9672) );
  INV_X1 U10832 ( .A(n9655), .ZN(n9667) );
  AOI21_X1 U10833 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9659) );
  NAND2_X1 U10834 ( .A1(n9660), .A2(n9659), .ZN(n9666) );
  AOI21_X1 U10835 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9664) );
  NAND2_X1 U10836 ( .A1(n9716), .A2(n9664), .ZN(n9665) );
  OAI211_X1 U10837 ( .C1(n9668), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9669)
         );
  INV_X1 U10838 ( .A(n9669), .ZN(n9671) );
  NAND2_X1 U10839 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9670) );
  OAI211_X1 U10840 ( .C1(n9724), .C2(n9672), .A(n9671), .B(n9670), .ZN(
        P1_U3254) );
  INV_X1 U10841 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9684) );
  AOI211_X1 U10842 ( .C1(n9675), .C2(n9674), .A(n9709), .B(n9673), .ZN(n9680)
         );
  AOI211_X1 U10843 ( .C1(n9678), .C2(n9677), .A(n9700), .B(n9676), .ZN(n9679)
         );
  AOI211_X1 U10844 ( .C1(n9712), .C2(n9681), .A(n9680), .B(n9679), .ZN(n9683)
         );
  NAND2_X1 U10845 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9682) );
  OAI211_X1 U10846 ( .C1(n9724), .C2(n9684), .A(n9683), .B(n9682), .ZN(
        P1_U3256) );
  INV_X1 U10847 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9696) );
  AOI211_X1 U10848 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n9700), .ZN(n9692)
         );
  AOI211_X1 U10849 ( .C1(n9690), .C2(n9689), .A(n9709), .B(n9688), .ZN(n9691)
         );
  AOI211_X1 U10850 ( .C1(n9712), .C2(n9693), .A(n9692), .B(n9691), .ZN(n9695)
         );
  NAND2_X1 U10851 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9694) );
  OAI211_X1 U10852 ( .C1(n9724), .C2(n9696), .A(n9695), .B(n9694), .ZN(
        P1_U3257) );
  AOI211_X1 U10853 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9709), .ZN(n9705)
         );
  AOI211_X1 U10854 ( .C1(n9703), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9704)
         );
  AOI211_X1 U10855 ( .C1(n9712), .C2(n9706), .A(n9705), .B(n9704), .ZN(n9708)
         );
  NAND2_X1 U10856 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9707) );
  OAI211_X1 U10857 ( .C1(n9724), .C2(n10001), .A(n9708), .B(n9707), .ZN(
        P1_U3258) );
  AOI21_X1 U10858 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9715) );
  AOI22_X1 U10859 ( .A1(n9715), .A2(n9714), .B1(n9713), .B2(n9712), .ZN(n9721)
         );
  OAI211_X1 U10860 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9720)
         );
  AND2_X1 U10861 ( .A1(n9721), .A2(n9720), .ZN(n9723) );
  NAND2_X1 U10862 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9722) );
  OAI211_X1 U10863 ( .C1(n9724), .C2(n9944), .A(n9723), .B(n9722), .ZN(
        P1_U3261) );
  XNOR2_X1 U10864 ( .A(n9726), .B(n9725), .ZN(n9730) );
  INV_X1 U10865 ( .A(n9727), .ZN(n9728) );
  AOI21_X1 U10866 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n9784) );
  AOI222_X1 U10867 ( .A1(n9785), .A2(n9745), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9767), .C1(n9756), .C2(n9731), .ZN(n9743) );
  NAND2_X1 U10868 ( .A1(n9733), .A2(n9732), .ZN(n9734) );
  AND2_X1 U10869 ( .A1(n9735), .A2(n9734), .ZN(n9792) );
  AOI21_X1 U10870 ( .B1(n9737), .B2(n9785), .A(n9736), .ZN(n9739) );
  NAND2_X1 U10871 ( .A1(n9739), .A2(n9738), .ZN(n9786) );
  NOR2_X1 U10872 ( .A1(n9786), .A2(n9740), .ZN(n9741) );
  AOI21_X1 U10873 ( .B1(n9792), .B2(n9764), .A(n9741), .ZN(n9742) );
  OAI211_X1 U10874 ( .C1(n9767), .C2(n9784), .A(n9743), .B(n9742), .ZN(
        P1_U3281) );
  AOI222_X1 U10875 ( .A1(n9746), .A2(n9745), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9767), .C1(n9756), .C2(n9744), .ZN(n9752) );
  INV_X1 U10876 ( .A(n9747), .ZN(n9748) );
  AOI22_X1 U10877 ( .A1(n9750), .A2(n9749), .B1(n9754), .B2(n9748), .ZN(n9751)
         );
  OAI211_X1 U10878 ( .C1(n9767), .C2(n9753), .A(n9752), .B(n9751), .ZN(
        P1_U3285) );
  NAND2_X1 U10879 ( .A1(n9755), .A2(n9754), .ZN(n9759) );
  AOI22_X1 U10880 ( .A1(n9767), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9757), .B2(
        n9756), .ZN(n9758) );
  OAI211_X1 U10881 ( .C1(n9761), .C2(n9760), .A(n9759), .B(n9758), .ZN(n9762)
         );
  AOI21_X1 U10882 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9765) );
  OAI21_X1 U10883 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(P1_U3288) );
  AND2_X1 U10884 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9972), .ZN(P1_U3294) );
  AND2_X1 U10885 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9972), .ZN(P1_U3295) );
  AND2_X1 U10886 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9972), .ZN(P1_U3296) );
  AND2_X1 U10887 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9972), .ZN(P1_U3297) );
  AND2_X1 U10888 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9972), .ZN(P1_U3298) );
  AND2_X1 U10889 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9972), .ZN(P1_U3299) );
  AND2_X1 U10890 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9972), .ZN(P1_U3300) );
  AND2_X1 U10891 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9972), .ZN(P1_U3301) );
  AND2_X1 U10892 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9972), .ZN(P1_U3303) );
  AND2_X1 U10893 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9972), .ZN(P1_U3304) );
  AND2_X1 U10894 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9972), .ZN(P1_U3305) );
  AND2_X1 U10895 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9972), .ZN(P1_U3306) );
  AND2_X1 U10896 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9972), .ZN(P1_U3307) );
  AND2_X1 U10897 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9972), .ZN(P1_U3308) );
  AND2_X1 U10898 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9972), .ZN(P1_U3309) );
  AND2_X1 U10899 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9972), .ZN(P1_U3310) );
  AND2_X1 U10900 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9972), .ZN(P1_U3311) );
  AND2_X1 U10901 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9972), .ZN(P1_U3312) );
  AND2_X1 U10902 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9972), .ZN(P1_U3313) );
  AND2_X1 U10903 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9972), .ZN(P1_U3314) );
  AND2_X1 U10904 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9972), .ZN(P1_U3315) );
  AND2_X1 U10905 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9972), .ZN(P1_U3316) );
  AND2_X1 U10906 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9972), .ZN(P1_U3317) );
  AND2_X1 U10907 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9972), .ZN(P1_U3318) );
  AND2_X1 U10908 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9972), .ZN(P1_U3319) );
  AND2_X1 U10909 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9972), .ZN(P1_U3320) );
  AND2_X1 U10910 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9972), .ZN(P1_U3321) );
  AND2_X1 U10911 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9972), .ZN(P1_U3322) );
  AND2_X1 U10912 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9972), .ZN(P1_U3323) );
  INV_X1 U10913 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9770) );
  OAI21_X1 U10914 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(P1_U3440) );
  OAI21_X1 U10915 ( .B1(n9773), .B2(n9787), .A(n9772), .ZN(n9775) );
  AOI211_X1 U10916 ( .C1(n9791), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9795)
         );
  INV_X1 U10917 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9777) );
  AOI22_X1 U10918 ( .A1(n9793), .A2(n9795), .B1(n9777), .B2(n6614), .ZN(
        P1_U3480) );
  OAI211_X1 U10919 ( .C1(n9780), .C2(n9787), .A(n9779), .B(n9778), .ZN(n9781)
         );
  AOI21_X1 U10920 ( .B1(n9782), .B2(n9791), .A(n9781), .ZN(n9796) );
  INV_X1 U10921 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9783) );
  AOI22_X1 U10922 ( .A1(n9793), .A2(n9796), .B1(n9783), .B2(n6614), .ZN(
        P1_U3483) );
  INV_X1 U10923 ( .A(n9784), .ZN(n9790) );
  INV_X1 U10924 ( .A(n9785), .ZN(n9788) );
  OAI21_X1 U10925 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(n9789) );
  AOI211_X1 U10926 ( .C1(n9792), .C2(n9791), .A(n9790), .B(n9789), .ZN(n9798)
         );
  AOI22_X1 U10927 ( .A1(n9793), .A2(n9798), .B1(n6212), .B2(n6614), .ZN(
        P1_U3489) );
  INV_X1 U10928 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U10929 ( .A1(n9799), .A2(n9795), .B1(n9794), .B2(n4846), .ZN(
        P1_U3531) );
  AOI22_X1 U10930 ( .A1(n9799), .A2(n9796), .B1(n6983), .B2(n4846), .ZN(
        P1_U3532) );
  AOI22_X1 U10931 ( .A1(n9799), .A2(n9798), .B1(n9797), .B2(n4846), .ZN(
        P1_U3534) );
  AOI21_X1 U10932 ( .B1(n9803), .B2(n9802), .A(n9801), .ZN(n9804) );
  OAI22_X1 U10933 ( .A1(n9805), .A2(n9974), .B1(n9844), .B2(n9804), .ZN(n9811)
         );
  AOI211_X1 U10934 ( .C1(n9809), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9810)
         );
  AOI211_X1 U10935 ( .C1(n9837), .C2(n4800), .A(n9811), .B(n9810), .ZN(n9817)
         );
  NAND2_X1 U10936 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  OAI211_X1 U10937 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6957), .A(n9817), .B(
        n9816), .ZN(P2_U3184) );
  AOI21_X1 U10938 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9822) );
  NOR2_X1 U10939 ( .A1(n9822), .A2(n9844), .ZN(n9823) );
  AOI211_X1 U10940 ( .C1(n9837), .C2(n9825), .A(n9824), .B(n9823), .ZN(n9826)
         );
  OAI21_X1 U10941 ( .B1(n9827), .B2(n9853), .A(n9826), .ZN(n9828) );
  INV_X1 U10942 ( .A(n9828), .ZN(n9834) );
  OAI21_X1 U10943 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9832) );
  AOI22_X1 U10944 ( .A1(n9835), .A2(P2_ADDR_REG_7__SCAN_IN), .B1(n9832), .B2(
        n9849), .ZN(n9833) );
  NAND2_X1 U10945 ( .A1(n9834), .A2(n9833), .ZN(P2_U3189) );
  AOI22_X1 U10946 ( .A1(n9837), .A2(n9836), .B1(n9835), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9857) );
  AOI21_X1 U10947 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9854) );
  AOI21_X1 U10948 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9845) );
  OR2_X1 U10949 ( .A1(n9845), .A2(n9844), .ZN(n9852) );
  OAI21_X1 U10950 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(n9850) );
  NAND2_X1 U10951 ( .A1(n9850), .A2(n9849), .ZN(n9851) );
  OAI211_X1 U10952 ( .C1(n9854), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9855)
         );
  INV_X1 U10953 ( .A(n9855), .ZN(n9856) );
  OAI211_X1 U10954 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5224), .A(n9857), .B(
        n9856), .ZN(P2_U3195) );
  AND2_X1 U10955 ( .A1(n9858), .A2(n9914), .ZN(n9859) );
  AOI21_X1 U10956 ( .B1(n9860), .B2(n9915), .A(n9859), .ZN(n9862) );
  AND2_X1 U10957 ( .A1(n9862), .A2(n9861), .ZN(n9923) );
  INV_X1 U10958 ( .A(n9923), .ZN(n9863) );
  OAI22_X1 U10959 ( .A1(n9919), .A2(P2_REG0_REG_2__SCAN_IN), .B1(n9863), .B2(
        n9921), .ZN(n9864) );
  INV_X1 U10960 ( .A(n9864), .ZN(P2_U3396) );
  INV_X1 U10961 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9869) );
  AOI22_X1 U10962 ( .A1(n9866), .A2(n9915), .B1(n9914), .B2(n9865), .ZN(n9867)
         );
  AND2_X1 U10963 ( .A1(n9868), .A2(n9867), .ZN(n9924) );
  AOI22_X1 U10964 ( .A1(n9921), .A2(n9869), .B1(n9924), .B2(n9919), .ZN(
        P2_U3399) );
  INV_X1 U10965 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9875) );
  INV_X1 U10966 ( .A(n9870), .ZN(n9874) );
  OAI21_X1 U10967 ( .B1(n9872), .B2(n9893), .A(n9871), .ZN(n9873) );
  AOI21_X1 U10968 ( .B1(n9874), .B2(n9915), .A(n9873), .ZN(n9925) );
  AOI22_X1 U10969 ( .A1(n9921), .A2(n9875), .B1(n9925), .B2(n9919), .ZN(
        P2_U3402) );
  INV_X1 U10970 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9881) );
  NOR2_X1 U10971 ( .A1(n9876), .A2(n9893), .ZN(n9878) );
  AOI211_X1 U10972 ( .C1(n9880), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9927)
         );
  AOI22_X1 U10973 ( .A1(n9921), .A2(n9881), .B1(n9927), .B2(n9919), .ZN(
        P2_U3405) );
  INV_X1 U10974 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9887) );
  OAI22_X1 U10975 ( .A1(n9883), .A2(n9902), .B1(n9882), .B2(n9893), .ZN(n9885)
         );
  NOR2_X1 U10976 ( .A1(n9883), .A2(n9901), .ZN(n9884) );
  NOR3_X1 U10977 ( .A1(n9886), .A2(n9885), .A3(n9884), .ZN(n9929) );
  AOI22_X1 U10978 ( .A1(n9921), .A2(n9887), .B1(n9929), .B2(n9919), .ZN(
        P2_U3411) );
  INV_X1 U10979 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9892) );
  OAI21_X1 U10980 ( .B1(n9889), .B2(n9893), .A(n9888), .ZN(n9890) );
  AOI21_X1 U10981 ( .B1(n9915), .B2(n9891), .A(n9890), .ZN(n9930) );
  AOI22_X1 U10982 ( .A1(n9921), .A2(n9892), .B1(n9930), .B2(n9919), .ZN(
        P2_U3414) );
  INV_X1 U10983 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10088) );
  OAI22_X1 U10984 ( .A1(n9895), .A2(n9902), .B1(n9894), .B2(n9893), .ZN(n9897)
         );
  AOI211_X1 U10985 ( .C1(n9899), .C2(n9898), .A(n9897), .B(n9896), .ZN(n9932)
         );
  AOI22_X1 U10986 ( .A1(n9921), .A2(n10088), .B1(n9932), .B2(n9919), .ZN(
        P2_U3417) );
  INV_X1 U10987 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9906) );
  AOI21_X1 U10988 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(n9904) );
  AOI211_X1 U10989 ( .C1(n9914), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9933)
         );
  AOI22_X1 U10990 ( .A1(n9921), .A2(n9906), .B1(n9933), .B2(n9919), .ZN(
        P2_U3420) );
  INV_X1 U10991 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U10992 ( .A1(n9907), .A2(n9915), .ZN(n9910) );
  NAND2_X1 U10993 ( .A1(n9908), .A2(n9914), .ZN(n9909) );
  AND3_X1 U10994 ( .A1(n9911), .A2(n9910), .A3(n9909), .ZN(n9934) );
  AOI22_X1 U10995 ( .A1(n9921), .A2(n9912), .B1(n9934), .B2(n9919), .ZN(
        P2_U3423) );
  INV_X1 U10996 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U10997 ( .A1(n9916), .A2(n9915), .B1(n9914), .B2(n9913), .ZN(n9918)
         );
  AND2_X1 U10998 ( .A1(n9918), .A2(n9917), .ZN(n9937) );
  AOI22_X1 U10999 ( .A1(n9921), .A2(n9920), .B1(n9937), .B2(n9919), .ZN(
        P2_U3426) );
  AOI22_X1 U11000 ( .A1(n9938), .A2(n9923), .B1(n9922), .B2(n9935), .ZN(
        P2_U3461) );
  AOI22_X1 U11001 ( .A1(n9938), .A2(n9924), .B1(n4824), .B2(n9935), .ZN(
        P2_U3462) );
  AOI22_X1 U11002 ( .A1(n9938), .A2(n9925), .B1(n5950), .B2(n9935), .ZN(
        P2_U3463) );
  INV_X1 U11003 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U11004 ( .A1(n9938), .A2(n9927), .B1(n9926), .B2(n9935), .ZN(
        P2_U3464) );
  AOI22_X1 U11005 ( .A1(n9938), .A2(n9929), .B1(n9928), .B2(n9935), .ZN(
        P2_U3466) );
  AOI22_X1 U11006 ( .A1(n9938), .A2(n9930), .B1(n5990), .B2(n9935), .ZN(
        P2_U3467) );
  AOI22_X1 U11007 ( .A1(n9938), .A2(n9932), .B1(n9931), .B2(n9935), .ZN(
        P2_U3468) );
  AOI22_X1 U11008 ( .A1(n9938), .A2(n9933), .B1(n5955), .B2(n9935), .ZN(
        P2_U3469) );
  AOI22_X1 U11009 ( .A1(n9938), .A2(n9934), .B1(n4818), .B2(n9935), .ZN(
        P2_U3470) );
  INV_X1 U11010 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9936) );
  AOI22_X1 U11011 ( .A1(n9938), .A2(n9937), .B1(n9936), .B2(n9935), .ZN(
        P2_U3471) );
  OAI222_X1 U11012 ( .A1(n6670), .A2(n9942), .B1(n6670), .B2(n9941), .C1(n9940), .C2(n9939), .ZN(ADD_1068_U5) );
  XOR2_X1 U11013 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11014 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9947) );
  XOR2_X1 U11015 ( .A(n9947), .B(n9946), .Z(ADD_1068_U55) );
  OAI21_X1 U11016 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(ADD_1068_U56) );
  OAI21_X1 U11017 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(ADD_1068_U57) );
  OAI21_X1 U11018 ( .B1(n9956), .B2(n9955), .A(n9954), .ZN(ADD_1068_U58) );
  OAI21_X1 U11019 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(ADD_1068_U59) );
  OAI21_X1 U11020 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(ADD_1068_U60) );
  OAI21_X1 U11021 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(ADD_1068_U61) );
  OAI21_X1 U11022 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(ADD_1068_U62) );
  OAI21_X1 U11023 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(ADD_1068_U63) );
  NAND2_X1 U11024 ( .A1(n9972), .A2(P1_D_REG_23__SCAN_IN), .ZN(n10164) );
  INV_X1 U11025 ( .A(SI_13_), .ZN(n9975) );
  INV_X1 U11026 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11027 ( .A1(n9975), .A2(keyinput101), .B1(keyinput94), .B2(n9974), 
        .ZN(n9973) );
  OAI221_X1 U11028 ( .B1(n9975), .B2(keyinput101), .C1(n9974), .C2(keyinput94), 
        .A(n9973), .ZN(n9984) );
  AOI22_X1 U11029 ( .A1(n10114), .A2(keyinput108), .B1(keyinput126), .B2(n9977), .ZN(n9976) );
  OAI221_X1 U11030 ( .B1(n10114), .B2(keyinput108), .C1(n9977), .C2(
        keyinput126), .A(n9976), .ZN(n9983) );
  INV_X1 U11031 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U11032 ( .A1(n10088), .A2(keyinput122), .B1(n10104), .B2(
        keyinput103), .ZN(n9978) );
  OAI221_X1 U11033 ( .B1(n10088), .B2(keyinput122), .C1(n10104), .C2(
        keyinput103), .A(n9978), .ZN(n9982) );
  XNOR2_X1 U11034 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(keyinput124), .ZN(n9980)
         );
  XNOR2_X1 U11035 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput82), .ZN(n9979) );
  NAND2_X1 U11036 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NOR4_X1 U11037 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(n10025)
         );
  AOI22_X1 U11038 ( .A1(n10102), .A2(keyinput114), .B1(n6498), .B2(keyinput95), 
        .ZN(n9985) );
  OAI221_X1 U11039 ( .B1(n10102), .B2(keyinput114), .C1(n6498), .C2(keyinput95), .A(n9985), .ZN(n9995) );
  AOI22_X1 U11040 ( .A1(n9988), .A2(keyinput68), .B1(n9987), .B2(keyinput125), 
        .ZN(n9986) );
  OAI221_X1 U11041 ( .B1(n9988), .B2(keyinput68), .C1(n9987), .C2(keyinput125), 
        .A(n9986), .ZN(n9994) );
  XNOR2_X1 U11042 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput65), .ZN(n9992)
         );
  XNOR2_X1 U11043 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput85), .ZN(n9991) );
  XNOR2_X1 U11044 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput111), .ZN(n9990) );
  XNOR2_X1 U11045 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput80), .ZN(n9989) );
  NAND4_X1 U11046 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), .ZN(n9993)
         );
  NOR3_X1 U11047 ( .A1(n9995), .A2(n9994), .A3(n9993), .ZN(n10024) );
  INV_X1 U11048 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9997) );
  INV_X1 U11049 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U11050 ( .A1(n9997), .A2(keyinput76), .B1(keyinput97), .B2(n10118), 
        .ZN(n9996) );
  OAI221_X1 U11051 ( .B1(n9997), .B2(keyinput76), .C1(n10118), .C2(keyinput97), 
        .A(n9996), .ZN(n10008) );
  INV_X1 U11052 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U11053 ( .A1(n10000), .A2(keyinput99), .B1(keyinput118), .B2(n9999), 
        .ZN(n9998) );
  OAI221_X1 U11054 ( .B1(n10000), .B2(keyinput99), .C1(n9999), .C2(keyinput118), .A(n9998), .ZN(n10007) );
  XNOR2_X1 U11055 ( .A(n10001), .B(keyinput77), .ZN(n10006) );
  XNOR2_X1 U11056 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput119), .ZN(n10004) );
  XNOR2_X1 U11057 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput75), .ZN(n10003) );
  XNOR2_X1 U11058 ( .A(P2_REG1_REG_28__SCAN_IN), .B(keyinput113), .ZN(n10002)
         );
  NAND3_X1 U11059 ( .A1(n10004), .A2(n10003), .A3(n10002), .ZN(n10005) );
  NOR4_X1 U11060 ( .A1(n10008), .A2(n10007), .A3(n10006), .A4(n10005), .ZN(
        n10023) );
  INV_X1 U11061 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10011) );
  INV_X1 U11062 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11063 ( .A1(n10011), .A2(keyinput73), .B1(n10010), .B2(keyinput91), 
        .ZN(n10009) );
  OAI221_X1 U11064 ( .B1(n10011), .B2(keyinput73), .C1(n10010), .C2(keyinput91), .A(n10009), .ZN(n10021) );
  INV_X1 U11065 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11066 ( .A1(n10133), .A2(keyinput100), .B1(n10013), .B2(keyinput86), .ZN(n10012) );
  OAI221_X1 U11067 ( .B1(n10133), .B2(keyinput100), .C1(n10013), .C2(
        keyinput86), .A(n10012), .ZN(n10020) );
  INV_X1 U11068 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10014) );
  XOR2_X1 U11069 ( .A(n10014), .B(keyinput72), .Z(n10018) );
  XNOR2_X1 U11070 ( .A(SI_4_), .B(keyinput69), .ZN(n10017) );
  XNOR2_X1 U11071 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput96), .ZN(n10016)
         );
  XNOR2_X1 U11072 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput71), .ZN(n10015) );
  NAND4_X1 U11073 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        n10019) );
  NOR3_X1 U11074 ( .A1(n10021), .A2(n10020), .A3(n10019), .ZN(n10022) );
  AND4_X1 U11075 ( .A1(n10025), .A2(n10024), .A3(n10023), .A4(n10022), .ZN(
        n10162) );
  OAI22_X1 U11076 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(keyinput112), .B1(
        keyinput92), .B2(P2_REG1_REG_6__SCAN_IN), .ZN(n10026) );
  AOI221_X1 U11077 ( .B1(P1_DATAO_REG_18__SCAN_IN), .B2(keyinput112), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput92), .A(n10026), .ZN(n10033) );
  OAI22_X1 U11078 ( .A1(P2_D_REG_4__SCAN_IN), .A2(keyinput98), .B1(keyinput127), .B2(P2_REG0_REG_26__SCAN_IN), .ZN(n10027) );
  AOI221_X1 U11079 ( .B1(P2_D_REG_4__SCAN_IN), .B2(keyinput98), .C1(
        P2_REG0_REG_26__SCAN_IN), .C2(keyinput127), .A(n10027), .ZN(n10032) );
  OAI22_X1 U11080 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(keyinput102), .B1(
        P2_D_REG_22__SCAN_IN), .B2(keyinput104), .ZN(n10028) );
  AOI221_X1 U11081 ( .B1(P1_REG0_REG_17__SCAN_IN), .B2(keyinput102), .C1(
        keyinput104), .C2(P2_D_REG_22__SCAN_IN), .A(n10028), .ZN(n10031) );
  OAI22_X1 U11082 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput78), .B1(
        keyinput107), .B2(SI_17_), .ZN(n10029) );
  AOI221_X1 U11083 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput78), .C1(SI_17_), 
        .C2(keyinput107), .A(n10029), .ZN(n10030) );
  NAND4_X1 U11084 ( .A1(n10033), .A2(n10032), .A3(n10031), .A4(n10030), .ZN(
        n10061) );
  OAI22_X1 U11085 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput67), .B1(
        P1_REG2_REG_18__SCAN_IN), .B2(keyinput70), .ZN(n10034) );
  AOI221_X1 U11086 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput67), .C1(
        keyinput70), .C2(P1_REG2_REG_18__SCAN_IN), .A(n10034), .ZN(n10041) );
  OAI22_X1 U11087 ( .A1(P1_REG0_REG_12__SCAN_IN), .A2(keyinput110), .B1(
        keyinput64), .B2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10035) );
  AOI221_X1 U11088 ( .B1(P1_REG0_REG_12__SCAN_IN), .B2(keyinput110), .C1(
        P1_ADDR_REG_6__SCAN_IN), .C2(keyinput64), .A(n10035), .ZN(n10040) );
  OAI22_X1 U11089 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput79), .B1(keyinput106), .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n10036) );
  AOI221_X1 U11090 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput79), .C1(
        P2_REG0_REG_16__SCAN_IN), .C2(keyinput106), .A(n10036), .ZN(n10039) );
  OAI22_X1 U11091 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput123), .B1(
        P1_REG2_REG_17__SCAN_IN), .B2(keyinput83), .ZN(n10037) );
  AOI221_X1 U11092 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput123), .C1(
        keyinput83), .C2(P1_REG2_REG_17__SCAN_IN), .A(n10037), .ZN(n10038) );
  NAND4_X1 U11093 ( .A1(n10041), .A2(n10040), .A3(n10039), .A4(n10038), .ZN(
        n10060) );
  OAI22_X1 U11094 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(keyinput117), .B1(
        keyinput121), .B2(P2_REG2_REG_29__SCAN_IN), .ZN(n10042) );
  AOI221_X1 U11095 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(keyinput117), .C1(
        P2_REG2_REG_29__SCAN_IN), .C2(keyinput121), .A(n10042), .ZN(n10049) );
  OAI22_X1 U11096 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(keyinput88), .B1(
        keyinput93), .B2(SI_31_), .ZN(n10043) );
  AOI221_X1 U11097 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(keyinput88), .C1(SI_31_), .C2(keyinput93), .A(n10043), .ZN(n10048) );
  OAI22_X1 U11098 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput74), .B1(
        P2_IR_REG_11__SCAN_IN), .B2(keyinput116), .ZN(n10044) );
  AOI221_X1 U11099 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput74), .C1(
        keyinput116), .C2(P2_IR_REG_11__SCAN_IN), .A(n10044), .ZN(n10047) );
  OAI22_X1 U11100 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput87), .B1(
        keyinput109), .B2(P2_REG2_REG_2__SCAN_IN), .ZN(n10045) );
  AOI221_X1 U11101 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG2_REG_2__SCAN_IN), .C2(keyinput109), .A(n10045), .ZN(n10046) );
  NAND4_X1 U11102 ( .A1(n10049), .A2(n10048), .A3(n10047), .A4(n10046), .ZN(
        n10059) );
  OAI22_X1 U11103 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput105), .B1(
        P1_REG0_REG_21__SCAN_IN), .B2(keyinput120), .ZN(n10050) );
  AOI221_X1 U11104 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput105), .C1(
        keyinput120), .C2(P1_REG0_REG_21__SCAN_IN), .A(n10050), .ZN(n10057) );
  OAI22_X1 U11105 ( .A1(P1_REG0_REG_6__SCAN_IN), .A2(keyinput66), .B1(
        P2_REG0_REG_18__SCAN_IN), .B2(keyinput84), .ZN(n10051) );
  AOI221_X1 U11106 ( .B1(P1_REG0_REG_6__SCAN_IN), .B2(keyinput66), .C1(
        keyinput84), .C2(P2_REG0_REG_18__SCAN_IN), .A(n10051), .ZN(n10056) );
  OAI22_X1 U11107 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(keyinput90), .B1(
        keyinput89), .B2(P1_REG3_REG_11__SCAN_IN), .ZN(n10052) );
  AOI221_X1 U11108 ( .B1(P1_DATAO_REG_12__SCAN_IN), .B2(keyinput90), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput89), .A(n10052), .ZN(n10055) );
  OAI22_X1 U11109 ( .A1(SI_3_), .A2(keyinput81), .B1(keyinput115), .B2(
        P2_IR_REG_1__SCAN_IN), .ZN(n10053) );
  AOI221_X1 U11110 ( .B1(SI_3_), .B2(keyinput81), .C1(P2_IR_REG_1__SCAN_IN), 
        .C2(keyinput115), .A(n10053), .ZN(n10054) );
  NAND4_X1 U11111 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10058) );
  NOR4_X1 U11112 ( .A1(n10061), .A2(n10060), .A3(n10059), .A4(n10058), .ZN(
        n10161) );
  AOI22_X1 U11113 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput13), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput61), .ZN(n10062) );
  OAI221_X1 U11114 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput13), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput61), .A(n10062), .ZN(n10069) );
  AOI22_X1 U11115 ( .A1(SI_31_), .A2(keyinput29), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(keyinput8), .ZN(n10063) );
  OAI221_X1 U11116 ( .B1(SI_31_), .B2(keyinput29), .C1(P1_REG2_REG_16__SCAN_IN), .C2(keyinput8), .A(n10063), .ZN(n10068) );
  AOI22_X1 U11117 ( .A1(P1_REG0_REG_6__SCAN_IN), .A2(keyinput2), .B1(
        P1_REG1_REG_25__SCAN_IN), .B2(keyinput22), .ZN(n10064) );
  OAI221_X1 U11118 ( .B1(P1_REG0_REG_6__SCAN_IN), .B2(keyinput2), .C1(
        P1_REG1_REG_25__SCAN_IN), .C2(keyinput22), .A(n10064), .ZN(n10067) );
  AOI22_X1 U11119 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(keyinput53), .B1(
        P1_REG0_REG_12__SCAN_IN), .B2(keyinput46), .ZN(n10065) );
  OAI221_X1 U11120 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(keyinput53), .C1(
        P1_REG0_REG_12__SCAN_IN), .C2(keyinput46), .A(n10065), .ZN(n10066) );
  NOR4_X1 U11121 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10100) );
  AOI22_X1 U11122 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(keyinput25), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput16), .ZN(n10070) );
  OAI221_X1 U11123 ( .B1(P1_REG3_REG_11__SCAN_IN), .B2(keyinput25), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput16), .A(n10070), .ZN(n10077) );
  AOI22_X1 U11124 ( .A1(P2_D_REG_7__SCAN_IN), .A2(keyinput4), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput10), .ZN(n10071) );
  OAI221_X1 U11125 ( .B1(P2_D_REG_7__SCAN_IN), .B2(keyinput4), .C1(
        P1_DATAO_REG_21__SCAN_IN), .C2(keyinput10), .A(n10071), .ZN(n10076) );
  AOI22_X1 U11126 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(keyinput62), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput28), .ZN(n10072) );
  OAI221_X1 U11127 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(keyinput62), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput28), .A(n10072), .ZN(n10075) );
  AOI22_X1 U11128 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput0), .B1(
        P1_REG2_REG_14__SCAN_IN), .B2(keyinput12), .ZN(n10073) );
  OAI221_X1 U11129 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput0), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(keyinput12), .A(n10073), .ZN(n10074) );
  NOR4_X1 U11130 ( .A1(n10077), .A2(n10076), .A3(n10075), .A4(n10074), .ZN(
        n10099) );
  AOI22_X1 U11131 ( .A1(P2_REG1_REG_20__SCAN_IN), .A2(keyinput35), .B1(
        P2_REG0_REG_26__SCAN_IN), .B2(keyinput63), .ZN(n10078) );
  OAI221_X1 U11132 ( .B1(P2_REG1_REG_20__SCAN_IN), .B2(keyinput35), .C1(
        P2_REG0_REG_26__SCAN_IN), .C2(keyinput63), .A(n10078), .ZN(n10085) );
  AOI22_X1 U11133 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(keyinput30), .B1(SI_4_), 
        .B2(keyinput5), .ZN(n10079) );
  OAI221_X1 U11134 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(keyinput30), .C1(SI_4_), 
        .C2(keyinput5), .A(n10079), .ZN(n10084) );
  AOI22_X1 U11135 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput32), .B1(
        P2_D_REG_4__SCAN_IN), .B2(keyinput34), .ZN(n10080) );
  OAI221_X1 U11136 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput32), .C1(
        P2_D_REG_4__SCAN_IN), .C2(keyinput34), .A(n10080), .ZN(n10083) );
  AOI22_X1 U11137 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(keyinput7), .B1(
        P1_REG3_REG_10__SCAN_IN), .B2(keyinput27), .ZN(n10081) );
  OAI221_X1 U11138 ( .B1(P2_IR_REG_28__SCAN_IN), .B2(keyinput7), .C1(
        P1_REG3_REG_10__SCAN_IN), .C2(keyinput27), .A(n10081), .ZN(n10082) );
  NOR4_X1 U11139 ( .A1(n10085), .A2(n10084), .A3(n10083), .A4(n10082), .ZN(
        n10098) );
  AOI22_X1 U11140 ( .A1(n10088), .A2(keyinput58), .B1(n10087), .B2(keyinput48), 
        .ZN(n10086) );
  OAI221_X1 U11141 ( .B1(n10088), .B2(keyinput58), .C1(n10087), .C2(keyinput48), .A(n10086), .ZN(n10096) );
  AOI22_X1 U11142 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(keyinput38), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(keyinput60), .ZN(n10089) );
  OAI221_X1 U11143 ( .B1(P1_REG0_REG_17__SCAN_IN), .B2(keyinput38), .C1(
        P1_DATAO_REG_27__SCAN_IN), .C2(keyinput60), .A(n10089), .ZN(n10095) );
  AOI22_X1 U11144 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(keyinput54), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(keyinput47), .ZN(n10090) );
  OAI221_X1 U11145 ( .B1(P2_REG0_REG_13__SCAN_IN), .B2(keyinput54), .C1(
        P1_REG2_REG_0__SCAN_IN), .C2(keyinput47), .A(n10090), .ZN(n10094) );
  XNOR2_X1 U11146 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput9), .ZN(n10092) );
  XNOR2_X1 U11147 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput18), .ZN(n10091)
         );
  NAND2_X1 U11148 ( .A1(n10092), .A2(n10091), .ZN(n10093) );
  NOR4_X1 U11149 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10097) );
  NAND4_X1 U11150 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10160) );
  AOI22_X1 U11151 ( .A1(n10102), .A2(keyinput50), .B1(keyinput45), .B2(n4799), 
        .ZN(n10101) );
  OAI221_X1 U11152 ( .B1(n10102), .B2(keyinput50), .C1(n4799), .C2(keyinput45), 
        .A(n10101), .ZN(n10112) );
  AOI22_X1 U11153 ( .A1(n10105), .A2(keyinput26), .B1(keyinput39), .B2(n10104), 
        .ZN(n10103) );
  OAI221_X1 U11154 ( .B1(n10105), .B2(keyinput26), .C1(n10104), .C2(keyinput39), .A(n10103), .ZN(n10111) );
  XNOR2_X1 U11155 ( .A(SI_3_), .B(keyinput17), .ZN(n10109) );
  XNOR2_X1 U11156 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput51), .ZN(n10108) );
  XNOR2_X1 U11157 ( .A(P2_REG1_REG_28__SCAN_IN), .B(keyinput49), .ZN(n10107)
         );
  XNOR2_X1 U11158 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput59), .ZN(n10106) );
  NAND4_X1 U11159 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10110) );
  NOR3_X1 U11160 ( .A1(n10112), .A2(n10111), .A3(n10110), .ZN(n10158) );
  AOI22_X1 U11161 ( .A1(n10115), .A2(keyinput20), .B1(n10114), .B2(keyinput44), 
        .ZN(n10113) );
  OAI221_X1 U11162 ( .B1(n10115), .B2(keyinput20), .C1(n10114), .C2(keyinput44), .A(n10113), .ZN(n10127) );
  AOI22_X1 U11163 ( .A1(n10118), .A2(keyinput33), .B1(n10117), .B2(keyinput14), 
        .ZN(n10116) );
  OAI221_X1 U11164 ( .B1(n10118), .B2(keyinput33), .C1(n10117), .C2(keyinput14), .A(n10116), .ZN(n10126) );
  AOI22_X1 U11165 ( .A1(n10121), .A2(keyinput24), .B1(n10120), .B2(keyinput23), 
        .ZN(n10119) );
  OAI221_X1 U11166 ( .B1(n10121), .B2(keyinput24), .C1(n10120), .C2(keyinput23), .A(n10119), .ZN(n10125) );
  XNOR2_X1 U11167 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput11), .ZN(n10123) );
  XNOR2_X1 U11168 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput3), .ZN(n10122)
         );
  NAND2_X1 U11169 ( .A1(n10123), .A2(n10122), .ZN(n10124) );
  NOR4_X1 U11170 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n10157) );
  AOI22_X1 U11171 ( .A1(n10130), .A2(keyinput15), .B1(n10129), .B2(keyinput43), 
        .ZN(n10128) );
  OAI221_X1 U11172 ( .B1(n10130), .B2(keyinput15), .C1(n10129), .C2(keyinput43), .A(n10128), .ZN(n10140) );
  INV_X1 U11173 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U11174 ( .A1(n10133), .A2(keyinput36), .B1(n10132), .B2(keyinput6), 
        .ZN(n10131) );
  OAI221_X1 U11175 ( .B1(n10133), .B2(keyinput36), .C1(n10132), .C2(keyinput6), 
        .A(n10131), .ZN(n10139) );
  XNOR2_X1 U11176 ( .A(P1_REG0_REG_28__SCAN_IN), .B(keyinput31), .ZN(n10137)
         );
  XNOR2_X1 U11177 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput52), .ZN(n10136) );
  XNOR2_X1 U11178 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput55), .ZN(n10135) );
  XNOR2_X1 U11179 ( .A(SI_13_), .B(keyinput37), .ZN(n10134) );
  NAND4_X1 U11180 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10138) );
  NOR3_X1 U11181 ( .A1(n10140), .A2(n10139), .A3(n10138), .ZN(n10156) );
  INV_X1 U11182 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U11183 ( .A1(n10143), .A2(keyinput56), .B1(keyinput19), .B2(n10142), 
        .ZN(n10141) );
  OAI221_X1 U11184 ( .B1(n10143), .B2(keyinput56), .C1(n10142), .C2(keyinput19), .A(n10141), .ZN(n10154) );
  INV_X1 U11185 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11186 ( .A1(n10146), .A2(keyinput1), .B1(keyinput42), .B2(n10145), 
        .ZN(n10144) );
  OAI221_X1 U11187 ( .B1(n10146), .B2(keyinput1), .C1(n10145), .C2(keyinput42), 
        .A(n10144), .ZN(n10153) );
  XNOR2_X1 U11188 ( .A(n10147), .B(keyinput40), .ZN(n10152) );
  XNOR2_X1 U11189 ( .A(P2_REG2_REG_29__SCAN_IN), .B(keyinput57), .ZN(n10150)
         );
  XNOR2_X1 U11190 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput41), .ZN(n10149) );
  XNOR2_X1 U11191 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput21), .ZN(n10148) );
  NAND3_X1 U11192 ( .A1(n10150), .A2(n10149), .A3(n10148), .ZN(n10151) );
  NOR4_X1 U11193 ( .A1(n10154), .A2(n10153), .A3(n10152), .A4(n10151), .ZN(
        n10155) );
  NAND4_X1 U11194 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10159) );
  AOI211_X1 U11195 ( .C1(n10162), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        n10163) );
  XNOR2_X1 U11196 ( .A(n10164), .B(n10163), .ZN(P1_U3302) );
  OAI21_X1 U11197 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(ADD_1068_U51) );
  OAI21_X1 U11198 ( .B1(n10170), .B2(n10169), .A(n10168), .ZN(ADD_1068_U47) );
  OAI21_X1 U11199 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(ADD_1068_U49) );
  OAI21_X1 U11200 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(ADD_1068_U48) );
  OAI21_X1 U11201 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(ADD_1068_U50) );
  AOI21_X1 U11202 ( .B1(n10182), .B2(n10181), .A(n10180), .ZN(ADD_1068_U54) );
  AOI21_X1 U11203 ( .B1(n10185), .B2(n10184), .A(n10183), .ZN(ADD_1068_U53) );
  OAI21_X1 U11204 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4845 ( .A(n5812), .Z(n5824) );
  CLKBUF_X2 U4870 ( .A(n4997), .Z(n6562) );
  XNOR2_X1 U4996 ( .A(n6416), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9109) );
endmodule

