

module b22_C_gen_AntiSAT_k_128_7 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222;

  CLKBUF_X2 U7214 ( .A(n11584), .Z(n11633) );
  CLKBUF_X2 U7215 ( .A(n6510), .Z(n8605) );
  CLKBUF_X2 U7216 ( .A(n8646), .Z(n6470) );
  XNOR2_X1 U7217 ( .A(n6468), .B(n10358), .ZN(n13020) );
  CLKBUF_X2 U7218 ( .A(n8535), .Z(n6509) );
  INV_X2 U7219 ( .A(n11835), .ZN(n11952) );
  OR2_X2 U7220 ( .A1(n10148), .A2(n7102), .ZN(n10353) );
  CLKBUF_X3 U7221 ( .A(n8891), .Z(n9723) );
  NAND2_X1 U7222 ( .A1(n12038), .A2(n8270), .ZN(n8290) );
  AND2_X1 U7223 ( .A1(n13676), .A2(n13680), .ZN(n7815) );
  AND2_X2 U7224 ( .A1(n13676), .A2(n7500), .ZN(n8138) );
  AND2_X2 U7225 ( .A1(n7499), .A2(n7500), .ZN(n8050) );
  NOR2_X2 U7226 ( .A1(n11235), .A2(n8205), .ZN(n10147) );
  NAND2_X1 U7227 ( .A1(n7494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7513) );
  NOR2_X1 U7228 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6658) );
  INV_X2 U7229 ( .A(n7773), .ZN(n8148) );
  AND2_X1 U7230 ( .A1(n12522), .A2(n9238), .ZN(n7440) );
  NOR2_X1 U7231 ( .A1(n12292), .A2(n8831), .ZN(n8832) );
  NOR2_X1 U7232 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7466) );
  OR2_X1 U7233 ( .A1(n9230), .A2(n9229), .ZN(n9231) );
  AND4_X1 U7234 ( .A1(n8799), .A2(n8798), .A3(n8797), .A4(n8978), .ZN(n8800)
         );
  NAND2_X1 U7235 ( .A1(n8920), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8921) );
  OAI21_X1 U7236 ( .B1(n7914), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7469) );
  INV_X1 U7237 ( .A(n14359), .ZN(n8270) );
  AND2_X1 U7238 ( .A1(n8270), .A2(n8269), .ZN(n8323) );
  NOR2_X1 U7239 ( .A1(n12493), .A2(n6722), .ZN(n12401) );
  INV_X1 U7240 ( .A(n11132), .ZN(n9891) );
  NAND2_X1 U7241 ( .A1(n9848), .A2(n9917), .ZN(n9849) );
  MUX2_X1 U7242 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8812), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8814) );
  AND2_X2 U7243 ( .A1(n8800), .A2(n8801), .ZN(n7430) );
  INV_X1 U7244 ( .A(n7791), .ZN(n8158) );
  AND2_X1 U7245 ( .A1(n7843), .A2(n7842), .ZN(n13629) );
  AND2_X1 U7246 ( .A1(n10274), .A2(n11977), .ZN(n11584) );
  CLKBUF_X2 U7247 ( .A(n8325), .Z(n8570) );
  INV_X1 U7248 ( .A(n8290), .ZN(n8646) );
  AND2_X1 U7249 ( .A1(n10744), .A2(n10891), .ZN(n10825) );
  INV_X1 U7250 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6497) );
  OAI21_X1 U7251 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n9385), .A(n9384), .ZN(
        n9433) );
  NAND2_X1 U7252 ( .A1(n9193), .A2(n9192), .ZN(n12506) );
  NAND2_X1 U7253 ( .A1(n12157), .A2(n12158), .ZN(n12117) );
  AOI21_X1 U7254 ( .B1(n8817), .B2(n11282), .A(n6664), .ZN(n10165) );
  OAI21_X1 U7255 ( .B1(n6531), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8830) );
  INV_X1 U7256 ( .A(n9862), .ZN(n11084) );
  XNOR2_X1 U7257 ( .A(n13608), .B(n13270), .ZN(n13433) );
  NAND2_X1 U7258 ( .A1(n8651), .A2(n14362), .ZN(n8304) );
  AND2_X1 U7259 ( .A1(n11975), .A2(n11794), .ZN(n14302) );
  INV_X1 U7260 ( .A(n9961), .ZN(n9960) );
  XNOR2_X1 U7261 ( .A(n8830), .B(n6723), .ZN(n12105) );
  NAND4_X1 U7262 ( .A1(n7586), .A2(n7585), .A3(n7584), .A4(n7583), .ZN(n13153)
         );
  NAND2_X1 U7263 ( .A1(n8268), .A2(n14352), .ZN(n14359) );
  INV_X1 U7264 ( .A(n14106), .ZN(n6857) );
  XOR2_X1 U7265 ( .A(n13585), .B(n10851), .Z(n6466) );
  XNOR2_X1 U7266 ( .A(n7469), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10148) );
  INV_X2 U7268 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9436) );
  NAND2_X2 U7269 ( .A1(n12792), .A2(n9694), .ZN(n12779) );
  XNOR2_X2 U7270 ( .A(n11665), .B(n11666), .ZN(n13131) );
  NAND2_X4 U7271 ( .A1(n7937), .A2(n7936), .ZN(n13608) );
  AND3_X2 U7272 ( .A1(n7467), .A2(n6658), .A3(n7466), .ZN(n7488) );
  INV_X1 U7273 ( .A(n10776), .ZN(n6467) );
  AOI21_X2 U7274 ( .B1(n13459), .B2(n6761), .A(n6759), .ZN(n13405) );
  NOR2_X4 U7275 ( .A1(n13460), .A2(n13464), .ZN(n13459) );
  NAND2_X2 U7276 ( .A1(n12148), .A2(n12147), .ZN(n12143) );
  NAND2_X2 U7277 ( .A1(n12057), .A2(n11663), .ZN(n11665) );
  NAND2_X2 U7278 ( .A1(n9762), .A2(n12184), .ZN(n11424) );
  XNOR2_X2 U7279 ( .A(n9390), .B(n9389), .ZN(n9431) );
  NAND2_X2 U7280 ( .A1(n6724), .A2(n9388), .ZN(n9390) );
  NAND2_X2 U7281 ( .A1(n13002), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7428) );
  AND2_X2 U7283 ( .A1(n7386), .A2(n7383), .ZN(n12698) );
  NAND2_X2 U7284 ( .A1(n6663), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8806) );
  CLKBUF_X2 U7285 ( .A(n10357), .Z(n6468) );
  INV_X2 U7286 ( .A(n8841), .ZN(n8839) );
  XNOR2_X2 U7287 ( .A(n7428), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8841) );
  XNOR2_X2 U7288 ( .A(n9849), .B(n14408), .ZN(n14401) );
  OAI222_X1 U7289 ( .A1(n9336), .A2(P3_U3151), .B1(n13004), .B2(n12321), .C1(
        n12387), .C2(n12320), .ZN(P3_U3267) );
  NAND2_X1 U7290 ( .A1(n9336), .A2(n9885), .ZN(n6501) );
  XNOR2_X2 U7291 ( .A(n13513), .B(n13261), .ZN(n13508) );
  INV_X2 U7292 ( .A(n13629), .ZN(n13513) );
  XNOR2_X2 U7293 ( .A(n9394), .B(n9393), .ZN(n9429) );
  NAND2_X2 U7294 ( .A1(n9391), .A2(n9392), .ZN(n9394) );
  XNOR2_X2 U7295 ( .A(n8921), .B(n8796), .ZN(n9862) );
  XNOR2_X2 U7296 ( .A(n8901), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U7297 ( .A1(n12706), .A2(n9776), .ZN(n11774) );
  OR2_X1 U7298 ( .A1(n13095), .A2(n6466), .ZN(n6799) );
  NAND2_X1 U7299 ( .A1(n14133), .A2(n14144), .ZN(n14132) );
  AND2_X1 U7300 ( .A1(n13396), .A2(n6602), .ZN(n13334) );
  NAND2_X1 U7301 ( .A1(n14505), .A2(n11886), .ZN(n14224) );
  INV_X1 U7302 ( .A(n11659), .ZN(n11418) );
  NAND2_X1 U7303 ( .A1(n8547), .A2(n8546), .ZN(n14160) );
  NAND2_X1 U7304 ( .A1(n8473), .A2(n8472), .ZN(n14513) );
  INV_X2 U7305 ( .A(n12143), .ZN(n15104) );
  CLKBUF_X1 U7306 ( .A(n10293), .Z(n14248) );
  NOR2_X1 U7307 ( .A1(n14641), .A2(n14240), .ZN(n14242) );
  NAND2_X1 U7308 ( .A1(n8839), .A2(n8846), .ZN(n8892) );
  INV_X1 U7310 ( .A(n8304), .ZN(n8535) );
  INV_X1 U7311 ( .A(n8312), .ZN(n9970) );
  INV_X1 U7312 ( .A(n10354), .ZN(n10338) );
  INV_X2 U7313 ( .A(n10150), .ZN(n10144) );
  MUX2_X1 U7314 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8266), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8268) );
  NAND2_X2 U7315 ( .A1(n8240), .A2(n10155), .ZN(n7161) );
  CLKBUF_X2 U7316 ( .A(n11027), .Z(n6500) );
  NOR2_X2 U7317 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8314) );
  AOI211_X1 U7318 ( .C1(n8213), .C2(n10269), .A(n8237), .B(n8204), .ZN(n8222)
         );
  AOI21_X1 U7319 ( .B1(n8185), .B2(n8184), .A(n8183), .ZN(n8213) );
  AOI21_X1 U7320 ( .B1(n9668), .B2(n14698), .A(n9667), .ZN(n9669) );
  NOR2_X1 U7321 ( .A1(n12299), .A2(n7065), .ZN(n9821) );
  AND2_X1 U7322 ( .A1(n12860), .A2(n15182), .ZN(n6671) );
  OR2_X1 U7323 ( .A1(n11772), .A2(n11778), .ZN(n12860) );
  OR2_X1 U7324 ( .A1(n9814), .A2(n12981), .ZN(n9820) );
  NAND2_X1 U7325 ( .A1(n6687), .A2(n6482), .ZN(n6481) );
  NAND2_X1 U7326 ( .A1(n6862), .A2(n6860), .ZN(n12101) );
  AOI21_X1 U7327 ( .B1(n6483), .B2(n12016), .A(n14672), .ZN(n6482) );
  NAND2_X1 U7328 ( .A1(n9374), .A2(n8629), .ZN(n6483) );
  OR2_X1 U7329 ( .A1(n9369), .A2(n12014), .ZN(n9374) );
  OAI21_X1 U7330 ( .B1(n11947), .B2(n7366), .A(n7367), .ZN(n11951) );
  OR2_X1 U7331 ( .A1(n14061), .A2(n14060), .ZN(n14063) );
  AND2_X1 U7332 ( .A1(n7440), .A2(n12400), .ZN(n6722) );
  NAND2_X1 U7333 ( .A1(n13763), .A2(n12351), .ZN(n13842) );
  AOI21_X1 U7334 ( .B1(n13302), .B2(n13301), .A(n13300), .ZN(n13557) );
  NOR2_X1 U7335 ( .A1(n14028), .A2(n14644), .ZN(n14265) );
  NAND2_X1 U7336 ( .A1(n14075), .A2(n7149), .ZN(n14068) );
  NAND2_X1 U7337 ( .A1(n14102), .A2(n6478), .ZN(n14075) );
  NAND2_X1 U7338 ( .A1(n14102), .A2(n8588), .ZN(n14077) );
  AND2_X1 U7339 ( .A1(n12277), .A2(n9709), .ZN(n12651) );
  AND2_X1 U7340 ( .A1(n9351), .A2(n9350), .ZN(n12303) );
  OAI21_X1 U7341 ( .B1(n14143), .B2(n14144), .A(n8565), .ZN(n14121) );
  NAND2_X1 U7342 ( .A1(n14164), .A2(n8555), .ZN(n14143) );
  INV_X1 U7343 ( .A(n13677), .ZN(n6486) );
  NAND2_X1 U7344 ( .A1(n14162), .A2(n14161), .ZN(n14164) );
  OR2_X1 U7345 ( .A1(n6965), .A2(n14033), .ZN(n9377) );
  AOI211_X1 U7346 ( .C1(n7243), .C2(n6511), .A(n13344), .B(n13281), .ZN(n6895)
         );
  NOR2_X1 U7347 ( .A1(n6472), .A2(n8545), .ZN(n14162) );
  OAI21_X1 U7348 ( .B1(n13700), .B2(n14316), .A(n9666), .ZN(n9667) );
  AOI21_X1 U7349 ( .B1(n14187), .B2(n8530), .A(n6473), .ZN(n6472) );
  AND2_X1 U7350 ( .A1(n12013), .A2(n8588), .ZN(n6478) );
  NAND2_X1 U7351 ( .A1(n8264), .A2(n8263), .ZN(n12382) );
  OAI21_X1 U7352 ( .B1(n14187), .B2(n8529), .A(n8530), .ZN(n14167) );
  NAND2_X1 U7353 ( .A1(n14225), .A2(n8505), .ZN(n14202) );
  XNOR2_X1 U7354 ( .A(n8122), .B(n8121), .ZN(n12036) );
  NAND2_X1 U7355 ( .A1(n6902), .A2(n6901), .ZN(n13428) );
  NOR2_X2 U7356 ( .A1(n13411), .A2(n13591), .ZN(n13396) );
  NAND2_X1 U7357 ( .A1(n14226), .A2(n14227), .ZN(n14225) );
  AND2_X1 U7358 ( .A1(n6479), .A2(n7446), .ZN(n14226) );
  OR2_X1 U7359 ( .A1(n13703), .A2(n13704), .ZN(n13701) );
  AND2_X1 U7360 ( .A1(n14554), .A2(n9472), .ZN(n9476) );
  NAND2_X1 U7361 ( .A1(n11385), .A2(n8469), .ZN(n11516) );
  NAND2_X1 U7362 ( .A1(n6751), .A2(n6752), .ZN(n13703) );
  NAND2_X1 U7363 ( .A1(n8557), .A2(n8556), .ZN(n14301) );
  NAND2_X1 U7364 ( .A1(n8022), .A2(n8021), .ZN(n13383) );
  NAND2_X1 U7365 ( .A1(n11386), .A2(n12004), .ZN(n11385) );
  NAND2_X1 U7366 ( .A1(n13131), .A2(n11664), .ZN(n13141) );
  OR2_X1 U7367 ( .A1(n11551), .A2(n7324), .ZN(n6751) );
  NAND2_X1 U7368 ( .A1(n7144), .A2(n7145), .ZN(n11386) );
  NAND2_X1 U7369 ( .A1(n8005), .A2(n8004), .ZN(n13591) );
  NOR2_X1 U7370 ( .A1(n11528), .A2(n11527), .ZN(n11529) );
  OR2_X1 U7371 ( .A1(n8492), .A2(n11482), .ZN(n7446) );
  NAND2_X1 U7372 ( .A1(n6474), .A2(n14168), .ZN(n6473) );
  INV_X1 U7373 ( .A(n9357), .ZN(n6480) );
  NAND2_X1 U7374 ( .A1(n8426), .A2(n8425), .ZN(n11352) );
  AND2_X1 U7375 ( .A1(n11986), .A2(n11481), .ZN(n11482) );
  NAND2_X1 U7376 ( .A1(n11886), .A2(n11881), .ZN(n11986) );
  OR2_X1 U7377 ( .A1(n11583), .A2(n14511), .ZN(n11886) );
  CLKBUF_X1 U7378 ( .A(n11583), .Z(n6670) );
  NAND2_X1 U7379 ( .A1(n8529), .A2(n8530), .ZN(n6474) );
  NAND2_X1 U7380 ( .A1(n8537), .A2(n8536), .ZN(n8544) );
  NAND2_X1 U7381 ( .A1(n6685), .A2(n8483), .ZN(n11583) );
  NAND2_X1 U7382 ( .A1(n10866), .A2(n10865), .ZN(n10995) );
  XNOR2_X1 U7383 ( .A(n7839), .B(n7838), .ZN(n10451) );
  NAND2_X1 U7384 ( .A1(n11140), .A2(n11996), .ZN(n8398) );
  OAI21_X1 U7385 ( .B1(n8371), .B2(n6476), .A(n6475), .ZN(n11140) );
  NAND2_X1 U7386 ( .A1(n8371), .A2(n8370), .ZN(n10832) );
  OR2_X1 U7387 ( .A1(n7929), .A2(n7191), .ZN(n6953) );
  XNOR2_X1 U7388 ( .A(n7835), .B(n7858), .ZN(n10420) );
  XNOR2_X1 U7389 ( .A(n7931), .B(SI_18_), .ZN(n7929) );
  NAND2_X1 U7390 ( .A1(n7806), .A2(n7805), .ZN(n13641) );
  XNOR2_X1 U7391 ( .A(n7857), .B(SI_14_), .ZN(n7835) );
  OAI21_X1 U7392 ( .B1(n7913), .B2(n7912), .A(n7911), .ZN(n7931) );
  OAI21_X1 U7393 ( .B1(n11199), .B2(n7339), .A(n7337), .ZN(n11327) );
  NAND2_X1 U7394 ( .A1(n7219), .A2(n7224), .ZN(n7857) );
  NAND2_X1 U7395 ( .A1(n8444), .A2(n8443), .ZN(n11866) );
  NAND2_X1 U7396 ( .A1(n8340), .A2(n8339), .ZN(n6489) );
  NAND2_X1 U7397 ( .A1(n7794), .A2(n7793), .ZN(n7819) );
  NAND2_X1 U7398 ( .A1(n13519), .A2(n10606), .ZN(n10633) );
  NAND2_X1 U7399 ( .A1(n8388), .A2(n8387), .ZN(n14668) );
  INV_X1 U7400 ( .A(n11997), .ZN(n6476) );
  NAND2_X1 U7401 ( .A1(n7705), .A2(n7704), .ZN(n11703) );
  NOR2_X1 U7402 ( .A1(n11839), .A2(n13880), .ZN(n8385) );
  NAND2_X1 U7403 ( .A1(n8377), .A2(n8376), .ZN(n11839) );
  NAND2_X1 U7404 ( .A1(n7661), .A2(n7660), .ZN(n14919) );
  CLKBUF_X1 U7405 ( .A(n12798), .Z(n12813) );
  INV_X1 U7406 ( .A(n8370), .ZN(n6477) );
  NAND2_X1 U7407 ( .A1(n7720), .A2(n7719), .ZN(n7723) );
  NOR2_X1 U7408 ( .A1(n11089), .A2(n9838), .ZN(n9839) );
  NAND2_X1 U7409 ( .A1(n6484), .A2(n8306), .ZN(n10519) );
  NAND2_X1 U7410 ( .A1(n15209), .A2(n9446), .ZN(n9451) );
  NAND2_X1 U7411 ( .A1(n12166), .A2(n12162), .ZN(n12112) );
  NAND2_X1 U7412 ( .A1(n10234), .A2(n10235), .ZN(n10509) );
  NAND2_X1 U7413 ( .A1(n11987), .A2(n14255), .ZN(n6484) );
  NAND2_X1 U7414 ( .A1(n7619), .A2(n7618), .ZN(n14904) );
  AND2_X1 U7415 ( .A1(n11818), .A2(n11817), .ZN(n11812) );
  NAND2_X1 U7416 ( .A1(n8346), .A2(n8345), .ZN(n11829) );
  NAND2_X1 U7417 ( .A1(n15211), .A2(n15210), .ZN(n15209) );
  XNOR2_X1 U7418 ( .A(n6725), .B(n9444), .ZN(n15211) );
  CLKBUF_X1 U7419 ( .A(n9675), .Z(n12606) );
  NAND2_X1 U7420 ( .A1(n10436), .A2(n10232), .ZN(n10235) );
  NAND2_X1 U7421 ( .A1(n11800), .A2(n11802), .ZN(n11987) );
  INV_X1 U7422 ( .A(n11801), .ZN(n11990) );
  NAND4_X2 U7423 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n12605)
         );
  NAND2_X1 U7424 ( .A1(n10463), .A2(n14641), .ZN(n11802) );
  NAND2_X1 U7425 ( .A1(n7595), .A2(n6810), .ZN(n13076) );
  NAND2_X1 U7426 ( .A1(n8285), .A2(n6537), .ZN(n13884) );
  INV_X1 U7427 ( .A(n10464), .ZN(n13885) );
  NOR2_X1 U7428 ( .A1(n11073), .A2(n7445), .ZN(n9836) );
  NAND2_X1 U7429 ( .A1(n8305), .A2(n10293), .ZN(n11800) );
  INV_X1 U7430 ( .A(n10293), .ZN(n10463) );
  AND2_X1 U7431 ( .A1(n8330), .A2(n8329), .ZN(n10464) );
  BUF_X2 U7432 ( .A(n10602), .Z(n13470) );
  AND3_X1 U7433 ( .A1(n8328), .A2(n8327), .A3(n8326), .ZN(n8329) );
  CLKBUF_X3 U7434 ( .A(n8892), .Z(n12085) );
  OAI211_X2 U7435 ( .C1(n8356), .C2(n9999), .A(n8335), .B(n8334), .ZN(n10714)
         );
  NAND2_X1 U7436 ( .A1(n7153), .A2(n7152), .ZN(n10491) );
  AND3_X1 U7437 ( .A1(n8309), .A2(n8308), .A3(n8307), .ZN(n8311) );
  NAND4_X1 U7438 ( .A1(n8294), .A2(n8293), .A3(n8292), .A4(n8291), .ZN(n10293)
         );
  AND2_X1 U7439 ( .A1(n8839), .A2(n8840), .ZN(n6504) );
  INV_X2 U7440 ( .A(n8356), .ZN(n11972) );
  BUF_X2 U7441 ( .A(n8331), .Z(n11971) );
  NAND2_X1 U7442 ( .A1(n8331), .A2(n8295), .ZN(n7134) );
  BUF_X2 U7443 ( .A(n8323), .Z(n6510) );
  OR2_X1 U7444 ( .A1(n9834), .A2(n9891), .ZN(n6727) );
  INV_X1 U7445 ( .A(n8290), .ZN(n6471) );
  NAND2_X1 U7446 ( .A1(n8325), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8293) );
  AND2_X1 U7447 ( .A1(n6505), .A2(n9961), .ZN(n8313) );
  NAND2_X1 U7448 ( .A1(n8707), .A2(n8706), .ZN(n14367) );
  XNOR2_X1 U7449 ( .A(n8838), .B(n8837), .ZN(n8840) );
  NAND2_X2 U7450 ( .A1(n6492), .A2(P2_U3088), .ZN(n13685) );
  NAND2_X1 U7451 ( .A1(n11017), .A2(n11016), .ZN(n11015) );
  NAND2_X2 U7452 ( .A1(n6492), .A2(P1_U3086), .ZN(n14363) );
  XNOR2_X1 U7453 ( .A(n7493), .B(n6659), .ZN(n13676) );
  NAND2_X2 U7454 ( .A1(n8262), .A2(n8261), .ZN(n14362) );
  XNOR2_X1 U7455 ( .A(n7590), .B(SI_3_), .ZN(n7587) );
  NAND2_X1 U7456 ( .A1(n7479), .A2(n7478), .ZN(n11235) );
  NAND2_X1 U7457 ( .A1(n7479), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7475) );
  MUX2_X1 U7458 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8260), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8262) );
  NAND2_X1 U7459 ( .A1(n8261), .A2(n7063), .ZN(n7062) );
  OR2_X1 U7460 ( .A1(n8808), .A2(n8807), .ZN(n8809) );
  NAND2_X1 U7461 ( .A1(n7524), .A2(SI_0_), .ZN(n7542) );
  NOR2_X1 U7462 ( .A1(n9114), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n9132) );
  XNOR2_X1 U7463 ( .A(n7480), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8205) );
  AND2_X1 U7464 ( .A1(n7677), .A2(n7306), .ZN(n7866) );
  XNOR2_X1 U7465 ( .A(n8886), .B(P3_IR_REG_2__SCAN_IN), .ZN(n11027) );
  AND2_X1 U7466 ( .A1(n8256), .A2(n7151), .ZN(n7150) );
  NOR2_X1 U7467 ( .A1(n7484), .A2(n8214), .ZN(n7490) );
  AND3_X1 U7468 ( .A1(n6990), .A2(n6989), .A3(n6995), .ZN(n6988) );
  NOR2_X1 U7469 ( .A1(n7487), .A2(n7486), .ZN(n7489) );
  AND2_X1 U7470 ( .A1(n8257), .A2(n8258), .ZN(n7381) );
  AND2_X1 U7471 ( .A1(n8250), .A2(n8251), .ZN(n7357) );
  AND2_X1 U7472 ( .A1(n6992), .A2(n7429), .ZN(n6989) );
  AND2_X1 U7473 ( .A1(n6994), .A2(n6993), .ZN(n6990) );
  INV_X1 U7474 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8829) );
  INV_X1 U7475 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6993) );
  NOR2_X1 U7476 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8798) );
  INV_X1 U7477 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8372) );
  INV_X1 U7478 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8796) );
  INV_X1 U7479 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n6994) );
  INV_X1 U7480 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n6995) );
  INV_X4 U7481 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7482 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8343) );
  INV_X1 U7483 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8978) );
  INV_X1 U7484 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8250) );
  INV_X1 U7485 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9115) );
  NOR2_X1 U7486 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8427) );
  NOR2_X1 U7487 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8246) );
  NOR2_X1 U7488 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n8245) );
  NOR2_X1 U7489 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7467) );
  INV_X1 U7490 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6488) );
  INV_X1 U7491 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6487) );
  INV_X1 U7492 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7429) );
  NOR2_X1 U7493 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8799) );
  NOR2_X1 U7494 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7470) );
  NOR2_X1 U7495 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7471) );
  NOR2_X1 U7496 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7472) );
  INV_X1 U7497 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8226) );
  INV_X4 U7498 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X4 U7499 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  AND2_X1 U7500 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n7063) );
  INV_X1 U7501 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7482) );
  INV_X1 U7502 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8224) );
  NOR2_X1 U7503 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7461) );
  NOR2_X1 U7504 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7462) );
  XNOR2_X1 U7505 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n9434) );
  INV_X1 U7506 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8825) );
  AOI21_X1 U7507 ( .B1(n11997), .B2(n6477), .A(n8385), .ZN(n6475) );
  NAND3_X1 U7508 ( .A1(n11385), .A2(n8469), .A3(n8493), .ZN(n6479) );
  NAND3_X1 U7509 ( .A1(n6481), .A2(n9358), .A3(n6480), .ZN(n12299) );
  NAND2_X1 U7510 ( .A1(n8312), .A2(n8331), .ZN(n6485) );
  NAND3_X1 U7511 ( .A1(n8317), .A2(n6485), .A3(n8318), .ZN(n11809) );
  NAND2_X1 U7512 ( .A1(n6486), .A2(n8331), .ZN(n11956) );
  AND2_X2 U7513 ( .A1(n6506), .A2(n9960), .ZN(n8331) );
  NAND4_X1 U7514 ( .A1(n8372), .A2(n8343), .A3(n6488), .A4(n6487), .ZN(n8247)
         );
  NAND2_X1 U7515 ( .A1(n6489), .A2(n10701), .ZN(n8355) );
  XNOR2_X1 U7516 ( .A(n6489), .B(n10701), .ZN(n10702) );
  NAND2_X1 U7517 ( .A1(n8702), .A2(n7381), .ZN(n8261) );
  NOR2_X1 U7518 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6490) );
  INV_X1 U7519 ( .A(n11516), .ZN(n6491) );
  INV_X1 U7520 ( .A(n9960), .ZN(n6492) );
  INV_X4 U7521 ( .A(n7547), .ZN(n9961) );
  NAND2_X1 U7522 ( .A1(n12837), .A2(n6496), .ZN(n6493) );
  AND2_X1 U7523 ( .A1(n6493), .A2(n6494), .ZN(n12816) );
  OR2_X1 U7524 ( .A1(n6495), .A2(n12824), .ZN(n6494) );
  INV_X1 U7525 ( .A(n12205), .ZN(n6495) );
  AND2_X1 U7526 ( .A1(n12201), .A2(n12205), .ZN(n6496) );
  NOR2_X2 U7527 ( .A1(n14397), .A2(n14398), .ZN(n14396) );
  INV_X1 U7528 ( .A(n10714), .ZN(n10558) );
  NAND4_X4 U7529 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n9672)
         );
  NOR2_X1 U7530 ( .A1(n12859), .A2(n6671), .ZN(n12929) );
  NAND2_X1 U7531 ( .A1(n8321), .A2(n8320), .ZN(n10548) );
  XNOR2_X2 U7532 ( .A(n6498), .B(n6497), .ZN(n8269) );
  NOR2_X1 U7533 ( .A1(n8267), .A2(n14351), .ZN(n6498) );
  XNOR2_X1 U7534 ( .A(n11849), .B(n13878), .ZN(n11999) );
  NAND2_X1 U7535 ( .A1(n9754), .A2(n12140), .ZN(n10775) );
  XNOR2_X1 U7536 ( .A(n13884), .B(n14652), .ZN(n11991) );
  NAND2_X4 U7537 ( .A1(n8311), .A2(n8310), .ZN(n8319) );
  INV_X2 U7538 ( .A(n7161), .ZN(n6499) );
  NAND2_X1 U7539 ( .A1(n6471), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8294) );
  OAI222_X1 U7540 ( .A1(P1_U3086), .A2(n12038), .B1(n14366), .B2(n13677), .C1(
        n12077), .C2(n14363), .ZN(P1_U3325) );
  NOR2_X2 U7541 ( .A1(n10637), .A2(n14919), .ZN(n6984) );
  NAND2_X1 U7542 ( .A1(n9336), .A2(n9885), .ZN(n6502) );
  NAND2_X2 U7543 ( .A1(n14132), .A2(n8684), .ZN(n14118) );
  AND2_X1 U7544 ( .A1(n8839), .A2(n8840), .ZN(n6503) );
  AND2_X1 U7545 ( .A1(n8839), .A2(n8840), .ZN(n12083) );
  NAND2_X1 U7546 ( .A1(n9336), .A2(n9885), .ZN(n6507) );
  INV_X1 U7547 ( .A(n8269), .ZN(n12038) );
  AND2_X1 U7548 ( .A1(n8269), .A2(n14359), .ZN(n8324) );
  NAND2_X1 U7549 ( .A1(n8651), .A2(n14362), .ZN(n6505) );
  NAND2_X1 U7550 ( .A1(n8651), .A2(n14362), .ZN(n6506) );
  OAI222_X1 U7551 ( .A1(n8651), .A2(P1_U3086), .B1(n14366), .B2(n13686), .C1(
        n12037), .C2(n14363), .ZN(P1_U3327) );
  NAND2_X1 U7552 ( .A1(n8841), .A2(n8846), .ZN(n8891) );
  NAND2_X1 U7553 ( .A1(n8841), .A2(n8840), .ZN(n8913) );
  NAND2_X1 U7554 ( .A1(n9336), .A2(n9885), .ZN(n9855) );
  INV_X4 U7555 ( .A(n13510), .ZN(n10602) );
  AND2_X4 U7556 ( .A1(n10267), .A2(n11012), .ZN(n13510) );
  NAND3_X2 U7557 ( .A1(n8297), .A2(n7134), .A3(n8298), .ZN(n14641) );
  XNOR2_X2 U7558 ( .A(n10623), .B(n8193), .ZN(n10227) );
  INV_X2 U7559 ( .A(n13018), .ZN(n10623) );
  AND3_X4 U7560 ( .A1(n8341), .A2(n8481), .A3(n8249), .ZN(n8533) );
  NAND2_X2 U7561 ( .A1(n9336), .A2(n9885), .ZN(n6508) );
  NOR2_X2 U7562 ( .A1(n13471), .A2(n13612), .ZN(n6978) );
  INV_X1 U7563 ( .A(n6674), .ZN(n6673) );
  AND3_X2 U7564 ( .A1(n7357), .A2(n8314), .A3(n6811), .ZN(n8341) );
  AND2_X2 U7565 ( .A1(n8533), .A2(n7150), .ZN(n8702) );
  OAI21_X2 U7566 ( .B1(n10518), .B2(n11990), .A(n8655), .ZN(n7057) );
  NAND2_X1 U7567 ( .A1(n8660), .A2(n8659), .ZN(n10817) );
  INV_X1 U7568 ( .A(n14641), .ZN(n8305) );
  OR2_X1 U7569 ( .A1(n12315), .A2(n14219), .ZN(n6694) );
  OAI21_X2 U7570 ( .B1(n14202), .B2(n8517), .A(n8678), .ZN(n14187) );
  AOI21_X1 U7571 ( .B1(n7217), .B2(n6940), .A(n6939), .ZN(n6938) );
  INV_X1 U7572 ( .A(n7880), .ZN(n6939) );
  INV_X1 U7573 ( .A(n7220), .ZN(n6940) );
  AOI21_X1 U7574 ( .B1(n11779), .B2(n7402), .A(n7455), .ZN(n7398) );
  NAND2_X1 U7575 ( .A1(n12950), .A2(n12589), .ZN(n7394) );
  OR2_X1 U7576 ( .A1(n12956), .A2(n12551), .ZN(n12239) );
  INV_X1 U7577 ( .A(n12370), .ZN(n12343) );
  INV_X1 U7578 ( .A(n14204), .ZN(n7088) );
  XNOR2_X1 U7579 ( .A(n12858), .B(n12585), .ZN(n12261) );
  NOR2_X1 U7580 ( .A1(n13239), .A2(n7182), .ZN(n7181) );
  INV_X1 U7581 ( .A(n7184), .ZN(n7182) );
  AOI21_X1 U7582 ( .B1(n7230), .B2(n7228), .A(n6558), .ZN(n7227) );
  INV_X1 U7583 ( .A(n7234), .ZN(n7228) );
  OAI211_X1 U7584 ( .C1(n12136), .C2(n12139), .A(n9754), .B(n12276), .ZN(n6709) );
  NAND2_X1 U7585 ( .A1(n7291), .A2(n7290), .ZN(n7824) );
  NAND2_X1 U7586 ( .A1(n7808), .A2(n7810), .ZN(n7290) );
  NAND2_X1 U7587 ( .A1(n6831), .A2(n11928), .ZN(n6830) );
  NAND2_X1 U7588 ( .A1(n7359), .A2(n7358), .ZN(n6831) );
  NAND2_X1 U7589 ( .A1(n6812), .A2(n11918), .ZN(n11922) );
  NAND2_X1 U7590 ( .A1(n6815), .A2(n11916), .ZN(n11920) );
  AOI21_X1 U7591 ( .B1(n12301), .B2(n11952), .A(n6689), .ZN(n6841) );
  AND2_X1 U7592 ( .A1(n13696), .A2(n11835), .ZN(n6689) );
  AOI21_X1 U7593 ( .B1(n6891), .B2(n6893), .A(n7260), .ZN(n6890) );
  AND2_X1 U7594 ( .A1(n7464), .A2(n7465), .ZN(n7309) );
  INV_X1 U7595 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U7596 ( .A1(n8040), .A2(n8039), .ZN(n6917) );
  AND2_X1 U7597 ( .A1(n7344), .A2(n7343), .ZN(n7342) );
  INV_X1 U7598 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7343) );
  NAND2_X1 U7599 ( .A1(n7929), .A2(n6952), .ZN(n6954) );
  AND2_X1 U7600 ( .A1(n7932), .A2(n6958), .ZN(n6952) );
  INV_X1 U7601 ( .A(n7954), .ZN(n6958) );
  INV_X1 U7602 ( .A(n7217), .ZN(n6941) );
  INV_X1 U7603 ( .A(n7762), .ZN(n6920) );
  NAND2_X1 U7604 ( .A1(n7765), .A2(n9967), .ZN(n7793) );
  OR2_X1 U7605 ( .A1(n9919), .A2(n14408), .ZN(n9921) );
  NAND2_X1 U7606 ( .A1(n7404), .A2(n7406), .ZN(n7403) );
  INV_X1 U7607 ( .A(n7408), .ZN(n7404) );
  NAND2_X1 U7608 ( .A1(n12663), .A2(n7406), .ZN(n7405) );
  INV_X1 U7609 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n6991) );
  INV_X1 U7610 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U7611 ( .A1(n8980), .A2(n8755), .ZN(n7273) );
  INV_X1 U7612 ( .A(n13455), .ZN(n7247) );
  NAND2_X1 U7613 ( .A1(n13612), .A2(n13462), .ZN(n7189) );
  NOR2_X1 U7614 ( .A1(n7231), .A2(n10989), .ZN(n7230) );
  INV_X1 U7615 ( .A(n7233), .ZN(n7231) );
  INV_X1 U7616 ( .A(n10233), .ZN(n10234) );
  AOI21_X1 U7617 ( .B1(n7177), .B2(n13247), .A(n6596), .ZN(n7175) );
  INV_X1 U7618 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7516) );
  AND2_X1 U7619 ( .A1(n7488), .A2(n7309), .ZN(n7308) );
  OR2_X1 U7620 ( .A1(n11559), .A2(n7326), .ZN(n7325) );
  INV_X1 U7621 ( .A(n11338), .ZN(n6734) );
  NOR2_X1 U7622 ( .A1(n11326), .A2(n7341), .ZN(n6738) );
  NOR2_X1 U7623 ( .A1(n6563), .A2(n6520), .ZN(n7068) );
  AND2_X1 U7624 ( .A1(n14060), .A2(n8600), .ZN(n7149) );
  AND2_X1 U7625 ( .A1(n11791), .A2(n11120), .ZN(n11975) );
  OAI21_X1 U7626 ( .B1(n8080), .B2(n6632), .A(n6926), .ZN(n8111) );
  AND2_X1 U7627 ( .A1(n6929), .A2(n6927), .ZN(n6926) );
  NAND2_X1 U7628 ( .A1(n6934), .A2(n6930), .ZN(n6929) );
  NAND2_X1 U7629 ( .A1(n8040), .A2(n6527), .ZN(n7202) );
  AND2_X1 U7630 ( .A1(n7221), .A2(n7856), .ZN(n7220) );
  NAND2_X1 U7631 ( .A1(n7222), .A2(n7224), .ZN(n7221) );
  XNOR2_X1 U7632 ( .A(n7613), .B(SI_4_), .ZN(n7610) );
  NAND2_X1 U7633 ( .A1(n7592), .A2(n7591), .ZN(n7612) );
  INV_X1 U7634 ( .A(n7587), .ZN(n7588) );
  AOI21_X1 U7635 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n10323), .A(n9411), .ZN(
        n9474) );
  NOR2_X1 U7636 ( .A1(n9422), .A2(n9423), .ZN(n9411) );
  NAND2_X1 U7637 ( .A1(n9784), .A2(n12278), .ZN(n12425) );
  NAND2_X1 U7638 ( .A1(n8928), .A2(n6538), .ZN(n11061) );
  AND2_X1 U7639 ( .A1(n12287), .A2(n12630), .ZN(n12103) );
  AND4_X1 U7640 ( .A1(n9286), .A2(n9285), .A3(n9284), .A4(n9283), .ZN(n12269)
         );
  NOR2_X1 U7641 ( .A1(n8818), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n8808) );
  NOR2_X1 U7642 ( .A1(n6779), .A2(n15022), .ZN(n6778) );
  INV_X1 U7643 ( .A(n6781), .ZN(n6779) );
  NAND2_X1 U7644 ( .A1(n15057), .A2(n6765), .ZN(n15074) );
  OR2_X1 U7645 ( .A1(n9910), .A2(n9911), .ZN(n6765) );
  INV_X1 U7646 ( .A(n7384), .ZN(n7383) );
  OAI21_X1 U7647 ( .B1(n7389), .B2(n7385), .A(n12109), .ZN(n7384) );
  NAND2_X1 U7648 ( .A1(n6865), .A2(n12277), .ZN(n6864) );
  NAND2_X1 U7649 ( .A1(n6867), .A2(n12651), .ZN(n6865) );
  INV_X1 U7650 ( .A(n12425), .ZN(n12640) );
  AND2_X1 U7651 ( .A1(n12858), .A2(n12265), .ZN(n9783) );
  OR2_X1 U7652 ( .A1(n11779), .A2(n11776), .ZN(n9781) );
  INV_X1 U7653 ( .A(n12082), .ZN(n12098) );
  INV_X1 U7654 ( .A(n12236), .ZN(n6721) );
  INV_X1 U7655 ( .A(n12105), .ZN(n12614) );
  OAI22_X1 U7656 ( .A1(n12081), .A2(n12080), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n13679), .ZN(n12092) );
  OAI21_X1 U7657 ( .B1(n9711), .B2(n9710), .A(n9712), .ZN(n9719) );
  OAI21_X1 U7658 ( .B1(n9248), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7280), .ZN(
        n9263) );
  INV_X1 U7659 ( .A(n7254), .ZN(n7253) );
  OAI21_X1 U7660 ( .B1(n9110), .B2(n7255), .A(n9128), .ZN(n7254) );
  NAND2_X1 U7661 ( .A1(n11733), .A2(n6541), .ZN(n7106) );
  XNOR2_X1 U7662 ( .A(n13076), .B(n10851), .ZN(n10408) );
  XNOR2_X1 U7663 ( .A(n13543), .B(n13226), .ZN(n8203) );
  INV_X1 U7664 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7463) );
  OAI21_X1 U7665 ( .B1(n13677), .B2(n8169), .A(n8168), .ZN(n13229) );
  XNOR2_X1 U7666 ( .A(n13561), .B(n13284), .ZN(n13312) );
  AOI21_X1 U7667 ( .B1(n7242), .B2(n7241), .A(n6578), .ZN(n7240) );
  XNOR2_X1 U7668 ( .A(n13578), .B(n13347), .ZN(n13363) );
  AOI21_X1 U7669 ( .B1(n7181), .B2(n7180), .A(n6595), .ZN(n7179) );
  INV_X1 U7670 ( .A(n7185), .ZN(n7180) );
  OR2_X1 U7671 ( .A1(n11003), .A2(n14459), .ZN(n10980) );
  NOR2_X1 U7672 ( .A1(n10879), .A2(n7235), .ZN(n7234) );
  INV_X1 U7673 ( .A(n10791), .ZN(n7235) );
  OR2_X1 U7674 ( .A1(n14937), .A2(n13147), .ZN(n7233) );
  AND2_X1 U7675 ( .A1(n7175), .A2(n7178), .ZN(n7174) );
  INV_X1 U7676 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7797) );
  AND2_X1 U7677 ( .A1(n13792), .A2(n12331), .ZN(n13713) );
  AOI21_X1 U7678 ( .B1(n11586), .B2(n13854), .A(n6747), .ZN(n6746) );
  INV_X1 U7679 ( .A(n7328), .ZN(n6747) );
  NAND2_X1 U7680 ( .A1(n13851), .A2(n11586), .ZN(n13773) );
  NAND3_X1 U7681 ( .A1(n14057), .A2(n13700), .A3(n6962), .ZN(n9351) );
  NOR2_X1 U7682 ( .A1(n12382), .A2(n6963), .ZN(n6962) );
  INV_X1 U7683 ( .A(n6964), .ZN(n6963) );
  NAND2_X1 U7684 ( .A1(n8521), .A2(n8520), .ZN(n14182) );
  AOI21_X1 U7685 ( .B1(n7084), .B2(n14227), .A(n6577), .ZN(n7083) );
  AOI21_X1 U7686 ( .B1(n7147), .B2(n8441), .A(n7146), .ZN(n7145) );
  INV_X1 U7687 ( .A(n8454), .ZN(n7146) );
  NAND2_X1 U7688 ( .A1(n8631), .A2(n8630), .ZN(n12308) );
  AND2_X1 U7689 ( .A1(n8883), .A2(n8866), .ZN(n10780) );
  AND2_X1 U7690 ( .A1(n12666), .A2(n12665), .ZN(n12667) );
  AOI22_X1 U7691 ( .A1(n13297), .A2(n13298), .B1(n13555), .B2(n13285), .ZN(
        n13288) );
  NAND2_X1 U7692 ( .A1(n13252), .A2(n13526), .ZN(n6950) );
  NAND2_X1 U7693 ( .A1(n7030), .A2(n7027), .ZN(n7028) );
  INV_X1 U7694 ( .A(n7032), .ZN(n7031) );
  OR2_X1 U7695 ( .A1(n7622), .A2(n7620), .ZN(n7299) );
  NAND2_X1 U7696 ( .A1(n11848), .A2(n11846), .ZN(n7369) );
  NAND2_X1 U7697 ( .A1(n11850), .A2(n11853), .ZN(n6850) );
  NAND2_X1 U7698 ( .A1(n6709), .A2(n6706), .ZN(n12146) );
  INV_X1 U7699 ( .A(n7823), .ZN(n6657) );
  NOR2_X1 U7700 ( .A1(n11873), .A2(n7376), .ZN(n7371) );
  INV_X1 U7701 ( .A(n7377), .ZN(n7376) );
  OAI22_X1 U7702 ( .A1(n11873), .A2(n7375), .B1(n11952), .B2(n11872), .ZN(
        n7373) );
  NAND2_X1 U7703 ( .A1(n7379), .A2(n7377), .ZN(n7375) );
  NAND2_X1 U7704 ( .A1(n11893), .A2(n6560), .ZN(n6817) );
  OAI22_X1 U7705 ( .A1(n11930), .A2(n7364), .B1(n11931), .B2(n7365), .ZN(
        n11934) );
  AND2_X1 U7706 ( .A1(n11931), .A2(n7365), .ZN(n7364) );
  INV_X1 U7707 ( .A(n11929), .ZN(n7365) );
  AOI211_X1 U7708 ( .C1(n12249), .C2(n12720), .A(n12248), .B(n12247), .ZN(
        n12253) );
  NAND2_X1 U7709 ( .A1(n6847), .A2(n6841), .ZN(n6846) );
  NOR2_X1 U7710 ( .A1(n6822), .A2(n6624), .ZN(n6819) );
  NAND2_X1 U7711 ( .A1(n11943), .A2(n11945), .ZN(n6820) );
  OR2_X1 U7712 ( .A1(n6841), .A2(n6840), .ZN(n6839) );
  NAND2_X1 U7713 ( .A1(n11954), .A2(n11950), .ZN(n6840) );
  NAND2_X1 U7714 ( .A1(n11954), .A2(n6834), .ZN(n6838) );
  NOR2_X1 U7715 ( .A1(n7999), .A2(SI_21_), .ZN(n7998) );
  NOR2_X1 U7716 ( .A1(n12663), .A2(n9777), .ZN(n12259) );
  OAI21_X1 U7717 ( .B1(n8118), .B2(n6684), .A(n6683), .ZN(n6682) );
  NAND2_X1 U7718 ( .A1(n8152), .A2(n8153), .ZN(n6683) );
  INV_X1 U7719 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7481) );
  NOR2_X1 U7720 ( .A1(n8121), .A2(n7216), .ZN(n7215) );
  INV_X1 U7721 ( .A(n8109), .ZN(n7216) );
  AOI21_X1 U7722 ( .B1(n7932), .B2(n6957), .A(n6956), .ZN(n6955) );
  INV_X1 U7723 ( .A(n7953), .ZN(n6956) );
  NOR2_X1 U7724 ( .A1(n7954), .A2(n7930), .ZN(n6957) );
  NAND2_X1 U7725 ( .A1(n7226), .A2(SI_13_), .ZN(n7225) );
  INV_X1 U7726 ( .A(n7818), .ZN(n7226) );
  NAND2_X1 U7727 ( .A1(n7818), .A2(n10007), .ZN(n7224) );
  INV_X1 U7728 ( .A(n7763), .ZN(n6923) );
  AND2_X1 U7729 ( .A1(n7744), .A2(n6923), .ZN(n6921) );
  INV_X1 U7730 ( .A(SI_11_), .ZN(n7747) );
  INV_X1 U7731 ( .A(n7022), .ZN(n7021) );
  OAI21_X1 U7732 ( .B1(n6512), .B2(n7024), .A(n7023), .ZN(n7022) );
  INV_X1 U7733 ( .A(n9073), .ZN(n7023) );
  OAI21_X1 U7734 ( .B1(n12506), .B2(n7007), .A(n7004), .ZN(n9230) );
  INV_X1 U7735 ( .A(n7008), .ZN(n7007) );
  AOI21_X1 U7736 ( .B1(n7008), .B2(n7006), .A(n7005), .ZN(n7004) );
  INV_X1 U7737 ( .A(n9224), .ZN(n7005) );
  AOI21_X1 U7738 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n10089), .A(n14428), .ZN(
        n9851) );
  INV_X1 U7739 ( .A(n9925), .ZN(n6791) );
  NAND2_X1 U7740 ( .A1(n6787), .A2(n6528), .ZN(n6786) );
  INV_X1 U7741 ( .A(n14437), .ZN(n6789) );
  NOR2_X1 U7742 ( .A1(n9704), .A2(n7409), .ZN(n7408) );
  INV_X1 U7743 ( .A(n9701), .ZN(n7409) );
  NAND2_X1 U7744 ( .A1(n7407), .A2(n7410), .ZN(n7406) );
  OR2_X1 U7745 ( .A1(n12660), .A2(n9780), .ZN(n11775) );
  INV_X1 U7746 ( .A(n12110), .ZN(n12660) );
  OR2_X1 U7747 ( .A1(n12873), .A2(n12524), .ZN(n12110) );
  NAND2_X1 U7748 ( .A1(n7394), .A2(n7392), .ZN(n7390) );
  OR2_X1 U7749 ( .A1(n12597), .A2(n12993), .ZN(n12205) );
  INV_X1 U7750 ( .A(n9687), .ZN(n7425) );
  OR2_X1 U7751 ( .A1(n12603), .A2(n15158), .ZN(n12163) );
  NAND2_X1 U7752 ( .A1(n12603), .A2(n15158), .ZN(n12165) );
  NAND2_X1 U7753 ( .A1(n7436), .A2(n7435), .ZN(n12162) );
  INV_X1 U7754 ( .A(n12604), .ZN(n7436) );
  OR2_X1 U7755 ( .A1(n12605), .A2(n15147), .ZN(n12157) );
  NAND2_X1 U7756 ( .A1(n7421), .A2(n7423), .ZN(n7419) );
  NAND2_X1 U7757 ( .A1(n12649), .A2(n7422), .ZN(n7421) );
  NAND2_X1 U7758 ( .A1(n9708), .A2(n9707), .ZN(n7422) );
  NAND2_X1 U7759 ( .A1(n7423), .A2(n9707), .ZN(n7420) );
  OR2_X1 U7760 ( .A1(n12877), .A2(n12507), .ZN(n11773) );
  AND2_X1 U7761 ( .A1(n12109), .A2(n12108), .ZN(n12248) );
  NAND2_X1 U7762 ( .A1(n7012), .A2(n8825), .ZN(n7011) );
  INV_X1 U7763 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7012) );
  INV_X1 U7764 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8804) );
  OAI21_X1 U7765 ( .B1(n9226), .B2(n6872), .A(n6870), .ZN(n8788) );
  AOI21_X1 U7766 ( .B1(n6873), .B2(n6871), .A(n6642), .ZN(n6870) );
  INV_X1 U7767 ( .A(n6873), .ZN(n6872) );
  OR2_X1 U7768 ( .A1(n8788), .A2(n11441), .ZN(n7280) );
  INV_X1 U7769 ( .A(n6892), .ZN(n6891) );
  INV_X1 U7770 ( .A(n9145), .ZN(n6893) );
  NAND2_X1 U7771 ( .A1(n9059), .A2(n8767), .ZN(n8768) );
  NAND2_X1 U7772 ( .A1(n8768), .A2(n10243), .ZN(n7279) );
  INV_X1 U7773 ( .A(n13676), .ZN(n7499) );
  AOI21_X1 U7774 ( .B1(n7245), .B2(n6904), .A(n6588), .ZN(n6903) );
  INV_X1 U7775 ( .A(n13464), .ZN(n6904) );
  OR2_X1 U7776 ( .A1(n7167), .A2(n11264), .ZN(n7166) );
  NAND2_X1 U7777 ( .A1(n7227), .A2(n6536), .ZN(n6910) );
  INV_X1 U7778 ( .A(n6911), .ZN(n6905) );
  AND2_X1 U7779 ( .A1(n7165), .A2(n10733), .ZN(n7164) );
  NAND2_X1 U7780 ( .A1(n10144), .A2(n11235), .ZN(n10348) );
  NOR2_X1 U7781 ( .A1(n6565), .A2(n13312), .ZN(n7177) );
  INV_X1 U7782 ( .A(n11550), .ZN(n6755) );
  INV_X1 U7783 ( .A(n6530), .ZN(n7326) );
  AOI21_X1 U7784 ( .B1(n6732), .B2(n6731), .A(n6730), .ZN(n6729) );
  INV_X1 U7785 ( .A(n11496), .ZN(n6730) );
  INV_X1 U7786 ( .A(n6737), .ZN(n6731) );
  AND2_X1 U7787 ( .A1(n6691), .A2(n6690), .ZN(n11965) );
  AOI21_X1 U7788 ( .B1(n6842), .B2(n6835), .A(n6832), .ZN(n6690) );
  OAI21_X1 U7789 ( .B1(n6842), .B2(n6845), .A(n11951), .ZN(n6691) );
  OR2_X1 U7790 ( .A1(n11792), .A2(n11794), .ZN(n6856) );
  NAND2_X1 U7791 ( .A1(n6855), .A2(n11960), .ZN(n6854) );
  NAND2_X1 U7792 ( .A1(n6598), .A2(n7096), .ZN(n7094) );
  NAND2_X1 U7793 ( .A1(n14120), .A2(n8685), .ZN(n7095) );
  NOR2_X1 U7794 ( .A1(n8687), .A2(n7093), .ZN(n7092) );
  INV_X1 U7795 ( .A(n8685), .ZN(n7093) );
  OR2_X1 U7796 ( .A1(n14513), .A2(n14523), .ZN(n11871) );
  OR2_X1 U7797 ( .A1(n11352), .A2(n8441), .ZN(n7148) );
  OR2_X1 U7798 ( .A1(n6969), .A2(n11854), .ZN(n6968) );
  NAND2_X1 U7799 ( .A1(n14531), .A2(n6970), .ZN(n6969) );
  INV_X1 U7800 ( .A(n11141), .ZN(n7077) );
  OR2_X1 U7801 ( .A1(n14668), .A2(n11185), .ZN(n7078) );
  NOR2_X1 U7802 ( .A1(n8666), .A2(n7075), .ZN(n7074) );
  INV_X1 U7803 ( .A(n7078), .ZN(n7075) );
  NAND2_X1 U7804 ( .A1(n14302), .A2(n14106), .ZN(n10286) );
  INV_X1 U7805 ( .A(n14295), .ZN(n14123) );
  INV_X1 U7806 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U7807 ( .A1(n8059), .A2(n8058), .ZN(n8080) );
  INV_X1 U7808 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U7809 ( .A1(n7204), .A2(SI_24_), .ZN(n7203) );
  INV_X1 U7810 ( .A(n8042), .ZN(n7204) );
  NAND2_X1 U7811 ( .A1(n8019), .A2(n8018), .ZN(n8040) );
  NAND2_X1 U7812 ( .A1(n8003), .A2(n8002), .ZN(n8017) );
  NAND2_X1 U7813 ( .A1(n6955), .A2(n6954), .ZN(n7995) );
  AOI21_X1 U7814 ( .B1(n6938), .B2(n6941), .A(n6633), .ZN(n6936) );
  INV_X1 U7815 ( .A(n6925), .ZN(n6924) );
  OAI21_X1 U7816 ( .B1(n7744), .B2(n7722), .A(n7746), .ZN(n6925) );
  AOI21_X1 U7817 ( .B1(n7698), .B2(n7199), .A(n6586), .ZN(n7198) );
  NAND2_X1 U7818 ( .A1(n7570), .A2(n7569), .ZN(n7589) );
  NAND2_X1 U7819 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n9387), .ZN(n9388) );
  INV_X1 U7820 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9387) );
  AOI22_X1 U7821 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n9447), .B1(n9448), .B2(
        n9400), .ZN(n9402) );
  OR2_X1 U7822 ( .A1(n9447), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n9400) );
  OAI21_X1 U7823 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n13950), .A(n9405), .ZN(
        n9427) );
  OAI22_X1 U7824 ( .A1(n9474), .A2(n9413), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n9412), .ZN(n9478) );
  OR2_X1 U7825 ( .A1(n8931), .A2(n11151), .ZN(n11060) );
  NAND2_X1 U7826 ( .A1(n9230), .A2(n9229), .ZN(n9238) );
  AND2_X1 U7827 ( .A1(n11154), .A2(n11150), .ZN(n11151) );
  NAND2_X1 U7828 ( .A1(n14977), .A2(n14976), .ZN(n14975) );
  AND4_X1 U7829 ( .A1(n9257), .A2(n9256), .A3(n9255), .A4(n9254), .ZN(n12403)
         );
  INV_X1 U7830 ( .A(n12085), .ZN(n9731) );
  NAND4_X1 U7831 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n9675)
         );
  OR2_X1 U7832 ( .A1(n9723), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U7833 ( .A1(n7117), .A2(n7115), .ZN(n11073) );
  NAND2_X1 U7834 ( .A1(n9835), .A2(n7118), .ZN(n7117) );
  OR2_X1 U7835 ( .A1(n11124), .A2(n7116), .ZN(n7115) );
  OAI21_X1 U7836 ( .B1(n11048), .B2(n7126), .A(n7125), .ZN(n11089) );
  NAND2_X1 U7837 ( .A1(n7129), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7126) );
  INV_X1 U7838 ( .A(n11090), .ZN(n7129) );
  OR2_X1 U7839 ( .A1(n11048), .A2(n11259), .ZN(n7128) );
  XNOR2_X1 U7840 ( .A(n7113), .B(n9950), .ZN(n14999) );
  OR2_X1 U7841 ( .A1(n10910), .A2(n7114), .ZN(n7113) );
  NOR2_X1 U7842 ( .A1(n9900), .A2(n8997), .ZN(n7114) );
  NAND2_X1 U7843 ( .A1(n6782), .A2(n6649), .ZN(n6781) );
  INV_X1 U7844 ( .A(n14994), .ZN(n6782) );
  NAND2_X1 U7845 ( .A1(n10913), .A2(n6525), .ZN(n6780) );
  INV_X1 U7846 ( .A(n6783), .ZN(n6777) );
  OR2_X1 U7847 ( .A1(n15013), .A2(n7121), .ZN(n7120) );
  AND2_X1 U7848 ( .A1(n15021), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7121) );
  AOI21_X1 U7849 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n15054), .A(n15046), .ZN(
        n9845) );
  NOR2_X1 U7850 ( .A1(n15074), .A2(n15075), .ZN(n15073) );
  AND2_X1 U7851 ( .A1(n9921), .A2(n9920), .ZN(n14412) );
  OAI21_X1 U7852 ( .B1(n14401), .B2(n7131), .A(n7130), .ZN(n14428) );
  NAND2_X1 U7853 ( .A1(n7132), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7131) );
  NAND2_X1 U7854 ( .A1(n9850), .A2(n7132), .ZN(n7130) );
  INV_X1 U7855 ( .A(n14427), .ZN(n7132) );
  NAND2_X1 U7856 ( .A1(n9923), .A2(n6647), .ZN(n6787) );
  INV_X1 U7857 ( .A(n6786), .ZN(n6788) );
  NAND2_X1 U7858 ( .A1(n14414), .A2(n6647), .ZN(n6790) );
  OR2_X1 U7859 ( .A1(n14442), .A2(n14443), .ZN(n7124) );
  NAND2_X1 U7860 ( .A1(n7123), .A2(n7122), .ZN(n12610) );
  INV_X1 U7861 ( .A(n9858), .ZN(n7122) );
  NAND2_X1 U7862 ( .A1(n9252), .A2(n8843), .ZN(n9282) );
  NOR2_X1 U7863 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n9282), .ZN(n9281) );
  INV_X1 U7864 ( .A(n7398), .ZN(n7397) );
  NAND2_X1 U7865 ( .A1(n6597), .A2(n7394), .ZN(n7389) );
  NAND2_X1 U7866 ( .A1(n7392), .A2(n12758), .ZN(n7391) );
  OR2_X1 U7867 ( .A1(n12759), .A2(n7390), .ZN(n7382) );
  INV_X1 U7868 ( .A(n12139), .ZN(n9797) );
  AND2_X1 U7869 ( .A1(n12297), .A2(n9797), .ZN(n12286) );
  OAI21_X1 U7870 ( .B1(n6864), .B2(n6861), .A(n9784), .ZN(n6860) );
  NAND2_X1 U7871 ( .A1(n11772), .A2(n6574), .ZN(n6862) );
  INV_X1 U7872 ( .A(n12278), .ZN(n6861) );
  AOI21_X1 U7873 ( .B1(n11756), .B2(n7416), .A(n7412), .ZN(n7411) );
  NAND2_X1 U7874 ( .A1(n7413), .A2(n7459), .ZN(n7412) );
  OR2_X1 U7875 ( .A1(n9717), .A2(n9738), .ZN(n7459) );
  NAND2_X1 U7876 ( .A1(n7416), .A2(n7418), .ZN(n7413) );
  AND2_X1 U7877 ( .A1(n7417), .A2(n12425), .ZN(n7416) );
  NAND2_X1 U7878 ( .A1(n7419), .A2(n7420), .ZN(n7417) );
  INV_X1 U7879 ( .A(n7419), .ZN(n7418) );
  INV_X1 U7880 ( .A(n7420), .ZN(n7415) );
  INV_X1 U7881 ( .A(n9783), .ZN(n6868) );
  INV_X1 U7882 ( .A(n12248), .ZN(n12707) );
  OR2_X1 U7883 ( .A1(n12962), .A2(n12487), .ZN(n12729) );
  NAND2_X1 U7884 ( .A1(n12729), .A2(n12237), .ZN(n12747) );
  NAND2_X1 U7885 ( .A1(n12137), .A2(n12139), .ZN(n15185) );
  AND2_X1 U7886 ( .A1(n12292), .A2(n12286), .ZN(n10678) );
  OAI21_X1 U7887 ( .B1(n9719), .B2(n9718), .A(n9721), .ZN(n12081) );
  AND2_X1 U7888 ( .A1(n7432), .A2(n8834), .ZN(n7431) );
  INV_X1 U7889 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U7890 ( .A1(n7281), .A2(n8794), .ZN(n9711) );
  OR2_X1 U7891 ( .A1(n9277), .A2(n8793), .ZN(n7281) );
  XNOR2_X1 U7892 ( .A(n8816), .B(P3_IR_REG_25__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U7893 ( .A1(n9211), .A2(n8785), .ZN(n9226) );
  NAND2_X1 U7894 ( .A1(n9209), .A2(n9208), .ZN(n9211) );
  NOR2_X1 U7895 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8803) );
  NAND2_X1 U7896 ( .A1(n6888), .A2(n6887), .ZN(n9196) );
  AND2_X1 U7897 ( .A1(n8780), .A2(n8779), .ZN(n9177) );
  INV_X1 U7898 ( .A(n8778), .ZN(n7261) );
  AND2_X1 U7899 ( .A1(n8778), .A2(n8777), .ZN(n9162) );
  NAND2_X1 U7900 ( .A1(n9163), .A2(n9162), .ZN(n9165) );
  OAI21_X1 U7901 ( .B1(n7252), .B2(n6893), .A(n6891), .ZN(n9163) );
  NAND2_X1 U7902 ( .A1(n9111), .A2(n7253), .ZN(n7252) );
  INV_X1 U7903 ( .A(n8772), .ZN(n7255) );
  AND2_X1 U7904 ( .A1(n8772), .A2(n8771), .ZN(n9110) );
  NAND2_X1 U7905 ( .A1(n9095), .A2(n8770), .ZN(n9111) );
  NAND2_X1 U7906 ( .A1(n9111), .A2(n9110), .ZN(n9113) );
  OR2_X1 U7907 ( .A1(n6516), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U7908 ( .A1(n9093), .A2(n9092), .ZN(n9095) );
  INV_X1 U7909 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8801) );
  OAI21_X1 U7910 ( .B1(n8768), .B2(n10243), .A(n7279), .ZN(n9082) );
  AND2_X1 U7911 ( .A1(n6876), .A2(n7262), .ZN(n6875) );
  AOI21_X1 U7912 ( .B1(n7265), .B2(n7267), .A(n7263), .ZN(n7262) );
  NAND2_X1 U7913 ( .A1(n9057), .A2(n9056), .ZN(n9059) );
  AND2_X1 U7914 ( .A1(n8932), .A2(n8800), .ZN(n9060) );
  NAND2_X1 U7915 ( .A1(n9013), .A2(n8759), .ZN(n9027) );
  NAND2_X1 U7916 ( .A1(n9011), .A2(n9010), .ZN(n9013) );
  OR2_X1 U7917 ( .A1(n8981), .A2(n8980), .ZN(n8983) );
  NAND2_X1 U7918 ( .A1(n8884), .A2(n7427), .ZN(n8920) );
  NAND2_X1 U7919 ( .A1(n8737), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8876) );
  AND2_X1 U7920 ( .A1(n7097), .A2(n6794), .ZN(n6793) );
  NAND2_X1 U7921 ( .A1(n11004), .A2(n6795), .ZN(n6794) );
  NOR2_X1 U7922 ( .A1(n11420), .A2(n7098), .ZN(n7097) );
  AND2_X1 U7923 ( .A1(n8237), .A2(n10150), .ZN(n10335) );
  INV_X1 U7924 ( .A(n11235), .ZN(n8237) );
  XNOR2_X1 U7925 ( .A(n13229), .B(n13254), .ZN(n7193) );
  NOR2_X1 U7926 ( .A1(n13312), .A2(n8202), .ZN(n7194) );
  AND4_X1 U7927 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(n13284)
         );
  NAND2_X1 U7928 ( .A1(n8157), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7585) );
  INV_X1 U7929 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U7930 ( .A1(n14845), .A2(n14844), .ZN(n14843) );
  NAND2_X1 U7931 ( .A1(n13321), .A2(n6985), .ZN(n13231) );
  NOR2_X1 U7932 ( .A1(n6519), .A2(n13555), .ZN(n6985) );
  NAND2_X1 U7933 ( .A1(n13306), .A2(n13550), .ZN(n13289) );
  INV_X1 U7934 ( .A(n13363), .ZN(n6899) );
  OR2_X1 U7935 ( .A1(n13277), .A2(n7243), .ZN(n6900) );
  NAND2_X1 U7936 ( .A1(n13277), .A2(n13388), .ZN(n13393) );
  OR2_X1 U7937 ( .A1(n13602), .A2(n13271), .ZN(n13272) );
  NOR2_X1 U7938 ( .A1(n7186), .A2(n7188), .ZN(n7185) );
  INV_X1 U7939 ( .A(n7189), .ZN(n7186) );
  NAND2_X1 U7940 ( .A1(n6581), .A2(n7189), .ZN(n7184) );
  NAND2_X1 U7941 ( .A1(n13463), .A2(n7245), .ZN(n13452) );
  INV_X1 U7942 ( .A(n13618), .ZN(n13221) );
  NAND2_X1 U7943 ( .A1(n13465), .A2(n13464), .ZN(n13463) );
  AND2_X1 U7944 ( .A1(n13259), .A2(n13258), .ZN(n7452) );
  NOR2_X1 U7945 ( .A1(n11265), .A2(n7171), .ZN(n7170) );
  INV_X1 U7946 ( .A(n7438), .ZN(n7171) );
  AND2_X1 U7947 ( .A1(n11264), .A2(n8188), .ZN(n10991) );
  OR2_X1 U7948 ( .A1(n14473), .A2(n13146), .ZN(n7438) );
  NOR2_X1 U7949 ( .A1(n6912), .A2(n7229), .ZN(n6911) );
  INV_X1 U7950 ( .A(n10794), .ZN(n6912) );
  INV_X1 U7951 ( .A(n7230), .ZN(n7229) );
  NAND2_X1 U7952 ( .A1(n10790), .A2(n10794), .ZN(n10792) );
  NAND2_X1 U7953 ( .A1(n7728), .A2(n7727), .ZN(n10856) );
  XNOR2_X1 U7954 ( .A(n10856), .B(n14456), .ZN(n10794) );
  NAND2_X1 U7955 ( .A1(n10595), .A2(n10594), .ZN(n7237) );
  NOR2_X1 U7956 ( .A1(n7158), .A2(n7159), .ZN(n7155) );
  NAND2_X1 U7957 ( .A1(n6980), .A2(n6979), .ZN(n10504) );
  XNOR2_X1 U7958 ( .A(n10476), .B(n10491), .ZN(n10233) );
  NAND2_X1 U7959 ( .A1(n10229), .A2(n10233), .ZN(n10470) );
  AND2_X1 U7960 ( .A1(n8192), .A2(n10232), .ZN(n10438) );
  INV_X1 U7961 ( .A(n10348), .ZN(n10267) );
  NAND2_X1 U7962 ( .A1(n8099), .A2(n8098), .ZN(n13561) );
  NAND2_X1 U7963 ( .A1(n8083), .A2(n8082), .ZN(n13566) );
  NAND2_X1 U7964 ( .A1(n7974), .A2(n7973), .ZN(n13597) );
  INV_X1 U7965 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7497) );
  AND2_X1 U7966 ( .A1(n8225), .A2(n8224), .ZN(n8229) );
  INV_X1 U7967 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U7968 ( .A1(n7677), .A2(n7308), .ZN(n7882) );
  NOR2_X1 U7969 ( .A1(n7329), .A2(n6580), .ZN(n7328) );
  NOR2_X1 U7970 ( .A1(n13774), .A2(n13781), .ZN(n7329) );
  AND2_X1 U7971 ( .A1(n7321), .A2(n13693), .ZN(n7320) );
  OR2_X1 U7972 ( .A1(n13843), .A2(n12359), .ZN(n7321) );
  NAND2_X1 U7973 ( .A1(n11327), .A2(n6737), .ZN(n6735) );
  AND2_X1 U7974 ( .A1(n13762), .A2(n7312), .ZN(n7311) );
  NAND2_X1 U7975 ( .A1(n7314), .A2(n7317), .ZN(n7312) );
  AND2_X1 U7976 ( .A1(n13761), .A2(n12340), .ZN(n13793) );
  NAND2_X1 U7977 ( .A1(n11648), .A2(n11647), .ZN(n12322) );
  INV_X1 U7978 ( .A(n7334), .ZN(n7333) );
  AOI21_X1 U7979 ( .B1(n7334), .B2(n7332), .A(n7331), .ZN(n7330) );
  NOR2_X1 U7980 ( .A1(n11198), .A2(n11203), .ZN(n7338) );
  AND2_X1 U7981 ( .A1(n11580), .A2(n11579), .ZN(n11586) );
  NAND2_X1 U7982 ( .A1(n6751), .A2(n6750), .ZN(n11580) );
  NOR2_X1 U7983 ( .A1(n11576), .A2(n6753), .ZN(n6750) );
  CLKBUF_X1 U7984 ( .A(n8290), .Z(n8574) );
  NAND2_X1 U7985 ( .A1(n8613), .A2(n8612), .ZN(n14046) );
  XNOR2_X1 U7986 ( .A(n14046), .B(n13871), .ZN(n14043) );
  NAND2_X1 U7987 ( .A1(n8511), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U7988 ( .A1(n14224), .A2(n7084), .ZN(n7080) );
  AOI21_X1 U7989 ( .B1(n7083), .B2(n7085), .A(n14186), .ZN(n7081) );
  INV_X1 U7990 ( .A(n7083), .ZN(n7082) );
  INV_X1 U7991 ( .A(n14224), .ZN(n7087) );
  NAND2_X1 U7992 ( .A1(n8432), .A2(n8431), .ZN(n11857) );
  NOR2_X1 U7993 ( .A1(n6968), .A2(n11190), .ZN(n11380) );
  NAND2_X1 U7994 ( .A1(n11974), .A2(n11973), .ZN(n14019) );
  NAND2_X1 U7995 ( .A1(n11956), .A2(n11955), .ZN(n11985) );
  NAND2_X1 U7996 ( .A1(n8590), .A2(n8589), .ZN(n14087) );
  NAND2_X1 U7997 ( .A1(n11976), .A2(n8651), .ZN(n14522) );
  INV_X1 U7998 ( .A(n14676), .ZN(n14661) );
  AND2_X1 U7999 ( .A1(n10274), .A2(n10290), .ZN(n10295) );
  AND2_X1 U8000 ( .A1(n8710), .A2(n8709), .ZN(n10281) );
  NAND2_X1 U8001 ( .A1(n8145), .A2(n8144), .ZN(n8127) );
  OR2_X1 U8002 ( .A1(n8164), .A2(n8163), .ZN(n8166) );
  INV_X1 U8003 ( .A(n8265), .ZN(n7061) );
  NOR2_X1 U8004 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n7060) );
  OAI21_X1 U8005 ( .B1(n6852), .B2(n7345), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8639) );
  NAND2_X1 U8006 ( .A1(n6937), .A2(n7217), .ZN(n7881) );
  NAND2_X1 U8007 ( .A1(n7819), .A2(n7220), .ZN(n6937) );
  AND2_X1 U8008 ( .A1(n8470), .A2(n8460), .ZN(n10385) );
  OR2_X1 U8009 ( .A1(n8374), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8386) );
  OR2_X1 U8010 ( .A1(n8359), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8374) );
  INV_X1 U8011 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6811) );
  XNOR2_X1 U8012 ( .A(n9434), .B(n9435), .ZN(n9437) );
  NOR2_X1 U8013 ( .A1(n15206), .A2(n9441), .ZN(n9445) );
  NAND2_X1 U8014 ( .A1(n7056), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8015 ( .A1(n7044), .A2(n7046), .ZN(n7043) );
  INV_X1 U8016 ( .A(n7047), .ZN(n7044) );
  AOI21_X1 U8017 ( .B1(n7050), .B2(n7048), .A(P2_ADDR_REG_16__SCAN_IN), .ZN(
        n7047) );
  INV_X1 U8018 ( .A(n7055), .ZN(n7048) );
  AOI21_X1 U8019 ( .B1(n6999), .B2(n7001), .A(n6628), .ZN(n6997) );
  OR2_X1 U8020 ( .A1(n12608), .A2(n10685), .ZN(n15116) );
  NOR2_X1 U8021 ( .A1(n7003), .A2(n11172), .ZN(n7002) );
  INV_X1 U8022 ( .A(n8951), .ZN(n7003) );
  OAI21_X1 U8023 ( .B1(n6883), .B2(n6884), .A(n12298), .ZN(n6711) );
  NAND2_X1 U8024 ( .A1(n12290), .A2(n6885), .ZN(n6884) );
  OAI21_X1 U8025 ( .B1(n6700), .B2(n6699), .A(n6698), .ZN(n12291) );
  INV_X1 U8026 ( .A(n15122), .ZN(n6699) );
  NAND2_X1 U8027 ( .A1(n6700), .A2(n12292), .ZN(n6698) );
  OR2_X1 U8028 ( .A1(n12289), .A2(n12288), .ZN(n6700) );
  NOR4_X1 U8029 ( .A1(n12287), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12131) );
  OR2_X1 U8030 ( .A1(n8892), .A2(n9863), .ZN(n8893) );
  OR2_X1 U8031 ( .A1(n8892), .A2(n11107), .ZN(n8853) );
  XNOR2_X1 U8032 ( .A(n8955), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11100) );
  XNOR2_X1 U8033 ( .A(n7120), .B(n15036), .ZN(n15031) );
  NOR2_X1 U8034 ( .A1(n15064), .A2(n9076), .ZN(n15063) );
  AOI21_X1 U8035 ( .B1(n12628), .B2(n15094), .A(n12627), .ZN(n6769) );
  XNOR2_X1 U8036 ( .A(n12624), .B(n12623), .ZN(n6770) );
  NAND2_X1 U8037 ( .A1(n12610), .A2(n6696), .ZN(n6695) );
  OR2_X1 U8038 ( .A1(n12617), .A2(n12751), .ZN(n6696) );
  OR2_X1 U8039 ( .A1(n9814), .A2(n12802), .ZN(n9802) );
  NAND2_X1 U8040 ( .A1(n9279), .A2(n9278), .ZN(n12559) );
  OR2_X1 U8041 ( .A1(n9714), .A2(n11349), .ZN(n9278) );
  NAND2_X1 U8042 ( .A1(n11783), .A2(n6672), .ZN(n12859) );
  NAND2_X1 U8043 ( .A1(n6522), .A2(n12804), .ZN(n6672) );
  NAND2_X1 U8044 ( .A1(n9265), .A2(n9264), .ZN(n12858) );
  OR2_X1 U8045 ( .A1(n9714), .A2(n11281), .ZN(n9264) );
  NAND2_X1 U8046 ( .A1(n6662), .A2(n6660), .ZN(n12863) );
  INV_X1 U8047 ( .A(n6661), .ZN(n6660) );
  NAND2_X1 U8048 ( .A1(n12864), .A2(n15175), .ZN(n6662) );
  OAI21_X1 U8049 ( .B1(n12672), .B2(n15117), .A(n12671), .ZN(n6661) );
  NAND2_X1 U8050 ( .A1(n9702), .A2(n9701), .ZN(n12684) );
  NAND2_X1 U8051 ( .A1(n9242), .A2(n9241), .ZN(n12691) );
  OR2_X1 U8052 ( .A1(n9714), .A2(n10847), .ZN(n9241) );
  AND3_X1 U8053 ( .A1(n8995), .A2(n8994), .A3(n8993), .ZN(n15170) );
  AND2_X1 U8054 ( .A1(n12614), .A2(n10579), .ZN(n15122) );
  AOI21_X1 U8055 ( .B1(n13008), .B2(n12098), .A(n12097), .ZN(n12914) );
  NOR2_X1 U8056 ( .A1(n12931), .A2(n12998), .ZN(n6714) );
  OR2_X1 U8057 ( .A1(n9714), .A2(n11137), .ZN(n9249) );
  NAND2_X1 U8058 ( .A1(n9184), .A2(n9183), .ZN(n12956) );
  NAND2_X1 U8059 ( .A1(n9135), .A2(n9134), .ZN(n12974) );
  NOR2_X1 U8060 ( .A1(n15191), .A2(n15185), .ZN(n12985) );
  INV_X1 U8061 ( .A(n13561), .ZN(n13319) );
  NAND2_X1 U8062 ( .A1(n7105), .A2(n7103), .ZN(n13010) );
  AND2_X1 U8063 ( .A1(n13011), .A2(n7104), .ZN(n7103) );
  NAND2_X1 U8064 ( .A1(n7106), .A2(n7107), .ZN(n7104) );
  AND2_X1 U8065 ( .A1(n11719), .A2(n11713), .ZN(n7111) );
  NAND2_X1 U8066 ( .A1(n13093), .A2(n11713), .ZN(n13027) );
  NAND2_X1 U8067 ( .A1(n7772), .A2(n7771), .ZN(n11003) );
  NAND2_X1 U8068 ( .A1(n13070), .A2(n10405), .ZN(n10406) );
  NAND2_X1 U8069 ( .A1(n6546), .A2(n11698), .ZN(n6804) );
  AND2_X1 U8070 ( .A1(n11698), .A2(n10848), .ZN(n6805) );
  NAND2_X1 U8071 ( .A1(n7754), .A2(n7753), .ZN(n14937) );
  NAND2_X1 U8072 ( .A1(n10374), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14470) );
  NAND2_X1 U8073 ( .A1(n7917), .A2(n7916), .ZN(n13612) );
  INV_X2 U8074 ( .A(n13126), .ZN(n14462) );
  OAI21_X1 U8075 ( .B1(n13366), .B2(n8139), .A(n8037), .ZN(n13347) );
  NOR2_X1 U8076 ( .A1(n14741), .A2(n14740), .ZN(n14739) );
  NAND2_X1 U8077 ( .A1(n8134), .A2(n8133), .ZN(n13543) );
  OAI21_X1 U8078 ( .B1(n13554), .B2(n14942), .A(n6946), .ZN(n6943) );
  AND2_X1 U8079 ( .A1(n6947), .A2(n6639), .ZN(n6946) );
  OR2_X1 U8080 ( .A1(n6625), .A2(n6948), .ZN(n6947) );
  OAI21_X1 U8081 ( .B1(n13329), .B2(n6763), .A(n6762), .ZN(n13251) );
  INV_X1 U8082 ( .A(n7174), .ZN(n6763) );
  AND2_X1 U8083 ( .A1(n6959), .A2(n13250), .ZN(n6762) );
  AOI21_X1 U8084 ( .B1(n11327), .B2(n11326), .A(n7341), .ZN(n11401) );
  NOR2_X1 U8085 ( .A1(n10939), .A2(n10940), .ZN(n11195) );
  INV_X1 U8086 ( .A(n11857), .ZN(n14531) );
  OR2_X1 U8087 ( .A1(n12018), .A2(n7140), .ZN(n7139) );
  OAI21_X1 U8088 ( .B1(n12018), .B2(n7138), .A(n7137), .ZN(n7136) );
  AND2_X1 U8089 ( .A1(n13869), .A2(n14498), .ZN(n8695) );
  NOR2_X1 U8090 ( .A1(n9376), .A2(n9375), .ZN(n14039) );
  NAND2_X1 U8091 ( .A1(n6667), .A2(n6665), .ZN(n9376) );
  NAND2_X1 U8092 ( .A1(n9372), .A2(n6666), .ZN(n6665) );
  NAND2_X2 U8093 ( .A1(n8289), .A2(n8288), .ZN(n14652) );
  NAND2_X1 U8094 ( .A1(n8313), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8318) );
  NOR2_X1 U8095 ( .A1(n7066), .A2(n14644), .ZN(n7065) );
  INV_X1 U8096 ( .A(n12303), .ZN(n7066) );
  NAND2_X1 U8097 ( .A1(n14687), .A2(n14669), .ZN(n14348) );
  XNOR2_X1 U8098 ( .A(n9437), .B(n7038), .ZN(n15221) );
  NOR2_X1 U8099 ( .A1(n14384), .A2(n6518), .ZN(n7033) );
  NOR2_X1 U8100 ( .A1(n7051), .A2(n14571), .ZN(n7050) );
  NAND2_X1 U8101 ( .A1(n14567), .A2(n7055), .ZN(n7052) );
  INV_X1 U8102 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7054) );
  OAI21_X1 U8103 ( .B1(n14371), .B2(n14372), .A(n7037), .ZN(n7036) );
  INV_X1 U8104 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7037) );
  OR2_X1 U8105 ( .A1(n7302), .A2(n7621), .ZN(n7300) );
  OR2_X1 U8106 ( .A1(n7664), .A2(n7662), .ZN(n7296) );
  AND2_X1 U8107 ( .A1(n11816), .A2(n11815), .ZN(n11820) );
  NAND2_X1 U8108 ( .A1(n7706), .A2(n7708), .ZN(n7284) );
  NAND2_X1 U8109 ( .A1(n7755), .A2(n7757), .ZN(n7287) );
  INV_X1 U8110 ( .A(n11838), .ZN(n7353) );
  INV_X1 U8111 ( .A(n11837), .ZN(n7348) );
  NAND2_X1 U8112 ( .A1(n7356), .A2(n11837), .ZN(n7355) );
  NAND2_X1 U8113 ( .A1(n6708), .A2(n6707), .ZN(n6706) );
  NOR2_X1 U8114 ( .A1(n12136), .A2(n12137), .ZN(n6708) );
  INV_X1 U8115 ( .A(n10775), .ZN(n6707) );
  NAND2_X1 U8116 ( .A1(n6849), .A2(n6848), .ZN(n11860) );
  AOI21_X1 U8117 ( .B1(n6517), .B2(n6851), .A(n6593), .ZN(n6848) );
  NOR2_X1 U8118 ( .A1(n11853), .A2(n11850), .ZN(n6851) );
  AND2_X1 U8119 ( .A1(n7920), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U8120 ( .A1(n7378), .A2(n11867), .ZN(n7377) );
  NOR2_X1 U8121 ( .A1(n7378), .A2(n11867), .ZN(n7379) );
  NOR4_X1 U8122 ( .A1(n12189), .A2(n12188), .A3(n12192), .A4(n12187), .ZN(
        n12199) );
  NAND2_X1 U8123 ( .A1(n7958), .A2(n7960), .ZN(n7293) );
  INV_X1 U8124 ( .A(n7373), .ZN(n7372) );
  AND2_X1 U8125 ( .A1(n11893), .A2(n11883), .ZN(n6818) );
  NAND2_X1 U8126 ( .A1(n6813), .A2(n6815), .ZN(n6812) );
  AND2_X1 U8127 ( .A1(n6814), .A2(n11916), .ZN(n6813) );
  NAND2_X1 U8128 ( .A1(n8006), .A2(n8008), .ZN(n7295) );
  AND2_X1 U8129 ( .A1(n11925), .A2(n7360), .ZN(n7359) );
  INV_X1 U8130 ( .A(n11923), .ZN(n7360) );
  OAI211_X1 U8131 ( .C1(n11924), .C2(n6830), .A(n6826), .B(n11927), .ZN(n6825)
         );
  NAND2_X1 U8132 ( .A1(n6829), .A2(n6828), .ZN(n6826) );
  INV_X1 U8133 ( .A(n6830), .ZN(n6829) );
  OAI21_X1 U8134 ( .B1(n11924), .B2(n7359), .A(n6827), .ZN(n6824) );
  NOR2_X1 U8135 ( .A1(n11928), .A2(n6828), .ZN(n6827) );
  NAND2_X1 U8136 ( .A1(n8045), .A2(n8047), .ZN(n7294) );
  NAND2_X1 U8137 ( .A1(n6705), .A2(n7407), .ZN(n6704) );
  INV_X1 U8138 ( .A(n12255), .ZN(n6705) );
  INV_X1 U8139 ( .A(n11940), .ZN(n7361) );
  AND2_X1 U8140 ( .A1(n11944), .A2(n6823), .ZN(n6822) );
  NAND2_X1 U8141 ( .A1(n6702), .A2(n6701), .ZN(n12264) );
  AND2_X1 U8142 ( .A1(n12261), .A2(n12669), .ZN(n6701) );
  OAI22_X1 U8143 ( .A1(n12254), .A2(n6704), .B1(n12939), .B2(n6703), .ZN(n6702) );
  NAND2_X1 U8144 ( .A1(n12526), .A2(n12286), .ZN(n6703) );
  NAND2_X1 U8145 ( .A1(n8084), .A2(n7305), .ZN(n7304) );
  AND2_X1 U8146 ( .A1(n10148), .A2(n8208), .ZN(n7807) );
  NAND2_X1 U8147 ( .A1(n6846), .A2(n6834), .ZN(n6833) );
  AND2_X1 U8148 ( .A1(n8078), .A2(SI_26_), .ZN(n6933) );
  INV_X1 U8149 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7505) );
  INV_X1 U8150 ( .A(n12505), .ZN(n7006) );
  AOI21_X1 U8151 ( .B1(n9225), .B2(n8786), .A(n6874), .ZN(n6873) );
  INV_X1 U8152 ( .A(n9239), .ZN(n6874) );
  INV_X1 U8153 ( .A(n8786), .ZN(n6871) );
  INV_X1 U8154 ( .A(n13268), .ZN(n7244) );
  NOR2_X1 U8155 ( .A1(n13578), .A2(n13383), .ZN(n6976) );
  NAND2_X1 U8156 ( .A1(n11946), .A2(n11949), .ZN(n7367) );
  NOR2_X1 U8157 ( .A1(n11949), .A2(n11946), .ZN(n7366) );
  NAND2_X1 U8158 ( .A1(n6821), .A2(n6820), .ZN(n11947) );
  NAND2_X1 U8159 ( .A1(n6836), .A2(n6569), .ZN(n6842) );
  OR2_X1 U8160 ( .A1(n6844), .A2(n6843), .ZN(n6836) );
  INV_X1 U8161 ( .A(n11793), .ZN(n6855) );
  AOI21_X1 U8162 ( .B1(n8079), .B2(n6933), .A(n6932), .ZN(n6931) );
  INV_X1 U8163 ( .A(n8093), .ZN(n6932) );
  AOI21_X1 U8164 ( .B1(n8079), .B2(n8078), .A(SI_26_), .ZN(n6934) );
  INV_X1 U8165 ( .A(n8078), .ZN(n6930) );
  NAND2_X1 U8166 ( .A1(n6931), .A2(n6928), .ZN(n6927) );
  INV_X1 U8167 ( .A(n6933), .ZN(n6928) );
  AND2_X1 U8168 ( .A1(n7210), .A2(n8016), .ZN(n7205) );
  NAND2_X1 U8169 ( .A1(n6954), .A2(n6688), .ZN(n8003) );
  AND2_X1 U8170 ( .A1(n6955), .A2(n6636), .ZN(n6688) );
  NAND2_X1 U8171 ( .A1(n7933), .A2(n10330), .ZN(n7953) );
  INV_X1 U8172 ( .A(n7909), .ZN(n7910) );
  INV_X1 U8173 ( .A(n7225), .ZN(n7222) );
  NOR2_X1 U8174 ( .A1(n7697), .A2(n7672), .ZN(n7197) );
  INV_X1 U8175 ( .A(n7676), .ZN(n7199) );
  AND2_X1 U8176 ( .A1(n6611), .A2(n9004), .ZN(n7024) );
  NAND2_X1 U8177 ( .A1(n7278), .A2(n12285), .ZN(n7275) );
  NOR2_X1 U8178 ( .A1(n12288), .A2(n6551), .ZN(n12107) );
  NAND2_X1 U8179 ( .A1(n8884), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9831) );
  OR2_X1 U8180 ( .A1(n11074), .A2(n10957), .ZN(n7116) );
  INV_X1 U8181 ( .A(n11074), .ZN(n7118) );
  NAND2_X1 U8182 ( .A1(n11076), .A2(n6557), .ZN(n9869) );
  OAI21_X1 U8183 ( .B1(n9900), .B2(n8996), .A(n10917), .ZN(n9873) );
  NAND2_X1 U8184 ( .A1(n9905), .A2(n9986), .ZN(n6783) );
  OAI21_X1 U8185 ( .B1(n9986), .B2(n9030), .A(n15016), .ZN(n9875) );
  OAI21_X1 U8186 ( .B1(n9911), .B2(n9861), .A(n15049), .ZN(n9877) );
  NAND2_X1 U8187 ( .A1(n15084), .A2(n9916), .ZN(n9879) );
  NAND2_X1 U8188 ( .A1(n14422), .A2(n6720), .ZN(n9881) );
  OR2_X1 U8189 ( .A1(n14418), .A2(n12892), .ZN(n6720) );
  INV_X1 U8190 ( .A(n7405), .ZN(n7399) );
  AND2_X1 U8191 ( .A1(n7407), .A2(n12680), .ZN(n12661) );
  INV_X1 U8192 ( .A(n12108), .ZN(n7385) );
  NAND2_X1 U8193 ( .A1(n7388), .A2(n12108), .ZN(n7387) );
  INV_X1 U8194 ( .A(n7390), .ZN(n7388) );
  AND2_X1 U8195 ( .A1(n12747), .A2(n12719), .ZN(n7395) );
  OR2_X1 U8196 ( .A1(n12601), .A2(n15170), .ZN(n12184) );
  INV_X1 U8197 ( .A(n12112), .ZN(n12160) );
  NAND2_X1 U8198 ( .A1(n12152), .A2(n12151), .ZN(n12115) );
  AND2_X1 U8199 ( .A1(n9815), .A2(n9728), .ZN(n12099) );
  INV_X1 U8200 ( .A(n12588), .ZN(n12507) );
  OR2_X1 U8201 ( .A1(n12595), .A2(n12389), .ZN(n12214) );
  AND2_X1 U8202 ( .A1(n6775), .A2(n8804), .ZN(n6772) );
  NAND2_X1 U8203 ( .A1(n7015), .A2(n7014), .ZN(n7013) );
  INV_X1 U8204 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7015) );
  INV_X1 U8205 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U8206 ( .A1(n7430), .A2(n6775), .ZN(n6774) );
  NOR2_X1 U8207 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8802) );
  AOI21_X1 U8208 ( .B1(n7259), .B2(n7261), .A(n7257), .ZN(n7256) );
  INV_X1 U8209 ( .A(n8780), .ZN(n7257) );
  NAND2_X1 U8210 ( .A1(n8781), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8783) );
  INV_X1 U8211 ( .A(n7266), .ZN(n7265) );
  OAI21_X1 U8212 ( .B1(n8761), .B2(n7267), .A(n8764), .ZN(n7266) );
  INV_X1 U8213 ( .A(n8762), .ZN(n7267) );
  INV_X1 U8214 ( .A(n8765), .ZN(n7263) );
  AND2_X1 U8215 ( .A1(n7265), .A2(n6879), .ZN(n6878) );
  NAND2_X1 U8216 ( .A1(n6880), .A2(n8759), .ZN(n6879) );
  INV_X1 U8217 ( .A(n9010), .ZN(n6880) );
  NAND2_X1 U8218 ( .A1(n6878), .A2(n6881), .ZN(n6876) );
  INV_X1 U8219 ( .A(n8759), .ZN(n6881) );
  OR2_X1 U8220 ( .A1(n8991), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9005) );
  AND2_X1 U8221 ( .A1(n6995), .A2(n6994), .ZN(n7427) );
  INV_X1 U8222 ( .A(n11416), .ZN(n7098) );
  INV_X1 U8223 ( .A(n10998), .ZN(n6795) );
  NOR2_X1 U8224 ( .A1(n7691), .A2(n7690), .ZN(n7710) );
  NOR2_X1 U8225 ( .A1(n13572), .A2(n6975), .ZN(n6974) );
  INV_X1 U8226 ( .A(n6976), .ZN(n6975) );
  NOR2_X1 U8227 ( .A1(n7827), .A2(n7826), .ZN(n7847) );
  NOR2_X1 U8228 ( .A1(n7758), .A2(n10999), .ZN(n7782) );
  NOR2_X1 U8229 ( .A1(n10883), .A2(n11003), .ZN(n6982) );
  NAND2_X1 U8230 ( .A1(n14904), .A2(n10543), .ZN(n10604) );
  OR2_X1 U8231 ( .A1(n14904), .A2(n10543), .ZN(n7160) );
  INV_X1 U8232 ( .A(n10507), .ZN(n7159) );
  INV_X1 U8233 ( .A(n10479), .ZN(n10481) );
  AND2_X1 U8234 ( .A1(n7160), .A2(n10604), .ZN(n10479) );
  NAND2_X1 U8235 ( .A1(n13396), .A2(n13585), .ZN(n13382) );
  NOR2_X1 U8236 ( .A1(n8217), .A2(n8216), .ZN(n8225) );
  NAND2_X1 U8237 ( .A1(n7110), .A2(n7488), .ZN(n8217) );
  INV_X1 U8238 ( .A(n13793), .ZN(n7317) );
  AOI21_X1 U8239 ( .B1(n13793), .B2(n7316), .A(n7315), .ZN(n7314) );
  NAND2_X1 U8240 ( .A1(n11960), .A2(n11120), .ZN(n10273) );
  INV_X1 U8241 ( .A(n13801), .ZN(n7332) );
  INV_X1 U8242 ( .A(n11585), .ZN(n12364) );
  INV_X1 U8243 ( .A(n10273), .ZN(n11977) );
  NAND2_X1 U8244 ( .A1(n12382), .A2(n13869), .ZN(n7143) );
  AND2_X1 U8245 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n8614), .ZN(n8272) );
  NOR2_X1 U8246 ( .A1(n12016), .A2(n7142), .ZN(n7141) );
  INV_X1 U8247 ( .A(n8629), .ZN(n7142) );
  NOR2_X1 U8248 ( .A1(n14046), .A2(n14058), .ZN(n6964) );
  NOR2_X1 U8249 ( .A1(n14160), .A2(n14170), .ZN(n6961) );
  AND2_X1 U8250 ( .A1(n8453), .A2(n8440), .ZN(n7147) );
  NAND2_X1 U8251 ( .A1(n10464), .A2(n10714), .ZN(n11818) );
  NAND2_X1 U8252 ( .A1(n14249), .A2(n14240), .ZN(n11796) );
  NAND2_X1 U8253 ( .A1(n14057), .A2(n8653), .ZN(n14045) );
  NAND2_X1 U8254 ( .A1(n14116), .A2(n8685), .ZN(n14096) );
  NOR2_X1 U8255 ( .A1(n14137), .A2(n14123), .ZN(n14122) );
  NAND2_X1 U8256 ( .A1(n7214), .A2(n7212), .ZN(n8145) );
  AOI21_X1 U8257 ( .B1(n7215), .B2(n8110), .A(n7213), .ZN(n7212) );
  INV_X1 U8258 ( .A(n8123), .ZN(n7213) );
  INV_X1 U8259 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8257) );
  OR2_X1 U8260 ( .A1(n8002), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U8261 ( .A1(n8003), .A2(n7209), .ZN(n7208) );
  AND2_X1 U8262 ( .A1(n8002), .A2(n7211), .ZN(n7209) );
  INV_X1 U8263 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U8264 ( .A1(n8643), .A2(n7342), .ZN(n8713) );
  AND2_X1 U8265 ( .A1(n8532), .A2(n6757), .ZN(n6756) );
  INV_X1 U8266 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6757) );
  AOI21_X1 U8267 ( .B1(n7220), .B2(n7223), .A(n7218), .ZN(n7217) );
  INV_X1 U8268 ( .A(n7224), .ZN(n7223) );
  INV_X1 U8269 ( .A(n7863), .ZN(n7218) );
  NAND2_X1 U8270 ( .A1(n7819), .A2(n7225), .ZN(n7219) );
  AOI21_X1 U8271 ( .B1(n6924), .B2(n6921), .A(n6920), .ZN(n6919) );
  NAND2_X1 U8272 ( .A1(n6924), .A2(n6923), .ZN(n6922) );
  INV_X1 U8273 ( .A(n7614), .ZN(n7195) );
  INV_X1 U8274 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9430) );
  AOI21_X1 U8275 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n9407), .A(n9406), .ZN(
        n9424) );
  OAI21_X1 U8276 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n13986), .A(n9410), .ZN(
        n9422) );
  NAND2_X1 U8277 ( .A1(n8900), .A2(n8899), .ZN(n12409) );
  AND2_X1 U8278 ( .A1(n12546), .A2(n7000), .ZN(n6999) );
  OR2_X1 U8279 ( .A1(n12484), .A2(n7001), .ZN(n7000) );
  INV_X1 U8280 ( .A(n9161), .ZN(n7001) );
  AND2_X1 U8281 ( .A1(n8861), .A2(n8860), .ZN(n7026) );
  OR2_X1 U8282 ( .A1(n12082), .A2(n9947), .ZN(n7025) );
  AND2_X1 U8283 ( .A1(n7009), .A2(n9207), .ZN(n7008) );
  INV_X1 U8284 ( .A(n12442), .ZN(n7009) );
  NAND2_X1 U8285 ( .A1(n12506), .A2(n12505), .ZN(n7010) );
  AOI21_X1 U8286 ( .B1(n14975), .B2(n7024), .A(n6512), .ZN(n12452) );
  INV_X1 U8287 ( .A(n9267), .ZN(n9252) );
  INV_X1 U8288 ( .A(n12138), .ZN(n10777) );
  AOI21_X1 U8289 ( .B1(n7021), .B2(n6512), .A(n6591), .ZN(n7020) );
  INV_X1 U8290 ( .A(n12550), .ZN(n12573) );
  AND2_X1 U8291 ( .A1(n11454), .A2(n12286), .ZN(n12572) );
  INV_X1 U8292 ( .A(n12134), .ZN(n6885) );
  AOI21_X1 U8293 ( .B1(n7276), .B2(n7274), .A(n12287), .ZN(n12289) );
  AOI21_X1 U8294 ( .B1(n7278), .B2(n7277), .A(n6551), .ZN(n7276) );
  NAND2_X1 U8295 ( .A1(n7275), .A2(n12286), .ZN(n7274) );
  NOR2_X1 U8296 ( .A1(n12076), .A2(n12286), .ZN(n7277) );
  AND2_X1 U8297 ( .A1(n12914), .A2(n12633), .ZN(n12288) );
  AND4_X1 U8298 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n12427)
         );
  AND4_X1 U8299 ( .A1(n9204), .A2(n9203), .A3(n9202), .A4(n9201), .ZN(n12443)
         );
  AND4_X1 U8300 ( .A1(n9190), .A2(n9189), .A3(n9188), .A4(n9187), .ZN(n12551)
         );
  AND4_X1 U8301 ( .A1(n9175), .A2(n9174), .A3(n9173), .A4(n9172), .ZN(n12487)
         );
  AND4_X1 U8302 ( .A1(n9159), .A2(n9158), .A3(n9157), .A4(n9156), .ZN(n12549)
         );
  AND4_X1 U8303 ( .A1(n9125), .A2(n9124), .A3(n9123), .A4(n9122), .ZN(n12477)
         );
  INV_X1 U8304 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9393) );
  OR2_X1 U8305 ( .A1(n11124), .A2(n10957), .ZN(n7119) );
  XNOR2_X1 U8306 ( .A(n9869), .B(n11057), .ZN(n11050) );
  XNOR2_X1 U8307 ( .A(n9871), .B(n9977), .ZN(n11036) );
  NAND2_X1 U8308 ( .A1(n11036), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11035) );
  INV_X1 U8309 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15087) );
  XNOR2_X1 U8310 ( .A(n9879), .B(n9117), .ZN(n14404) );
  NAND2_X1 U8311 ( .A1(n14423), .A2(n14424), .ZN(n14422) );
  NAND2_X1 U8312 ( .A1(n7124), .A2(n6562), .ZN(n7123) );
  NAND2_X1 U8313 ( .A1(n6785), .A2(n6784), .ZN(n12618) );
  NAND2_X1 U8314 ( .A1(n6786), .A2(n6529), .ZN(n6784) );
  NOR2_X1 U8315 ( .A1(n9706), .A2(n12269), .ZN(n9708) );
  OR2_X1 U8316 ( .A1(n12559), .A2(n12584), .ZN(n9707) );
  OAI21_X1 U8317 ( .B1(n9702), .B2(n7405), .A(n7401), .ZN(n11780) );
  AND2_X1 U8318 ( .A1(n12257), .A2(n12665), .ZN(n11776) );
  NAND2_X1 U8319 ( .A1(n7400), .A2(n7406), .ZN(n12670) );
  NAND2_X1 U8320 ( .A1(n9702), .A2(n7408), .ZN(n7400) );
  OR2_X1 U8321 ( .A1(n12676), .A2(n12403), .ZN(n6894) );
  OR2_X1 U8322 ( .A1(n9780), .A2(n12661), .ZN(n12665) );
  NAND2_X1 U8323 ( .A1(n6719), .A2(n6718), .ZN(n12666) );
  INV_X1 U8324 ( .A(n11775), .ZN(n6718) );
  OR2_X1 U8325 ( .A1(n12691), .A2(n12526), .ZN(n12662) );
  NOR2_X1 U8326 ( .A1(n9243), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U8327 ( .A1(n12529), .A2(n9232), .ZN(n9243) );
  AND2_X1 U8328 ( .A1(n9215), .A2(n9214), .ZN(n9232) );
  NOR2_X1 U8329 ( .A1(n9199), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U8330 ( .A1(n9170), .A2(n9169), .ZN(n9185) );
  OR2_X1 U8331 ( .A1(n9185), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9199) );
  NOR2_X1 U8332 ( .A1(n9136), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9154) );
  INV_X1 U8333 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9554) );
  OR2_X1 U8334 ( .A1(n9044), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9065) );
  OR2_X1 U8335 ( .A1(n9065), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9074) );
  NOR2_X1 U8336 ( .A1(n7425), .A2(n6587), .ZN(n7424) );
  INV_X1 U8337 ( .A(n12113), .ZN(n12824) );
  NAND2_X1 U8338 ( .A1(n11452), .A2(n12192), .ZN(n7426) );
  AND2_X1 U8339 ( .A1(n9017), .A2(n8842), .ZN(n9032) );
  INV_X1 U8340 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n9031) );
  AOI21_X1 U8341 ( .B1(n11256), .B2(n6564), .A(n6515), .ZN(n11284) );
  INV_X1 U8342 ( .A(n9680), .ZN(n7437) );
  NAND2_X1 U8343 ( .A1(n11284), .A2(n12172), .ZN(n11362) );
  AND2_X1 U8344 ( .A1(n12114), .A2(n11306), .ZN(n11307) );
  NAND2_X1 U8345 ( .A1(n12163), .A2(n12165), .ZN(n12114) );
  INV_X1 U8346 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9564) );
  INV_X1 U8347 ( .A(n11255), .ZN(n11256) );
  AND2_X1 U8348 ( .A1(n12293), .A2(n15167), .ZN(n9325) );
  OR2_X1 U8349 ( .A1(n11454), .A2(n12276), .ZN(n12550) );
  AND2_X1 U8350 ( .A1(n12633), .A2(n12632), .ZN(n12912) );
  AND4_X1 U8351 ( .A1(n9343), .A2(n9342), .A3(n9341), .A4(n9340), .ZN(n9738)
         );
  NOR2_X1 U8352 ( .A1(n12076), .A2(n12099), .ZN(n12281) );
  INV_X1 U8353 ( .A(n12572), .ZN(n12548) );
  AND2_X1 U8354 ( .A1(n7393), .A2(n6555), .ZN(n12748) );
  NAND2_X1 U8355 ( .A1(n12759), .A2(n12231), .ZN(n7393) );
  INV_X1 U8356 ( .A(n12747), .ZN(n6716) );
  AND2_X1 U8357 ( .A1(n12224), .A2(n12220), .ZN(n12768) );
  INV_X1 U8358 ( .A(n12788), .ZN(n9769) );
  NAND2_X1 U8359 ( .A1(n9786), .A2(n9785), .ZN(n15175) );
  NOR2_X1 U8360 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(n7433), .ZN(n7432) );
  NAND2_X1 U8361 ( .A1(n8804), .A2(n7434), .ZN(n7433) );
  INV_X1 U8362 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U8363 ( .A1(n8792), .A2(n8791), .ZN(n9277) );
  NAND2_X1 U8364 ( .A1(n9263), .A2(n8790), .ZN(n8792) );
  NAND2_X1 U8365 ( .A1(n7280), .A2(n8789), .ZN(n9248) );
  NAND2_X1 U8366 ( .A1(n8782), .A2(n8783), .ZN(n9194) );
  OR2_X1 U8367 ( .A1(n8781), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8782) );
  AOI21_X1 U8368 ( .B1(n7253), .B2(n7255), .A(n7251), .ZN(n7250) );
  INV_X1 U8369 ( .A(n8774), .ZN(n7251) );
  AND2_X1 U8370 ( .A1(n8776), .A2(n8775), .ZN(n9145) );
  AND2_X1 U8371 ( .A1(n8770), .A2(n8769), .ZN(n9092) );
  AND2_X1 U8372 ( .A1(n6995), .A2(n6992), .ZN(n6986) );
  NAND2_X1 U8373 ( .A1(n6869), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9084) );
  AOI21_X1 U8374 ( .B1(n7271), .B2(n7270), .A(n7269), .ZN(n7268) );
  INV_X1 U8375 ( .A(n8757), .ZN(n7269) );
  INV_X1 U8376 ( .A(n8755), .ZN(n7270) );
  AND2_X1 U8377 ( .A1(n8747), .A2(n8746), .ZN(n8922) );
  XNOR2_X1 U8378 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8857) );
  INV_X1 U8379 ( .A(n8100), .ZN(n8102) );
  OR2_X1 U8380 ( .A1(n7812), .A2(n7811), .ZN(n7827) );
  NAND2_X1 U8381 ( .A1(n6803), .A2(n6802), .ZN(n10863) );
  AND2_X1 U8382 ( .A1(n6804), .A2(n10855), .ZN(n6802) );
  NAND2_X1 U8383 ( .A1(n6541), .A2(n7108), .ZN(n7107) );
  INV_X1 U8384 ( .A(n13037), .ZN(n7108) );
  OR2_X1 U8385 ( .A1(n7666), .A2(n7665), .ZN(n7691) );
  OR2_X1 U8386 ( .A1(n7647), .A2(n7646), .ZN(n7666) );
  AND2_X1 U8387 ( .A1(n8009), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U8388 ( .A1(n7101), .A2(n10593), .ZN(n13071) );
  AND2_X1 U8389 ( .A1(n10370), .A2(n10365), .ZN(n7101) );
  OR2_X1 U8390 ( .A1(n7946), .A2(n13083), .ZN(n7985) );
  OR2_X1 U8391 ( .A1(n7738), .A2(n7737), .ZN(n7758) );
  XNOR2_X1 U8392 ( .A(n11742), .B(n10623), .ZN(n10357) );
  NAND2_X1 U8393 ( .A1(n6809), .A2(n11680), .ZN(n13109) );
  INV_X1 U8394 ( .A(n13112), .ZN(n6809) );
  OR2_X1 U8395 ( .A1(n13120), .A2(n11732), .ZN(n11733) );
  AND4_X1 U8396 ( .A1(n8107), .A2(n8106), .A3(n8105), .A4(n8104), .ZN(n11740)
         );
  INV_X1 U8397 ( .A(n8050), .ZN(n8139) );
  NOR2_X1 U8398 ( .A1(n13159), .A2(n13160), .ZN(n13158) );
  NOR2_X1 U8399 ( .A1(n14717), .A2(n14716), .ZN(n14715) );
  INV_X1 U8400 ( .A(n7109), .ZN(n8215) );
  NAND2_X1 U8401 ( .A1(n14789), .A2(n6631), .ZN(n14803) );
  AOI21_X1 U8402 ( .B1(n13198), .B2(n14796), .A(n14802), .ZN(n14816) );
  OAI21_X1 U8403 ( .B1(n13202), .B2(n13201), .A(n14826), .ZN(n13204) );
  NAND2_X1 U8404 ( .A1(n14843), .A2(n6646), .ZN(n14861) );
  OAI21_X1 U8405 ( .B1(n14865), .B2(n13207), .A(n14860), .ZN(n13208) );
  AOI21_X1 U8406 ( .B1(n6913), .B2(n7238), .A(n6575), .ZN(n13318) );
  NAND2_X1 U8407 ( .A1(n6973), .A2(n13283), .ZN(n7238) );
  NAND2_X1 U8408 ( .A1(n13349), .A2(n7239), .ZN(n13339) );
  OR2_X1 U8409 ( .A1(n13572), .A2(n13282), .ZN(n7239) );
  NAND2_X1 U8410 ( .A1(n13396), .A2(n6974), .ZN(n13352) );
  AND2_X1 U8411 ( .A1(n13248), .A2(n13246), .ZN(n13338) );
  NAND2_X1 U8412 ( .A1(n13410), .A2(n13222), .ZN(n13411) );
  AND2_X1 U8413 ( .A1(n7181), .A2(n13427), .ZN(n6761) );
  OAI21_X1 U8414 ( .B1(n7179), .B2(n6760), .A(n6583), .ZN(n6759) );
  AOI21_X1 U8415 ( .B1(n6903), .B2(n7246), .A(n6523), .ZN(n6901) );
  NAND2_X1 U8416 ( .A1(n6978), .A2(n6977), .ZN(n13437) );
  NAND2_X1 U8417 ( .A1(n13511), .A2(n13629), .ZN(n13509) );
  NAND2_X1 U8418 ( .A1(n7166), .A2(n6521), .ZN(n7169) );
  NOR2_X1 U8419 ( .A1(n11271), .A2(n13636), .ZN(n13511) );
  INV_X1 U8420 ( .A(n6908), .ZN(n11270) );
  OAI211_X1 U8421 ( .C1(n10790), .C2(n6910), .A(n6907), .B(n6542), .ZN(n6908)
         );
  NAND2_X1 U8422 ( .A1(n6982), .A2(n6981), .ZN(n11271) );
  INV_X1 U8423 ( .A(n6982), .ZN(n10986) );
  NAND2_X1 U8424 ( .A1(n7163), .A2(n6573), .ZN(n10797) );
  NOR2_X1 U8425 ( .A1(n6571), .A2(n10794), .ZN(n6764) );
  OAI21_X1 U8426 ( .B1(n10756), .B2(n6543), .A(n10733), .ZN(n10796) );
  NOR2_X1 U8427 ( .A1(n10764), .A2(n11703), .ZN(n10763) );
  NAND2_X1 U8428 ( .A1(n6984), .A2(n6983), .ZN(n10764) );
  NAND2_X1 U8429 ( .A1(n7157), .A2(n10477), .ZN(n10511) );
  NAND2_X1 U8430 ( .A1(n10509), .A2(n10507), .ZN(n7157) );
  NAND2_X1 U8431 ( .A1(n9943), .A2(n7571), .ZN(n7153) );
  AOI22_X1 U8432 ( .A1(n8167), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n7572), .B2(
        n14699), .ZN(n7152) );
  AND2_X1 U8433 ( .A1(n10335), .A2(n10154), .ZN(n13523) );
  NAND2_X1 U8434 ( .A1(n6469), .A2(n11012), .ZN(n10265) );
  NAND2_X1 U8435 ( .A1(n6949), .A2(n14944), .ZN(n6948) );
  INV_X1 U8436 ( .A(n13256), .ZN(n6949) );
  INV_X1 U8437 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U8438 ( .A1(n7174), .A2(n7173), .ZN(n6959) );
  INV_X1 U8439 ( .A(n7177), .ZN(n7173) );
  NAND2_X1 U8440 ( .A1(n7176), .A2(n7174), .ZN(n13301) );
  NAND4_X1 U8441 ( .A1(n7236), .A2(n7490), .A3(n7489), .A4(n7109), .ZN(n7494)
         );
  AND2_X1 U8442 ( .A1(n7488), .A2(n8234), .ZN(n7236) );
  INV_X1 U8443 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7514) );
  AND2_X1 U8444 ( .A1(n7308), .A2(n7307), .ZN(n7306) );
  INV_X1 U8445 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7307) );
  AOI21_X1 U8446 ( .B1(n7323), .B2(n7326), .A(n6590), .ZN(n7322) );
  NAND2_X1 U8447 ( .A1(n7323), .A2(n6755), .ZN(n6754) );
  NAND2_X1 U8448 ( .A1(n8568), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8581) );
  OR2_X1 U8449 ( .A1(n8539), .A2(n8538), .ZN(n8548) );
  NOR2_X1 U8450 ( .A1(n11638), .A2(n14302), .ZN(n12372) );
  AOI21_X1 U8451 ( .B1(n6737), .B2(n7341), .A(n6592), .ZN(n6736) );
  INV_X1 U8452 ( .A(n11331), .ZN(n6740) );
  INV_X1 U8453 ( .A(n11330), .ZN(n6741) );
  NOR2_X1 U8454 ( .A1(n13742), .A2(n7335), .ZN(n7334) );
  INV_X1 U8455 ( .A(n11628), .ZN(n7335) );
  NAND2_X1 U8456 ( .A1(n13802), .A2(n13801), .ZN(n7336) );
  AND2_X1 U8457 ( .A1(n13752), .A2(n13750), .ZN(n11559) );
  INV_X1 U8458 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8445) );
  AND2_X1 U8459 ( .A1(n12351), .A2(n12350), .ZN(n13762) );
  AND2_X1 U8460 ( .A1(n8499), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U8461 ( .A1(n13772), .A2(n11594), .ZN(n13723) );
  NAND2_X1 U8462 ( .A1(n13773), .A2(n13774), .ZN(n13772) );
  INV_X1 U8463 ( .A(n8604), .ZN(n8591) );
  NOR2_X1 U8464 ( .A1(n8406), .A2(n11501), .ZN(n8418) );
  NOR2_X1 U8465 ( .A1(n8446), .A2(n8445), .ZN(n8463) );
  AND2_X1 U8466 ( .A1(n13712), .A2(n11645), .ZN(n11647) );
  INV_X1 U8467 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8433) );
  OR2_X1 U8468 ( .A1(n8434), .A2(n8433), .ZN(n8446) );
  NAND2_X1 U8469 ( .A1(n13842), .A2(n13843), .ZN(n13841) );
  OR2_X1 U8470 ( .A1(n13853), .A2(n13854), .ZN(n13851) );
  INV_X1 U8471 ( .A(n12372), .ZN(n11585) );
  OR2_X1 U8472 ( .A1(n8475), .A2(n8474), .ZN(n8485) );
  NOR2_X1 U8473 ( .A1(n8485), .A2(n8484), .ZN(n8499) );
  AOI22_X1 U8474 ( .A1(n11970), .A2(n11969), .B1(n11968), .B2(n11967), .ZN(
        n11984) );
  INV_X1 U8475 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11501) );
  NAND2_X1 U8476 ( .A1(n12018), .A2(n7143), .ZN(n7137) );
  NOR2_X1 U8477 ( .A1(n7141), .A2(n7140), .ZN(n7138) );
  INV_X1 U8478 ( .A(n7143), .ZN(n7140) );
  AND2_X1 U8479 ( .A1(n14033), .A2(n9356), .ZN(n7067) );
  INV_X1 U8480 ( .A(n12014), .ZN(n6666) );
  NAND2_X1 U8481 ( .A1(n6668), .A2(n12014), .ZN(n6667) );
  NAND2_X1 U8482 ( .A1(n9370), .A2(n9371), .ZN(n6668) );
  NOR2_X1 U8483 ( .A1(n12013), .A2(n7094), .ZN(n7090) );
  AND2_X1 U8484 ( .A1(n14081), .A2(n7092), .ZN(n7091) );
  NAND2_X1 U8485 ( .A1(n7089), .A2(n7094), .ZN(n14082) );
  NAND2_X1 U8486 ( .A1(n14118), .A2(n7092), .ZN(n7089) );
  INV_X1 U8487 ( .A(n12011), .ZN(n14120) );
  OR2_X1 U8488 ( .A1(n14118), .A2(n14120), .ZN(n14116) );
  NAND2_X1 U8489 ( .A1(n6961), .A2(n6960), .ZN(n14137) );
  INV_X1 U8490 ( .A(n6961), .ZN(n14156) );
  NAND2_X1 U8491 ( .A1(n7070), .A2(n7069), .ZN(n14148) );
  NOR2_X1 U8492 ( .A1(n14161), .A2(n8681), .ZN(n7069) );
  NAND2_X1 U8493 ( .A1(n14185), .A2(n14320), .ZN(n14170) );
  OR2_X1 U8494 ( .A1(n8523), .A2(n8522), .ZN(n8539) );
  NAND2_X1 U8495 ( .A1(n8510), .A2(n8509), .ZN(n14213) );
  AND2_X1 U8496 ( .A1(n11870), .A2(n8491), .ZN(n8493) );
  INV_X1 U8497 ( .A(n11871), .ZN(n7064) );
  NAND2_X1 U8498 ( .A1(n10451), .A2(n11971), .ZN(n6685) );
  NOR2_X1 U8499 ( .A1(n6968), .A2(n11866), .ZN(n6967) );
  NAND2_X1 U8500 ( .A1(n7148), .A2(n8440), .ZN(n11373) );
  NAND2_X1 U8501 ( .A1(n7148), .A2(n7147), .ZN(n11375) );
  AOI21_X1 U8502 ( .B1(n11996), .B2(n7074), .A(n6552), .ZN(n7072) );
  NAND2_X1 U8503 ( .A1(n7076), .A2(n7074), .ZN(n11184) );
  NAND2_X1 U8504 ( .A1(n7077), .A2(n7079), .ZN(n7076) );
  NOR2_X1 U8505 ( .A1(n11190), .A2(n11849), .ZN(n11296) );
  INV_X1 U8506 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8389) );
  OR2_X1 U8507 ( .A1(n8390), .A2(n8389), .ZN(n8406) );
  INV_X1 U8508 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8378) );
  OR2_X1 U8509 ( .A1(n8379), .A2(n8378), .ZN(n8390) );
  NAND2_X1 U8510 ( .A1(n8337), .A2(n8336), .ZN(n7133) );
  INV_X1 U8511 ( .A(n12317), .ZN(n6972) );
  NAND2_X1 U8512 ( .A1(n14075), .A2(n8600), .ZN(n14066) );
  NAND2_X1 U8513 ( .A1(n8579), .A2(n8578), .ZN(n14289) );
  INV_X1 U8514 ( .A(n14522), .ZN(n14642) );
  INV_X1 U8515 ( .A(n14680), .ZN(n14669) );
  AND2_X1 U8516 ( .A1(n8702), .A2(n6615), .ZN(n8267) );
  INV_X1 U8517 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7380) );
  XNOR2_X1 U8518 ( .A(n8132), .B(n8131), .ZN(n13670) );
  NAND2_X1 U8519 ( .A1(n8166), .A2(n8129), .ZN(n8132) );
  XNOR2_X1 U8520 ( .A(n8145), .B(n8144), .ZN(n13678) );
  OAI21_X1 U8521 ( .B1(n8111), .B2(n8110), .A(n8109), .ZN(n8122) );
  XNOR2_X1 U8522 ( .A(n8111), .B(n8096), .ZN(n11655) );
  NAND3_X1 U8523 ( .A1(n8533), .A2(n8257), .A3(n7150), .ZN(n8706) );
  OAI21_X1 U8524 ( .B1(n8080), .B2(n8079), .A(n8078), .ZN(n8094) );
  XNOR2_X1 U8525 ( .A(n8080), .B(n8079), .ZN(n11475) );
  AND2_X1 U8526 ( .A1(n8699), .A2(n8698), .ZN(n8712) );
  XNOR2_X1 U8527 ( .A(n8055), .B(n8056), .ZN(n11439) );
  XNOR2_X1 U8528 ( .A(n7972), .B(n7971), .ZN(n11234) );
  INV_X1 U8529 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8638) );
  OAI21_X1 U8530 ( .B1(n7723), .B2(n7744), .A(n6924), .ZN(n7764) );
  NAND2_X1 U8531 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  NAND2_X1 U8532 ( .A1(n7200), .A2(n7676), .ZN(n7699) );
  INV_X1 U8533 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n9385) );
  INV_X1 U8534 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9386) );
  INV_X1 U8535 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9389) );
  INV_X1 U8536 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13916) );
  NAND2_X1 U8537 ( .A1(n9399), .A2(n9398), .ZN(n9448) );
  NAND2_X1 U8538 ( .A1(n14550), .A2(n6680), .ZN(n9471) );
  OAI21_X1 U8539 ( .B1(n14551), .B2(n14552), .A(n6681), .ZN(n6680) );
  INV_X1 U8540 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6681) );
  AOI21_X1 U8541 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9415), .A(n9414), .ZN(
        n9421) );
  AND2_X1 U8542 ( .A1(n8881), .A2(n15116), .ZN(n8882) );
  NAND2_X1 U8543 ( .A1(n7010), .A2(n9207), .ZN(n12441) );
  NAND2_X1 U8544 ( .A1(n7017), .A2(n6540), .ZN(n7016) );
  OAI22_X1 U8545 ( .A1(n12082), .A2(n9982), .B1(n6500), .B2(n9855), .ZN(n6674)
         );
  NAND2_X1 U8546 ( .A1(n6998), .A2(n9161), .ZN(n12547) );
  NAND2_X1 U8547 ( .A1(n12485), .A2(n12484), .ZN(n6998) );
  NAND2_X1 U8548 ( .A1(n8952), .A2(n8951), .ZN(n11173) );
  INV_X1 U8549 ( .A(n12530), .ZN(n14982) );
  NAND2_X1 U8550 ( .A1(n9322), .A2(n9321), .ZN(n14974) );
  AND2_X1 U8551 ( .A1(n9335), .A2(n9334), .ZN(n14985) );
  INV_X1 U8552 ( .A(n14973), .ZN(n12577) );
  AND4_X1 U8553 ( .A1(n12090), .A2(n9735), .A3(n9734), .A4(n9733), .ZN(n12102)
         );
  NAND4_X1 U8554 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n12585)
         );
  INV_X1 U8555 ( .A(n12443), .ZN(n12589) );
  NAND4_X1 U8556 ( .A1(n8947), .A2(n8946), .A3(n8945), .A4(n8944), .ZN(n12604)
         );
  OR2_X1 U8557 ( .A1(n9723), .A2(n11168), .ZN(n8917) );
  INV_X1 U8558 ( .A(P3_U3897), .ZN(n12607) );
  CLKBUF_X1 U8559 ( .A(n8880), .Z(n12608) );
  AND2_X1 U8560 ( .A1(n9833), .A2(n7119), .ZN(n11075) );
  INV_X1 U8561 ( .A(n7128), .ZN(n11047) );
  INV_X1 U8562 ( .A(n9837), .ZN(n7127) );
  NOR2_X1 U8563 ( .A1(n11032), .A2(n9840), .ZN(n10912) );
  NAND2_X1 U8564 ( .A1(n10913), .A2(n9902), .ZN(n14996) );
  INV_X1 U8565 ( .A(n7113), .ZN(n9841) );
  NAND2_X1 U8566 ( .A1(n6780), .A2(n6781), .ZN(n15023) );
  INV_X1 U8567 ( .A(n7120), .ZN(n9843) );
  NOR2_X1 U8568 ( .A1(n15039), .A2(n6766), .ZN(n15059) );
  AND2_X1 U8569 ( .A1(n9907), .A2(n9908), .ZN(n6766) );
  NAND2_X1 U8570 ( .A1(n15059), .A2(n15058), .ZN(n15057) );
  NOR2_X1 U8571 ( .A1(n15063), .A2(n9846), .ZN(n15083) );
  NOR2_X1 U8572 ( .A1(n15083), .A2(n15082), .ZN(n15081) );
  AOI21_X1 U8573 ( .B1(n9914), .B2(n9913), .A(n15073), .ZN(n15099) );
  NOR2_X1 U8574 ( .A1(n14401), .A2(n14402), .ZN(n14400) );
  NOR2_X1 U8575 ( .A1(n14414), .A2(n9923), .ZN(n14421) );
  NAND2_X1 U8576 ( .A1(n6790), .A2(n6526), .ZN(n14438) );
  AND2_X1 U8577 ( .A1(n6788), .A2(n6790), .ZN(n14436) );
  INV_X1 U8578 ( .A(n7124), .ZN(n14444) );
  AND2_X1 U8579 ( .A1(n9934), .A2(n9933), .ZN(n15089) );
  NAND2_X1 U8580 ( .A1(n6652), .A2(n14441), .ZN(n9938) );
  NAND2_X1 U8581 ( .A1(n6653), .A2(n12610), .ZN(n6652) );
  NAND2_X1 U8582 ( .A1(n9859), .A2(n9858), .ZN(n6653) );
  INV_X1 U8583 ( .A(n7123), .ZN(n9859) );
  AND2_X1 U8584 ( .A1(n9800), .A2(n9339), .ZN(n12645) );
  AND2_X1 U8585 ( .A1(n9338), .A2(n8845), .ZN(n12655) );
  NAND2_X1 U8586 ( .A1(n8811), .A2(n8810), .ZN(n12855) );
  OR2_X1 U8587 ( .A1(n9714), .A2(n7211), .ZN(n9227) );
  NAND2_X1 U8588 ( .A1(n7382), .A2(n7389), .ZN(n12708) );
  NAND2_X1 U8589 ( .A1(n9213), .A2(n9212), .ZN(n12877) );
  OR2_X1 U8590 ( .A1(n9714), .A2(n10683), .ZN(n9212) );
  NAND2_X1 U8591 ( .A1(n9119), .A2(n9118), .ZN(n12896) );
  NOR3_X1 U8592 ( .A1(n9799), .A2(n15122), .A3(n15185), .ZN(n12798) );
  AND3_X1 U8593 ( .A1(n8958), .A2(n8957), .A3(n8956), .ZN(n15158) );
  AND2_X1 U8594 ( .A1(n12694), .A2(n9798), .ZN(n12802) );
  INV_X1 U8595 ( .A(n15175), .ZN(n15164) );
  NAND2_X1 U8596 ( .A1(n9325), .A2(n15122), .ZN(n15121) );
  AND2_X1 U8597 ( .A1(n9799), .A2(n15121), .ZN(n15128) );
  OR2_X1 U8598 ( .A1(n12082), .A2(n9959), .ZN(n8877) );
  OR2_X1 U8599 ( .A1(n8984), .A2(n9958), .ZN(n8873) );
  INV_X1 U8600 ( .A(n15205), .ZN(n15203) );
  OAI22_X1 U8601 ( .A1(n12307), .A2(n12082), .B1(n12306), .B2(n9714), .ZN(
        n12915) );
  NAND2_X1 U8602 ( .A1(n9716), .A2(n9715), .ZN(n12921) );
  OAI21_X1 U8603 ( .B1(n11756), .B2(n7418), .A(n7416), .ZN(n12641) );
  AOI21_X1 U8604 ( .B1(n11772), .B2(n6539), .A(n6864), .ZN(n12639) );
  NAND2_X1 U8605 ( .A1(n6863), .A2(n6866), .ZN(n12650) );
  NAND2_X1 U8606 ( .A1(n11772), .A2(n11754), .ZN(n6863) );
  NOR2_X1 U8607 ( .A1(n11772), .A2(n9783), .ZN(n11755) );
  INV_X1 U8608 ( .A(n12691), .ZN(n12939) );
  NAND2_X1 U8609 ( .A1(n9198), .A2(n9197), .ZN(n12950) );
  OR2_X1 U8610 ( .A1(n9714), .A2(n10578), .ZN(n9197) );
  NAND2_X1 U8611 ( .A1(n9168), .A2(n9167), .ZN(n12962) );
  NAND2_X1 U8612 ( .A1(n9153), .A2(n9152), .ZN(n12968) );
  AND3_X1 U8613 ( .A1(n9064), .A2(n9063), .A3(n9062), .ZN(n12993) );
  INV_X1 U8614 ( .A(n10618), .ZN(n10685) );
  AND2_X1 U8615 ( .A1(n9294), .A2(n9293), .ZN(n12999) );
  INV_X1 U8616 ( .A(n9318), .ZN(n13001) );
  NAND2_X1 U8617 ( .A1(n9856), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13000) );
  XNOR2_X1 U8618 ( .A(n12096), .B(n12095), .ZN(n13008) );
  OR2_X1 U8619 ( .A1(n12092), .A2(n12091), .ZN(n12094) );
  XNOR2_X1 U8620 ( .A(n12092), .B(n6669), .ZN(n12307) );
  INV_X1 U8621 ( .A(n12091), .ZN(n6669) );
  NAND2_X1 U8622 ( .A1(n8836), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8838) );
  INV_X1 U8623 ( .A(SI_25_), .ZN(n11281) );
  OAI21_X1 U8624 ( .B1(n9226), .B2(n9225), .A(n8786), .ZN(n9240) );
  AND2_X1 U8625 ( .A1(n9313), .A2(n6513), .ZN(n12297) );
  XNOR2_X1 U8626 ( .A(n8826), .B(n8825), .ZN(n12139) );
  INV_X1 U8627 ( .A(SI_20_), .ZN(n10578) );
  XNOR2_X1 U8628 ( .A(n8828), .B(n6775), .ZN(n10579) );
  INV_X1 U8629 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n6723) );
  OAI21_X1 U8630 ( .B1(n9163), .B2(n7261), .A(n7259), .ZN(n9180) );
  NAND2_X1 U8631 ( .A1(n9165), .A2(n8778), .ZN(n9178) );
  INV_X1 U8632 ( .A(SI_16_), .ZN(n10088) );
  OAI21_X1 U8633 ( .B1(n9111), .B2(n7255), .A(n7253), .ZN(n9131) );
  NAND2_X1 U8634 ( .A1(n9113), .A2(n8772), .ZN(n9129) );
  INV_X1 U8635 ( .A(SI_15_), .ZN(n10058) );
  INV_X1 U8636 ( .A(SI_12_), .ZN(n9967) );
  NAND2_X1 U8637 ( .A1(n7264), .A2(n8762), .ZN(n9053) );
  NAND2_X1 U8638 ( .A1(n9027), .A2(n8761), .ZN(n7264) );
  NAND2_X1 U8639 ( .A1(n8983), .A2(n8755), .ZN(n8990) );
  NOR2_X1 U8640 ( .A1(n6492), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14381) );
  AND2_X1 U8641 ( .A1(n12052), .A2(n11657), .ZN(n11658) );
  INV_X1 U8642 ( .A(n10856), .ZN(n14928) );
  NAND2_X1 U8643 ( .A1(n10593), .A2(n10365), .ZN(n10373) );
  AND2_X1 U8644 ( .A1(n12066), .A2(n10848), .ZN(n6806) );
  NAND2_X1 U8645 ( .A1(n6792), .A2(n11004), .ZN(n11417) );
  NAND2_X1 U8646 ( .A1(n14464), .A2(n10998), .ZN(n6792) );
  INV_X1 U8647 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10999) );
  OR2_X1 U8648 ( .A1(n11727), .A2(n11728), .ZN(n6801) );
  NAND2_X1 U8649 ( .A1(n13141), .A2(n11668), .ZN(n13043) );
  NAND2_X1 U8650 ( .A1(n7885), .A2(n7884), .ZN(n13485) );
  NAND2_X1 U8651 ( .A1(n13141), .A2(n7099), .ZN(n13057) );
  AND2_X1 U8652 ( .A1(n11668), .A2(n7100), .ZN(n7099) );
  INV_X1 U8653 ( .A(n13044), .ZN(n7100) );
  NAND2_X1 U8654 ( .A1(n9945), .A2(n8097), .ZN(n6810) );
  AND4_X2 U8655 ( .A1(n7532), .A2(n7531), .A3(n7530), .A4(n7529), .ZN(n8193)
         );
  NAND2_X1 U8656 ( .A1(n11709), .A2(n13086), .ZN(n13093) );
  AOI21_X1 U8657 ( .B1(n11682), .B2(n13111), .A(n6589), .ZN(n6808) );
  NOR2_X1 U8658 ( .A1(n10349), .A2(n10334), .ZN(n13122) );
  NAND2_X1 U8659 ( .A1(n13109), .A2(n11682), .ZN(n13090) );
  NAND2_X1 U8660 ( .A1(n11417), .A2(n11416), .ZN(n11419) );
  NAND2_X1 U8661 ( .A1(n10995), .A2(n10994), .ZN(n14461) );
  NAND2_X1 U8662 ( .A1(n10534), .A2(n7112), .ZN(n10666) );
  AND2_X1 U8663 ( .A1(n10541), .A2(n10533), .ZN(n7112) );
  NAND2_X1 U8664 ( .A1(n10534), .A2(n10533), .ZN(n10539) );
  NOR2_X1 U8665 ( .A1(n13119), .A2(n11733), .ZN(n13127) );
  OR2_X1 U8666 ( .A1(n14462), .A2(n13510), .ZN(n13132) );
  XNOR2_X1 U8667 ( .A(n7192), .B(n13216), .ZN(n8204) );
  NAND2_X1 U8668 ( .A1(n8203), .A2(n6550), .ZN(n7192) );
  INV_X1 U8669 ( .A(n11740), .ZN(n13285) );
  NAND4_X1 U8670 ( .A1(n7541), .A2(n7540), .A3(n7539), .A4(n7538), .ZN(n13155)
         );
  INV_X1 U8671 ( .A(n8193), .ZN(n13156) );
  NOR2_X1 U8672 ( .A1(n10081), .A2(n10080), .ZN(n10079) );
  NAND2_X1 U8673 ( .A1(n13190), .A2(n6629), .ZN(n14754) );
  NAND2_X1 U8674 ( .A1(n14754), .A2(n14753), .ZN(n14752) );
  AND2_X1 U8675 ( .A1(n7703), .A2(n7725), .ZN(n14759) );
  AOI21_X1 U8676 ( .B1(n13195), .B2(n13194), .A(n14764), .ZN(n14775) );
  NAND2_X1 U8677 ( .A1(n14791), .A2(n14790), .ZN(n14789) );
  AND2_X1 U8678 ( .A1(n7803), .A2(n7840), .ZN(n14817) );
  INV_X1 U8679 ( .A(n13231), .ZN(n13230) );
  OR2_X1 U8680 ( .A1(n13306), .A2(n13550), .ZN(n6692) );
  OR3_X1 U8681 ( .A1(n13321), .A2(n13320), .A3(n10602), .ZN(n13559) );
  AND2_X1 U8682 ( .A1(n6898), .A2(n6897), .ZN(n13351) );
  NAND2_X1 U8683 ( .A1(n6900), .A2(n7240), .ZN(n13364) );
  NAND2_X1 U8684 ( .A1(n13393), .A2(n7242), .ZN(n13380) );
  NAND2_X1 U8685 ( .A1(n6758), .A2(n7179), .ZN(n13419) );
  NAND2_X1 U8686 ( .A1(n13459), .A2(n7181), .ZN(n6758) );
  NAND2_X1 U8687 ( .A1(n7183), .A2(n7184), .ZN(n13434) );
  NAND2_X1 U8688 ( .A1(n7187), .A2(n7185), .ZN(n7183) );
  NAND2_X1 U8689 ( .A1(n13452), .A2(n13268), .ZN(n13432) );
  NAND2_X1 U8690 ( .A1(n13463), .A2(n13266), .ZN(n13454) );
  NAND2_X1 U8691 ( .A1(n7873), .A2(n7872), .ZN(n13618) );
  NAND2_X1 U8692 ( .A1(n7168), .A2(n11264), .ZN(n13237) );
  NAND2_X1 U8693 ( .A1(n7172), .A2(n7170), .ZN(n7168) );
  NAND2_X1 U8694 ( .A1(n7172), .A2(n7438), .ZN(n11266) );
  NAND2_X1 U8695 ( .A1(n10790), .A2(n6911), .ZN(n6909) );
  NAND2_X1 U8696 ( .A1(n7232), .A2(n7233), .ZN(n10990) );
  NAND2_X1 U8697 ( .A1(n10792), .A2(n7234), .ZN(n7232) );
  NAND2_X1 U8698 ( .A1(n10792), .A2(n10791), .ZN(n10880) );
  INV_X1 U8699 ( .A(n13533), .ZN(n10597) );
  AND2_X1 U8700 ( .A1(n13527), .A2(n10500), .ZN(n13534) );
  OAI21_X1 U8701 ( .B1(n7870), .B2(n9942), .A(n7249), .ZN(n7248) );
  AND2_X1 U8702 ( .A1(n13527), .A2(n10428), .ZN(n13530) );
  INV_X1 U8703 ( .A(n13530), .ZN(n13489) );
  INV_X1 U8704 ( .A(n13515), .ZN(n13538) );
  INV_X2 U8705 ( .A(n14957), .ZN(n14960) );
  INV_X1 U8706 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U8707 ( .A1(n13672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7493) );
  XNOR2_X1 U8708 ( .A(n8235), .B(n8234), .ZN(n13690) );
  NAND2_X1 U8709 ( .A1(n8233), .A2(n8232), .ZN(n11440) );
  INV_X1 U8710 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10789) );
  INV_X1 U8711 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10446) );
  INV_X1 U8712 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10401) );
  INV_X1 U8713 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10452) );
  INV_X1 U8714 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10421) );
  INV_X1 U8715 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10097) );
  INV_X1 U8716 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10070) );
  INV_X1 U8717 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10047) );
  INV_X1 U8718 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10039) );
  INV_X1 U8719 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10006) );
  INV_X1 U8720 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9990) );
  INV_X1 U8721 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9972) );
  INV_X1 U8722 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9966) );
  INV_X1 U8723 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9946) );
  INV_X1 U8724 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U8725 ( .A1(n13692), .A2(n6748), .ZN(n13694) );
  OAI21_X1 U8726 ( .B1(n13842), .B2(n12359), .A(n7320), .ZN(n13692) );
  NAND2_X1 U8727 ( .A1(n13841), .A2(n6749), .ZN(n6748) );
  NOR2_X1 U8728 ( .A1(n13693), .A2(n12359), .ZN(n6749) );
  AOI21_X1 U8729 ( .B1(n7328), .B2(n13781), .A(n6579), .ZN(n7327) );
  AOI21_X1 U8730 ( .B1(n7320), .B2(n12359), .A(n12369), .ZN(n7319) );
  NAND2_X1 U8731 ( .A1(n6735), .A2(n6736), .ZN(n11339) );
  NAND2_X1 U8732 ( .A1(n7336), .A2(n11628), .ZN(n13743) );
  NAND2_X1 U8733 ( .A1(n13749), .A2(n11559), .ZN(n13751) );
  AND2_X1 U8734 ( .A1(n11199), .A2(n11198), .ZN(n11246) );
  INV_X1 U8735 ( .A(n14213), .ZN(n14488) );
  NAND2_X1 U8736 ( .A1(n13716), .A2(n13792), .ZN(n7313) );
  NOR2_X1 U8737 ( .A1(n13847), .A2(n14522), .ZN(n13825) );
  INV_X1 U8738 ( .A(n13877), .ZN(n13827) );
  OAI21_X2 U8739 ( .B1(n10296), .B2(n10650), .A(n14206), .ZN(n13817) );
  NOR2_X1 U8740 ( .A1(n11244), .A2(n11243), .ZN(n7339) );
  AOI21_X1 U8741 ( .B1(n7340), .B2(n11244), .A(n7338), .ZN(n7337) );
  NAND2_X1 U8742 ( .A1(n11198), .A2(n11203), .ZN(n7340) );
  OR2_X1 U8743 ( .A1(n10292), .A2(n12031), .ZN(n13847) );
  NAND2_X1 U8744 ( .A1(n10285), .A2(n10284), .ZN(n13864) );
  NAND4_X1 U8745 ( .A1(n8619), .A2(n8618), .A3(n8617), .A4(n8616), .ZN(n13871)
         );
  OAI21_X1 U8746 ( .B1(n14139), .B2(n8543), .A(n8564), .ZN(n14152) );
  NAND2_X1 U8747 ( .A1(n8554), .A2(n8553), .ZN(n14317) );
  OR2_X1 U8748 ( .A1(n8516), .A2(n8515), .ZN(n13872) );
  NAND2_X1 U8749 ( .A1(n8533), .A2(n8532), .ZN(n8637) );
  INV_X1 U8750 ( .A(n14289), .ZN(n14115) );
  NAND2_X1 U8751 ( .A1(n14368), .A2(n8304), .ZN(n14295) );
  NAND2_X1 U8752 ( .A1(n7080), .A2(n7083), .ZN(n14190) );
  NAND2_X1 U8753 ( .A1(n7087), .A2(n12005), .ZN(n7086) );
  NAND2_X1 U8754 ( .A1(n8498), .A2(n8497), .ZN(n14236) );
  NAND2_X1 U8755 ( .A1(n8462), .A2(n8461), .ZN(n14525) );
  NOR3_X1 U8756 ( .A1(n11190), .A2(n11854), .A3(n11849), .ZN(n11354) );
  NAND2_X1 U8757 ( .A1(n10295), .A2(n10294), .ZN(n14206) );
  INV_X1 U8758 ( .A(n14206), .ZN(n14243) );
  INV_X1 U8759 ( .A(n14019), .ZN(n14329) );
  INV_X1 U8760 ( .A(n11985), .ZN(n14333) );
  INV_X1 U8761 ( .A(n14087), .ZN(n14341) );
  NAND2_X1 U8762 ( .A1(n10048), .A2(n10295), .ZN(n14639) );
  NAND2_X1 U8763 ( .A1(n8166), .A2(n8165), .ZN(n13677) );
  NOR2_X1 U8764 ( .A1(n7061), .A2(n7060), .ZN(n7059) );
  INV_X1 U8765 ( .A(n8712), .ZN(n11542) );
  INV_X1 U8766 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10787) );
  INV_X1 U8767 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10449) );
  INV_X1 U8768 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10422) );
  INV_X1 U8769 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10453) );
  INV_X1 U8770 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10447) );
  INV_X1 U8771 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10243) );
  INV_X1 U8772 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10092) );
  INV_X1 U8773 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10045) );
  INV_X1 U8774 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10040) );
  INV_X1 U8775 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10003) );
  INV_X1 U8776 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9991) );
  AND2_X1 U8777 ( .A1(n8375), .A2(n8386), .ZN(n13939) );
  INV_X1 U8778 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U8779 ( .A1(n7357), .A2(n8314), .ZN(n8286) );
  XNOR2_X1 U8780 ( .A(n8296), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13888) );
  NOR2_X1 U8781 ( .A1(n15220), .A2(n9438), .ZN(n14377) );
  NAND2_X1 U8782 ( .A1(n14376), .A2(n7039), .ZN(n15217) );
  OAI21_X1 U8783 ( .B1(n14377), .B2(n14378), .A(n7040), .ZN(n7039) );
  INV_X1 U8784 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7040) );
  NOR2_X1 U8785 ( .A1(n15217), .A2(n15218), .ZN(n15216) );
  INV_X1 U8786 ( .A(n9445), .ZN(n6725) );
  INV_X1 U8787 ( .A(n9457), .ZN(n9458) );
  XNOR2_X1 U8788 ( .A(n9471), .B(n9470), .ZN(n14556) );
  INV_X1 U8789 ( .A(n9469), .ZN(n9470) );
  NAND2_X1 U8790 ( .A1(n7042), .A2(n7041), .ZN(n14397) );
  AOI22_X1 U8791 ( .A1(n7047), .A2(n7049), .B1(n7045), .B2(n7051), .ZN(n7041)
         );
  INV_X1 U8792 ( .A(n7050), .ZN(n7049) );
  INV_X1 U8793 ( .A(n6711), .ZN(n6710) );
  XNOR2_X1 U8794 ( .A(n6695), .B(n12619), .ZN(n12629) );
  NAND2_X1 U8795 ( .A1(n12676), .A2(n12901), .ZN(n6679) );
  NOR2_X1 U8796 ( .A1(n6714), .A2(n6713), .ZN(n6712) );
  NOR2_X1 U8797 ( .A1(n15193), .A2(n12930), .ZN(n6713) );
  NAND2_X1 U8798 ( .A1(n12676), .A2(n12985), .ZN(n6678) );
  AND2_X1 U8799 ( .A1(n6803), .A2(n6804), .ZN(n11705) );
  NAND2_X1 U8800 ( .A1(n13554), .A2(n13553), .ZN(n13651) );
  INV_X1 U8801 ( .A(n6943), .ZN(n6942) );
  NOR2_X1 U8802 ( .A1(n6625), .A2(n14942), .ZN(n6945) );
  AOI21_X1 U8803 ( .B1(n12317), .B2(n14124), .A(n12316), .ZN(n6693) );
  NOR2_X1 U8804 ( .A1(n9359), .A2(n9361), .ZN(n9362) );
  NOR2_X1 U8805 ( .A1(n12301), .A2(n14348), .ZN(n9359) );
  AOI21_X1 U8806 ( .B1(n9668), .B2(n14687), .A(n9381), .ZN(n9382) );
  NAND2_X1 U8807 ( .A1(n6626), .A2(n9380), .ZN(n9381) );
  NAND2_X1 U8808 ( .A1(n7030), .A2(n7029), .ZN(n15214) );
  INV_X1 U8809 ( .A(n7028), .ZN(n15213) );
  NAND2_X1 U8810 ( .A1(n7052), .A2(n7053), .ZN(n14572) );
  AND2_X1 U8811 ( .A1(n7052), .A2(n7050), .ZN(n14570) );
  XNOR2_X1 U8812 ( .A(n9665), .B(n9494), .ZN(n7034) );
  NAND2_X1 U8813 ( .A1(n10274), .A2(n10273), .ZN(n11638) );
  INV_X1 U8814 ( .A(n7523), .ZN(n7547) );
  AND2_X1 U8815 ( .A1(n7240), .A2(n6899), .ZN(n6511) );
  CLKBUF_X3 U8816 ( .A(n7807), .Z(n7773) );
  NAND3_X2 U8817 ( .A1(n6856), .A2(n6854), .A3(n6853), .ZN(n11835) );
  INV_X1 U8818 ( .A(n13388), .ZN(n7241) );
  AND3_X1 U8819 ( .A1(n6610), .A2(n6990), .A3(n6986), .ZN(n8932) );
  NOR2_X1 U8820 ( .A1(n9042), .A2(n11465), .ZN(n6512) );
  OR2_X1 U8821 ( .A1(n9311), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8822 ( .A1(n7088), .A2(n6547), .ZN(n7085) );
  NOR2_X1 U8823 ( .A1(n7013), .A2(n7011), .ZN(n6514) );
  NOR2_X1 U8824 ( .A1(n9680), .A2(n11307), .ZN(n6515) );
  INV_X1 U8825 ( .A(n11954), .ZN(n6843) );
  NAND3_X1 U8826 ( .A1(n8932), .A2(n7430), .A3(n7429), .ZN(n6516) );
  INV_X1 U8827 ( .A(n12231), .ZN(n12758) );
  INV_X1 U8828 ( .A(n7243), .ZN(n7242) );
  NAND2_X1 U8829 ( .A1(n13381), .A2(n13279), .ZN(n7243) );
  AND2_X1 U8830 ( .A1(n6594), .A2(n6850), .ZN(n6517) );
  INV_X1 U8831 ( .A(n11996), .ZN(n7079) );
  OR2_X1 U8832 ( .A1(n12921), .A2(n9738), .ZN(n9784) );
  OR2_X1 U8833 ( .A1(n9452), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6518) );
  OR2_X1 U8834 ( .A1(n13229), .A2(n13293), .ZN(n6519) );
  AND2_X1 U8835 ( .A1(n14046), .A2(n8690), .ZN(n6520) );
  NAND2_X1 U8836 ( .A1(n11923), .A2(n11926), .ZN(n7358) );
  INV_X1 U8837 ( .A(n7358), .ZN(n6828) );
  OR2_X1 U8838 ( .A1(n13636), .A2(n13504), .ZN(n6521) );
  XOR2_X1 U8839 ( .A(n11780), .B(n11779), .Z(n6522) );
  AND2_X1 U8840 ( .A1(n13608), .A2(n13270), .ZN(n6523) );
  AND2_X1 U8841 ( .A1(n10471), .A2(n8190), .ZN(n10508) );
  AND4_X1 U8842 ( .A1(n9247), .A2(n9246), .A3(n9245), .A4(n9244), .ZN(n12526)
         );
  INV_X1 U8843 ( .A(n11960), .ZN(n11794) );
  XNOR2_X1 U8844 ( .A(n8642), .B(P1_IR_REG_21__SCAN_IN), .ZN(n11960) );
  INV_X1 U8845 ( .A(n14168), .ZN(n7071) );
  AND2_X1 U8846 ( .A1(n13263), .A2(n13262), .ZN(n6524) );
  INV_X1 U8847 ( .A(n13792), .ZN(n7316) );
  AND2_X1 U8848 ( .A1(n6649), .A2(n9902), .ZN(n6525) );
  AND2_X1 U8849 ( .A1(n6787), .A2(n14419), .ZN(n6526) );
  NAND2_X1 U8850 ( .A1(n9250), .A2(n9249), .ZN(n12676) );
  NAND2_X1 U8851 ( .A1(n13618), .A2(n13238), .ZN(n7190) );
  XNOR2_X1 U8852 ( .A(n8534), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14106) );
  AND2_X1 U8853 ( .A1(n8039), .A2(SI_24_), .ZN(n6527) );
  AND2_X1 U8854 ( .A1(n6789), .A2(n14419), .ZN(n6528) );
  OR2_X1 U8855 ( .A1(n6791), .A2(n14433), .ZN(n6529) );
  INV_X1 U8856 ( .A(n13076), .ZN(n6979) );
  NOR2_X1 U8857 ( .A1(n11400), .A2(n6738), .ZN(n6737) );
  INV_X2 U8858 ( .A(n9883), .ZN(n9922) );
  OR2_X1 U8859 ( .A1(n11562), .A2(n11561), .ZN(n6530) );
  OR2_X1 U8860 ( .A1(n9149), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6531) );
  INV_X1 U8861 ( .A(n15154), .ZN(n7435) );
  INV_X1 U8862 ( .A(n8913), .ZN(n9732) );
  INV_X1 U8863 ( .A(n11027), .ZN(n6656) );
  AND2_X1 U8864 ( .A1(n7677), .A2(n7309), .ZN(n7702) );
  AND2_X1 U8865 ( .A1(n7336), .A2(n7334), .ZN(n6532) );
  NAND2_X1 U8866 ( .A1(n8712), .A2(n8711), .ZN(n10274) );
  NAND2_X1 U8867 ( .A1(n6728), .A2(n13713), .ZN(n13716) );
  AND2_X1 U8868 ( .A1(n7313), .A2(n13793), .ZN(n6533) );
  OR2_X1 U8869 ( .A1(n9311), .A2(n7013), .ZN(n6534) );
  AND2_X1 U8870 ( .A1(n7026), .A2(n7025), .ZN(n6535) );
  INV_X1 U8871 ( .A(n11754), .ZN(n12266) );
  OR2_X1 U8872 ( .A1(n12559), .A2(n12269), .ZN(n11754) );
  INV_X1 U8873 ( .A(n12005), .ZN(n14227) );
  NAND2_X1 U8874 ( .A1(n13641), .A2(n13145), .ZN(n6536) );
  AND3_X1 U8875 ( .A1(n8284), .A2(n8283), .A3(n8282), .ZN(n6537) );
  NOR2_X1 U8876 ( .A1(n12408), .A2(n8931), .ZN(n6538) );
  AND2_X1 U8877 ( .A1(n12651), .A2(n11754), .ZN(n6539) );
  NOR2_X1 U8878 ( .A1(n12495), .A2(n7447), .ZN(n6540) );
  NAND2_X1 U8879 ( .A1(n11735), .A2(n11734), .ZN(n6541) );
  OR2_X1 U8880 ( .A1(n13641), .A2(n13145), .ZN(n6542) );
  AND2_X1 U8881 ( .A1(n11703), .A2(n10868), .ZN(n6543) );
  NOR2_X1 U8882 ( .A1(n12601), .A2(n9682), .ZN(n6544) );
  NAND2_X1 U8883 ( .A1(n13396), .A2(n6976), .ZN(n6545) );
  AND2_X1 U8884 ( .A1(n10850), .A2(n10849), .ZN(n6546) );
  OR2_X1 U8885 ( .A1(n14494), .A2(n14500), .ZN(n6547) );
  NAND3_X1 U8886 ( .A1(n7528), .A2(n7527), .A3(n7526), .ZN(n13018) );
  XNOR2_X1 U8887 ( .A(n7612), .B(n7610), .ZN(n9945) );
  NAND2_X1 U8888 ( .A1(n8417), .A2(n8416), .ZN(n11854) );
  INV_X1 U8889 ( .A(n14568), .ZN(n7056) );
  AND2_X1 U8890 ( .A1(n7187), .A2(n7190), .ZN(n6548) );
  INV_X1 U8891 ( .A(n13608), .ZN(n6977) );
  AND2_X1 U8892 ( .A1(n7381), .A2(n8259), .ZN(n6549) );
  AND4_X1 U8893 ( .A1(n13286), .A2(n7194), .A3(n7193), .A4(n7178), .ZN(n6550)
         );
  INV_X1 U8894 ( .A(n13566), .ZN(n6973) );
  INV_X1 U8895 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13003) );
  AND2_X1 U8896 ( .A1(n12915), .A2(n12102), .ZN(n6551) );
  AND2_X1 U8897 ( .A1(n6950), .A2(n13256), .ZN(n13553) );
  INV_X1 U8898 ( .A(n12256), .ZN(n7407) );
  AND2_X1 U8899 ( .A1(n11849), .A2(n11535), .ZN(n6552) );
  INV_X1 U8900 ( .A(n11953), .ZN(n6834) );
  NOR2_X1 U8901 ( .A1(n13543), .A2(n13226), .ZN(n6553) );
  OR2_X1 U8902 ( .A1(n13223), .A2(n13282), .ZN(n6554) );
  INV_X1 U8903 ( .A(n8085), .ZN(n7305) );
  INV_X1 U8904 ( .A(n11856), .ZN(n7370) );
  NAND2_X1 U8905 ( .A1(n12968), .A2(n12592), .ZN(n6555) );
  NOR2_X1 U8906 ( .A1(n14095), .A2(n14087), .ZN(n14057) );
  AND2_X1 U8907 ( .A1(n7170), .A2(n13236), .ZN(n6556) );
  OR2_X1 U8908 ( .A1(n11084), .A2(n8915), .ZN(n6557) );
  AND2_X1 U8909 ( .A1(n11003), .A2(n13146), .ZN(n6558) );
  AND3_X1 U8910 ( .A1(n6799), .A2(n6798), .A3(n6797), .ZN(n6559) );
  INV_X1 U8911 ( .A(n7402), .ZN(n7401) );
  OAI22_X1 U8912 ( .A1(n12669), .A2(n7403), .B1(n12935), .B2(n12403), .ZN(
        n7402) );
  NAND2_X1 U8913 ( .A1(n8064), .A2(n8063), .ZN(n13572) );
  NOR2_X1 U8914 ( .A1(n11886), .A2(n11961), .ZN(n6560) );
  NAND2_X1 U8915 ( .A1(n6987), .A2(n7430), .ZN(n8827) );
  NAND2_X1 U8916 ( .A1(n8314), .A2(n8250), .ZN(n8332) );
  AND2_X1 U8917 ( .A1(n11725), .A2(n13095), .ZN(n6561) );
  OR2_X1 U8918 ( .A1(n14433), .A2(n9851), .ZN(n6562) );
  INV_X1 U8919 ( .A(n8117), .ZN(n6684) );
  NOR2_X1 U8920 ( .A1(n14040), .A2(n14042), .ZN(n6563) );
  AND2_X1 U8921 ( .A1(n7437), .A2(n12112), .ZN(n6564) );
  NAND2_X1 U8922 ( .A1(n14568), .A2(n7054), .ZN(n7053) );
  INV_X1 U8923 ( .A(n7053), .ZN(n7051) );
  INV_X1 U8924 ( .A(n14058), .ZN(n8653) );
  NAND2_X1 U8925 ( .A1(n8602), .A2(n8601), .ZN(n14058) );
  NOR2_X1 U8926 ( .A1(n13247), .A2(n13248), .ZN(n6565) );
  NAND2_X1 U8927 ( .A1(n6561), .A2(n6466), .ZN(n6566) );
  INV_X1 U8928 ( .A(n7246), .ZN(n7245) );
  NAND2_X1 U8929 ( .A1(n7247), .A2(n13266), .ZN(n7246) );
  NOR2_X1 U8930 ( .A1(n14567), .A2(n14568), .ZN(n6567) );
  INV_X1 U8931 ( .A(n10795), .ZN(n7165) );
  NAND2_X1 U8932 ( .A1(n6627), .A2(n7071), .ZN(n7070) );
  AND2_X1 U8933 ( .A1(n8116), .A2(n8115), .ZN(n13308) );
  INV_X1 U8934 ( .A(n13308), .ZN(n13555) );
  INV_X1 U8935 ( .A(n11866), .ZN(n13760) );
  INV_X1 U8936 ( .A(n13383), .ZN(n13585) );
  INV_X1 U8937 ( .A(n11869), .ZN(n7378) );
  INV_X1 U8938 ( .A(n12013), .ZN(n14081) );
  INV_X1 U8939 ( .A(n7046), .ZN(n7045) );
  OAI21_X1 U8940 ( .B1(n7051), .B2(n7055), .A(n14571), .ZN(n7046) );
  AND2_X1 U8941 ( .A1(n8147), .A2(n8146), .ZN(n13550) );
  INV_X1 U8942 ( .A(n13550), .ZN(n13293) );
  NOR2_X1 U8943 ( .A1(n12133), .A2(n12132), .ZN(n6568) );
  AND2_X1 U8944 ( .A1(n6839), .A2(n6838), .ZN(n6569) );
  INV_X1 U8945 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7038) );
  NOR2_X1 U8946 ( .A1(n14400), .A2(n9850), .ZN(n6570) );
  AOI21_X1 U8947 ( .B1(n12308), .B2(n14669), .A(n12310), .ZN(n6971) );
  AND2_X1 U8948 ( .A1(n6543), .A2(n10733), .ZN(n6571) );
  OR3_X1 U8949 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6572) );
  OR2_X1 U8950 ( .A1(n10795), .A2(n6764), .ZN(n6573) );
  AND2_X1 U8951 ( .A1(n6539), .A2(n9784), .ZN(n6574) );
  NAND2_X1 U8952 ( .A1(n14057), .A2(n6964), .ZN(n6965) );
  INV_X1 U8953 ( .A(n6739), .ZN(n11520) );
  AND2_X1 U8954 ( .A1(n13566), .A2(n13346), .ZN(n6575) );
  AND2_X1 U8955 ( .A1(n7010), .A2(n7008), .ZN(n6576) );
  INV_X1 U8956 ( .A(n6852), .ZN(n8643) );
  NOR2_X1 U8957 ( .A1(n14213), .A2(n14233), .ZN(n6577) );
  NOR2_X1 U8958 ( .A1(n13383), .A2(n13280), .ZN(n6578) );
  NOR2_X1 U8959 ( .A1(n11616), .A2(n11615), .ZN(n6579) );
  INV_X1 U8960 ( .A(n8687), .ZN(n7096) );
  INV_X1 U8961 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U8962 ( .A1(n13780), .A2(n11613), .ZN(n6580) );
  AND2_X1 U8963 ( .A1(n7395), .A2(n6555), .ZN(n7392) );
  AND2_X1 U8964 ( .A1(n13451), .A2(n13267), .ZN(n6581) );
  INV_X1 U8965 ( .A(n13281), .ZN(n6897) );
  AND2_X1 U8966 ( .A1(n13578), .A2(n13347), .ZN(n13281) );
  INV_X1 U8967 ( .A(n9704), .ZN(n7410) );
  AND2_X1 U8968 ( .A1(n12691), .A2(n12587), .ZN(n9704) );
  NAND2_X1 U8969 ( .A1(n8862), .A2(n10783), .ZN(n9754) );
  INV_X1 U8970 ( .A(n7190), .ZN(n7188) );
  AND2_X1 U8971 ( .A1(n7350), .A2(n7355), .ZN(n6582) );
  NAND2_X1 U8972 ( .A1(n13602), .A2(n13240), .ZN(n6583) );
  NAND3_X1 U8973 ( .A1(n7109), .A2(n7488), .A3(n7110), .ZN(n6584) );
  AND2_X1 U8974 ( .A1(n6773), .A2(n6987), .ZN(n8823) );
  NAND2_X1 U8975 ( .A1(n7677), .A2(n7464), .ZN(n6585) );
  INV_X1 U8976 ( .A(n6753), .ZN(n6752) );
  NAND2_X1 U8977 ( .A1(n7322), .A2(n6754), .ZN(n6753) );
  AND2_X1 U8978 ( .A1(n7700), .A2(SI_8_), .ZN(n6586) );
  AND2_X1 U8979 ( .A1(n12598), .A2(n9688), .ZN(n6587) );
  OR2_X1 U8980 ( .A1(n13269), .A2(n7244), .ZN(n6588) );
  AND2_X1 U8981 ( .A1(n13087), .A2(n11707), .ZN(n6589) );
  INV_X1 U8982 ( .A(n6898), .ZN(n13582) );
  NAND2_X1 U8983 ( .A1(n6900), .A2(n6511), .ZN(n6898) );
  AND2_X1 U8984 ( .A1(n11568), .A2(n11567), .ZN(n6590) );
  NAND2_X1 U8985 ( .A1(n9072), .A2(n12453), .ZN(n6591) );
  INV_X1 U8986 ( .A(n7345), .ZN(n7344) );
  NAND2_X1 U8987 ( .A1(n8638), .A2(n7346), .ZN(n7345) );
  INV_X1 U8988 ( .A(n12663), .ZN(n12669) );
  NAND2_X1 U8989 ( .A1(n12257), .A2(n6894), .ZN(n12663) );
  AND2_X1 U8990 ( .A1(n6741), .A2(n6740), .ZN(n6592) );
  NAND2_X1 U8991 ( .A1(n8533), .A2(n8256), .ZN(n8698) );
  INV_X1 U8992 ( .A(n6867), .ZN(n6866) );
  OAI21_X1 U8993 ( .B1(n12266), .B2(n6868), .A(n11753), .ZN(n6867) );
  AND2_X1 U8994 ( .A1(n11855), .A2(n7370), .ZN(n6593) );
  OR2_X1 U8995 ( .A1(n7370), .A2(n11855), .ZN(n6594) );
  NOR2_X1 U8996 ( .A1(n6977), .A2(n13270), .ZN(n6595) );
  NOR2_X1 U8997 ( .A1(n13319), .A2(n13249), .ZN(n6596) );
  INV_X1 U8998 ( .A(n11950), .ZN(n6847) );
  NAND2_X1 U8999 ( .A1(n9699), .A2(n7391), .ZN(n6597) );
  NAND2_X1 U9000 ( .A1(n7095), .A2(n14099), .ZN(n6598) );
  XNOR2_X1 U9001 ( .A(n8644), .B(n8638), .ZN(n11120) );
  OR2_X1 U9002 ( .A1(n9454), .A2(n9453), .ZN(n6599) );
  AND2_X1 U9003 ( .A1(n7441), .A2(n14189), .ZN(n6600) );
  NAND2_X1 U9004 ( .A1(n13250), .A2(n8186), .ZN(n13298) );
  INV_X1 U9005 ( .A(n13298), .ZN(n7178) );
  AND2_X1 U9006 ( .A1(n11779), .A2(n7399), .ZN(n6601) );
  INV_X1 U9007 ( .A(n14033), .ZN(n13700) );
  NAND2_X1 U9008 ( .A1(n8623), .A2(n8622), .ZN(n14033) );
  AND2_X1 U9009 ( .A1(n6974), .A2(n6973), .ZN(n6602) );
  AND2_X1 U9010 ( .A1(n12018), .A2(n7141), .ZN(n6603) );
  NAND2_X1 U9011 ( .A1(n9228), .A2(n9227), .ZN(n12873) );
  AND2_X1 U9012 ( .A1(n7634), .A2(SI_5_), .ZN(n6604) );
  AND2_X1 U9013 ( .A1(n10996), .A2(n10994), .ZN(n6605) );
  AND2_X1 U9014 ( .A1(n13393), .A2(n13279), .ZN(n6606) );
  AND2_X1 U9015 ( .A1(n6540), .A2(n12524), .ZN(n6607) );
  AND2_X1 U9016 ( .A1(n6694), .A2(n6693), .ZN(n6608) );
  OR2_X1 U9017 ( .A1(n8047), .A2(n8045), .ZN(n6609) );
  AND2_X1 U9018 ( .A1(n6991), .A2(n8796), .ZN(n6610) );
  NOR2_X1 U9019 ( .A1(n11444), .A2(n9042), .ZN(n6611) );
  OR2_X1 U9020 ( .A1(n8006), .A2(n8008), .ZN(n6612) );
  OR2_X1 U9021 ( .A1(n7958), .A2(n7960), .ZN(n6613) );
  OR2_X1 U9022 ( .A1(n11848), .A2(n11846), .ZN(n6614) );
  AND2_X1 U9023 ( .A1(n6549), .A2(n7380), .ZN(n6615) );
  INV_X1 U9024 ( .A(n10480), .ZN(n7158) );
  AND2_X1 U9025 ( .A1(n7342), .A2(n7347), .ZN(n6616) );
  OR2_X1 U9026 ( .A1(n8084), .A2(n7305), .ZN(n6617) );
  AND2_X1 U9027 ( .A1(n6756), .A2(n8638), .ZN(n6618) );
  INV_X1 U9028 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8234) );
  OR2_X1 U9029 ( .A1(n7663), .A2(n7298), .ZN(n6619) );
  AND2_X1 U9030 ( .A1(n6972), .A2(n6971), .ZN(n6620) );
  INV_X1 U9031 ( .A(n7324), .ZN(n7323) );
  NAND2_X1 U9032 ( .A1(n13813), .A2(n7325), .ZN(n7324) );
  INV_X1 U9033 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U9034 ( .A1(n7707), .A2(n7286), .ZN(n6621) );
  NAND2_X1 U9035 ( .A1(n7756), .A2(n7289), .ZN(n6622) );
  NAND2_X1 U9036 ( .A1(n7809), .A2(n7292), .ZN(n6623) );
  OR2_X1 U9037 ( .A1(n13555), .A2(n11740), .ZN(n13250) );
  OR2_X1 U9038 ( .A1(n6841), .A2(n6847), .ZN(n6837) );
  AND2_X1 U9039 ( .A1(n11942), .A2(n11940), .ZN(n6624) );
  INV_X1 U9040 ( .A(n6733), .ZN(n6732) );
  NAND2_X1 U9041 ( .A1(n6736), .A2(n6734), .ZN(n6733) );
  INV_X1 U9042 ( .A(n7272), .ZN(n7271) );
  NAND2_X1 U9043 ( .A1(n7273), .A2(n8989), .ZN(n7272) );
  INV_X1 U9044 ( .A(n11730), .ZN(n11708) );
  AND4_X1 U9045 ( .A1(n9237), .A2(n9236), .A3(n9235), .A4(n9234), .ZN(n12524)
         );
  AND2_X1 U9046 ( .A1(n13256), .A2(n13500), .ZN(n6625) );
  NAND2_X1 U9047 ( .A1(n14975), .A2(n9004), .ZN(n11442) );
  NAND2_X1 U9048 ( .A1(n11551), .A2(n11550), .ZN(n13749) );
  OR2_X1 U9049 ( .A1(n13700), .A2(n14348), .ZN(n6626) );
  NAND2_X1 U9050 ( .A1(n7426), .A2(n9687), .ZN(n12832) );
  NAND2_X1 U9051 ( .A1(n13751), .A2(n6530), .ZN(n13812) );
  INV_X1 U9052 ( .A(n14301), .ZN(n6960) );
  INV_X1 U9053 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n6775) );
  INV_X1 U9054 ( .A(n13761), .ZN(n7315) );
  INV_X1 U9055 ( .A(n11646), .ZN(n7331) );
  NAND2_X1 U9056 ( .A1(n7452), .A2(n13508), .ZN(n13507) );
  AND2_X1 U9057 ( .A1(n14188), .A2(n8680), .ZN(n6627) );
  NAND2_X1 U9058 ( .A1(n13507), .A2(n13262), .ZN(n13493) );
  NAND2_X1 U9059 ( .A1(n8932), .A2(n7430), .ZN(n9085) );
  AND2_X1 U9060 ( .A1(n9176), .A2(n12591), .ZN(n6628) );
  NOR2_X1 U9061 ( .A1(n13437), .A2(n13602), .ZN(n13410) );
  INV_X1 U9062 ( .A(n6978), .ZN(n13447) );
  INV_X1 U9063 ( .A(n8324), .ZN(n8363) );
  OR2_X1 U9064 ( .A1(n13191), .A2(n14953), .ZN(n6629) );
  AND2_X1 U9065 ( .A1(n7086), .A2(n7084), .ZN(n6630) );
  INV_X1 U9066 ( .A(SI_13_), .ZN(n10007) );
  OR2_X1 U9067 ( .A1(n13197), .A2(n14958), .ZN(n6631) );
  INV_X1 U9068 ( .A(n7085), .ZN(n7084) );
  NOR2_X1 U9069 ( .A1(n6934), .A2(n6931), .ZN(n6632) );
  INV_X1 U9070 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10224) );
  INV_X1 U9071 ( .A(n7930), .ZN(n7191) );
  AND2_X1 U9072 ( .A1(n7864), .A2(n10088), .ZN(n6633) );
  INV_X1 U9073 ( .A(n7260), .ZN(n7259) );
  OAI21_X1 U9074 ( .B1(n9162), .B2(n7261), .A(n9177), .ZN(n7260) );
  INV_X1 U9075 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9942) );
  OR2_X1 U9076 ( .A1(n12931), .A2(n12911), .ZN(n6634) );
  NOR2_X1 U9077 ( .A1(n13065), .A2(n13510), .ZN(n6635) );
  NOR2_X1 U9078 ( .A1(n7994), .A2(n7998), .ZN(n6636) );
  OR2_X1 U9079 ( .A1(n6778), .A2(n6777), .ZN(n6637) );
  AND2_X1 U9080 ( .A1(n6525), .A2(n6783), .ZN(n6638) );
  NAND2_X2 U9081 ( .A1(n10264), .A2(n13466), .ZN(n13527) );
  INV_X1 U9082 ( .A(n9885), .ZN(n9883) );
  INV_X1 U9083 ( .A(n11004), .ZN(n6796) );
  NAND2_X1 U9084 ( .A1(n8640), .A2(n8713), .ZN(n11791) );
  NOR2_X1 U9085 ( .A1(n7484), .A2(n7487), .ZN(n7110) );
  AND2_X1 U9086 ( .A1(n15205), .A2(n15167), .ZN(n12901) );
  AOI21_X1 U9087 ( .B1(n11362), .B2(n9683), .A(n6544), .ZN(n11425) );
  INV_X1 U9088 ( .A(n13641), .ZN(n6981) );
  OR2_X1 U9089 ( .A1(n14944), .A2(n6951), .ZN(n6639) );
  OR2_X1 U9090 ( .A1(n11145), .A2(n14668), .ZN(n11190) );
  NAND2_X1 U9091 ( .A1(n7237), .A2(n10596), .ZN(n13532) );
  INV_X1 U9092 ( .A(n6984), .ZN(n10636) );
  AND2_X1 U9093 ( .A1(n7076), .A2(n7078), .ZN(n6640) );
  AOI21_X1 U9094 ( .B1(n12143), .B2(n15109), .A(n9674), .ZN(n10951) );
  AND2_X1 U9095 ( .A1(n6780), .A2(n6778), .ZN(n6641) );
  AND2_X1 U9096 ( .A1(n8787), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6642) );
  AND2_X1 U9097 ( .A1(n8042), .A2(n11137), .ZN(n6643) );
  AND2_X1 U9098 ( .A1(n6735), .A2(n6732), .ZN(n6644) );
  AND2_X1 U9099 ( .A1(n7203), .A2(n8056), .ZN(n6645) );
  NAND2_X1 U9100 ( .A1(n9730), .A2(n12134), .ZN(n12804) );
  INV_X1 U9101 ( .A(n11849), .ZN(n6970) );
  INV_X1 U9102 ( .A(SI_22_), .ZN(n7211) );
  NAND2_X1 U9103 ( .A1(n6858), .A2(n6857), .ZN(n11793) );
  NAND2_X1 U9104 ( .A1(n10283), .A2(n12370), .ZN(n14672) );
  INV_X1 U9105 ( .A(n6469), .ZN(n13216) );
  NAND2_X1 U9106 ( .A1(n7681), .A2(n7680), .ZN(n12070) );
  INV_X1 U9107 ( .A(n12070), .ZN(n6983) );
  INV_X1 U9108 ( .A(n10503), .ZN(n6980) );
  OR2_X1 U9109 ( .A1(n14856), .A2(n13206), .ZN(n6646) );
  NAND2_X1 U9110 ( .A1(n9884), .A2(n10089), .ZN(n6647) );
  AND2_X1 U9111 ( .A1(n7128), .A2(n7127), .ZN(n6648) );
  NAND2_X1 U9112 ( .A1(n9903), .A2(n15003), .ZN(n6649) );
  AND2_X1 U9113 ( .A1(n11793), .A2(n11792), .ZN(n6650) );
  INV_X1 U9114 ( .A(n14433), .ZN(n10093) );
  INV_X1 U9115 ( .A(SI_26_), .ZN(n11349) );
  AND2_X1 U9116 ( .A1(n6647), .A2(n6529), .ZN(n6651) );
  XNOR2_X1 U9117 ( .A(n8819), .B(P3_IR_REG_26__SCAN_IN), .ZN(n11346) );
  INV_X1 U9118 ( .A(n11346), .ZN(n6664) );
  INV_X1 U9119 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6887) );
  NAND2_X2 U9120 ( .A1(n6492), .A2(P3_U3151), .ZN(n13004) );
  NAND2_X1 U9121 ( .A1(n9827), .A2(n6654), .ZN(n11017) );
  NAND2_X1 U9122 ( .A1(n6656), .A2(n6655), .ZN(n6654) );
  INV_X1 U9123 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U9124 ( .A1(n9836), .A2(n11057), .ZN(n9837) );
  NAND2_X1 U9125 ( .A1(n8885), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U9126 ( .A1(n6992), .A2(n6993), .ZN(n8885) );
  NOR2_X1 U9127 ( .A1(n15031), .A2(n12839), .ZN(n15030) );
  AOI22_X2 U9128 ( .A1(n13389), .A2(n7241), .B1(n13243), .B2(n13278), .ZN(
        n13374) );
  NAND4_X1 U9129 ( .A1(n7490), .A2(n7489), .A3(n7109), .A4(n7488), .ZN(n8223)
         );
  AND3_X2 U9130 ( .A1(n7462), .A2(n7548), .A3(n7461), .ZN(n7109) );
  NAND2_X1 U9131 ( .A1(n10797), .A2(n10798), .ZN(n10875) );
  NAND2_X1 U9132 ( .A1(n7176), .A2(n7175), .ZN(n13299) );
  INV_X1 U9133 ( .A(n7248), .ZN(n7550) );
  NAND2_X1 U9134 ( .A1(n10756), .A2(n7164), .ZN(n7163) );
  NAND2_X1 U9135 ( .A1(n10981), .A2(n10980), .ZN(n7172) );
  INV_X4 U9136 ( .A(n7161), .ZN(n7572) );
  AOI21_X1 U9137 ( .B1(n7824), .B2(n7825), .A(n6657), .ZN(n7453) );
  MUX2_X1 U9138 ( .A(n13157), .B(n8170), .S(n10354), .Z(n7519) );
  NAND2_X1 U9139 ( .A1(n7303), .A2(n7304), .ZN(n8118) );
  NAND2_X1 U9140 ( .A1(n7559), .A2(n7558), .ZN(n7577) );
  OAI22_X1 U9141 ( .A1(n7919), .A2(n7282), .B1(n7920), .B2(n7283), .ZN(n7940)
         );
  NAND2_X1 U9142 ( .A1(n7521), .A2(n7520), .ZN(n7535) );
  OAI21_X1 U9143 ( .B1(n7824), .B2(n7825), .A(n7890), .ZN(n7899) );
  OAI21_X2 U9144 ( .B1(n11424), .B2(n9763), .A(n12190), .ZN(n11459) );
  NAND2_X1 U9145 ( .A1(n8813), .A2(n7432), .ZN(n6663) );
  XNOR2_X1 U9146 ( .A(n7525), .B(P2_IR_REG_1__SCAN_IN), .ZN(n13162) );
  NAND2_X1 U9147 ( .A1(n8822), .A2(n8821), .ZN(n9318) );
  NAND2_X4 U9148 ( .A1(n8833), .A2(n8832), .ZN(n10776) );
  NAND2_X1 U9149 ( .A1(n11174), .A2(n8968), .ZN(n14965) );
  NAND2_X1 U9150 ( .A1(n7206), .A2(SI_22_), .ZN(n7207) );
  OAI21_X1 U9151 ( .B1(n12476), .B2(n9144), .A(n9143), .ZN(n12485) );
  NAND2_X1 U9152 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  NAND2_X1 U9153 ( .A1(n9196), .A2(n8783), .ZN(n9209) );
  NAND2_X1 U9154 ( .A1(n9084), .A2(n7279), .ZN(n9093) );
  INV_X1 U9155 ( .A(n9082), .ZN(n6869) );
  INV_X1 U9156 ( .A(n9194), .ZN(n6888) );
  NAND2_X1 U9157 ( .A1(n6697), .A2(n14684), .ZN(n6686) );
  NAND2_X1 U9158 ( .A1(n7258), .A2(n7256), .ZN(n8781) );
  NAND2_X1 U9159 ( .A1(n6859), .A2(n8747), .ZN(n8938) );
  NAND2_X1 U9160 ( .A1(n8905), .A2(n8745), .ZN(n8923) );
  NAND2_X1 U9161 ( .A1(n9011), .A2(n6878), .ZN(n6877) );
  NAND2_X1 U9162 ( .A1(n6877), .A2(n6875), .ZN(n9057) );
  OAI211_X1 U9163 ( .C1(n6886), .C2(n12296), .A(n6882), .B(n6710), .ZN(
        P3_U3296) );
  AND2_X2 U9164 ( .A1(n10618), .A2(n8880), .ZN(n12138) );
  NAND2_X2 U9165 ( .A1(n6717), .A2(n6716), .ZN(n12744) );
  AOI21_X2 U9166 ( .B1(n9768), .B2(n12209), .A(n9767), .ZN(n12787) );
  NAND2_X1 U9167 ( .A1(n12668), .A2(n12667), .ZN(n12864) );
  NAND2_X1 U9168 ( .A1(n12825), .A2(n12824), .ZN(n12823) );
  NAND2_X1 U9169 ( .A1(n11303), .A2(n11305), .ZN(n11304) );
  NAND2_X1 U9170 ( .A1(n7439), .A2(n12720), .ZN(n12716) );
  MUX2_X1 U9171 ( .A(n12861), .B(n12929), .S(n15205), .Z(n12862) );
  NAND2_X1 U9172 ( .A1(n12787), .A2(n9769), .ZN(n12786) );
  AOI21_X1 U9173 ( .B1(n12744), .B2(n9774), .A(n6721), .ZN(n7439) );
  NAND2_X1 U9174 ( .A1(n10950), .A2(n10948), .ZN(n10949) );
  NOR2_X1 U9175 ( .A1(n11777), .A2(n12261), .ZN(n11778) );
  NAND2_X2 U9176 ( .A1(n6673), .A2(n8890), .ZN(n15106) );
  AOI21_X1 U9177 ( .B1(n12860), .B2(n15175), .A(n12468), .ZN(n11783) );
  NAND2_X1 U9178 ( .A1(n6675), .A2(n7294), .ZN(n8067) );
  NAND3_X1 U9179 ( .A1(n8030), .A2(n8029), .A3(n6609), .ZN(n6675) );
  NAND2_X1 U9180 ( .A1(n6676), .A2(n7295), .ZN(n8025) );
  NAND3_X1 U9181 ( .A1(n7982), .A2(n7981), .A3(n6612), .ZN(n6676) );
  NAND2_X1 U9182 ( .A1(n6677), .A2(n7293), .ZN(n7977) );
  NAND3_X1 U9183 ( .A1(n7945), .A2(n7944), .A3(n6613), .ZN(n6677) );
  INV_X1 U9184 ( .A(n12315), .ZN(n6697) );
  NAND2_X1 U9185 ( .A1(n7612), .A2(n7611), .ZN(n7615) );
  INV_X1 U9186 ( .A(n6682), .ZN(n8151) );
  NOR2_X1 U9187 ( .A1(n8872), .A2(n8871), .ZN(n8880) );
  NAND2_X2 U9188 ( .A1(n8878), .A2(n8877), .ZN(n10618) );
  NAND2_X1 U9189 ( .A1(n12716), .A2(n9775), .ZN(n12706) );
  NAND2_X1 U9190 ( .A1(n12838), .A2(n9766), .ZN(n12837) );
  NAND2_X1 U9191 ( .A1(n12934), .A2(n6678), .ZN(P3_U3451) );
  NAND2_X1 U9192 ( .A1(n12866), .A2(n6679), .ZN(P3_U3483) );
  INV_X1 U9193 ( .A(n7918), .ZN(n7283) );
  NOR2_X1 U9194 ( .A1(n14395), .A2(n14394), .ZN(n14393) );
  XNOR2_X1 U9195 ( .A(n9464), .B(n9465), .ZN(n14395) );
  NAND2_X1 U9196 ( .A1(n14565), .A2(n14566), .ZN(n14562) );
  NAND2_X1 U9197 ( .A1(n14371), .A2(n14372), .ZN(n14370) );
  NAND2_X1 U9198 ( .A1(n14556), .A2(n14555), .ZN(n14554) );
  XOR2_X2 U9199 ( .A(n9451), .B(P2_ADDR_REG_6__SCAN_IN), .Z(n14386) );
  XNOR2_X1 U9200 ( .A(n9443), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U9201 ( .A1(n7285), .A2(n7284), .ZN(n7731) );
  NAND2_X1 U9202 ( .A1(n7288), .A2(n7287), .ZN(n7776) );
  NAND2_X1 U9203 ( .A1(n7297), .A2(n6619), .ZN(n7684) );
  NAND2_X1 U9204 ( .A1(n7301), .A2(n7300), .ZN(n7640) );
  NAND2_X1 U9205 ( .A1(n14068), .A2(n8611), .ZN(n14041) );
  INV_X1 U9206 ( .A(n9382), .ZN(P1_U3523) );
  NAND2_X1 U9207 ( .A1(n7196), .A2(n7198), .ZN(n7720) );
  NAND3_X1 U9208 ( .A1(n6686), .A2(n12318), .A3(n6620), .ZN(n9365) );
  OAI21_X1 U9209 ( .B1(n9821), .B2(n14695), .A(n9825), .ZN(P1_U3556) );
  NAND2_X1 U9210 ( .A1(n9374), .A2(n7141), .ZN(n6687) );
  AOI21_X2 U9211 ( .B1(n8696), .B2(n14676), .A(n8695), .ZN(n12318) );
  AOI21_X1 U9212 ( .B1(n9368), .B2(n12014), .A(n7067), .ZN(n9353) );
  NAND3_X1 U9213 ( .A1(n12061), .A2(n6805), .A3(n12066), .ZN(n6803) );
  NAND2_X1 U9214 ( .A1(n11659), .A2(n11658), .ZN(n12057) );
  NAND2_X2 U9215 ( .A1(n8677), .A2(n12008), .ZN(n14505) );
  INV_X1 U9216 ( .A(n8003), .ZN(n7206) );
  NOR3_X1 U9217 ( .A1(n12030), .A2(n12029), .A3(n12028), .ZN(n12035) );
  NAND2_X1 U9218 ( .A1(n13469), .A2(n13221), .ZN(n13471) );
  NAND2_X1 U9219 ( .A1(n10763), .A2(n14928), .ZN(n10802) );
  NAND2_X1 U9220 ( .A1(n10377), .A2(n10431), .ZN(n10503) );
  NAND3_X1 U9221 ( .A1(n13289), .A2(n6692), .A3(n13510), .ZN(n13549) );
  XNOR2_X1 U9222 ( .A(n9845), .B(n9914), .ZN(n15064) );
  OAI21_X1 U9223 ( .B1(n12283), .B2(n12282), .A(n12281), .ZN(n7278) );
  INV_X1 U9224 ( .A(n13339), .ZN(n6913) );
  OAI21_X1 U9225 ( .B1(n6918), .B2(n6922), .A(n6919), .ZN(n7792) );
  OAI22_X1 U9226 ( .A1(n13318), .A2(n13317), .B1(n13284), .B2(n13319), .ZN(
        n13297) );
  NAND2_X1 U9227 ( .A1(n6896), .A2(n6895), .ZN(n13349) );
  NAND2_X1 U9228 ( .A1(n6715), .A2(n6712), .ZN(P3_U3452) );
  OR2_X1 U9229 ( .A1(n12929), .A2(n15191), .ZN(n6715) );
  INV_X1 U9230 ( .A(n12743), .ZN(n6717) );
  AND3_X2 U9231 ( .A1(n6988), .A2(n7450), .A3(n6610), .ZN(n6987) );
  NAND2_X1 U9232 ( .A1(n12862), .A2(n6634), .ZN(P3_U3484) );
  INV_X1 U9233 ( .A(n12696), .ZN(n6719) );
  NAND2_X1 U9234 ( .A1(n6916), .A2(n7657), .ZN(n7674) );
  NAND2_X1 U9235 ( .A1(n12140), .A2(n12138), .ZN(n9755) );
  NAND2_X2 U9236 ( .A1(n11774), .A2(n11773), .ZN(n12696) );
  OAI21_X1 U9237 ( .B1(n6770), .B2(n15076), .A(n6769), .ZN(n6768) );
  INV_X1 U9238 ( .A(n6768), .ZN(n6767) );
  INV_X1 U9239 ( .A(n8885), .ZN(n8884) );
  OAI21_X1 U9240 ( .B1(n12571), .B2(n12568), .A(n12567), .ZN(n12476) );
  NAND2_X1 U9241 ( .A1(n9107), .A2(n9106), .ZN(n12393) );
  INV_X2 U9242 ( .A(n10776), .ZN(n8926) );
  AND2_X2 U9243 ( .A1(n12105), .A2(n10579), .ZN(n12292) );
  NAND2_X1 U9244 ( .A1(n9433), .A2(n9432), .ZN(n6724) );
  NAND2_X2 U9245 ( .A1(n14564), .A2(n14562), .ZN(n14567) );
  NOR2_X1 U9246 ( .A1(n14390), .A2(n9463), .ZN(n9464) );
  NAND2_X1 U9247 ( .A1(n9434), .A2(n9383), .ZN(n9384) );
  NOR2_X2 U9248 ( .A1(n14386), .A2(n14385), .ZN(n14384) );
  NAND2_X1 U9249 ( .A1(n14370), .A2(n7036), .ZN(n7035) );
  XNOR2_X1 U9250 ( .A(n7035), .B(n7034), .ZN(SUB_1596_U4) );
  NAND2_X1 U9251 ( .A1(n6726), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7511) );
  NAND3_X1 U9252 ( .A1(n14018), .A2(n7505), .A3(n7506), .ZN(n6726) );
  INV_X1 U9253 ( .A(n7074), .ZN(n7073) );
  AOI21_X2 U9254 ( .B1(n14118), .B2(n7091), .A(n7090), .ZN(n14080) );
  NAND2_X1 U9255 ( .A1(n14148), .A2(n8682), .ZN(n14133) );
  NAND2_X1 U9256 ( .A1(n8676), .A2(n8675), .ZN(n11507) );
  NAND2_X1 U9257 ( .A1(n11293), .A2(n8669), .ZN(n11350) );
  OAI21_X2 U9258 ( .B1(n14224), .B2(n7082), .A(n7081), .ZN(n14188) );
  NAND2_X1 U9259 ( .A1(n7058), .A2(n8671), .ZN(n11371) );
  NAND2_X1 U9260 ( .A1(n9365), .A2(n14698), .ZN(n9367) );
  INV_X1 U9261 ( .A(n11295), .ZN(n8668) );
  OAI21_X2 U9262 ( .B1(n14061), .B2(n8689), .A(n7068), .ZN(n9368) );
  NOR2_X1 U9263 ( .A1(n11033), .A2(n8971), .ZN(n11032) );
  XNOR2_X1 U9264 ( .A(n9839), .B(n9977), .ZN(n11033) );
  NAND2_X1 U9265 ( .A1(n9833), .A2(n6727), .ZN(n11124) );
  NAND2_X1 U9266 ( .A1(n9834), .A2(n9891), .ZN(n9833) );
  OAI21_X1 U9267 ( .B1(n12629), .B2(n15102), .A(n6767), .ZN(P3_U3201) );
  NOR2_X1 U9268 ( .A1(n14999), .A2(n9016), .ZN(n14998) );
  NOR2_X1 U9269 ( .A1(n10912), .A2(n10911), .ZN(n10910) );
  NOR2_X1 U9270 ( .A1(n15015), .A2(n15014), .ZN(n15013) );
  XNOR2_X1 U9271 ( .A(n9851), .B(n14433), .ZN(n14442) );
  NAND2_X1 U9272 ( .A1(n13716), .A2(n7314), .ZN(n7310) );
  NAND2_X1 U9273 ( .A1(n12322), .A2(n13712), .ZN(n6728) );
  OAI21_X1 U9274 ( .B1(n11327), .B2(n6733), .A(n6729), .ZN(n6739) );
  NAND3_X1 U9275 ( .A1(n6744), .A2(n7327), .A3(n6742), .ZN(n13728) );
  NAND2_X1 U9276 ( .A1(n6746), .A2(n6743), .ZN(n6742) );
  INV_X1 U9277 ( .A(n11586), .ZN(n6743) );
  NAND2_X1 U9278 ( .A1(n6745), .A2(n6746), .ZN(n6744) );
  INV_X1 U9279 ( .A(n13853), .ZN(n6745) );
  NAND2_X2 U9280 ( .A1(n11793), .A2(n10273), .ZN(n12370) );
  NAND2_X1 U9281 ( .A1(n8533), .A2(n6618), .ZN(n8641) );
  NAND2_X1 U9282 ( .A1(n8533), .A2(n6756), .ZN(n6852) );
  INV_X1 U9283 ( .A(n13427), .ZN(n6760) );
  NAND2_X2 U9284 ( .A1(n13343), .A2(n6554), .ZN(n13329) );
  INV_X1 U9285 ( .A(n7610), .ZN(n7611) );
  MUX2_X1 U9286 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7547), .Z(n7613) );
  NOR2_X2 U9287 ( .A1(n6771), .A2(n6774), .ZN(n8813) );
  NAND2_X1 U9288 ( .A1(n6514), .A2(n6987), .ZN(n6771) );
  NAND4_X1 U9289 ( .A1(n6514), .A2(n6987), .A3(n6772), .A4(n7430), .ZN(n8818)
         );
  INV_X1 U9290 ( .A(n6774), .ZN(n6773) );
  NAND2_X1 U9291 ( .A1(n10913), .A2(n6638), .ZN(n6776) );
  NAND2_X1 U9292 ( .A1(n6776), .A2(n6637), .ZN(n15041) );
  NAND2_X1 U9293 ( .A1(n14414), .A2(n6651), .ZN(n6785) );
  NAND3_X1 U9294 ( .A1(n13071), .A2(n10402), .A3(n13078), .ZN(n13070) );
  XNOR2_X1 U9295 ( .A(n10408), .B(n10403), .ZN(n13078) );
  OAI21_X2 U9296 ( .B1(n14464), .B2(n6796), .A(n6793), .ZN(n11659) );
  AND2_X2 U9297 ( .A1(n6566), .A2(n6800), .ZN(n13063) );
  NAND4_X1 U9298 ( .A1(n6797), .A2(n6799), .A3(n6798), .A4(n6635), .ZN(n6800)
         );
  OR2_X1 U9299 ( .A1(n11725), .A2(n6466), .ZN(n6797) );
  NAND3_X1 U9300 ( .A1(n11725), .A2(n13095), .A3(n6466), .ZN(n6798) );
  INV_X1 U9301 ( .A(n6800), .ZN(n12039) );
  NOR2_X2 U9302 ( .A1(n13036), .A2(n13037), .ZN(n13119) );
  NAND2_X2 U9303 ( .A1(n13061), .A2(n6801), .ZN(n13036) );
  NAND2_X1 U9304 ( .A1(n6806), .A2(n12061), .ZN(n12072) );
  NAND2_X1 U9305 ( .A1(n13112), .A2(n11682), .ZN(n6807) );
  NAND2_X1 U9306 ( .A1(n6807), .A2(n6808), .ZN(n11709) );
  INV_X1 U9307 ( .A(n11919), .ZN(n6814) );
  NAND3_X1 U9308 ( .A1(n6816), .A2(n6817), .A3(n6600), .ZN(n6815) );
  NAND3_X1 U9309 ( .A1(n11884), .A2(n6818), .A3(n11885), .ZN(n6816) );
  NAND2_X1 U9310 ( .A1(n7362), .A2(n6819), .ZN(n6821) );
  INV_X1 U9311 ( .A(n11943), .ZN(n6823) );
  NAND2_X1 U9312 ( .A1(n6825), .A2(n6824), .ZN(n11930) );
  INV_X1 U9313 ( .A(n6833), .ZN(n6845) );
  NOR2_X1 U9314 ( .A1(n6837), .A2(n6833), .ZN(n6832) );
  NAND2_X1 U9315 ( .A1(n6837), .A2(n11953), .ZN(n6835) );
  INV_X1 U9316 ( .A(n6846), .ZN(n6844) );
  NAND2_X1 U9317 ( .A1(n11851), .A2(n6517), .ZN(n6849) );
  NAND3_X1 U9318 ( .A1(n11793), .A2(n11120), .A3(n11792), .ZN(n6853) );
  INV_X1 U9319 ( .A(n11791), .ZN(n6858) );
  MUX2_X1 U9320 ( .A(n11836), .B(n13882), .S(n11835), .Z(n7349) );
  NAND2_X1 U9321 ( .A1(n8938), .A2(n8937), .ZN(n8750) );
  NAND2_X1 U9322 ( .A1(n8923), .A2(n8922), .ZN(n6859) );
  XNOR2_X1 U9323 ( .A(n12106), .B(n12614), .ZN(n6883) );
  NAND2_X1 U9324 ( .A1(n6568), .A2(n12290), .ZN(n6882) );
  INV_X1 U9325 ( .A(n12291), .ZN(n6886) );
  NAND2_X1 U9326 ( .A1(n7252), .A2(n6891), .ZN(n6889) );
  NAND2_X1 U9327 ( .A1(n6889), .A2(n6890), .ZN(n7258) );
  OAI21_X1 U9328 ( .B1(n7250), .B2(n6893), .A(n8776), .ZN(n6892) );
  NAND2_X1 U9329 ( .A1(n9146), .A2(n9145), .ZN(n9148) );
  NAND2_X1 U9330 ( .A1(n7252), .A2(n7250), .ZN(n9146) );
  NAND2_X1 U9331 ( .A1(n13277), .A2(n6511), .ZN(n6896) );
  NAND2_X1 U9332 ( .A1(n13465), .A2(n6903), .ZN(n6902) );
  INV_X1 U9333 ( .A(n6910), .ZN(n6906) );
  NAND2_X1 U9334 ( .A1(n6906), .A2(n6905), .ZN(n6907) );
  NAND2_X1 U9335 ( .A1(n6909), .A2(n7227), .ZN(n11268) );
  XNOR2_X1 U9336 ( .A(n7589), .B(n7587), .ZN(n9943) );
  AOI21_X2 U9337 ( .B1(n13552), .B2(n14934), .A(n13551), .ZN(n13554) );
  NAND2_X1 U9338 ( .A1(n6915), .A2(n6914), .ZN(n7655) );
  AOI21_X1 U9339 ( .B1(n7632), .B2(n7195), .A(n6604), .ZN(n6914) );
  NAND3_X1 U9340 ( .A1(n7612), .A2(n7611), .A3(n7632), .ZN(n6915) );
  NAND2_X1 U9341 ( .A1(n7655), .A2(n7654), .ZN(n6916) );
  NAND2_X1 U9342 ( .A1(n6917), .A2(n6643), .ZN(n7201) );
  NAND2_X1 U9343 ( .A1(n6917), .A2(n8042), .ZN(n8057) );
  INV_X1 U9344 ( .A(n7723), .ZN(n6918) );
  NAND2_X1 U9345 ( .A1(n7819), .A2(n6938), .ZN(n6935) );
  NAND2_X1 U9346 ( .A1(n6935), .A2(n6936), .ZN(n7913) );
  NAND2_X1 U9347 ( .A1(n13252), .A2(n6945), .ZN(n6944) );
  NAND2_X1 U9348 ( .A1(n6944), .A2(n6942), .ZN(P2_U3496) );
  NAND2_X1 U9349 ( .A1(n6953), .A2(n7932), .ZN(n7955) );
  NAND2_X1 U9350 ( .A1(n8702), .A2(n6549), .ZN(n8265) );
  NOR2_X2 U9351 ( .A1(n14205), .A2(n14182), .ZN(n14185) );
  INV_X1 U9352 ( .A(n6965), .ZN(n14049) );
  INV_X1 U9353 ( .A(n11190), .ZN(n6966) );
  NAND2_X1 U9354 ( .A1(n6967), .A2(n6966), .ZN(n11391) );
  NOR2_X2 U9355 ( .A1(n10504), .A2(n14904), .ZN(n13535) );
  NOR2_X2 U9356 ( .A1(n10430), .A2(n10591), .ZN(n10431) );
  NAND2_X2 U9357 ( .A1(n7161), .A2(n9961), .ZN(n8169) );
  XNOR2_X2 U9358 ( .A(n7162), .B(n7516), .ZN(n10155) );
  XNOR2_X2 U9359 ( .A(n7513), .B(n7514), .ZN(n8240) );
  AND2_X2 U9360 ( .A1(n13321), .A2(n13308), .ZN(n13306) );
  INV_X2 U9361 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6992) );
  NAND3_X1 U9362 ( .A1(n8884), .A2(n7427), .A3(n8796), .ZN(n8933) );
  NAND2_X1 U9363 ( .A1(n12485), .A2(n6999), .ZN(n6996) );
  NAND2_X1 U9364 ( .A1(n6996), .A2(n6997), .ZN(n12418) );
  NAND2_X1 U9365 ( .A1(n8952), .A2(n7002), .ZN(n11174) );
  NAND2_X1 U9366 ( .A1(n8823), .A2(n8825), .ZN(n9311) );
  NAND2_X1 U9367 ( .A1(n12523), .A2(n6607), .ZN(n7018) );
  NAND2_X1 U9368 ( .A1(n12523), .A2(n12524), .ZN(n12522) );
  NAND2_X1 U9369 ( .A1(n7018), .A2(n7016), .ZN(n12463) );
  NAND2_X1 U9370 ( .A1(n9238), .A2(n9260), .ZN(n7017) );
  OAI21_X2 U9371 ( .B1(n12463), .B2(n12465), .A(n12464), .ZN(n12462) );
  NAND2_X1 U9372 ( .A1(n14975), .A2(n7021), .ZN(n7019) );
  NAND2_X1 U9373 ( .A1(n7019), .A2(n7020), .ZN(n12514) );
  NAND2_X4 U9374 ( .A1(n6501), .A2(n9960), .ZN(n12082) );
  AOI21_X1 U9375 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(n14384), .A(n7031), .ZN(
        n7027) );
  AND2_X2 U9376 ( .A1(n6599), .A2(n7028), .ZN(n9459) );
  OAI21_X1 U9377 ( .B1(n14384), .B2(n9452), .A(P2_ADDR_REG_7__SCAN_IN), .ZN(
        n7029) );
  INV_X1 U9378 ( .A(n7033), .ZN(n7030) );
  AOI21_X1 U9379 ( .B1(n9452), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n15215), .ZN(
        n7032) );
  NOR2_X1 U9380 ( .A1(n14384), .A2(n9452), .ZN(n9454) );
  NAND2_X1 U9381 ( .A1(n14567), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U9382 ( .A1(n7057), .A2(n11812), .ZN(n8656) );
  XNOR2_X1 U9383 ( .A(n11989), .B(n7057), .ZN(n10552) );
  NAND2_X1 U9384 ( .A1(n11371), .A2(n12002), .ZN(n8673) );
  NAND2_X1 U9385 ( .A1(n11350), .A2(n8670), .ZN(n7058) );
  NAND2_X2 U9386 ( .A1(n7062), .A2(n7059), .ZN(n8651) );
  OAI21_X2 U9387 ( .B1(n11507), .B2(n7064), .A(n11880), .ZN(n11491) );
  INV_X1 U9388 ( .A(n7070), .ZN(n14169) );
  NOR2_X1 U9389 ( .A1(n14169), .A2(n8681), .ZN(n14150) );
  OAI21_X2 U9390 ( .B1(n7077), .B2(n7073), .A(n7072), .ZN(n11295) );
  NAND2_X1 U9391 ( .A1(n7086), .A2(n6547), .ZN(n14203) );
  OAI22_X1 U9392 ( .A1(n10817), .A2(n8662), .B1(n8661), .B2(n11836), .ZN(
        n10830) );
  NAND2_X1 U9393 ( .A1(n8673), .A2(n8672), .ZN(n11384) );
  NAND2_X1 U9394 ( .A1(n8668), .A2(n8667), .ZN(n11293) );
  NAND2_X1 U9395 ( .A1(n8331), .A2(n9943), .ZN(n8335) );
  NAND2_X1 U9396 ( .A1(n13885), .A2(n10558), .ZN(n11817) );
  XNOR2_X1 U9397 ( .A(n10147), .B(n10150), .ZN(n7102) );
  AND2_X2 U9398 ( .A1(n10353), .A2(n10352), .ZN(n11730) );
  NAND2_X1 U9399 ( .A1(n13036), .A2(n7106), .ZN(n7105) );
  OAI21_X1 U9400 ( .B1(n13036), .B2(n7107), .A(n7106), .ZN(n13012) );
  NAND4_X1 U9401 ( .A1(n7109), .A2(n7488), .A3(n7110), .A4(n7483), .ZN(n7476)
         );
  NAND2_X1 U9402 ( .A1(n13093), .A2(n7111), .ZN(n13028) );
  NAND2_X1 U9403 ( .A1(n10995), .A2(n6605), .ZN(n14464) );
  NAND2_X1 U9404 ( .A1(n10406), .A2(n10407), .ZN(n10534) );
  INV_X1 U9405 ( .A(n7119), .ZN(n11123) );
  NAND2_X1 U9406 ( .A1(n9837), .A2(n7129), .ZN(n7125) );
  NAND2_X1 U9407 ( .A1(n7133), .A2(n8338), .ZN(n8340) );
  XNOR2_X1 U9408 ( .A(n7133), .B(n11991), .ZN(n14654) );
  NAND2_X1 U9409 ( .A1(n9374), .A2(n6603), .ZN(n7135) );
  OAI211_X1 U9410 ( .C1(n9374), .C2(n7139), .A(n7136), .B(n7135), .ZN(n12315)
         );
  NAND2_X1 U9411 ( .A1(n11352), .A2(n7147), .ZN(n7144) );
  NAND2_X1 U9412 ( .A1(n10509), .A2(n7155), .ZN(n7154) );
  NAND2_X1 U9413 ( .A1(n10508), .A2(n10480), .ZN(n7156) );
  NAND4_X1 U9414 ( .A1(n7154), .A2(n7160), .A3(n7156), .A4(n10604), .ZN(n10605) );
  NAND2_X2 U9415 ( .A1(n7161), .A2(n9960), .ZN(n7870) );
  OAI21_X2 U9416 ( .B1(n8223), .B2(n7515), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7162) );
  INV_X1 U9417 ( .A(n13236), .ZN(n7167) );
  AOI21_X2 U9418 ( .B1(n7172), .B2(n6556), .A(n7169), .ZN(n13499) );
  NAND2_X1 U9419 ( .A1(n13329), .A2(n7177), .ZN(n7176) );
  AOI21_X1 U9420 ( .B1(n13329), .B2(n13248), .A(n13247), .ZN(n13313) );
  INV_X1 U9421 ( .A(n13459), .ZN(n7187) );
  MUX2_X1 U9422 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7547), .Z(n7590) );
  NAND2_X1 U9423 ( .A1(n7615), .A2(n7614), .ZN(n7633) );
  NAND2_X1 U9424 ( .A1(n7674), .A2(n7197), .ZN(n7196) );
  NAND2_X1 U9425 ( .A1(n7674), .A2(n7673), .ZN(n7200) );
  NAND3_X1 U9426 ( .A1(n7202), .A2(n6645), .A3(n7201), .ZN(n8059) );
  NAND3_X1 U9427 ( .A1(n7202), .A2(n7203), .A3(n7201), .ZN(n8055) );
  NAND3_X1 U9428 ( .A1(n7207), .A2(n7205), .A3(n7208), .ZN(n8019) );
  NAND3_X1 U9429 ( .A1(n7208), .A2(n7210), .A3(n7207), .ZN(n8566) );
  NAND2_X1 U9430 ( .A1(n8111), .A2(n7215), .ZN(n7214) );
  NAND3_X1 U9431 ( .A1(n7237), .A2(n10597), .A3(n10596), .ZN(n13531) );
  NAND2_X1 U9432 ( .A1(n13507), .A2(n6524), .ZN(n13492) );
  INV_X2 U9433 ( .A(n7870), .ZN(n8167) );
  NAND2_X1 U9434 ( .A1(n7572), .A2(n10074), .ZN(n7249) );
  OAI21_X1 U9435 ( .B1(n8981), .B2(n7272), .A(n7268), .ZN(n9011) );
  NOR2_X2 U9436 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7548) );
  NAND2_X1 U9437 ( .A1(n7940), .A2(n7941), .ZN(n7939) );
  NAND3_X1 U9438 ( .A1(n7689), .A2(n7688), .A3(n6621), .ZN(n7285) );
  INV_X1 U9439 ( .A(n7706), .ZN(n7286) );
  NAND3_X1 U9440 ( .A1(n7736), .A2(n7735), .A3(n6622), .ZN(n7288) );
  INV_X1 U9441 ( .A(n7755), .ZN(n7289) );
  NAND3_X1 U9442 ( .A1(n7781), .A2(n7780), .A3(n6623), .ZN(n7291) );
  INV_X1 U9443 ( .A(n7808), .ZN(n7292) );
  NAND3_X1 U9444 ( .A1(n7645), .A2(n7644), .A3(n7296), .ZN(n7297) );
  INV_X1 U9445 ( .A(n7662), .ZN(n7298) );
  NAND3_X1 U9446 ( .A1(n7603), .A2(n7602), .A3(n7299), .ZN(n7301) );
  INV_X1 U9447 ( .A(n7620), .ZN(n7302) );
  NAND3_X1 U9448 ( .A1(n8072), .A2(n6617), .A3(n8071), .ZN(n7303) );
  NAND2_X1 U9449 ( .A1(n7310), .A2(n7311), .ZN(n13763) );
  NAND2_X1 U9450 ( .A1(n7318), .A2(n7319), .ZN(n12376) );
  NAND2_X1 U9451 ( .A1(n13842), .A2(n7320), .ZN(n7318) );
  OAI21_X1 U9452 ( .B1(n13802), .B2(n7333), .A(n7330), .ZN(n11648) );
  AND2_X1 U9453 ( .A1(n11324), .A2(n11325), .ZN(n7341) );
  NAND2_X1 U9454 ( .A1(n8643), .A2(n6616), .ZN(n8715) );
  NAND2_X1 U9455 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  NAND2_X1 U9456 ( .A1(n7349), .A2(n7348), .ZN(n7354) );
  INV_X1 U9457 ( .A(n7349), .ZN(n7356) );
  NAND2_X1 U9458 ( .A1(n7354), .A2(n7353), .ZN(n7350) );
  OAI211_X1 U9459 ( .C1(n7354), .C2(n7352), .A(n7351), .B(n11842), .ZN(n11841)
         );
  NAND2_X1 U9460 ( .A1(n11838), .A2(n7355), .ZN(n7351) );
  INV_X1 U9461 ( .A(n7355), .ZN(n7352) );
  NAND2_X1 U9462 ( .A1(n11941), .A2(n7361), .ZN(n7363) );
  NAND3_X1 U9463 ( .A1(n11939), .A2(n11938), .A3(n7363), .ZN(n7362) );
  NAND2_X1 U9464 ( .A1(n11934), .A2(n11935), .ZN(n11933) );
  NAND3_X1 U9465 ( .A1(n11845), .A2(n11844), .A3(n6614), .ZN(n7368) );
  NAND2_X1 U9466 ( .A1(n7368), .A2(n7369), .ZN(n11851) );
  NAND2_X1 U9467 ( .A1(n11868), .A2(n7371), .ZN(n7374) );
  OAI21_X1 U9468 ( .B1(n11868), .B2(n7379), .A(n7377), .ZN(n11876) );
  NAND2_X1 U9469 ( .A1(n7374), .A2(n7372), .ZN(n11874) );
  OR2_X1 U9470 ( .A1(n12759), .A2(n7387), .ZN(n7386) );
  INV_X1 U9471 ( .A(n9702), .ZN(n7396) );
  AOI21_X1 U9472 ( .B1(n7396), .B2(n6601), .A(n7397), .ZN(n9705) );
  INV_X1 U9473 ( .A(n7411), .ZN(n9729) );
  AOI21_X1 U9474 ( .B1(n11756), .B2(n7415), .A(n7418), .ZN(n7414) );
  OAI21_X1 U9475 ( .B1(n11756), .B2(n9708), .A(n9707), .ZN(n12652) );
  NAND2_X1 U9476 ( .A1(n12273), .A2(n12427), .ZN(n7423) );
  NAND2_X1 U9477 ( .A1(n7426), .A2(n7424), .ZN(n9690) );
  NAND2_X1 U9478 ( .A1(n8813), .A2(n7431), .ZN(n8836) );
  OR2_X1 U9479 ( .A1(n7870), .A2(n8739), .ZN(n7527) );
  OAI21_X1 U9480 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7537) );
  INV_X1 U9481 ( .A(n12299), .ZN(n12305) );
  NAND2_X1 U9482 ( .A1(n9365), .A2(n14687), .ZN(n8736) );
  OR2_X1 U9483 ( .A1(n8215), .A2(n8214), .ZN(n8216) );
  AND2_X1 U9484 ( .A1(n8203), .A2(n8155), .ZN(n8149) );
  OR2_X1 U9485 ( .A1(n8913), .A2(n6655), .ZN(n8894) );
  INV_X1 U9486 ( .A(n7866), .ZN(n7867) );
  NAND2_X1 U9487 ( .A1(n11530), .A2(n11529), .ZN(n11551) );
  INV_X1 U9488 ( .A(n11526), .ZN(n11528) );
  NAND2_X1 U9489 ( .A1(n8646), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8299) );
  OAI21_X1 U9490 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8244) );
  INV_X1 U9491 ( .A(n8840), .ZN(n8846) );
  OAI21_X1 U9492 ( .B1(n9821), .B2(n14685), .A(n9362), .ZN(P1_U3524) );
  AND3_X1 U9493 ( .A1(n11984), .A2(n11983), .A3(n7451), .ZN(n12029) );
  NAND2_X1 U9494 ( .A1(n8646), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8310) );
  XNOR2_X1 U9495 ( .A(n11197), .B(n10938), .ZN(n10939) );
  NAND2_X1 U9496 ( .A1(n10937), .A2(n10936), .ZN(n11197) );
  NAND2_X1 U9497 ( .A1(n8665), .A2(n8664), .ZN(n11141) );
  NAND2_X1 U9498 ( .A1(n13736), .A2(n13735), .ZN(n13734) );
  NOR3_X1 U9499 ( .A1(n14168), .A2(n11907), .A3(n11906), .ZN(n7441) );
  OR2_X1 U9500 ( .A1(n11839), .A2(n11142), .ZN(n7442) );
  INV_X1 U9501 ( .A(n12195), .ZN(n9764) );
  INV_X2 U9502 ( .A(n15128), .ZN(n15126) );
  INV_X1 U9503 ( .A(n12389), .ZN(n9693) );
  NOR2_X1 U9504 ( .A1(n8511), .A2(n8500), .ZN(n7443) );
  OR2_X1 U9505 ( .A1(n6507), .A2(n6992), .ZN(n7444) );
  AND2_X1 U9506 ( .A1(n9862), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7445) );
  INV_X1 U9507 ( .A(n11100), .ZN(n9955) );
  AND2_X1 U9508 ( .A1(n12400), .A2(n12587), .ZN(n7447) );
  OR2_X1 U9509 ( .A1(n12301), .A2(n13869), .ZN(n7448) );
  INV_X1 U9510 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9453) );
  INV_X1 U9511 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7506) );
  INV_X1 U9512 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9442) );
  AND2_X1 U9513 ( .A1(n7793), .A2(n7767), .ZN(n7449) );
  XNOR2_X1 U9514 ( .A(n12950), .B(n12589), .ZN(n12720) );
  AND4_X1 U9515 ( .A1(n8803), .A2(n8802), .A3(n8829), .A4(n9115), .ZN(n7450)
         );
  INV_X1 U9516 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11689) );
  NAND2_X1 U9517 ( .A1(n14698), .A2(n14669), .ZN(n14316) );
  INV_X1 U9518 ( .A(n14316), .ZN(n9824) );
  AND2_X2 U9519 ( .A1(n8733), .A2(n9363), .ZN(n14687) );
  AND2_X1 U9520 ( .A1(n12024), .A2(n12026), .ZN(n7451) );
  NOR2_X1 U9521 ( .A1(n9232), .A2(n9216), .ZN(n7454) );
  AND2_X1 U9522 ( .A1(n12858), .A2(n12585), .ZN(n7455) );
  NAND2_X2 U9523 ( .A1(n10647), .A2(n14206), .ZN(n14253) );
  AND2_X2 U9524 ( .A1(n9364), .A2(n9363), .ZN(n14698) );
  INV_X2 U9525 ( .A(n14698), .ZN(n14695) );
  AND2_X1 U9526 ( .A1(n9820), .A2(n9819), .ZN(n7456) );
  AND2_X1 U9527 ( .A1(n9802), .A2(n9801), .ZN(n7457) );
  AND2_X1 U9528 ( .A1(n9788), .A2(n9787), .ZN(n7458) );
  INV_X1 U9529 ( .A(n14043), .ZN(n14040) );
  NOR3_X1 U9530 ( .A1(n13306), .A2(n13305), .A3(n10602), .ZN(n7460) );
  INV_X1 U9531 ( .A(n12382), .ZN(n12301) );
  INV_X1 U9532 ( .A(n13597), .ZN(n13222) );
  OR2_X1 U9533 ( .A1(n11800), .A2(n11835), .ZN(n11805) );
  AND2_X1 U9534 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  MUX2_X1 U9535 ( .A(n11818), .B(n11817), .S(n11952), .Z(n11819) );
  MUX2_X1 U9536 ( .A(n13883), .B(n11829), .S(n11835), .Z(n11828) );
  NAND2_X1 U9537 ( .A1(n11827), .A2(n11826), .ZN(n11832) );
  NAND2_X1 U9538 ( .A1(n7779), .A2(n7778), .ZN(n7780) );
  NAND2_X1 U9539 ( .A1(n11865), .A2(n11864), .ZN(n11868) );
  AND2_X1 U9540 ( .A1(n7889), .A2(n7896), .ZN(n7890) );
  INV_X1 U9541 ( .A(n11910), .ZN(n11915) );
  NOR2_X1 U9542 ( .A1(n11915), .A2(n11914), .ZN(n11916) );
  NAND2_X1 U9543 ( .A1(n7943), .A2(n7942), .ZN(n7944) );
  INV_X1 U9544 ( .A(n12165), .ZN(n12171) );
  NAND2_X1 U9545 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  INV_X1 U9546 ( .A(n11986), .ZN(n12008) );
  NOR3_X1 U9547 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .A3(
        P1_IR_REG_16__SCAN_IN), .ZN(n8249) );
  OR4_X1 U9548 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10135) );
  INV_X1 U9549 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U9550 ( .A1(n6500), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9827) );
  OR2_X1 U9551 ( .A1(n14033), .A2(n13870), .ZN(n8629) );
  AND4_X1 U9552 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n8256)
         );
  INV_X1 U9553 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8251) );
  INV_X1 U9554 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7508) );
  AND2_X1 U9555 ( .A1(n11060), .A2(n11062), .ZN(n8948) );
  INV_X1 U9556 ( .A(n9833), .ZN(n9835) );
  NOR2_X1 U9557 ( .A1(n11100), .A2(n8959), .ZN(n9838) );
  NAND2_X1 U9558 ( .A1(n12595), .A2(n9693), .ZN(n9694) );
  NAND2_X1 U9559 ( .A1(n12596), .A2(n14450), .ZN(n12210) );
  AND2_X1 U9560 ( .A1(n7847), .A2(n7846), .ZN(n7900) );
  AND2_X1 U9561 ( .A1(n8086), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8100) );
  INV_X1 U9562 ( .A(n13572), .ZN(n13223) );
  INV_X1 U9563 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9564 ( .A1(n10935), .A2(n10934), .ZN(n10936) );
  INV_X2 U9565 ( .A(n11638), .ZN(n12360) );
  INV_X1 U9566 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8347) );
  INV_X1 U9567 ( .A(n11998), .ZN(n8667) );
  INV_X1 U9568 ( .A(n12016), .ZN(n9352) );
  INV_X1 U9569 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8259) );
  INV_X1 U9570 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U9571 ( .A1(n7523), .A2(n8739), .ZN(n7522) );
  NOR2_X1 U9572 ( .A1(n9427), .A2(n9426), .ZN(n9406) );
  INV_X1 U9573 ( .A(n12396), .ZN(n9106) );
  INV_X1 U9574 ( .A(n10579), .ZN(n9746) );
  AND2_X1 U9575 ( .A1(n6504), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U9576 ( .A1(n9919), .A2(n14408), .ZN(n9920) );
  INV_X1 U9577 ( .A(n9921), .ZN(n9923) );
  INV_X1 U9578 ( .A(n12261), .ZN(n11779) );
  OR2_X1 U9579 ( .A1(n9120), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9136) );
  INV_X1 U9580 ( .A(n12833), .ZN(n9766) );
  OAI21_X1 U9581 ( .B1(n9304), .B2(n9303), .A(n10165), .ZN(n9741) );
  INV_X1 U9582 ( .A(n9950), .ZN(n15003) );
  AND3_X1 U9583 ( .A1(n9318), .A2(n9317), .A3(n9741), .ZN(n9332) );
  AND2_X1 U9584 ( .A1(n8759), .A2(n8758), .ZN(n9010) );
  INV_X1 U9585 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10412) );
  INV_X1 U9586 ( .A(n10372), .ZN(n10370) );
  NOR2_X1 U9587 ( .A1(n8048), .A2(n8049), .ZN(n8073) );
  NOR2_X1 U9588 ( .A1(n7985), .A2(n7983), .ZN(n8009) );
  OR2_X1 U9589 ( .A1(n7921), .A2(n11689), .ZN(n7946) );
  NAND2_X1 U9590 ( .A1(n7900), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7921) );
  INV_X1 U9591 ( .A(n7814), .ZN(n7709) );
  INV_X1 U9592 ( .A(n13410), .ZN(n13422) );
  INV_X1 U9593 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8474) );
  INV_X1 U9594 ( .A(n10460), .ZN(n10457) );
  INV_X1 U9595 ( .A(n11196), .ZN(n10938) );
  AOI22_X1 U9596 ( .A1(n12372), .A2(n14248), .B1(n11584), .B2(n14641), .ZN(
        n10460) );
  INV_X1 U9597 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8484) );
  NOR2_X1 U9598 ( .A1(n8548), .A2(n13808), .ZN(n8558) );
  NAND2_X1 U9599 ( .A1(n12301), .A2(n13869), .ZN(n8691) );
  INV_X1 U9600 ( .A(n14057), .ZN(n14086) );
  INV_X1 U9601 ( .A(n11812), .ZN(n11989) );
  NAND2_X1 U9602 ( .A1(n7748), .A2(n7747), .ZN(n7762) );
  INV_X1 U9603 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9407) );
  OAI21_X1 U9604 ( .B1(P3_ADDR_REG_16__SCAN_IN), .B2(n9419), .A(n9418), .ZN(
        n9487) );
  NOR2_X1 U9605 ( .A1(n9074), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9100) );
  INV_X1 U9606 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12529) );
  OR2_X1 U9607 ( .A1(n9811), .A2(n9745), .ZN(n12530) );
  AND2_X1 U9608 ( .A1(n9826), .A2(n9309), .ZN(n12293) );
  INV_X1 U9609 ( .A(n12083), .ZN(n9280) );
  AOI22_X1 U9610 ( .A1(n11087), .A2(n11088), .B1(n11100), .B2(n9898), .ZN(
        n11031) );
  OR2_X1 U9611 ( .A1(n9714), .A2(n12074), .ZN(n8810) );
  AND2_X1 U9612 ( .A1(n9154), .A2(n9554), .ZN(n9170) );
  INV_X1 U9613 ( .A(n12122), .ZN(n12815) );
  OR2_X1 U9614 ( .A1(n9714), .A2(n12321), .ZN(n9715) );
  NAND2_X1 U9615 ( .A1(n12194), .A2(n12195), .ZN(n12192) );
  INV_X1 U9616 ( .A(n12297), .ZN(n12137) );
  INV_X1 U9617 ( .A(n12804), .ZN(n15117) );
  AND2_X1 U9618 ( .A1(n8774), .A2(n8773), .ZN(n9128) );
  AND2_X1 U9619 ( .A1(n8767), .A2(n8766), .ZN(n9056) );
  AND2_X1 U9620 ( .A1(n8749), .A2(n8748), .ZN(n8937) );
  INV_X1 U9621 ( .A(n10864), .ZN(n10865) );
  INV_X1 U9622 ( .A(n13111), .ZN(n11680) );
  INV_X1 U9623 ( .A(n13026), .ZN(n11719) );
  INV_X1 U9624 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13083) );
  INV_X1 U9625 ( .A(n10540), .ZN(n10541) );
  OR2_X1 U9626 ( .A1(n10343), .A2(n14889), .ZN(n10349) );
  NAND2_X1 U9627 ( .A1(n8031), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8048) );
  INV_X1 U9628 ( .A(n13286), .ZN(n13287) );
  OAI21_X1 U9629 ( .B1(n13242), .B2(n13597), .A(n13241), .ZN(n13389) );
  INV_X1 U9630 ( .A(n10793), .ZN(n10798) );
  OR2_X1 U9631 ( .A1(n10265), .A2(n10263), .ZN(n13466) );
  NAND2_X1 U9632 ( .A1(n13216), .A2(n11012), .ZN(n10334) );
  OAI21_X1 U9633 ( .B1(n13428), .B2(n13273), .A(n13272), .ZN(n13409) );
  INV_X1 U9634 ( .A(n13523), .ZN(n13505) );
  INV_X1 U9635 ( .A(n14927), .ZN(n14936) );
  OR2_X1 U9636 ( .A1(n7768), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n7796) );
  INV_X1 U9637 ( .A(n10295), .ZN(n10282) );
  INV_X1 U9638 ( .A(n8592), .ZN(n8580) );
  INV_X1 U9639 ( .A(n13884), .ZN(n10572) );
  AND2_X1 U9640 ( .A1(n13724), .A2(n11603), .ZN(n13780) );
  INV_X1 U9641 ( .A(n13825), .ZN(n13857) );
  AND2_X1 U9642 ( .A1(n6858), .A2(n11960), .ZN(n11976) );
  AND2_X1 U9643 ( .A1(n8632), .A2(n8275), .ZN(n12377) );
  AND2_X1 U9644 ( .A1(n8558), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8568) );
  INV_X1 U9645 ( .A(n8651), .ZN(n13896) );
  INV_X1 U9646 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n13950) );
  INV_X1 U9647 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n13986) );
  OR2_X1 U9648 ( .A1(n14059), .A2(n14644), .ZN(n14276) );
  INV_X1 U9649 ( .A(n11909), .ZN(n8681) );
  NAND2_X1 U9650 ( .A1(n11487), .A2(n14503), .ZN(n14220) );
  INV_X1 U9651 ( .A(n14499), .ZN(n14523) );
  INV_X1 U9652 ( .A(n13874), .ZN(n14510) );
  INV_X1 U9653 ( .A(n14520), .ZN(n14498) );
  NAND2_X1 U9654 ( .A1(n10646), .A2(n10645), .ZN(n10647) );
  AND2_X1 U9655 ( .A1(n8679), .A2(n8678), .ZN(n14204) );
  NAND2_X1 U9656 ( .A1(n11791), .A2(n8645), .ZN(n14680) );
  INV_X1 U9657 ( .A(n14302), .ZN(n14644) );
  AOI21_X1 U9658 ( .B1(n10281), .B2(n10050), .A(n10049), .ZN(n10644) );
  INV_X1 U9659 ( .A(n8533), .ZN(n8518) );
  INV_X1 U9660 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9447) );
  AOI21_X1 U9661 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n9409), .A(n9408), .ZN(
        n9468) );
  AND2_X1 U9662 ( .A1(n11135), .A2(n9305), .ZN(n9306) );
  OAI21_X1 U9663 ( .B1(n12273), .B2(n14973), .A(n9346), .ZN(n9347) );
  NOR2_X1 U9664 ( .A1(n8969), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9017) );
  INV_X1 U9665 ( .A(n14985), .ZN(n12532) );
  NAND2_X1 U9666 ( .A1(n9032), .A2(n9031), .ZN(n9044) );
  OR2_X1 U9667 ( .A1(n8960), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8969) );
  OR2_X1 U9668 ( .A1(n9723), .A2(n9800), .ZN(n12090) );
  AND4_X1 U9669 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n12486)
         );
  INV_X1 U9670 ( .A(n15092), .ZN(n15002) );
  NOR2_X1 U9671 ( .A1(n9743), .A2(n9742), .ZN(n9795) );
  INV_X1 U9672 ( .A(n12651), .ZN(n12649) );
  INV_X1 U9673 ( .A(n15185), .ZN(n15167) );
  OR2_X1 U9674 ( .A1(n15175), .A2(n15182), .ZN(n15190) );
  AND2_X1 U9675 ( .A1(n15122), .A2(n12137), .ZN(n15182) );
  NAND2_X1 U9676 ( .A1(n9308), .A2(n6534), .ZN(n9856) );
  AND2_X1 U9677 ( .A1(n8757), .A2(n8756), .ZN(n8989) );
  NOR2_X2 U9678 ( .A1(n10349), .A2(n10337), .ZN(n13126) );
  INV_X1 U9679 ( .A(n8138), .ZN(n8162) );
  AND2_X1 U9680 ( .A1(n7834), .A2(n7833), .ZN(n13261) );
  INV_X1 U9681 ( .A(n14873), .ZN(n14823) );
  INV_X1 U9682 ( .A(n14805), .ZN(n14877) );
  AOI21_X1 U9683 ( .B1(n13285), .B2(n13523), .A(n13255), .ZN(n13256) );
  INV_X1 U9684 ( .A(n13503), .ZN(n13521) );
  INV_X1 U9685 ( .A(n13466), .ZN(n13529) );
  NAND2_X1 U9686 ( .A1(n10334), .A2(n10267), .ZN(n14927) );
  INV_X1 U9687 ( .A(n13229), .ZN(n13548) );
  INV_X1 U9688 ( .A(n14934), .ZN(n14922) );
  NAND2_X1 U9689 ( .A1(n13648), .A2(n10353), .ZN(n14934) );
  INV_X1 U9690 ( .A(n14886), .ZN(n10333) );
  INV_X1 U9691 ( .A(n13864), .ZN(n13844) );
  NAND2_X1 U9692 ( .A1(n11976), .A2(n13896), .ZN(n14520) );
  AND2_X1 U9693 ( .A1(n8577), .A2(n8576), .ZN(n11637) );
  INV_X1 U9694 ( .A(n8605), .ZN(n8543) );
  INV_X1 U9695 ( .A(n14626), .ZN(n14600) );
  AND2_X1 U9696 ( .A1(n10108), .A2(n10107), .ZN(n14628) );
  INV_X1 U9697 ( .A(n11993), .ZN(n10819) );
  AND2_X1 U9698 ( .A1(n12311), .A2(n6857), .ZN(n14124) );
  INV_X1 U9699 ( .A(n14196), .ZN(n14246) );
  AND3_X1 U9700 ( .A1(n14313), .A2(n14312), .A3(n14311), .ZN(n14345) );
  NAND2_X1 U9701 ( .A1(n8694), .A2(n11963), .ZN(n14676) );
  AND3_X1 U9702 ( .A1(n10836), .A2(n10835), .A3(n10834), .ZN(n10905) );
  INV_X1 U9703 ( .A(n14672), .ZN(n14684) );
  AND2_X1 U9704 ( .A1(n8403), .A2(n8414), .ZN(n13972) );
  NAND2_X1 U9705 ( .A1(n11346), .A2(n9306), .ZN(n9826) );
  AND2_X1 U9706 ( .A1(n9326), .A2(n15121), .ZN(n14973) );
  INV_X1 U9707 ( .A(n14974), .ZN(n12579) );
  INV_X1 U9708 ( .A(n12269), .ZN(n12584) );
  OR2_X1 U9709 ( .A1(n9931), .A2(n9857), .ZN(n15102) );
  AND2_X1 U9710 ( .A1(n12810), .A2(n12809), .ZN(n14453) );
  OR2_X1 U9711 ( .A1(n15128), .A2(n15119), .ZN(n12694) );
  INV_X1 U9712 ( .A(n12901), .ZN(n12911) );
  AND2_X2 U9713 ( .A1(n9795), .A2(n9752), .ZN(n15205) );
  INV_X1 U9714 ( .A(n12676), .ZN(n12935) );
  NAND2_X1 U9715 ( .A1(n15193), .A2(n15190), .ZN(n12981) );
  AND3_X1 U9716 ( .A1(n14453), .A2(n14452), .A3(n14451), .ZN(n14455) );
  INV_X2 U9717 ( .A(n15191), .ZN(n15193) );
  AND2_X1 U9718 ( .A1(n9813), .A2(n9812), .ZN(n15191) );
  INV_X1 U9719 ( .A(SI_29_), .ZN(n12388) );
  INV_X1 U9720 ( .A(SI_23_), .ZN(n10847) );
  INV_X1 U9721 ( .A(SI_19_), .ZN(n10330) );
  INV_X1 U9722 ( .A(SI_14_), .ZN(n10042) );
  INV_X1 U9723 ( .A(n9900), .ZN(n10921) );
  INV_X1 U9724 ( .A(n14381), .ZN(n12387) );
  INV_X1 U9725 ( .A(n13136), .ZN(n14458) );
  INV_X1 U9726 ( .A(n14467), .ZN(n13139) );
  INV_X1 U9727 ( .A(n11746), .ZN(n13144) );
  OR2_X1 U9728 ( .A1(n7761), .A2(n7760), .ZN(n13146) );
  INV_X1 U9729 ( .A(n14851), .ZN(n14881) );
  NAND2_X1 U9730 ( .A1(n13527), .A2(n13216), .ZN(n13515) );
  INV_X1 U9731 ( .A(n13534), .ZN(n13475) );
  OR2_X1 U9732 ( .A1(n10161), .A2(n14886), .ZN(n14957) );
  OR2_X1 U9733 ( .A1(n10161), .A2(n10333), .ZN(n14942) );
  INV_X2 U9734 ( .A(n14942), .ZN(n14944) );
  OR2_X1 U9735 ( .A1(n14889), .A2(n14883), .ZN(n14884) );
  INV_X1 U9736 ( .A(n8205), .ZN(n11012) );
  INV_X1 U9737 ( .A(n14817), .ZN(n13200) );
  AND2_X1 U9738 ( .A1(n10064), .A2(n10062), .ZN(n14596) );
  INV_X1 U9739 ( .A(n8544), .ZN(n14320) );
  INV_X1 U9740 ( .A(n14236), .ZN(n14494) );
  INV_X1 U9741 ( .A(n13817), .ZN(n13858) );
  NAND4_X1 U9742 ( .A1(n8279), .A2(n8278), .A3(n8277), .A4(n8276), .ZN(n13869)
         );
  INV_X1 U9743 ( .A(n11637), .ZN(n14134) );
  CLKBUF_X1 U9744 ( .A(P1_U4016), .Z(n13881) );
  NAND2_X1 U9745 ( .A1(n10108), .A2(n8651), .ZN(n14618) );
  INV_X1 U9746 ( .A(n14596), .ZN(n14637) );
  NAND2_X1 U9747 ( .A1(n14253), .A2(n10651), .ZN(n14196) );
  NAND2_X1 U9748 ( .A1(n14253), .A2(n14684), .ZN(n14219) );
  INV_X1 U9749 ( .A(n14124), .ZN(n14239) );
  AOI21_X1 U9750 ( .B1(n12382), .B2(n9824), .A(n9823), .ZN(n9825) );
  AND3_X1 U9751 ( .A1(n14528), .A2(n14527), .A3(n14526), .ZN(n14547) );
  INV_X1 U9752 ( .A(n14687), .ZN(n14685) );
  AND2_X1 U9753 ( .A1(n14367), .A2(n11477), .ZN(n10279) );
  AND2_X1 U9754 ( .A1(n10060), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10290) );
  INV_X1 U9755 ( .A(n14003), .ZN(n13998) );
  INV_X1 U9756 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10072) );
  NOR2_X2 U9757 ( .A1(n9826), .A2(n13000), .ZN(P3_U3897) );
  AND2_X1 U9758 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9939), .ZN(P2_U3947) );
  INV_X1 U9759 ( .A(n9669), .ZN(P1_U3555) );
  NAND2_X1 U9760 ( .A1(n8736), .A2(n8735), .ZN(P1_U3525) );
  NAND2_X1 U9761 ( .A1(n7109), .A2(n7463), .ZN(n7658) );
  NOR2_X2 U9762 ( .A1(n7658), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U9763 ( .A1(n7866), .A2(n7468), .ZN(n7914) );
  NAND2_X1 U9764 ( .A1(n7471), .A2(n7470), .ZN(n7487) );
  NOR2_X1 U9765 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7473) );
  NAND2_X1 U9766 ( .A1(n7473), .A2(n7472), .ZN(n7484) );
  INV_X1 U9767 ( .A(n7476), .ZN(n7474) );
  NAND2_X1 U9768 ( .A1(n7474), .A2(n7482), .ZN(n7479) );
  XNOR2_X2 U9769 ( .A(n7475), .B(P2_IR_REG_22__SCAN_IN), .ZN(n10150) );
  NAND2_X1 U9770 ( .A1(n7476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7477) );
  MUX2_X1 U9771 ( .A(n7477), .B(P2_IR_REG_31__SCAN_IN), .S(n7482), .Z(n7478)
         );
  NAND2_X1 U9772 ( .A1(n6584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7480) );
  AND2_X1 U9773 ( .A1(n10144), .A2(n10147), .ZN(n8208) );
  INV_X2 U9774 ( .A(n7807), .ZN(n8170) );
  NAND3_X1 U9775 ( .A1(n7483), .A2(n7482), .A3(n7481), .ZN(n8214) );
  INV_X1 U9776 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7485) );
  NAND3_X1 U9777 ( .A1(n8224), .A2(n8226), .A3(n7485), .ZN(n7486) );
  INV_X1 U9778 ( .A(n7494), .ZN(n7492) );
  NAND2_X1 U9779 ( .A1(n7514), .A2(n7516), .ZN(n7495) );
  NOR2_X1 U9780 ( .A1(n7495), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7491) );
  NAND2_X1 U9781 ( .A1(n7492), .A2(n7491), .ZN(n13672) );
  NAND2_X1 U9782 ( .A1(n7495), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7496) );
  NAND2_X1 U9783 ( .A1(n7513), .A2(n7496), .ZN(n7498) );
  NAND2_X1 U9785 ( .A1(n8050), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7504) );
  INV_X1 U9786 ( .A(n7500), .ZN(n13680) );
  AND2_X2 U9787 ( .A1(n7499), .A2(n13680), .ZN(n7814) );
  NAND2_X1 U9788 ( .A1(n7814), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U9789 ( .A1(n7815), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7502) );
  NAND2_X1 U9790 ( .A1(n8138), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7501) );
  NAND4_X2 U9791 ( .A1(n7504), .A2(n7501), .A3(n7502), .A4(n7503), .ZN(n13157)
         );
  NAND2_X1 U9792 ( .A1(n8170), .A2(n13157), .ZN(n7518) );
  INV_X1 U9793 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14018) );
  INV_X1 U9794 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7507) );
  NAND3_X1 U9795 ( .A1(n7507), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U9796 ( .A1(n7509), .A2(n7508), .ZN(n7510) );
  NAND2_X2 U9797 ( .A1(n7511), .A2(n7510), .ZN(n7523) );
  NAND2_X1 U9798 ( .A1(n9961), .A2(SI_0_), .ZN(n7512) );
  XNOR2_X1 U9799 ( .A(n7512), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13691) );
  NAND2_X1 U9800 ( .A1(n8234), .A2(n7514), .ZN(n7515) );
  MUX2_X1 U9801 ( .A(n13691), .B(P2_IR_REG_0__SCAN_IN), .S(n6499), .Z(n10354)
         );
  INV_X1 U9802 ( .A(n10147), .ZN(n10352) );
  AOI21_X1 U9803 ( .B1(n6469), .B2(n10144), .A(n10352), .ZN(n7517) );
  OAI21_X1 U9804 ( .B1(n7518), .B2(n10354), .A(n7517), .ZN(n7521) );
  NAND2_X1 U9805 ( .A1(n7519), .A2(n7518), .ZN(n7520) );
  INV_X1 U9806 ( .A(n8169), .ZN(n7571) );
  INV_X1 U9807 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9962) );
  INV_X1 U9808 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8739) );
  OAI21_X2 U9809 ( .B1(n7523), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7522), .ZN(
        n7543) );
  XNOR2_X2 U9810 ( .A(n7543), .B(SI_1_), .ZN(n7545) );
  MUX2_X1 U9811 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n7523), .Z(n7524) );
  XNOR2_X1 U9812 ( .A(n7542), .B(n7545), .ZN(n8295) );
  NAND2_X1 U9813 ( .A1(n7571), .A2(n8295), .ZN(n7528) );
  NAND2_X1 U9814 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7525) );
  NAND2_X1 U9815 ( .A1(n7572), .A2(n13162), .ZN(n7526) );
  NAND2_X1 U9816 ( .A1(n8050), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7532) );
  NAND2_X1 U9817 ( .A1(n7815), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7531) );
  NAND2_X1 U9818 ( .A1(n8138), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7530) );
  NAND2_X1 U9819 ( .A1(n7814), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7529) );
  MUX2_X1 U9820 ( .A(n10623), .B(n8193), .S(n8170), .Z(n7534) );
  MUX2_X1 U9821 ( .A(n13156), .B(n13018), .S(n8170), .Z(n7533) );
  NAND2_X1 U9822 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  NAND2_X1 U9823 ( .A1(n7537), .A2(n7536), .ZN(n7554) );
  NAND2_X1 U9824 ( .A1(n7814), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U9825 ( .A1(n8050), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7540) );
  NAND2_X1 U9826 ( .A1(n7815), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U9827 ( .A1(n8138), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7538) );
  INV_X1 U9828 ( .A(n7542), .ZN(n7546) );
  INV_X1 U9829 ( .A(SI_1_), .ZN(n9948) );
  NOR2_X1 U9830 ( .A1(n7543), .A2(n9948), .ZN(n7544) );
  AOI21_X2 U9831 ( .B1(n7546), .B2(n7545), .A(n7544), .ZN(n7567) );
  XNOR2_X1 U9832 ( .A(n7567), .B(SI_2_), .ZN(n7566) );
  INV_X1 U9833 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9969) );
  MUX2_X1 U9834 ( .A(n9969), .B(n9942), .S(n9961), .Z(n7564) );
  XNOR2_X1 U9835 ( .A(n7566), .B(n7564), .ZN(n8312) );
  NAND2_X1 U9836 ( .A1(n8312), .A2(n7571), .ZN(n7551) );
  INV_X1 U9837 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13671) );
  OR2_X1 U9838 ( .A1(n7548), .A2(n13671), .ZN(n7549) );
  XNOR2_X1 U9839 ( .A(n7549), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10074) );
  NAND2_X2 U9840 ( .A1(n7551), .A2(n7550), .ZN(n10591) );
  MUX2_X1 U9841 ( .A(n13155), .B(n10591), .S(n8170), .Z(n7555) );
  NAND2_X1 U9842 ( .A1(n7554), .A2(n7555), .ZN(n7553) );
  MUX2_X1 U9843 ( .A(n10591), .B(n13155), .S(n8170), .Z(n7552) );
  NAND2_X1 U9844 ( .A1(n7553), .A2(n7552), .ZN(n7559) );
  INV_X1 U9845 ( .A(n7554), .ZN(n7557) );
  INV_X1 U9846 ( .A(n7555), .ZN(n7556) );
  NAND2_X1 U9847 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  NAND2_X1 U9848 ( .A1(n7814), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7563) );
  INV_X1 U9849 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U9850 ( .A1(n8050), .A2(n10490), .ZN(n7562) );
  NAND2_X1 U9851 ( .A1(n7815), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7561) );
  NAND2_X1 U9852 ( .A1(n8138), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7560) );
  NAND4_X1 U9853 ( .A1(n7563), .A2(n7562), .A3(n7561), .A4(n7560), .ZN(n13154)
         );
  INV_X1 U9854 ( .A(n7564), .ZN(n7565) );
  NAND2_X1 U9855 ( .A1(n7566), .A2(n7565), .ZN(n7570) );
  INV_X1 U9856 ( .A(n7567), .ZN(n7568) );
  NAND2_X1 U9857 ( .A1(n7568), .A2(SI_2_), .ZN(n7569) );
  INV_X1 U9858 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U9859 ( .A1(n7548), .A2(n7573), .ZN(n7593) );
  NAND2_X1 U9860 ( .A1(n7593), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7574) );
  XNOR2_X1 U9861 ( .A(n7574), .B(P2_IR_REG_3__SCAN_IN), .ZN(n14699) );
  MUX2_X1 U9862 ( .A(n13154), .B(n10491), .S(n7773), .Z(n7578) );
  NAND2_X1 U9863 ( .A1(n7577), .A2(n7578), .ZN(n7576) );
  MUX2_X1 U9864 ( .A(n13154), .B(n10491), .S(n8148), .Z(n7575) );
  NAND2_X1 U9865 ( .A1(n7576), .A2(n7575), .ZN(n7582) );
  INV_X1 U9866 ( .A(n7577), .ZN(n7580) );
  INV_X1 U9867 ( .A(n7578), .ZN(n7579) );
  NAND2_X1 U9868 ( .A1(n7580), .A2(n7579), .ZN(n7581) );
  NAND2_X1 U9869 ( .A1(n7582), .A2(n7581), .ZN(n7598) );
  NAND2_X1 U9870 ( .A1(n8138), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7586) );
  INV_X2 U9871 ( .A(n7709), .ZN(n8157) );
  NAND2_X1 U9872 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7604) );
  OAI21_X1 U9873 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n7604), .ZN(n13074) );
  INV_X1 U9874 ( .A(n13074), .ZN(n10505) );
  NAND2_X1 U9875 ( .A1(n8050), .A2(n10505), .ZN(n7584) );
  NAND2_X1 U9876 ( .A1(n7815), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U9877 ( .A1(n7589), .A2(n7588), .ZN(n7592) );
  NAND2_X1 U9878 ( .A1(n7590), .A2(SI_3_), .ZN(n7591) );
  INV_X2 U9879 ( .A(n8169), .ZN(n8097) );
  OR2_X1 U9880 ( .A1(n7593), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7616) );
  NAND2_X1 U9881 ( .A1(n7616), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7594) );
  XNOR2_X1 U9882 ( .A(n7594), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14711) );
  AOI22_X1 U9883 ( .A1(n8167), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7572), .B2(
        n14711), .ZN(n7595) );
  MUX2_X1 U9884 ( .A(n13153), .B(n13076), .S(n8170), .Z(n7599) );
  NAND2_X1 U9885 ( .A1(n7598), .A2(n7599), .ZN(n7597) );
  MUX2_X1 U9886 ( .A(n13153), .B(n13076), .S(n7773), .Z(n7596) );
  NAND2_X1 U9887 ( .A1(n7597), .A2(n7596), .ZN(n7603) );
  INV_X1 U9888 ( .A(n7598), .ZN(n7601) );
  INV_X1 U9889 ( .A(n7599), .ZN(n7600) );
  NAND2_X1 U9890 ( .A1(n7601), .A2(n7600), .ZN(n7602) );
  NAND2_X1 U9891 ( .A1(n8138), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9892 ( .A1(n7814), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7608) );
  NOR2_X1 U9893 ( .A1(n7604), .A2(n10412), .ZN(n7623) );
  INV_X1 U9894 ( .A(n7623), .ZN(n7625) );
  NAND2_X1 U9895 ( .A1(n7604), .A2(n10412), .ZN(n7605) );
  AND2_X1 U9896 ( .A1(n7625), .A2(n7605), .ZN(n10474) );
  NAND2_X1 U9897 ( .A1(n8050), .A2(n10474), .ZN(n7607) );
  NAND2_X1 U9898 ( .A1(n7815), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7606) );
  NAND4_X1 U9899 ( .A1(n7609), .A2(n7608), .A3(n7607), .A4(n7606), .ZN(n13524)
         );
  NAND2_X1 U9900 ( .A1(n7613), .A2(SI_4_), .ZN(n7614) );
  MUX2_X1 U9901 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9961), .Z(n7634) );
  XNOR2_X1 U9902 ( .A(n7634), .B(SI_5_), .ZN(n7631) );
  XNOR2_X1 U9903 ( .A(n7633), .B(n7631), .ZN(n9965) );
  NAND2_X1 U9904 ( .A1(n9965), .A2(n8097), .ZN(n7619) );
  OAI21_X1 U9905 ( .B1(n7616), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7617) );
  XNOR2_X1 U9906 ( .A(n7617), .B(P2_IR_REG_5__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U9907 ( .A1(n8167), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7572), .B2(
        n14723), .ZN(n7618) );
  MUX2_X1 U9908 ( .A(n13524), .B(n14904), .S(n7773), .Z(n7621) );
  MUX2_X1 U9909 ( .A(n13524), .B(n14904), .S(n8148), .Z(n7620) );
  INV_X1 U9910 ( .A(n7621), .ZN(n7622) );
  NAND2_X1 U9911 ( .A1(n8157), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7630) );
  NAND2_X1 U9912 ( .A1(n8158), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U9913 ( .A1(n7623), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7647) );
  INV_X1 U9914 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7624) );
  NAND2_X1 U9915 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  AND2_X1 U9916 ( .A1(n7647), .A2(n7626), .ZN(n13528) );
  NAND2_X1 U9917 ( .A1(n8050), .A2(n13528), .ZN(n7628) );
  NAND2_X1 U9918 ( .A1(n8138), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7627) );
  NAND4_X1 U9919 ( .A1(n7630), .A2(n7629), .A3(n7628), .A4(n7627), .ZN(n13152)
         );
  INV_X1 U9920 ( .A(n7631), .ZN(n7632) );
  MUX2_X1 U9921 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9961), .Z(n7656) );
  XNOR2_X1 U9922 ( .A(n7656), .B(SI_6_), .ZN(n7653) );
  XNOR2_X1 U9923 ( .A(n7655), .B(n7653), .ZN(n9971) );
  NAND2_X1 U9924 ( .A1(n9971), .A2(n8097), .ZN(n7637) );
  NAND2_X1 U9925 ( .A1(n8215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7635) );
  XNOR2_X1 U9926 ( .A(n7635), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U9927 ( .A1(n8167), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7572), .B2(
        n14735), .ZN(n7636) );
  NAND2_X1 U9928 ( .A1(n7637), .A2(n7636), .ZN(n14912) );
  MUX2_X1 U9929 ( .A(n13152), .B(n14912), .S(n8148), .Z(n7641) );
  NAND2_X1 U9930 ( .A1(n7640), .A2(n7641), .ZN(n7639) );
  MUX2_X1 U9931 ( .A(n13152), .B(n14912), .S(n7773), .Z(n7638) );
  NAND2_X1 U9932 ( .A1(n7639), .A2(n7638), .ZN(n7645) );
  INV_X1 U9933 ( .A(n7640), .ZN(n7643) );
  INV_X1 U9934 ( .A(n7641), .ZN(n7642) );
  NAND2_X1 U9935 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  NAND2_X1 U9936 ( .A1(n8157), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U9937 ( .A1(n8158), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7651) );
  INV_X1 U9938 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7646) );
  NAND2_X1 U9939 ( .A1(n7647), .A2(n7646), .ZN(n7648) );
  AND2_X1 U9940 ( .A1(n7666), .A2(n7648), .ZN(n10674) );
  NAND2_X1 U9941 ( .A1(n8050), .A2(n10674), .ZN(n7650) );
  NAND2_X1 U9942 ( .A1(n8138), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7649) );
  NAND4_X1 U9943 ( .A1(n7652), .A2(n7651), .A3(n7650), .A4(n7649), .ZN(n13522)
         );
  INV_X1 U9944 ( .A(n7653), .ZN(n7654) );
  NAND2_X1 U9945 ( .A1(n7656), .A2(SI_6_), .ZN(n7657) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9961), .Z(n7675) );
  XNOR2_X1 U9947 ( .A(n7675), .B(SI_7_), .ZN(n7672) );
  XNOR2_X1 U9948 ( .A(n7674), .B(n7672), .ZN(n9989) );
  NAND2_X1 U9949 ( .A1(n9989), .A2(n8097), .ZN(n7661) );
  NAND2_X1 U9950 ( .A1(n7658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7659) );
  XNOR2_X1 U9951 ( .A(n7659), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U9952 ( .A1(n8167), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6499), .B2(
        n13175), .ZN(n7660) );
  MUX2_X1 U9953 ( .A(n13522), .B(n14919), .S(n7773), .Z(n7663) );
  MUX2_X1 U9954 ( .A(n13522), .B(n14919), .S(n8148), .Z(n7662) );
  INV_X1 U9955 ( .A(n7663), .ZN(n7664) );
  NAND2_X1 U9956 ( .A1(n8138), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9957 ( .A1(n8157), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7670) );
  INV_X1 U9958 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7665) );
  NAND2_X1 U9959 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  NAND2_X1 U9960 ( .A1(n7691), .A2(n7667), .ZN(n12060) );
  INV_X1 U9961 ( .A(n12060), .ZN(n10689) );
  NAND2_X1 U9962 ( .A1(n8050), .A2(n10689), .ZN(n7669) );
  NAND2_X1 U9963 ( .A1(n7815), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7668) );
  NAND4_X1 U9964 ( .A1(n7671), .A2(n7670), .A3(n7669), .A4(n7668), .ZN(n13151)
         );
  INV_X1 U9965 ( .A(n7672), .ZN(n7673) );
  NAND2_X1 U9966 ( .A1(n7675), .A2(SI_7_), .ZN(n7676) );
  MUX2_X1 U9967 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9961), .Z(n7700) );
  XNOR2_X1 U9968 ( .A(n7700), .B(SI_8_), .ZN(n7697) );
  XNOR2_X1 U9969 ( .A(n7699), .B(n7697), .ZN(n10002) );
  NAND2_X1 U9970 ( .A1(n10002), .A2(n8097), .ZN(n7681) );
  INV_X1 U9971 ( .A(n7677), .ZN(n7678) );
  NAND2_X1 U9972 ( .A1(n7678), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7679) );
  XNOR2_X1 U9973 ( .A(n7679), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14747) );
  AOI22_X1 U9974 ( .A1(n8167), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7572), .B2(
        n14747), .ZN(n7680) );
  MUX2_X1 U9975 ( .A(n13151), .B(n12070), .S(n8170), .Z(n7685) );
  NAND2_X1 U9976 ( .A1(n7684), .A2(n7685), .ZN(n7683) );
  MUX2_X1 U9977 ( .A(n13151), .B(n12070), .S(n7773), .Z(n7682) );
  NAND2_X1 U9978 ( .A1(n7683), .A2(n7682), .ZN(n7689) );
  INV_X1 U9979 ( .A(n7684), .ZN(n7687) );
  INV_X1 U9980 ( .A(n7685), .ZN(n7686) );
  NAND2_X1 U9981 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  NAND2_X1 U9982 ( .A1(n8138), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U9983 ( .A1(n8157), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7695) );
  INV_X1 U9984 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7690) );
  INV_X1 U9985 ( .A(n7710), .ZN(n7712) );
  NAND2_X1 U9986 ( .A1(n7691), .A2(n7690), .ZN(n7692) );
  AND2_X1 U9987 ( .A1(n7712), .A2(n7692), .ZN(n11694) );
  NAND2_X1 U9988 ( .A1(n8050), .A2(n11694), .ZN(n7694) );
  NAND2_X1 U9989 ( .A1(n7815), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7693) );
  NAND4_X1 U9990 ( .A1(n7696), .A2(n7695), .A3(n7694), .A4(n7693), .ZN(n13149)
         );
  INV_X1 U9991 ( .A(n7697), .ZN(n7698) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9961), .Z(n7721) );
  XNOR2_X1 U9993 ( .A(n7721), .B(SI_9_), .ZN(n7718) );
  XNOR2_X1 U9994 ( .A(n7720), .B(n7718), .ZN(n10038) );
  NAND2_X1 U9995 ( .A1(n10038), .A2(n8097), .ZN(n7705) );
  NAND2_X1 U9996 ( .A1(n6585), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7701) );
  MUX2_X1 U9997 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7701), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7703) );
  INV_X1 U9998 ( .A(n7702), .ZN(n7725) );
  AOI22_X1 U9999 ( .A1(n8167), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6499), .B2(
        n14759), .ZN(n7704) );
  MUX2_X1 U10000 ( .A(n13149), .B(n11703), .S(n7773), .Z(n7707) );
  MUX2_X1 U10001 ( .A(n13149), .B(n11703), .S(n8148), .Z(n7706) );
  INV_X1 U10002 ( .A(n7707), .ZN(n7708) );
  NAND2_X1 U10003 ( .A1(n8138), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U10004 ( .A1(n8157), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U10005 ( .A1(n7710), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7738) );
  INV_X1 U10006 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U10007 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  AND2_X1 U10008 ( .A1(n7738), .A2(n7713), .ZN(n10871) );
  NAND2_X1 U10009 ( .A1(n8050), .A2(n10871), .ZN(n7715) );
  NAND2_X1 U10010 ( .A1(n7815), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7714) );
  NAND4_X1 U10011 ( .A1(n7717), .A2(n7716), .A3(n7715), .A4(n7714), .ZN(n13148) );
  INV_X1 U10012 ( .A(n7718), .ZN(n7719) );
  NAND2_X1 U10013 ( .A1(n7721), .A2(SI_9_), .ZN(n7722) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9961), .Z(n7745) );
  XNOR2_X1 U10015 ( .A(n7745), .B(SI_10_), .ZN(n7744) );
  XNOR2_X1 U10016 ( .A(n7724), .B(n7744), .ZN(n10044) );
  NAND2_X1 U10017 ( .A1(n10044), .A2(n8097), .ZN(n7728) );
  NAND2_X1 U10018 ( .A1(n7725), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7726) );
  XNOR2_X1 U10019 ( .A(n7726), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14772) );
  AOI22_X1 U10020 ( .A1(n8167), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7572), 
        .B2(n14772), .ZN(n7727) );
  MUX2_X1 U10021 ( .A(n13148), .B(n10856), .S(n8148), .Z(n7732) );
  NAND2_X1 U10022 ( .A1(n7731), .A2(n7732), .ZN(n7730) );
  MUX2_X1 U10023 ( .A(n13148), .B(n10856), .S(n7773), .Z(n7729) );
  NAND2_X1 U10024 ( .A1(n7730), .A2(n7729), .ZN(n7736) );
  INV_X1 U10025 ( .A(n7731), .ZN(n7734) );
  INV_X1 U10026 ( .A(n7732), .ZN(n7733) );
  NAND2_X1 U10027 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U10028 ( .A1(n8157), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7743) );
  INV_X1 U10029 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10030 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  NAND2_X1 U10031 ( .A1(n7758), .A2(n7739), .ZN(n14469) );
  INV_X1 U10032 ( .A(n14469), .ZN(n10804) );
  NAND2_X1 U10033 ( .A1(n8050), .A2(n10804), .ZN(n7742) );
  NAND2_X1 U10034 ( .A1(n7815), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U10035 ( .A1(n8138), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7740) );
  NAND4_X1 U10036 ( .A1(n7743), .A2(n7742), .A3(n7741), .A4(n7740), .ZN(n13147) );
  NAND2_X1 U10037 ( .A1(n7745), .A2(SI_10_), .ZN(n7746) );
  MUX2_X1 U10038 ( .A(n10072), .B(n10070), .S(n9961), .Z(n7748) );
  INV_X1 U10039 ( .A(n7748), .ZN(n7749) );
  NAND2_X1 U10040 ( .A1(n7749), .A2(SI_11_), .ZN(n7750) );
  NAND2_X1 U10041 ( .A1(n7762), .A2(n7750), .ZN(n7763) );
  XNOR2_X1 U10042 ( .A(n7764), .B(n7763), .ZN(n10069) );
  NAND2_X1 U10043 ( .A1(n10069), .A2(n8097), .ZN(n7754) );
  INV_X1 U10044 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U10045 ( .A1(n7702), .A2(n7751), .ZN(n7768) );
  NAND2_X1 U10046 ( .A1(n7768), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7752) );
  XNOR2_X1 U10047 ( .A(n7752), .B(P2_IR_REG_11__SCAN_IN), .ZN(n14784) );
  AOI22_X1 U10048 ( .A1(n8167), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n14784), 
        .B2(n6499), .ZN(n7753) );
  MUX2_X1 U10049 ( .A(n13147), .B(n14937), .S(n7773), .Z(n7756) );
  MUX2_X1 U10050 ( .A(n13147), .B(n14937), .S(n8148), .Z(n7755) );
  INV_X1 U10051 ( .A(n7756), .ZN(n7757) );
  INV_X1 U10052 ( .A(n7782), .ZN(n7784) );
  NAND2_X1 U10053 ( .A1(n7758), .A2(n10999), .ZN(n7759) );
  NAND2_X1 U10054 ( .A1(n7784), .A2(n7759), .ZN(n11000) );
  INV_X1 U10055 ( .A(n7815), .ZN(n7791) );
  OAI22_X1 U10056 ( .A1(n11000), .A2(n8139), .B1(n7791), .B2(n14477), .ZN(
        n7761) );
  INV_X1 U10057 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n13198) );
  INV_X1 U10058 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13180) );
  OAI22_X1 U10059 ( .A1(n8162), .A2(n13198), .B1(n7709), .B2(n13180), .ZN(
        n7760) );
  MUX2_X1 U10060 ( .A(n10092), .B(n10097), .S(n9961), .Z(n7765) );
  INV_X1 U10061 ( .A(n7765), .ZN(n7766) );
  NAND2_X1 U10062 ( .A1(n7766), .A2(SI_12_), .ZN(n7767) );
  XNOR2_X1 U10063 ( .A(n7792), .B(n7449), .ZN(n10091) );
  NAND2_X1 U10064 ( .A1(n10091), .A2(n8097), .ZN(n7772) );
  NAND2_X1 U10065 ( .A1(n7796), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7769) );
  XNOR2_X1 U10066 ( .A(n7769), .B(n7797), .ZN(n14796) );
  OAI22_X1 U10067 ( .A1(n14796), .A2(n7161), .B1(n7870), .B2(n10097), .ZN(
        n7770) );
  INV_X1 U10068 ( .A(n7770), .ZN(n7771) );
  MUX2_X1 U10069 ( .A(n13146), .B(n11003), .S(n8170), .Z(n7777) );
  NAND2_X1 U10070 ( .A1(n7776), .A2(n7777), .ZN(n7775) );
  MUX2_X1 U10071 ( .A(n13146), .B(n11003), .S(n7773), .Z(n7774) );
  NAND2_X1 U10072 ( .A1(n7775), .A2(n7774), .ZN(n7781) );
  INV_X1 U10073 ( .A(n7776), .ZN(n7779) );
  INV_X1 U10074 ( .A(n7777), .ZN(n7778) );
  INV_X1 U10075 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U10076 ( .A1(n7782), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7812) );
  INV_X1 U10077 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U10078 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  NAND2_X1 U10079 ( .A1(n7812), .A2(n7785), .ZN(n11408) );
  OR2_X1 U10080 ( .A1(n11408), .A2(n8139), .ZN(n7789) );
  NAND2_X1 U10081 ( .A1(n8157), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10082 ( .A1(n8138), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7786) );
  AND2_X1 U10083 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  OAI211_X1 U10084 ( .C1(n7791), .C2(n7790), .A(n7789), .B(n7788), .ZN(n13145)
         );
  NAND2_X1 U10085 ( .A1(n7792), .A2(n7449), .ZN(n7794) );
  MUX2_X1 U10086 ( .A(n10243), .B(n10224), .S(n9961), .Z(n7818) );
  XNOR2_X1 U10087 ( .A(n7818), .B(SI_13_), .ZN(n7795) );
  XNOR2_X1 U10088 ( .A(n7819), .B(n7795), .ZN(n10223) );
  NAND2_X1 U10089 ( .A1(n10223), .A2(n8097), .ZN(n7806) );
  INV_X1 U10090 ( .A(n7796), .ZN(n7798) );
  NAND2_X1 U10091 ( .A1(n7798), .A2(n7797), .ZN(n7800) );
  NAND2_X1 U10092 ( .A1(n7800), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7799) );
  MUX2_X1 U10093 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7799), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7803) );
  INV_X1 U10094 ( .A(n7800), .ZN(n7802) );
  INV_X1 U10095 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U10096 ( .A1(n7802), .A2(n7801), .ZN(n7840) );
  NOR2_X1 U10097 ( .A1(n7870), .A2(n10224), .ZN(n7804) );
  AOI21_X1 U10098 ( .B1(n14817), .B2(n7572), .A(n7804), .ZN(n7805) );
  MUX2_X1 U10099 ( .A(n13145), .B(n13641), .S(n7773), .Z(n7809) );
  MUX2_X1 U10100 ( .A(n13145), .B(n13641), .S(n8170), .Z(n7808) );
  INV_X1 U10101 ( .A(n7809), .ZN(n7810) );
  INV_X1 U10102 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U10103 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  NAND2_X1 U10104 ( .A1(n7827), .A2(n7813), .ZN(n12048) );
  AOI22_X1 U10105 ( .A1(n8138), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n8157), .B2(
        P2_REG2_REG_14__SCAN_IN), .ZN(n7817) );
  NAND2_X1 U10106 ( .A1(n8158), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7816) );
  OAI211_X1 U10107 ( .C1(n12048), .C2(n8139), .A(n7817), .B(n7816), .ZN(n13257) );
  MUX2_X1 U10108 ( .A(n10447), .B(n10421), .S(n9961), .Z(n7858) );
  NAND2_X1 U10109 ( .A1(n10420), .A2(n8097), .ZN(n7822) );
  NAND2_X1 U10110 ( .A1(n7840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7820) );
  XNOR2_X1 U10111 ( .A(n7820), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14822) );
  AOI22_X1 U10112 ( .A1(n14822), .A2(n7572), .B1(n8167), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n7821) );
  NAND2_X2 U10113 ( .A1(n7822), .A2(n7821), .ZN(n13636) );
  MUX2_X1 U10114 ( .A(n13257), .B(n13636), .S(n8148), .Z(n7825) );
  MUX2_X1 U10115 ( .A(n13257), .B(n13636), .S(n7773), .Z(n7823) );
  INV_X1 U10116 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7826) );
  INV_X1 U10117 ( .A(n7847), .ZN(n7874) );
  NAND2_X1 U10118 ( .A1(n7827), .A2(n7826), .ZN(n7828) );
  NAND2_X1 U10119 ( .A1(n7874), .A2(n7828), .ZN(n13498) );
  OR2_X1 U10120 ( .A1(n13498), .A2(n8139), .ZN(n7834) );
  INV_X1 U10121 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U10122 ( .A1(n8158), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10123 ( .A1(n8157), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7829) );
  OAI211_X1 U10124 ( .C1(n8162), .C2(n7831), .A(n7830), .B(n7829), .ZN(n7832)
         );
  INV_X1 U10125 ( .A(n7832), .ZN(n7833) );
  NAND2_X1 U10126 ( .A1(n7835), .A2(n7858), .ZN(n7837) );
  NAND2_X1 U10127 ( .A1(n7857), .A2(n10042), .ZN(n7836) );
  MUX2_X1 U10128 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9961), .Z(n7854) );
  INV_X1 U10129 ( .A(n7854), .ZN(n7860) );
  XNOR2_X1 U10130 ( .A(n7860), .B(SI_15_), .ZN(n7838) );
  NAND2_X1 U10131 ( .A1(n10451), .A2(n8097), .ZN(n7843) );
  OAI21_X1 U10132 ( .B1(n7840), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7841) );
  XNOR2_X1 U10133 ( .A(n7841), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13203) );
  AOI22_X1 U10134 ( .A1(n13203), .A2(n7572), .B1(n8167), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7842) );
  MUX2_X1 U10135 ( .A(n13261), .B(n13629), .S(n8148), .Z(n7892) );
  INV_X1 U10136 ( .A(n13261), .ZN(n13480) );
  MUX2_X1 U10137 ( .A(n13480), .B(n13513), .S(n7773), .Z(n7891) );
  NAND2_X1 U10138 ( .A1(n7892), .A2(n7891), .ZN(n7889) );
  INV_X1 U10139 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7845) );
  INV_X1 U10140 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7844) );
  OAI21_X1 U10141 ( .B1(n7874), .B2(n7845), .A(n7844), .ZN(n7848) );
  AND2_X1 U10142 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n7846) );
  INV_X1 U10143 ( .A(n7900), .ZN(n7901) );
  AND2_X1 U10144 ( .A1(n7848), .A2(n7901), .ZN(n13050) );
  NAND2_X1 U10145 ( .A1(n13050), .A2(n8050), .ZN(n7853) );
  INV_X1 U10146 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13207) );
  NAND2_X1 U10147 ( .A1(n8157), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10148 ( .A1(n8158), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7849) );
  OAI211_X1 U10149 ( .C1(n13207), .C2(n8162), .A(n7850), .B(n7849), .ZN(n7851)
         );
  INV_X1 U10150 ( .A(n7851), .ZN(n7852) );
  NAND2_X1 U10151 ( .A1(n7853), .A2(n7852), .ZN(n13481) );
  NAND2_X1 U10152 ( .A1(n7854), .A2(SI_15_), .ZN(n7861) );
  OAI21_X1 U10153 ( .B1(n10042), .B2(n7858), .A(n7861), .ZN(n7855) );
  INV_X1 U10154 ( .A(n7855), .ZN(n7856) );
  INV_X1 U10155 ( .A(n7858), .ZN(n7859) );
  NOR2_X1 U10156 ( .A1(n7859), .A2(SI_14_), .ZN(n7862) );
  AOI22_X1 U10157 ( .A1(n7862), .A2(n7861), .B1(n10058), .B2(n7860), .ZN(n7863) );
  MUX2_X1 U10158 ( .A(n10422), .B(n10401), .S(n9961), .Z(n7864) );
  XNOR2_X1 U10159 ( .A(n7864), .B(SI_16_), .ZN(n7880) );
  MUX2_X1 U10160 ( .A(n10449), .B(n10446), .S(n9961), .Z(n7909) );
  XNOR2_X1 U10161 ( .A(n7909), .B(SI_17_), .ZN(n7865) );
  XNOR2_X1 U10162 ( .A(n7913), .B(n7865), .ZN(n10445) );
  NAND2_X1 U10163 ( .A1(n10445), .A2(n8097), .ZN(n7873) );
  NAND2_X1 U10164 ( .A1(n7867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7868) );
  MUX2_X1 U10165 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7868), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7869) );
  NAND2_X1 U10166 ( .A1(n7869), .A2(n7914), .ZN(n14865) );
  OAI22_X1 U10167 ( .A1(n14865), .A2(n7161), .B1(n7870), .B2(n10446), .ZN(
        n7871) );
  INV_X1 U10168 ( .A(n7871), .ZN(n7872) );
  MUX2_X1 U10169 ( .A(n13481), .B(n13618), .S(n7773), .Z(n7894) );
  NAND2_X1 U10170 ( .A1(n13618), .A2(n13481), .ZN(n13266) );
  XNOR2_X1 U10171 ( .A(n7874), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n13484) );
  NAND2_X1 U10172 ( .A1(n13484), .A2(n8050), .ZN(n7879) );
  INV_X1 U10173 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13488) );
  NAND2_X1 U10174 ( .A1(n8138), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10175 ( .A1(n8158), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7875) );
  OAI211_X1 U10176 ( .C1(n7709), .C2(n13488), .A(n7876), .B(n7875), .ZN(n7877)
         );
  INV_X1 U10177 ( .A(n7877), .ZN(n7878) );
  NAND2_X1 U10178 ( .A1(n7879), .A2(n7878), .ZN(n13264) );
  AND2_X1 U10179 ( .A1(n13264), .A2(n8148), .ZN(n7887) );
  NOR2_X1 U10180 ( .A1(n13264), .A2(n8170), .ZN(n7886) );
  XNOR2_X1 U10181 ( .A(n7881), .B(n7880), .ZN(n10400) );
  NAND2_X1 U10182 ( .A1(n10400), .A2(n8097), .ZN(n7885) );
  NAND2_X1 U10183 ( .A1(n7882), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7883) );
  XNOR2_X1 U10184 ( .A(n7883), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13172) );
  AOI22_X1 U10185 ( .A1(n6499), .A2(n13172), .B1(n8167), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n7884) );
  MUX2_X1 U10186 ( .A(n7887), .B(n7886), .S(n13485), .Z(n7888) );
  AOI21_X1 U10187 ( .B1(n7894), .B2(n13266), .A(n7888), .ZN(n7896) );
  XNOR2_X1 U10188 ( .A(n13485), .B(n13264), .ZN(n13494) );
  OAI21_X1 U10189 ( .B1(n7892), .B2(n7891), .A(n13494), .ZN(n7897) );
  NOR2_X1 U10190 ( .A1(n13618), .A2(n13481), .ZN(n7893) );
  NOR2_X1 U10191 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  AOI21_X1 U10192 ( .B1(n7897), .B2(n7896), .A(n7895), .ZN(n7898) );
  OAI21_X1 U10193 ( .B1(n7453), .B2(n7899), .A(n7898), .ZN(n7919) );
  INV_X1 U10194 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n14871) );
  NAND2_X1 U10195 ( .A1(n7901), .A2(n14871), .ZN(n7902) );
  NAND2_X1 U10196 ( .A1(n7921), .A2(n7902), .ZN(n13448) );
  OR2_X1 U10197 ( .A1(n13448), .A2(n8139), .ZN(n7908) );
  INV_X1 U10198 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U10199 ( .A1(n8157), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10200 ( .A1(n8158), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7903) );
  OAI211_X1 U10201 ( .C1(n8162), .C2(n7905), .A(n7904), .B(n7903), .ZN(n7906)
         );
  INV_X1 U10202 ( .A(n7906), .ZN(n7907) );
  NAND2_X1 U10203 ( .A1(n7908), .A2(n7907), .ZN(n13267) );
  NOR2_X1 U10204 ( .A1(n7910), .A2(SI_17_), .ZN(n7912) );
  NAND2_X1 U10205 ( .A1(n7910), .A2(SI_17_), .ZN(n7911) );
  MUX2_X1 U10206 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9961), .Z(n7930) );
  XNOR2_X1 U10207 ( .A(n7929), .B(n7930), .ZN(n10718) );
  NAND2_X1 U10208 ( .A1(n10718), .A2(n8097), .ZN(n7917) );
  NAND2_X1 U10209 ( .A1(n7914), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7915) );
  XNOR2_X1 U10210 ( .A(n7915), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U10211 ( .A1(n13209), .A2(n7572), .B1(n8167), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n7916) );
  MUX2_X1 U10212 ( .A(n13267), .B(n13612), .S(n8170), .Z(n7920) );
  MUX2_X1 U10213 ( .A(n13267), .B(n13612), .S(n7773), .Z(n7918) );
  NAND2_X1 U10214 ( .A1(n7921), .A2(n11689), .ZN(n7922) );
  NAND2_X1 U10215 ( .A1(n7946), .A2(n7922), .ZN(n13439) );
  OR2_X1 U10216 ( .A1(n13439), .A2(n8139), .ZN(n7928) );
  INV_X1 U10217 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U10218 ( .A1(n8158), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U10219 ( .A1(n8157), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7923) );
  OAI211_X1 U10220 ( .C1(n8162), .C2(n7925), .A(n7924), .B(n7923), .ZN(n7926)
         );
  INV_X1 U10221 ( .A(n7926), .ZN(n7927) );
  NAND2_X1 U10222 ( .A1(n7928), .A2(n7927), .ZN(n13270) );
  NAND2_X1 U10223 ( .A1(n7931), .A2(SI_18_), .ZN(n7932) );
  MUX2_X1 U10224 ( .A(n10787), .B(n10789), .S(n9961), .Z(n7933) );
  INV_X1 U10225 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U10226 ( .A1(n7934), .A2(SI_19_), .ZN(n7935) );
  NAND2_X1 U10227 ( .A1(n7953), .A2(n7935), .ZN(n7954) );
  XNOR2_X1 U10228 ( .A(n7955), .B(n7954), .ZN(n8531) );
  INV_X1 U10229 ( .A(n8531), .ZN(n10788) );
  NAND2_X1 U10230 ( .A1(n8531), .A2(n8097), .ZN(n7937) );
  AOI22_X1 U10231 ( .A1(n6469), .A2(n6499), .B1(n8167), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n7936) );
  MUX2_X1 U10232 ( .A(n13270), .B(n13608), .S(n7773), .Z(n7941) );
  MUX2_X1 U10233 ( .A(n13270), .B(n13608), .S(n8170), .Z(n7938) );
  NAND2_X1 U10234 ( .A1(n7939), .A2(n7938), .ZN(n7945) );
  INV_X1 U10235 ( .A(n7940), .ZN(n7943) );
  INV_X1 U10236 ( .A(n7941), .ZN(n7942) );
  NAND2_X1 U10237 ( .A1(n7946), .A2(n13083), .ZN(n7947) );
  NAND2_X1 U10238 ( .A1(n7985), .A2(n7947), .ZN(n13423) );
  INV_X1 U10239 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10240 ( .A1(n8157), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10241 ( .A1(n8158), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7948) );
  OAI211_X1 U10242 ( .C1(n7950), .C2(n8162), .A(n7949), .B(n7948), .ZN(n7951)
         );
  INV_X1 U10243 ( .A(n7951), .ZN(n7952) );
  OAI21_X1 U10244 ( .B1(n13423), .B2(n8139), .A(n7952), .ZN(n13271) );
  XNOR2_X1 U10245 ( .A(n7995), .B(n10578), .ZN(n7967) );
  MUX2_X1 U10246 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9961), .Z(n7996) );
  XNOR2_X1 U10247 ( .A(n7967), .B(n7996), .ZN(n11010) );
  NAND2_X1 U10248 ( .A1(n11010), .A2(n8097), .ZN(n7957) );
  NAND2_X1 U10249 ( .A1(n8167), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7956) );
  NAND2_X2 U10250 ( .A1(n7957), .A2(n7956), .ZN(n13602) );
  MUX2_X1 U10251 ( .A(n13271), .B(n13602), .S(n8148), .Z(n7959) );
  MUX2_X1 U10252 ( .A(n13271), .B(n13602), .S(n7773), .Z(n7958) );
  INV_X1 U10253 ( .A(n7959), .ZN(n7960) );
  XNOR2_X1 U10254 ( .A(n7985), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n13413) );
  NAND2_X1 U10255 ( .A1(n13413), .A2(n8050), .ZN(n7966) );
  INV_X1 U10256 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10257 ( .A1(n8158), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U10258 ( .A1(n8157), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7961) );
  OAI211_X1 U10259 ( .C1(n8162), .C2(n7963), .A(n7962), .B(n7961), .ZN(n7964)
         );
  INV_X1 U10260 ( .A(n7964), .ZN(n7965) );
  NAND2_X1 U10261 ( .A1(n7966), .A2(n7965), .ZN(n13274) );
  INV_X1 U10262 ( .A(n7967), .ZN(n7968) );
  NAND2_X1 U10263 ( .A1(n7968), .A2(n7996), .ZN(n7970) );
  OR2_X1 U10264 ( .A1(n7995), .A2(n10578), .ZN(n7969) );
  NAND2_X1 U10265 ( .A1(n7970), .A2(n7969), .ZN(n7972) );
  MUX2_X1 U10266 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9961), .Z(n7999) );
  XNOR2_X1 U10267 ( .A(n7999), .B(SI_21_), .ZN(n7971) );
  NAND2_X1 U10268 ( .A1(n11234), .A2(n8097), .ZN(n7974) );
  NAND2_X1 U10269 ( .A1(n8167), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7973) );
  MUX2_X1 U10270 ( .A(n13274), .B(n13597), .S(n7773), .Z(n7978) );
  NAND2_X1 U10271 ( .A1(n7977), .A2(n7978), .ZN(n7976) );
  MUX2_X1 U10272 ( .A(n13274), .B(n13597), .S(n8148), .Z(n7975) );
  NAND2_X1 U10273 ( .A1(n7976), .A2(n7975), .ZN(n7982) );
  INV_X1 U10274 ( .A(n7977), .ZN(n7980) );
  INV_X1 U10275 ( .A(n7978), .ZN(n7979) );
  NAND2_X1 U10276 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  NAND2_X1 U10277 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n7983) );
  INV_X1 U10278 ( .A(n8009), .ZN(n7987) );
  INV_X1 U10279 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13031) );
  INV_X1 U10280 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7984) );
  OAI21_X1 U10281 ( .B1(n7985), .B2(n13031), .A(n7984), .ZN(n7986) );
  NAND2_X1 U10282 ( .A1(n7987), .A2(n7986), .ZN(n13400) );
  OR2_X1 U10283 ( .A1(n13400), .A2(n8139), .ZN(n7993) );
  INV_X1 U10284 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10285 ( .A1(n8158), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10286 ( .A1(n8157), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7988) );
  OAI211_X1 U10287 ( .C1(n8162), .C2(n7990), .A(n7989), .B(n7988), .ZN(n7991)
         );
  INV_X1 U10288 ( .A(n7991), .ZN(n7992) );
  NAND2_X1 U10289 ( .A1(n7993), .A2(n7992), .ZN(n13278) );
  NOR2_X1 U10290 ( .A1(n7996), .A2(SI_20_), .ZN(n7994) );
  INV_X1 U10291 ( .A(n7996), .ZN(n7997) );
  NOR2_X1 U10292 ( .A1(n7997), .A2(n10578), .ZN(n8001) );
  INV_X1 U10293 ( .A(n7998), .ZN(n8000) );
  AOI22_X1 U10294 ( .A1(n8001), .A2(n8000), .B1(n7999), .B2(SI_21_), .ZN(n8002) );
  MUX2_X1 U10295 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9961), .Z(n8016) );
  XNOR2_X1 U10296 ( .A(n8566), .B(n8016), .ZN(n11251) );
  NAND2_X1 U10297 ( .A1(n11251), .A2(n8097), .ZN(n8005) );
  NAND2_X1 U10298 ( .A1(n8167), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8004) );
  MUX2_X1 U10299 ( .A(n13278), .B(n13591), .S(n8148), .Z(n8007) );
  MUX2_X1 U10300 ( .A(n13278), .B(n13591), .S(n7773), .Z(n8006) );
  INV_X1 U10301 ( .A(n8007), .ZN(n8008) );
  NOR2_X1 U10302 ( .A1(n8009), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8010) );
  OR2_X1 U10303 ( .A1(n8031), .A2(n8010), .ZN(n12041) );
  INV_X1 U10304 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10305 ( .A1(n8158), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10306 ( .A1(n8157), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8011) );
  OAI211_X1 U10307 ( .C1(n8162), .C2(n8013), .A(n8012), .B(n8011), .ZN(n8014)
         );
  INV_X1 U10308 ( .A(n8014), .ZN(n8015) );
  OAI21_X1 U10309 ( .B1(n12041), .B2(n8139), .A(n8015), .ZN(n13280) );
  NAND2_X1 U10310 ( .A1(n8017), .A2(SI_22_), .ZN(n8018) );
  MUX2_X1 U10311 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9961), .Z(n8041) );
  XNOR2_X1 U10312 ( .A(n8041), .B(SI_23_), .ZN(n8020) );
  XNOR2_X1 U10313 ( .A(n8040), .B(n8020), .ZN(n11318) );
  NAND2_X1 U10314 ( .A1(n11318), .A2(n8097), .ZN(n8022) );
  NAND2_X1 U10315 ( .A1(n8167), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8021) );
  MUX2_X1 U10316 ( .A(n13280), .B(n13383), .S(n7773), .Z(n8026) );
  NAND2_X1 U10317 ( .A1(n8025), .A2(n8026), .ZN(n8024) );
  MUX2_X1 U10318 ( .A(n13280), .B(n13383), .S(n8170), .Z(n8023) );
  NAND2_X1 U10319 ( .A1(n8024), .A2(n8023), .ZN(n8030) );
  INV_X1 U10320 ( .A(n8025), .ZN(n8028) );
  INV_X1 U10321 ( .A(n8026), .ZN(n8027) );
  OR2_X1 U10322 ( .A1(n8031), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10323 ( .A1(n8032), .A2(n8048), .ZN(n13366) );
  INV_X1 U10324 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10325 ( .A1(n8158), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8034) );
  NAND2_X1 U10326 ( .A1(n8157), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8033) );
  OAI211_X1 U10327 ( .C1(n8162), .C2(n8035), .A(n8034), .B(n8033), .ZN(n8036)
         );
  INV_X1 U10328 ( .A(n8036), .ZN(n8037) );
  INV_X1 U10329 ( .A(n8041), .ZN(n8038) );
  NAND2_X1 U10330 ( .A1(n8038), .A2(n10847), .ZN(n8039) );
  NAND2_X1 U10331 ( .A1(n8041), .A2(SI_23_), .ZN(n8042) );
  MUX2_X1 U10332 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6492), .Z(n8056) );
  NAND2_X1 U10333 ( .A1(n11439), .A2(n8097), .ZN(n8044) );
  NAND2_X1 U10334 ( .A1(n8167), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8043) );
  NAND2_X2 U10335 ( .A1(n8044), .A2(n8043), .ZN(n13578) );
  MUX2_X1 U10336 ( .A(n13347), .B(n13578), .S(n8148), .Z(n8046) );
  MUX2_X1 U10337 ( .A(n13347), .B(n13578), .S(n7773), .Z(n8045) );
  INV_X1 U10338 ( .A(n8046), .ZN(n8047) );
  NAND2_X1 U10339 ( .A1(n8157), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U10340 ( .A1(n8138), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8053) );
  INV_X1 U10341 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8049) );
  AOI21_X1 U10342 ( .B1(n8049), .B2(n8048), .A(n8073), .ZN(n13354) );
  NAND2_X1 U10343 ( .A1(n8050), .A2(n13354), .ZN(n8052) );
  NAND2_X1 U10344 ( .A1(n8158), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8051) );
  NAND4_X1 U10345 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), .ZN(n13282) );
  NAND2_X1 U10346 ( .A1(n8057), .A2(SI_24_), .ZN(n8058) );
  INV_X1 U10347 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11476) );
  INV_X1 U10348 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11480) );
  MUX2_X1 U10349 ( .A(n11476), .B(n11480), .S(n9961), .Z(n8060) );
  NAND2_X1 U10350 ( .A1(n8060), .A2(n11281), .ZN(n8078) );
  INV_X1 U10351 ( .A(n8060), .ZN(n8061) );
  NAND2_X1 U10352 ( .A1(n8061), .A2(SI_25_), .ZN(n8062) );
  NAND2_X1 U10353 ( .A1(n8078), .A2(n8062), .ZN(n8079) );
  NAND2_X1 U10354 ( .A1(n11475), .A2(n8097), .ZN(n8064) );
  NAND2_X1 U10355 ( .A1(n8167), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8063) );
  MUX2_X1 U10356 ( .A(n13282), .B(n13572), .S(n7773), .Z(n8068) );
  NAND2_X1 U10357 ( .A1(n8067), .A2(n8068), .ZN(n8066) );
  MUX2_X1 U10358 ( .A(n13282), .B(n13572), .S(n8148), .Z(n8065) );
  NAND2_X1 U10359 ( .A1(n8066), .A2(n8065), .ZN(n8072) );
  INV_X1 U10360 ( .A(n8067), .ZN(n8070) );
  INV_X1 U10361 ( .A(n8068), .ZN(n8069) );
  NAND2_X1 U10362 ( .A1(n8070), .A2(n8069), .ZN(n8071) );
  NAND2_X1 U10363 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8073), .ZN(n8087) );
  OAI21_X1 U10364 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n8073), .A(n8087), .ZN(
        n13335) );
  OR2_X1 U10365 ( .A1(n8139), .A2(n13335), .ZN(n8077) );
  NAND2_X1 U10366 ( .A1(n8157), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10367 ( .A1(n8138), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U10368 ( .A1(n8158), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8074) );
  NAND4_X1 U10369 ( .A1(n8077), .A2(n8076), .A3(n8075), .A4(n8074), .ZN(n13346) );
  INV_X1 U10370 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14364) );
  INV_X1 U10371 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13689) );
  MUX2_X1 U10372 ( .A(n14364), .B(n13689), .S(n6492), .Z(n8093) );
  XNOR2_X1 U10373 ( .A(n8093), .B(SI_26_), .ZN(n8081) );
  XNOR2_X1 U10374 ( .A(n8094), .B(n8081), .ZN(n13687) );
  NAND2_X1 U10375 ( .A1(n13687), .A2(n8097), .ZN(n8083) );
  NAND2_X1 U10376 ( .A1(n8167), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8082) );
  MUX2_X1 U10377 ( .A(n13346), .B(n13566), .S(n8148), .Z(n8085) );
  MUX2_X1 U10378 ( .A(n13346), .B(n13566), .S(n7773), .Z(n8084) );
  NAND2_X1 U10379 ( .A1(n8157), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10380 ( .A1(n8138), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U10381 ( .A1(n8158), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8090) );
  INV_X1 U10382 ( .A(n8087), .ZN(n8086) );
  INV_X1 U10383 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U10384 ( .A1(n8087), .A2(n13013), .ZN(n8088) );
  NAND2_X1 U10385 ( .A1(n8102), .A2(n8088), .ZN(n13322) );
  OR2_X1 U10386 ( .A1(n8139), .A2(n13322), .ZN(n8089) );
  MUX2_X1 U10387 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6492), .Z(n8108) );
  INV_X1 U10388 ( .A(n8108), .ZN(n8095) );
  XNOR2_X1 U10389 ( .A(n8095), .B(SI_27_), .ZN(n8096) );
  NAND2_X1 U10390 ( .A1(n11655), .A2(n8097), .ZN(n8099) );
  NAND2_X1 U10391 ( .A1(n8167), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8098) );
  MUX2_X1 U10392 ( .A(n13284), .B(n13319), .S(n7773), .Z(n8117) );
  NAND2_X1 U10393 ( .A1(n8138), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U10394 ( .A1(n8157), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10395 ( .A1(n8158), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10396 ( .A1(n8100), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13290) );
  INV_X1 U10397 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U10398 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  NAND2_X1 U10399 ( .A1(n13290), .A2(n8103), .ZN(n13303) );
  OR2_X1 U10400 ( .A1(n8139), .A2(n13303), .ZN(n8104) );
  NOR2_X1 U10401 ( .A1(n8108), .A2(SI_27_), .ZN(n8110) );
  NAND2_X1 U10402 ( .A1(n8108), .A2(SI_27_), .ZN(n8109) );
  INV_X1 U10403 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12037) );
  INV_X1 U10404 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9720) );
  MUX2_X1 U10405 ( .A(n12037), .B(n9720), .S(n6492), .Z(n8112) );
  INV_X1 U10406 ( .A(SI_28_), .ZN(n12321) );
  NAND2_X1 U10407 ( .A1(n8112), .A2(n12321), .ZN(n8123) );
  INV_X1 U10408 ( .A(n8112), .ZN(n8113) );
  NAND2_X1 U10409 ( .A1(n8113), .A2(SI_28_), .ZN(n8114) );
  NAND2_X1 U10410 ( .A1(n8123), .A2(n8114), .ZN(n8121) );
  NAND2_X1 U10411 ( .A1(n12036), .A2(n8097), .ZN(n8116) );
  NAND2_X1 U10412 ( .A1(n8167), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8115) );
  MUX2_X1 U10413 ( .A(n11740), .B(n13308), .S(n7773), .Z(n8153) );
  MUX2_X1 U10414 ( .A(n13285), .B(n13555), .S(n8148), .Z(n8152) );
  NAND2_X1 U10415 ( .A1(n8118), .A2(n6684), .ZN(n8120) );
  INV_X1 U10416 ( .A(n13284), .ZN(n13249) );
  MUX2_X1 U10417 ( .A(n13249), .B(n13561), .S(n8148), .Z(n8119) );
  NAND2_X1 U10418 ( .A1(n8120), .A2(n8119), .ZN(n8150) );
  MUX2_X1 U10419 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6492), .Z(n8124) );
  XNOR2_X1 U10420 ( .A(n8124), .B(n12388), .ZN(n8144) );
  INV_X1 U10421 ( .A(n8124), .ZN(n8125) );
  NAND2_X1 U10422 ( .A1(n8125), .A2(n12388), .ZN(n8126) );
  NAND2_X1 U10423 ( .A1(n8127), .A2(n8126), .ZN(n8164) );
  MUX2_X1 U10424 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6492), .Z(n8128) );
  NAND2_X1 U10425 ( .A1(n8128), .A2(SI_30_), .ZN(n8129) );
  OAI21_X1 U10426 ( .B1(SI_30_), .B2(n8128), .A(n8129), .ZN(n8163) );
  MUX2_X1 U10427 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6492), .Z(n8130) );
  XNOR2_X1 U10428 ( .A(n8130), .B(SI_31_), .ZN(n8131) );
  NAND2_X1 U10429 ( .A1(n13670), .A2(n8097), .ZN(n8134) );
  NAND2_X1 U10430 ( .A1(n8167), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8133) );
  INV_X1 U10431 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10432 ( .A1(n8157), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10433 ( .A1(n8158), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8135) );
  OAI211_X1 U10434 ( .C1(n8162), .C2(n8137), .A(n8136), .B(n8135), .ZN(n13226)
         );
  NAND2_X1 U10435 ( .A1(n8157), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10436 ( .A1(n8158), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10437 ( .A1(n8138), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8141) );
  OR2_X1 U10438 ( .A1(n8139), .A2(n13290), .ZN(n8140) );
  AND4_X1 U10439 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n11746)
         );
  NAND2_X1 U10440 ( .A1(n13678), .A2(n8097), .ZN(n8147) );
  NAND2_X1 U10441 ( .A1(n8167), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8146) );
  MUX2_X1 U10442 ( .A(n11746), .B(n13550), .S(n7773), .Z(n8175) );
  MUX2_X1 U10443 ( .A(n13144), .B(n13293), .S(n8148), .Z(n8174) );
  NAND2_X1 U10444 ( .A1(n8175), .A2(n8174), .ZN(n8155) );
  NAND3_X1 U10445 ( .A1(n8151), .A2(n8150), .A3(n8149), .ZN(n8179) );
  INV_X1 U10446 ( .A(n8152), .ZN(n8156) );
  INV_X1 U10447 ( .A(n8153), .ZN(n8154) );
  NAND4_X1 U10448 ( .A1(n8203), .A2(n8156), .A3(n8155), .A4(n8154), .ZN(n8178)
         );
  INV_X1 U10449 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U10450 ( .A1(n8157), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U10451 ( .A1(n8158), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8159) );
  OAI211_X1 U10452 ( .C1(n8162), .C2(n8161), .A(n8160), .B(n8159), .ZN(n13254)
         );
  NAND2_X1 U10453 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  NAND2_X1 U10454 ( .A1(n8167), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8168) );
  MUX2_X1 U10455 ( .A(n13254), .B(n13229), .S(n8170), .Z(n8181) );
  OR2_X1 U10456 ( .A1(n10265), .A2(n10144), .ZN(n8206) );
  NAND2_X1 U10457 ( .A1(n8170), .A2(n13226), .ZN(n8171) );
  NAND4_X1 U10458 ( .A1(n8206), .A2(n8237), .A3(n10334), .A4(n8171), .ZN(n8172) );
  AND2_X1 U10459 ( .A1(n8172), .A2(n13254), .ZN(n8173) );
  AOI21_X1 U10460 ( .B1(n13229), .B2(n7773), .A(n8173), .ZN(n8180) );
  OAI22_X1 U10461 ( .A1(n8181), .A2(n8180), .B1(n8175), .B2(n8174), .ZN(n8176)
         );
  NAND2_X1 U10462 ( .A1(n8176), .A2(n8203), .ZN(n8177) );
  NAND3_X1 U10463 ( .A1(n8179), .A2(n8178), .A3(n8177), .ZN(n8185) );
  NAND2_X1 U10464 ( .A1(n8181), .A2(n8180), .ZN(n8184) );
  MUX2_X1 U10465 ( .A(n13226), .B(n13543), .S(n7773), .Z(n8182) );
  NOR2_X1 U10466 ( .A1(n6553), .A2(n8182), .ZN(n8183) );
  INV_X1 U10467 ( .A(n10265), .ZN(n10269) );
  NAND2_X1 U10468 ( .A1(n13555), .A2(n11740), .ZN(n8186) );
  INV_X1 U10469 ( .A(n13346), .ZN(n13283) );
  OR2_X1 U10470 ( .A1(n13566), .A2(n13283), .ZN(n13248) );
  NAND2_X1 U10471 ( .A1(n13566), .A2(n13283), .ZN(n13246) );
  INV_X1 U10472 ( .A(n13280), .ZN(n13065) );
  NAND2_X1 U10473 ( .A1(n13383), .A2(n13065), .ZN(n13244) );
  OR2_X1 U10474 ( .A1(n13383), .A2(n13065), .ZN(n8187) );
  NAND2_X1 U10475 ( .A1(n13244), .A2(n8187), .ZN(n13381) );
  INV_X1 U10476 ( .A(n13274), .ZN(n13242) );
  XNOR2_X1 U10477 ( .A(n13597), .B(n13242), .ZN(n13408) );
  INV_X1 U10478 ( .A(n13278), .ZN(n13030) );
  XNOR2_X1 U10479 ( .A(n13591), .B(n13030), .ZN(n13388) );
  XNOR2_X1 U10480 ( .A(n13602), .B(n13271), .ZN(n13427) );
  INV_X1 U10481 ( .A(n13257), .ZN(n13504) );
  XNOR2_X1 U10482 ( .A(n13636), .B(n13504), .ZN(n11269) );
  INV_X1 U10483 ( .A(n13481), .ZN(n13238) );
  XNOR2_X1 U10484 ( .A(n13618), .B(n13238), .ZN(n13464) );
  INV_X1 U10485 ( .A(n13145), .ZN(n12049) );
  OR2_X1 U10486 ( .A1(n13641), .A2(n12049), .ZN(n11264) );
  NAND2_X1 U10487 ( .A1(n13641), .A2(n12049), .ZN(n8188) );
  INV_X1 U10488 ( .A(n13147), .ZN(n11005) );
  NAND2_X1 U10489 ( .A1(n14937), .A2(n11005), .ZN(n10874) );
  OR2_X1 U10490 ( .A1(n14937), .A2(n11005), .ZN(n8189) );
  NAND2_X1 U10491 ( .A1(n10874), .A2(n8189), .ZN(n10793) );
  INV_X1 U10492 ( .A(n13148), .ZN(n14456) );
  INV_X1 U10493 ( .A(n13149), .ZN(n10868) );
  XNOR2_X1 U10494 ( .A(n11703), .B(n10868), .ZN(n10758) );
  XNOR2_X1 U10495 ( .A(n12070), .B(n13151), .ZN(n10729) );
  INV_X1 U10496 ( .A(n13524), .ZN(n10543) );
  OR2_X1 U10497 ( .A1(n13076), .A2(n13153), .ZN(n10471) );
  NAND2_X1 U10498 ( .A1(n13076), .A2(n13153), .ZN(n8190) );
  INV_X1 U10499 ( .A(n13154), .ZN(n10476) );
  INV_X1 U10500 ( .A(n13155), .ZN(n10236) );
  NAND2_X1 U10501 ( .A1(n10591), .A2(n10236), .ZN(n10232) );
  INV_X1 U10502 ( .A(n10591), .ZN(n8191) );
  NAND2_X1 U10503 ( .A1(n8191), .A2(n13155), .ZN(n8192) );
  NAND2_X1 U10504 ( .A1(n13157), .A2(n10354), .ZN(n10225) );
  OAI21_X1 U10505 ( .B1(n13157), .B2(n10354), .A(n10225), .ZN(n13647) );
  NAND4_X1 U10506 ( .A1(n10438), .A2(n8205), .A3(n10227), .A4(n13647), .ZN(
        n8194) );
  NOR4_X1 U10507 ( .A1(n10481), .A2(n10508), .A3(n10233), .A4(n8194), .ZN(
        n8195) );
  XNOR2_X1 U10508 ( .A(n14919), .B(n13522), .ZN(n10632) );
  XNOR2_X1 U10509 ( .A(n14912), .B(n13152), .ZN(n13533) );
  NAND4_X1 U10510 ( .A1(n10729), .A2(n8195), .A3(n10632), .A4(n13533), .ZN(
        n8196) );
  NOR4_X1 U10511 ( .A1(n10793), .A2(n10794), .A3(n10758), .A4(n8196), .ZN(
        n8197) );
  XNOR2_X1 U10512 ( .A(n11003), .B(n13146), .ZN(n10881) );
  NAND4_X1 U10513 ( .A1(n10991), .A2(n13494), .A3(n8197), .A4(n10881), .ZN(
        n8198) );
  NOR4_X1 U10514 ( .A1(n13508), .A2(n11269), .A3(n13464), .A4(n8198), .ZN(
        n8199) );
  XNOR2_X1 U10515 ( .A(n13612), .B(n13267), .ZN(n13455) );
  NAND4_X1 U10516 ( .A1(n13427), .A2(n8199), .A3(n13433), .A4(n13455), .ZN(
        n8200) );
  NOR4_X1 U10517 ( .A1(n13381), .A2(n13408), .A3(n13388), .A4(n8200), .ZN(
        n8201) );
  XNOR2_X1 U10518 ( .A(n13572), .B(n13282), .ZN(n13344) );
  NAND4_X1 U10519 ( .A1(n13338), .A2(n8201), .A3(n13344), .A4(n13363), .ZN(
        n8202) );
  XNOR2_X1 U10520 ( .A(n13293), .B(n13144), .ZN(n13286) );
  NAND2_X1 U10521 ( .A1(n8237), .A2(n8205), .ZN(n10151) );
  OAI21_X1 U10522 ( .B1(n10151), .B2(n13216), .A(n8206), .ZN(n8207) );
  INV_X1 U10523 ( .A(n8207), .ZN(n8212) );
  INV_X1 U10524 ( .A(n8208), .ZN(n8209) );
  OAI211_X1 U10525 ( .C1(n6469), .C2(n11235), .A(n10334), .B(n8209), .ZN(n8210) );
  NAND2_X1 U10526 ( .A1(n8213), .A2(n8210), .ZN(n8211) );
  OAI21_X1 U10527 ( .B1(n8213), .B2(n8212), .A(n8211), .ZN(n8221) );
  INV_X1 U10528 ( .A(n8225), .ZN(n8218) );
  NAND2_X1 U10529 ( .A1(n8218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8219) );
  XNOR2_X1 U10530 ( .A(n8219), .B(P2_IR_REG_23__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U10531 ( .A1(n8238), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11321) );
  INV_X1 U10532 ( .A(n11321), .ZN(n8220) );
  NAND2_X1 U10533 ( .A1(n8229), .A2(n8226), .ZN(n8232) );
  NAND2_X1 U10534 ( .A1(n8232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8227) );
  MUX2_X1 U10535 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8227), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8228) );
  AND2_X1 U10536 ( .A1(n8223), .A2(n8228), .ZN(n10126) );
  INV_X1 U10537 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U10538 ( .A1(n8230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8231) );
  MUX2_X1 U10539 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8231), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8233) );
  NAND2_X1 U10540 ( .A1(n8223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8235) );
  NOR2_X1 U10541 ( .A1(n11440), .A2(n13690), .ZN(n8236) );
  NAND2_X1 U10542 ( .A1(n10126), .A2(n8236), .ZN(n10143) );
  NOR2_X1 U10543 ( .A1(n10143), .A2(n8238), .ZN(n9939) );
  INV_X1 U10544 ( .A(n8238), .ZN(n10142) );
  AOI21_X1 U10545 ( .B1(n10335), .B2(n10142), .A(n7572), .ZN(n8239) );
  OR2_X1 U10546 ( .A1(n9939), .A2(n8239), .ZN(n10032) );
  NOR2_X2 U10547 ( .A1(n10032), .A2(P2_U3088), .ZN(n14849) );
  INV_X1 U10548 ( .A(n14849), .ZN(n10033) );
  NOR4_X1 U10549 ( .A1(n10033), .A2(n10334), .A3(n8240), .A4(n10155), .ZN(
        n8242) );
  OAI21_X1 U10550 ( .B1(n10150), .B2(n11321), .A(P2_B_REG_SCAN_IN), .ZN(n8241)
         );
  OR2_X1 U10551 ( .A1(n8242), .A2(n8241), .ZN(n8243) );
  NAND2_X1 U10552 ( .A1(n8244), .A2(n8243), .ZN(P2_U3328) );
  NAND3_X1 U10553 ( .A1(n8427), .A2(n8246), .A3(n8245), .ZN(n8248) );
  NOR2_X2 U10554 ( .A1(n8248), .A2(n8247), .ZN(n8481) );
  NOR2_X1 U10555 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n8255) );
  NOR2_X1 U10556 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8254) );
  NOR2_X1 U10557 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8253) );
  INV_X1 U10558 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10559 ( .A1(n8706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10560 ( .A1(n12036), .A2(n11971), .ZN(n8264) );
  INV_X1 U10561 ( .A(n8313), .ZN(n8356) );
  NAND2_X1 U10562 ( .A1(n11972), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10563 ( .A1(n8265), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8266) );
  INV_X1 U10564 ( .A(n8267), .ZN(n14352) );
  NAND2_X1 U10565 ( .A1(n6470), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8279) );
  INV_X4 U10566 ( .A(n8363), .ZN(n8647) );
  NAND2_X1 U10567 ( .A1(n8647), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U10568 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8348) );
  NOR2_X1 U10569 ( .A1(n8348), .A2(n8347), .ZN(n8364) );
  NAND2_X1 U10570 ( .A1(n8364), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U10571 ( .A1(n8418), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10572 ( .A1(n8463), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8475) );
  INV_X1 U10573 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8522) );
  INV_X1 U10574 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8538) );
  INV_X1 U10575 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13808) );
  INV_X1 U10576 ( .A(n8581), .ZN(n8271) );
  NAND2_X1 U10577 ( .A1(n8271), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U10578 ( .A1(n8580), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U10579 ( .A1(n8591), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8615) );
  INV_X1 U10580 ( .A(n8615), .ZN(n8603) );
  NAND2_X1 U10581 ( .A1(n8603), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8624) );
  INV_X1 U10582 ( .A(n8624), .ZN(n8614) );
  NAND2_X1 U10583 ( .A1(n8272), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8632) );
  INV_X1 U10584 ( .A(n8272), .ZN(n8274) );
  INV_X1 U10585 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10586 ( .A1(n8274), .A2(n8273), .ZN(n8275) );
  NAND2_X1 U10587 ( .A1(n8605), .A2(n12377), .ZN(n8277) );
  AND2_X2 U10588 ( .A1(n12038), .A2(n14359), .ZN(n8325) );
  NAND2_X1 U10589 ( .A1(n8570), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U10590 ( .A1(n8647), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8285) );
  INV_X1 U10591 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8322) );
  INV_X1 U10592 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U10593 ( .A1(n8322), .A2(n8280), .ZN(n8281) );
  AND2_X1 U10594 ( .A1(n8281), .A2(n8348), .ZN(n10927) );
  NAND2_X1 U10595 ( .A1(n6510), .A2(n10927), .ZN(n8284) );
  NAND2_X1 U10596 ( .A1(n8325), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10597 ( .A1(n8646), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U10598 ( .A1(n8286), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8287) );
  XNOR2_X1 U10599 ( .A(n8287), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14582) );
  AOI22_X1 U10600 ( .A1(n8313), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6509), .B2(
        n14582), .ZN(n8289) );
  NAND2_X1 U10601 ( .A1(n9945), .A2(n8331), .ZN(n8288) );
  INV_X1 U10602 ( .A(n11991), .ZN(n8338) );
  NAND2_X1 U10603 ( .A1(n8323), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10604 ( .A1(n8324), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8291) );
  INV_X1 U10605 ( .A(n8295), .ZN(n9963) );
  NAND2_X1 U10606 ( .A1(n8313), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U10607 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8296) );
  NAND2_X1 U10608 ( .A1(n8535), .A2(n13888), .ZN(n8297) );
  NAND2_X1 U10609 ( .A1(n6510), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10610 ( .A1(n8324), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10611 ( .A1(n8325), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8300) );
  NAND4_X2 U10612 ( .A1(n8302), .A2(n8301), .A3(n8300), .A4(n8299), .ZN(n10303) );
  INV_X1 U10613 ( .A(SI_0_), .ZN(n9958) );
  NOR2_X1 U10614 ( .A1(n9961), .A2(n9958), .ZN(n8303) );
  INV_X1 U10615 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8874) );
  XNOR2_X1 U10616 ( .A(n8303), .B(n8874), .ZN(n14369) );
  MUX2_X1 U10617 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14369), .S(n8304), .Z(n14240)
         );
  NAND2_X1 U10618 ( .A1(n10303), .A2(n14240), .ZN(n14255) );
  NAND2_X1 U10619 ( .A1(n10463), .A2(n8305), .ZN(n8306) );
  NAND2_X1 U10620 ( .A1(n8324), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10621 ( .A1(n8325), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U10622 ( .A1(n8323), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8307) );
  INV_X1 U10623 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14351) );
  OR2_X1 U10624 ( .A1(n8314), .A2(n14351), .ZN(n8315) );
  XNOR2_X1 U10625 ( .A(n8315), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13907) );
  INV_X1 U10626 ( .A(n13907), .ZN(n8316) );
  OR2_X1 U10627 ( .A1(n8304), .A2(n8316), .ZN(n8317) );
  XNOR2_X2 U10628 ( .A(n8319), .B(n11809), .ZN(n11801) );
  NAND2_X1 U10629 ( .A1(n10519), .A2(n11990), .ZN(n8321) );
  INV_X1 U10630 ( .A(n8319), .ZN(n11808) );
  INV_X1 U10631 ( .A(n11809), .ZN(n10653) );
  NAND2_X1 U10632 ( .A1(n11808), .A2(n10653), .ZN(n8320) );
  NAND2_X1 U10633 ( .A1(n6510), .A2(n8322), .ZN(n8330) );
  NAND2_X1 U10634 ( .A1(n6471), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10635 ( .A1(n8324), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10636 ( .A1(n8325), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8326) );
  INV_X1 U10637 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U10638 ( .A1(n8332), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8333) );
  XNOR2_X1 U10639 ( .A(n8333), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13924) );
  NAND2_X1 U10640 ( .A1(n8535), .A2(n13924), .ZN(n8334) );
  NAND2_X1 U10641 ( .A1(n10548), .A2(n11989), .ZN(n8337) );
  NAND2_X1 U10642 ( .A1(n10464), .A2(n10558), .ZN(n8336) );
  INV_X1 U10643 ( .A(n14652), .ZN(n11822) );
  NAND2_X1 U10644 ( .A1(n10572), .A2(n11822), .ZN(n8339) );
  NAND2_X1 U10645 ( .A1(n9965), .A2(n11971), .ZN(n8346) );
  NOR2_X1 U10646 ( .A1(n8341), .A2(n14351), .ZN(n8342) );
  MUX2_X1 U10647 ( .A(n14351), .B(n8342), .S(P1_IR_REG_5__SCAN_IN), .Z(n8344)
         );
  AND2_X1 U10648 ( .A1(n8341), .A2(n8343), .ZN(n8357) );
  OR2_X1 U10649 ( .A1(n8344), .A2(n8357), .ZN(n10125) );
  INV_X1 U10650 ( .A(n10125), .ZN(n10204) );
  AOI22_X1 U10651 ( .A1(n11972), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6509), 
        .B2(n10204), .ZN(n8345) );
  NAND2_X1 U10652 ( .A1(n8647), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10653 ( .A1(n6470), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8352) );
  AND2_X1 U10654 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  NOR2_X1 U10655 ( .A1(n8364), .A2(n8349), .ZN(n10890) );
  NAND2_X1 U10656 ( .A1(n8605), .A2(n10890), .ZN(n8351) );
  NAND2_X1 U10657 ( .A1(n8570), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8350) );
  NAND4_X1 U10658 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n13883) );
  XNOR2_X1 U10659 ( .A(n11829), .B(n13883), .ZN(n11992) );
  INV_X1 U10660 ( .A(n11992), .ZN(n10701) );
  OR2_X1 U10661 ( .A1(n13883), .A2(n11829), .ZN(n8354) );
  NAND2_X1 U10662 ( .A1(n8355), .A2(n8354), .ZN(n10818) );
  NAND2_X1 U10663 ( .A1(n9971), .A2(n11971), .ZN(n8362) );
  INV_X1 U10664 ( .A(n8357), .ZN(n8359) );
  NAND2_X1 U10665 ( .A1(n8359), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8358) );
  MUX2_X1 U10666 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8358), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n8360) );
  AND2_X1 U10667 ( .A1(n8360), .A2(n8374), .ZN(n10247) );
  AOI22_X1 U10668 ( .A1(n11972), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6509), 
        .B2(n10247), .ZN(n8361) );
  NAND2_X1 U10669 ( .A1(n8362), .A2(n8361), .ZN(n11836) );
  NAND2_X1 U10670 ( .A1(n8647), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U10671 ( .A1(n6470), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8368) );
  OR2_X1 U10672 ( .A1(n8364), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8365) );
  AND2_X1 U10673 ( .A1(n8379), .A2(n8365), .ZN(n11207) );
  NAND2_X1 U10674 ( .A1(n8605), .A2(n11207), .ZN(n8367) );
  NAND2_X1 U10675 ( .A1(n8570), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8366) );
  NAND4_X1 U10676 ( .A1(n8369), .A2(n8368), .A3(n8367), .A4(n8366), .ZN(n13882) );
  XNOR2_X1 U10677 ( .A(n11836), .B(n13882), .ZN(n11993) );
  NAND2_X1 U10678 ( .A1(n10818), .A2(n10819), .ZN(n8371) );
  OR2_X1 U10679 ( .A1(n11836), .A2(n13882), .ZN(n8370) );
  NAND2_X1 U10680 ( .A1(n9989), .A2(n11971), .ZN(n8377) );
  NAND2_X1 U10681 ( .A1(n8374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8373) );
  MUX2_X1 U10682 ( .A(n8373), .B(P1_IR_REG_31__SCAN_IN), .S(n8372), .Z(n8375)
         );
  AOI22_X1 U10683 ( .A1(n11972), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6509), 
        .B2(n13939), .ZN(n8376) );
  NAND2_X1 U10684 ( .A1(n8647), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10685 ( .A1(n8570), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10686 ( .A1(n8379), .A2(n8378), .ZN(n8380) );
  AND2_X1 U10687 ( .A1(n8390), .A2(n8380), .ZN(n11396) );
  NAND2_X1 U10688 ( .A1(n8605), .A2(n11396), .ZN(n8382) );
  NAND2_X1 U10689 ( .A1(n6470), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8381) );
  NAND4_X1 U10690 ( .A1(n8384), .A2(n8383), .A3(n8382), .A4(n8381), .ZN(n13880) );
  INV_X1 U10691 ( .A(n13880), .ZN(n11142) );
  XNOR2_X1 U10692 ( .A(n11839), .B(n11142), .ZN(n11997) );
  NAND2_X1 U10693 ( .A1(n10002), .A2(n11971), .ZN(n8388) );
  NAND2_X1 U10694 ( .A1(n8386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8400) );
  XNOR2_X1 U10695 ( .A(n8400), .B(P1_IR_REG_8__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U10696 ( .A1(n11972), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6509), 
        .B2(n13955), .ZN(n8387) );
  NAND2_X1 U10697 ( .A1(n8647), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10698 ( .A1(n8570), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10699 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  NAND2_X1 U10700 ( .A1(n8406), .A2(n8391), .ZN(n11342) );
  INV_X1 U10701 ( .A(n11342), .ZN(n8392) );
  NAND2_X1 U10702 ( .A1(n8605), .A2(n8392), .ZN(n8394) );
  NAND2_X1 U10703 ( .A1(n6470), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8393) );
  NAND4_X1 U10704 ( .A1(n8396), .A2(n8395), .A3(n8394), .A4(n8393), .ZN(n13879) );
  INV_X1 U10705 ( .A(n13879), .ZN(n11185) );
  XNOR2_X1 U10706 ( .A(n14668), .B(n11185), .ZN(n11996) );
  OR2_X1 U10707 ( .A1(n14668), .A2(n13879), .ZN(n8397) );
  NAND2_X1 U10708 ( .A1(n8398), .A2(n8397), .ZN(n11183) );
  NAND2_X1 U10709 ( .A1(n10038), .A2(n11971), .ZN(n8405) );
  INV_X1 U10710 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8399) );
  AOI21_X1 U10711 ( .B1(n8400), .B2(n8399), .A(n14351), .ZN(n8401) );
  NAND2_X1 U10712 ( .A1(n8401), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8403) );
  INV_X1 U10713 ( .A(n8401), .ZN(n8429) );
  INV_X1 U10714 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10715 ( .A1(n8429), .A2(n8402), .ZN(n8414) );
  AOI22_X1 U10716 ( .A1(n11972), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6509), 
        .B2(n13972), .ZN(n8404) );
  NAND2_X2 U10717 ( .A1(n8405), .A2(n8404), .ZN(n11849) );
  NAND2_X1 U10718 ( .A1(n6470), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U10719 ( .A1(n8647), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8410) );
  AND2_X1 U10720 ( .A1(n8406), .A2(n11501), .ZN(n8407) );
  NOR2_X1 U10721 ( .A1(n8418), .A2(n8407), .ZN(n11504) );
  NAND2_X1 U10722 ( .A1(n8605), .A2(n11504), .ZN(n8409) );
  NAND2_X1 U10723 ( .A1(n8570), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8408) );
  NAND4_X1 U10724 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n13878) );
  INV_X1 U10725 ( .A(n11999), .ZN(n8666) );
  NAND2_X1 U10726 ( .A1(n11183), .A2(n8666), .ZN(n8413) );
  OR2_X1 U10727 ( .A1(n11849), .A2(n13878), .ZN(n8412) );
  NAND2_X1 U10728 ( .A1(n8413), .A2(n8412), .ZN(n11292) );
  NAND2_X1 U10729 ( .A1(n10044), .A2(n11971), .ZN(n8417) );
  NAND2_X1 U10730 ( .A1(n8414), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8415) );
  XNOR2_X1 U10731 ( .A(n8415), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U10732 ( .A1(n11972), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6509), 
        .B2(n10317), .ZN(n8416) );
  NAND2_X1 U10733 ( .A1(n8647), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10734 ( .A1(n6470), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8422) );
  OR2_X1 U10735 ( .A1(n8418), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8419) );
  AND2_X1 U10736 ( .A1(n8419), .A2(n8434), .ZN(n11537) );
  NAND2_X1 U10737 ( .A1(n8605), .A2(n11537), .ZN(n8421) );
  NAND2_X1 U10738 ( .A1(n8570), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8420) );
  NAND4_X1 U10739 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n13877) );
  OR2_X1 U10740 ( .A1(n11854), .A2(n13827), .ZN(n8669) );
  NAND2_X1 U10741 ( .A1(n11854), .A2(n13827), .ZN(n8424) );
  NAND2_X1 U10742 ( .A1(n8669), .A2(n8424), .ZN(n11998) );
  NAND2_X1 U10743 ( .A1(n11292), .A2(n11998), .ZN(n8426) );
  OR2_X1 U10744 ( .A1(n11854), .A2(n13877), .ZN(n8425) );
  NAND2_X1 U10745 ( .A1(n10069), .A2(n11971), .ZN(n8432) );
  OR2_X1 U10746 ( .A1(n6490), .A2(n14351), .ZN(n8428) );
  NAND2_X1 U10747 ( .A1(n8429), .A2(n8428), .ZN(n8442) );
  INV_X1 U10748 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8430) );
  XNOR2_X1 U10749 ( .A(n8442), .B(n8430), .ZN(n13988) );
  AOI22_X1 U10750 ( .A1(n11972), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6509), 
        .B2(n13988), .ZN(n8431) );
  NAND2_X1 U10751 ( .A1(n6470), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10752 ( .A1(n8647), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10753 ( .A1(n8434), .A2(n8433), .ZN(n8435) );
  AND2_X1 U10754 ( .A1(n8446), .A2(n8435), .ZN(n13830) );
  NAND2_X1 U10755 ( .A1(n8605), .A2(n13830), .ZN(n8437) );
  NAND2_X1 U10756 ( .A1(n8570), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8436) );
  NAND4_X1 U10757 ( .A1(n8439), .A2(n8438), .A3(n8437), .A4(n8436), .ZN(n13876) );
  NOR2_X1 U10758 ( .A1(n11857), .A2(n13876), .ZN(n8441) );
  NAND2_X1 U10759 ( .A1(n11857), .A2(n13876), .ZN(n8440) );
  NAND2_X1 U10760 ( .A1(n10091), .A2(n11971), .ZN(n8444) );
  OAI21_X1 U10761 ( .B1(n8442), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8456) );
  XNOR2_X1 U10762 ( .A(n8456), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U10763 ( .A1(n11972), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10325), 
        .B2(n6509), .ZN(n8443) );
  NAND2_X1 U10764 ( .A1(n8647), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U10765 ( .A1(n6470), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8450) );
  AND2_X1 U10766 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  NOR2_X1 U10767 ( .A1(n8463), .A2(n8447), .ZN(n13757) );
  NAND2_X1 U10768 ( .A1(n6510), .A2(n13757), .ZN(n8449) );
  NAND2_X1 U10769 ( .A1(n8570), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8448) );
  NAND4_X1 U10770 ( .A1(n8451), .A2(n8450), .A3(n8449), .A4(n8448), .ZN(n13875) );
  OR2_X1 U10771 ( .A1(n11866), .A2(n13875), .ZN(n8454) );
  NAND2_X1 U10772 ( .A1(n11866), .A2(n13875), .ZN(n8452) );
  NAND2_X1 U10773 ( .A1(n8454), .A2(n8452), .ZN(n12002) );
  INV_X1 U10774 ( .A(n12002), .ZN(n8453) );
  NAND2_X1 U10775 ( .A1(n10223), .A2(n11971), .ZN(n8462) );
  INV_X1 U10776 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10777 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  NAND2_X1 U10778 ( .A1(n8457), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8459) );
  INV_X1 U10779 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U10780 ( .A1(n8459), .A2(n8458), .ZN(n8470) );
  OR2_X1 U10781 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  AOI22_X1 U10782 ( .A1(n10385), .A2(n6509), .B1(n11972), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8461) );
  NAND2_X1 U10783 ( .A1(n8647), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10784 ( .A1(n6470), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8467) );
  OR2_X1 U10785 ( .A1(n8463), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8464) );
  AND2_X1 U10786 ( .A1(n8475), .A2(n8464), .ZN(n13816) );
  NAND2_X1 U10787 ( .A1(n8605), .A2(n13816), .ZN(n8466) );
  NAND2_X1 U10788 ( .A1(n8570), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8465) );
  NAND4_X1 U10789 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n13874) );
  XNOR2_X1 U10790 ( .A(n14525), .B(n14510), .ZN(n12004) );
  OR2_X1 U10791 ( .A1(n14525), .A2(n13874), .ZN(n8469) );
  NAND2_X1 U10792 ( .A1(n10420), .A2(n11971), .ZN(n8473) );
  NAND2_X1 U10793 ( .A1(n8470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U10794 ( .A(n8471), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U10795 ( .A1(n10383), .A2(n6509), .B1(n11972), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U10796 ( .A1(n6470), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U10797 ( .A1(n8647), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10798 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  AND2_X1 U10799 ( .A1(n8485), .A2(n8476), .ZN(n13708) );
  NAND2_X1 U10800 ( .A1(n6510), .A2(n13708), .ZN(n8478) );
  NAND2_X1 U10801 ( .A1(n8570), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8477) );
  NAND4_X1 U10802 ( .A1(n8480), .A2(n8479), .A3(n8478), .A4(n8477), .ZN(n14499) );
  NAND2_X1 U10803 ( .A1(n14513), .A2(n14523), .ZN(n11880) );
  NAND2_X1 U10804 ( .A1(n11871), .A2(n11880), .ZN(n11870) );
  INV_X1 U10805 ( .A(n11870), .ZN(n12007) );
  AND2_X1 U10806 ( .A1(n8481), .A2(n8341), .ZN(n8495) );
  OR2_X1 U10807 ( .A1(n8495), .A2(n14351), .ZN(n8482) );
  XNOR2_X1 U10808 ( .A(n8482), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U10809 ( .A1(n11972), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6509), 
        .B2(n10969), .ZN(n8483) );
  NAND2_X1 U10810 ( .A1(n6470), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10811 ( .A1(n8647), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8489) );
  AND2_X1 U10812 ( .A1(n8485), .A2(n8484), .ZN(n8486) );
  NOR2_X1 U10813 ( .A1(n8499), .A2(n8486), .ZN(n13861) );
  NAND2_X1 U10814 ( .A1(n8605), .A2(n13861), .ZN(n8488) );
  NAND2_X1 U10815 ( .A1(n8570), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8487) );
  NAND4_X1 U10816 ( .A1(n8490), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n13873) );
  OR2_X1 U10817 ( .A1(n6670), .A2(n13873), .ZN(n8491) );
  INV_X1 U10818 ( .A(n8491), .ZN(n8492) );
  NAND2_X1 U10819 ( .A1(n14513), .A2(n14499), .ZN(n11481) );
  INV_X1 U10820 ( .A(n13873), .ZN(n14511) );
  NAND2_X1 U10821 ( .A1(n11583), .A2(n14511), .ZN(n11881) );
  NAND2_X1 U10822 ( .A1(n10400), .A2(n11971), .ZN(n8498) );
  INV_X1 U10823 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10824 ( .A1(n8495), .A2(n8494), .ZN(n8506) );
  NAND2_X1 U10825 ( .A1(n8506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8496) );
  XNOR2_X1 U10826 ( .A(n8496), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U10827 ( .A1(n11972), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6509), 
        .B2(n10973), .ZN(n8497) );
  NOR2_X1 U10828 ( .A1(n8499), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U10829 ( .A1(n7443), .A2(n8605), .ZN(n8504) );
  NAND2_X1 U10830 ( .A1(n6470), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10831 ( .A1(n8647), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U10832 ( .A1(n8570), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8501) );
  NAND4_X1 U10833 ( .A1(n8504), .A2(n8503), .A3(n8502), .A4(n8501), .ZN(n14500) );
  XNOR2_X1 U10834 ( .A(n14236), .B(n14500), .ZN(n12005) );
  OR2_X1 U10835 ( .A1(n14236), .A2(n14500), .ZN(n8505) );
  NAND2_X1 U10836 ( .A1(n10445), .A2(n11971), .ZN(n8510) );
  OAI21_X1 U10837 ( .B1(n8506), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8507) );
  MUX2_X1 U10838 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8507), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8508) );
  AND2_X1 U10839 ( .A1(n8508), .A2(n8518), .ZN(n14003) );
  AOI22_X1 U10840 ( .A1(n11972), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6509), 
        .B2(n14003), .ZN(n8509) );
  OR2_X1 U10841 ( .A1(n8511), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10842 ( .A1(n8523), .A2(n8512), .ZN(n14207) );
  INV_X1 U10843 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11224) );
  OAI22_X1 U10844 ( .A1(n14207), .A2(n8543), .B1(n8290), .B2(n11224), .ZN(
        n8516) );
  NAND2_X1 U10845 ( .A1(n8647), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U10846 ( .A1(n8570), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U10847 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  OR2_X1 U10848 ( .A1(n14213), .A2(n13872), .ZN(n8679) );
  INV_X1 U10849 ( .A(n8679), .ZN(n8517) );
  NAND2_X1 U10850 ( .A1(n14213), .A2(n13872), .ZN(n8678) );
  NAND2_X1 U10851 ( .A1(n10718), .A2(n11971), .ZN(n8521) );
  NAND2_X1 U10852 ( .A1(n8518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8519) );
  XNOR2_X1 U10853 ( .A(n8519), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14633) );
  AOI22_X1 U10854 ( .A1(n11972), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6509), 
        .B2(n14633), .ZN(n8520) );
  INV_X1 U10855 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14195) );
  NAND2_X1 U10856 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  NAND2_X1 U10857 ( .A1(n8539), .A2(n8524), .ZN(n14194) );
  OR2_X1 U10858 ( .A1(n14194), .A2(n8543), .ZN(n8528) );
  NAND2_X1 U10859 ( .A1(n8570), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10860 ( .A1(n6470), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8525) );
  AND2_X1 U10861 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  OAI211_X1 U10862 ( .C1(n8363), .C2(n14195), .A(n8528), .B(n8527), .ZN(n14485) );
  AND2_X1 U10863 ( .A1(n14182), .A2(n14485), .ZN(n8529) );
  OR2_X1 U10864 ( .A1(n14182), .A2(n14485), .ZN(n8530) );
  NAND2_X1 U10865 ( .A1(n8531), .A2(n11971), .ZN(n8537) );
  NAND2_X1 U10866 ( .A1(n8637), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8534) );
  AOI22_X1 U10867 ( .A1(n11972), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14106), 
        .B2(n6509), .ZN(n8536) );
  NAND2_X1 U10868 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  NAND2_X1 U10869 ( .A1(n8548), .A2(n8540), .ZN(n14171) );
  AOI22_X1 U10870 ( .A1(n6470), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8647), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U10871 ( .A1(n8570), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8541) );
  OAI211_X1 U10872 ( .C1(n14171), .C2(n8543), .A(n8542), .B(n8541), .ZN(n14199) );
  INV_X1 U10873 ( .A(n14199), .ZN(n14155) );
  OR2_X1 U10874 ( .A1(n8544), .A2(n14155), .ZN(n11908) );
  NAND2_X1 U10875 ( .A1(n8544), .A2(n14155), .ZN(n11909) );
  NAND2_X1 U10876 ( .A1(n11908), .A2(n11909), .ZN(n14168) );
  NOR2_X1 U10877 ( .A1(n8544), .A2(n14199), .ZN(n8545) );
  NAND2_X1 U10878 ( .A1(n11010), .A2(n11971), .ZN(n8547) );
  NAND2_X1 U10879 ( .A1(n11972), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8546) );
  AND2_X1 U10880 ( .A1(n8548), .A2(n13808), .ZN(n8549) );
  NOR2_X1 U10881 ( .A1(n8558), .A2(n8549), .ZN(n14151) );
  NAND2_X1 U10882 ( .A1(n14151), .A2(n8605), .ZN(n8554) );
  INV_X1 U10883 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U10884 ( .A1(n8647), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10885 ( .A1(n8570), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8550) );
  OAI211_X1 U10886 ( .C1(n14314), .C2(n8574), .A(n8551), .B(n8550), .ZN(n8552)
         );
  INV_X1 U10887 ( .A(n8552), .ZN(n8553) );
  INV_X1 U10888 ( .A(n14317), .ZN(n11917) );
  XNOR2_X1 U10889 ( .A(n14160), .B(n11917), .ZN(n14161) );
  NAND2_X1 U10890 ( .A1(n14160), .A2(n14317), .ZN(n8555) );
  NAND2_X1 U10891 ( .A1(n11234), .A2(n11971), .ZN(n8557) );
  NAND2_X1 U10892 ( .A1(n11972), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8556) );
  NOR2_X1 U10893 ( .A1(n8558), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8559) );
  OR2_X1 U10894 ( .A1(n8568), .A2(n8559), .ZN(n14139) );
  INV_X1 U10895 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U10896 ( .A1(n8570), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10897 ( .A1(n8647), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8560) );
  OAI211_X1 U10898 ( .C1(n8574), .C2(n8562), .A(n8561), .B(n8560), .ZN(n8563)
         );
  INV_X1 U10899 ( .A(n8563), .ZN(n8564) );
  XNOR2_X1 U10900 ( .A(n14301), .B(n14152), .ZN(n14144) );
  OR2_X1 U10901 ( .A1(n14301), .A2(n14152), .ZN(n8565) );
  OR2_X1 U10902 ( .A1(n8566), .A2(n6492), .ZN(n8567) );
  XNOR2_X1 U10903 ( .A(n8567), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14368) );
  OR2_X1 U10904 ( .A1(n8568), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10905 ( .A1(n8569), .A2(n8581), .ZN(n14125) );
  INV_X1 U10906 ( .A(n14125), .ZN(n11652) );
  NAND2_X1 U10907 ( .A1(n11652), .A2(n6510), .ZN(n8577) );
  INV_X1 U10908 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U10909 ( .A1(n8570), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U10910 ( .A1(n8647), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8571) );
  OAI211_X1 U10911 ( .C1(n8574), .C2(n8573), .A(n8572), .B(n8571), .ZN(n8575)
         );
  INV_X1 U10912 ( .A(n8575), .ZN(n8576) );
  XNOR2_X1 U10913 ( .A(n14295), .B(n11637), .ZN(n12011) );
  NAND2_X1 U10914 ( .A1(n14121), .A2(n14120), .ZN(n14119) );
  NAND2_X1 U10915 ( .A1(n11318), .A2(n11971), .ZN(n8579) );
  NAND2_X1 U10916 ( .A1(n11972), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U10917 ( .A1(n6470), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U10918 ( .A1(n8647), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8584) );
  INV_X1 U10919 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13719) );
  AOI21_X1 U10920 ( .B1(n13719), .B2(n8581), .A(n8580), .ZN(n14108) );
  NAND2_X1 U10921 ( .A1(n8605), .A2(n14108), .ZN(n8583) );
  NAND2_X1 U10922 ( .A1(n8570), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8582) );
  NAND4_X1 U10923 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n14079) );
  NAND2_X1 U10924 ( .A1(n14289), .A2(n14079), .ZN(n8588) );
  OR2_X1 U10925 ( .A1(n14289), .A2(n14079), .ZN(n8586) );
  NAND2_X1 U10926 ( .A1(n8588), .A2(n8586), .ZN(n14099) );
  AND2_X1 U10927 ( .A1(n14295), .A2(n11637), .ZN(n14097) );
  NOR2_X1 U10928 ( .A1(n14099), .A2(n14097), .ZN(n8587) );
  NAND2_X1 U10929 ( .A1(n14119), .A2(n8587), .ZN(n14102) );
  NAND2_X1 U10930 ( .A1(n11439), .A2(n11971), .ZN(n8590) );
  NAND2_X1 U10931 ( .A1(n11972), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U10932 ( .A1(n8647), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10933 ( .A1(n6470), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8596) );
  INV_X1 U10934 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8593) );
  AOI21_X1 U10935 ( .B1(n8593), .B2(n8592), .A(n8591), .ZN(n14088) );
  NAND2_X1 U10936 ( .A1(n8605), .A2(n14088), .ZN(n8595) );
  NAND2_X1 U10937 ( .A1(n8570), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8594) );
  NAND4_X1 U10938 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n14112) );
  INV_X1 U10939 ( .A(n14112), .ZN(n8598) );
  OR2_X1 U10940 ( .A1(n14087), .A2(n8598), .ZN(n8688) );
  NAND2_X1 U10941 ( .A1(n14087), .A2(n8598), .ZN(n8599) );
  NAND2_X1 U10942 ( .A1(n8688), .A2(n8599), .ZN(n12013) );
  OR2_X1 U10943 ( .A1(n14087), .A2(n14112), .ZN(n8600) );
  NAND2_X1 U10944 ( .A1(n11475), .A2(n11971), .ZN(n8602) );
  NAND2_X1 U10945 ( .A1(n11972), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U10946 ( .A1(n6470), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U10947 ( .A1(n8647), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8608) );
  INV_X1 U10948 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13768) );
  AOI21_X1 U10949 ( .B1(n13768), .B2(n8604), .A(n8603), .ZN(n14069) );
  NAND2_X1 U10950 ( .A1(n8605), .A2(n14069), .ZN(n8607) );
  NAND2_X1 U10951 ( .A1(n8570), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8606) );
  NAND4_X1 U10952 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n14078) );
  INV_X1 U10953 ( .A(n14078), .ZN(n13797) );
  NAND2_X1 U10954 ( .A1(n14058), .A2(n13797), .ZN(n14042) );
  OR2_X1 U10955 ( .A1(n14058), .A2(n13797), .ZN(n8610) );
  NAND2_X1 U10956 ( .A1(n14042), .A2(n8610), .ZN(n14060) );
  INV_X1 U10957 ( .A(n14060), .ZN(n14065) );
  NAND2_X1 U10958 ( .A1(n14058), .A2(n14078), .ZN(n8611) );
  NAND2_X1 U10959 ( .A1(n13687), .A2(n11971), .ZN(n8613) );
  NAND2_X1 U10960 ( .A1(n11972), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U10961 ( .A1(n8647), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U10962 ( .A1(n8570), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8618) );
  INV_X1 U10963 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13846) );
  AOI21_X1 U10964 ( .B1(n13846), .B2(n8615), .A(n8614), .ZN(n14050) );
  NAND2_X1 U10965 ( .A1(n6510), .A2(n14050), .ZN(n8617) );
  NAND2_X1 U10966 ( .A1(n6470), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10967 ( .A1(n14041), .A2(n14040), .ZN(n8621) );
  NAND2_X1 U10968 ( .A1(n14046), .A2(n13871), .ZN(n8620) );
  NAND2_X1 U10969 ( .A1(n8621), .A2(n8620), .ZN(n9369) );
  NAND2_X1 U10970 ( .A1(n11655), .A2(n11971), .ZN(n8623) );
  NAND2_X1 U10971 ( .A1(n11972), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U10972 ( .A1(n6470), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U10973 ( .A1(n8647), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8627) );
  XNOR2_X1 U10974 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n8624), .ZN(n14032) );
  NAND2_X1 U10975 ( .A1(n8605), .A2(n14032), .ZN(n8626) );
  NAND2_X1 U10976 ( .A1(n8570), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8625) );
  NAND4_X1 U10977 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n13870) );
  XNOR2_X1 U10978 ( .A(n14033), .B(n13870), .ZN(n12014) );
  XNOR2_X1 U10979 ( .A(n12382), .B(n13869), .ZN(n12016) );
  NAND2_X1 U10980 ( .A1(n13678), .A2(n11971), .ZN(n8631) );
  NAND2_X1 U10981 ( .A1(n11972), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U10982 ( .A1(n6470), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10983 ( .A1(n8647), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8635) );
  INV_X1 U10984 ( .A(n8632), .ZN(n12309) );
  NAND2_X1 U10985 ( .A1(n6510), .A2(n12309), .ZN(n8634) );
  NAND2_X1 U10986 ( .A1(n8570), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8633) );
  NAND4_X1 U10987 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .ZN(n13868) );
  INV_X1 U10988 ( .A(n13868), .ZN(n9355) );
  XNOR2_X1 U10989 ( .A(n12308), .B(n9355), .ZN(n12018) );
  MUX2_X1 U10990 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8639), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8640) );
  NAND2_X1 U10991 ( .A1(n8641), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8642) );
  INV_X1 U10992 ( .A(n11976), .ZN(n10283) );
  NAND2_X1 U10993 ( .A1(n6852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U10994 ( .A1(n11120), .A2(n6857), .ZN(n8717) );
  AND2_X1 U10995 ( .A1(n11794), .A2(n8717), .ZN(n8645) );
  NAND2_X1 U10996 ( .A1(n6470), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U10997 ( .A1(n8647), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U10998 ( .A1(n8570), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8648) );
  NAND3_X1 U10999 ( .A1(n8650), .A2(n8649), .A3(n8648), .ZN(n13867) );
  INV_X1 U11000 ( .A(P1_B_REG_SCAN_IN), .ZN(n8700) );
  NOR2_X1 U11001 ( .A1(n14362), .A2(n8700), .ZN(n8652) );
  NOR2_X1 U11002 ( .A1(n14522), .A2(n8652), .ZN(n14021) );
  AND2_X1 U11003 ( .A1(n13867), .A2(n14021), .ZN(n12310) );
  NAND2_X1 U11004 ( .A1(n14242), .A2(n10653), .ZN(n10553) );
  OR2_X1 U11005 ( .A1(n10553), .A2(n10714), .ZN(n10745) );
  NOR2_X2 U11006 ( .A1(n10745), .A2(n14652), .ZN(n10744) );
  INV_X1 U11007 ( .A(n11829), .ZN(n10891) );
  INV_X1 U11008 ( .A(n11836), .ZN(n14660) );
  NAND2_X1 U11009 ( .A1(n10825), .A2(n14660), .ZN(n10837) );
  OR2_X1 U11010 ( .A1(n10837), .A2(n11839), .ZN(n11145) );
  INV_X1 U11011 ( .A(n11854), .ZN(n14681) );
  OR2_X2 U11012 ( .A1(n11391), .A2(n14525), .ZN(n11508) );
  NOR2_X2 U11013 ( .A1(n11508), .A2(n14513), .ZN(n11487) );
  NOR2_X1 U11014 ( .A1(n14220), .A2(n14236), .ZN(n14221) );
  NAND2_X1 U11015 ( .A1(n14221), .A2(n14488), .ZN(n14205) );
  NAND2_X1 U11016 ( .A1(n14122), .A2(n14115), .ZN(n14095) );
  NOR2_X2 U11017 ( .A1(n12308), .A2(n9351), .ZN(n14027) );
  AOI211_X1 U11018 ( .C1(n12308), .C2(n9351), .A(n14644), .B(n14027), .ZN(
        n12317) );
  INV_X1 U11019 ( .A(n10303), .ZN(n14249) );
  NAND2_X1 U11020 ( .A1(n11802), .A2(n11796), .ZN(n8654) );
  NAND2_X1 U11021 ( .A1(n8654), .A2(n11800), .ZN(n10518) );
  NAND2_X1 U11022 ( .A1(n11808), .A2(n11809), .ZN(n8655) );
  NAND2_X1 U11023 ( .A1(n8656), .A2(n11818), .ZN(n10746) );
  NAND2_X1 U11024 ( .A1(n10746), .A2(n11991), .ZN(n8657) );
  NAND2_X1 U11025 ( .A1(n10572), .A2(n14652), .ZN(n11816) );
  NAND2_X1 U11026 ( .A1(n8657), .A2(n11816), .ZN(n10700) );
  NAND2_X1 U11027 ( .A1(n10700), .A2(n11992), .ZN(n8660) );
  INV_X1 U11028 ( .A(n13883), .ZN(n8658) );
  NAND2_X1 U11029 ( .A1(n8658), .A2(n11829), .ZN(n8659) );
  INV_X1 U11030 ( .A(n13882), .ZN(n8661) );
  AND2_X1 U11031 ( .A1(n11836), .A2(n8661), .ZN(n8662) );
  INV_X1 U11032 ( .A(n10830), .ZN(n8663) );
  NAND2_X1 U11033 ( .A1(n8663), .A2(n7442), .ZN(n8665) );
  NAND2_X1 U11034 ( .A1(n11839), .A2(n11142), .ZN(n8664) );
  INV_X1 U11035 ( .A(n13878), .ZN(n11535) );
  INV_X1 U11036 ( .A(n13876), .ZN(n11372) );
  NAND2_X1 U11037 ( .A1(n11857), .A2(n11372), .ZN(n8670) );
  OR2_X1 U11038 ( .A1(n11857), .A2(n11372), .ZN(n8671) );
  INV_X1 U11039 ( .A(n13875), .ZN(n14521) );
  OR2_X1 U11040 ( .A1(n11866), .A2(n14521), .ZN(n8672) );
  INV_X1 U11041 ( .A(n12004), .ZN(n8674) );
  NAND2_X1 U11042 ( .A1(n11384), .A2(n8674), .ZN(n8676) );
  OR2_X1 U11043 ( .A1(n14525), .A2(n14510), .ZN(n8675) );
  INV_X1 U11044 ( .A(n11491), .ZN(n8677) );
  INV_X1 U11045 ( .A(n13872), .ZN(n14233) );
  INV_X1 U11046 ( .A(n14485), .ZN(n14175) );
  XNOR2_X1 U11047 ( .A(n14182), .B(n14175), .ZN(n14186) );
  INV_X1 U11048 ( .A(n14186), .ZN(n14189) );
  OR2_X1 U11049 ( .A1(n14182), .A2(n14175), .ZN(n8680) );
  INV_X1 U11050 ( .A(n14161), .ZN(n14149) );
  OR2_X1 U11051 ( .A1(n14160), .A2(n11917), .ZN(n8682) );
  INV_X1 U11052 ( .A(n14152), .ZN(n8683) );
  OR2_X1 U11053 ( .A1(n14301), .A2(n8683), .ZN(n8684) );
  OR2_X1 U11054 ( .A1(n14295), .A2(n14134), .ZN(n8685) );
  INV_X1 U11055 ( .A(n14079), .ZN(n8686) );
  AND2_X1 U11056 ( .A1(n14289), .A2(n8686), .ZN(n8687) );
  NAND2_X1 U11057 ( .A1(n14080), .A2(n8688), .ZN(n14061) );
  OR2_X1 U11058 ( .A1(n14060), .A2(n14040), .ZN(n8689) );
  INV_X1 U11059 ( .A(n13871), .ZN(n8690) );
  INV_X1 U11060 ( .A(n13870), .ZN(n9356) );
  NAND2_X1 U11061 ( .A1(n9353), .A2(n7448), .ZN(n8692) );
  INV_X1 U11062 ( .A(n13869), .ZN(n13696) );
  NAND2_X1 U11063 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  XNOR2_X1 U11064 ( .A(n8693), .B(n12018), .ZN(n8696) );
  OR2_X1 U11065 ( .A1(n11791), .A2(n6857), .ZN(n8694) );
  INV_X1 U11066 ( .A(n11120), .ZN(n11795) );
  NAND2_X1 U11067 ( .A1(n11960), .A2(n11795), .ZN(n11963) );
  NAND2_X1 U11068 ( .A1(n8715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8697) );
  MUX2_X1 U11069 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8697), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8699) );
  NAND2_X1 U11070 ( .A1(n8712), .A2(n8700), .ZN(n8710) );
  NAND2_X1 U11071 ( .A1(n8698), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8701) );
  MUX2_X1 U11072 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8701), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8703) );
  INV_X1 U11073 ( .A(n8702), .ZN(n8704) );
  NAND2_X1 U11074 ( .A1(n8703), .A2(n8704), .ZN(n11477) );
  AND2_X1 U11075 ( .A1(n11477), .A2(P1_B_REG_SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11076 ( .A1(n8704), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8705) );
  MUX2_X1 U11077 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8705), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8707) );
  AOI21_X1 U11078 ( .B1(n11542), .B2(n8708), .A(n14367), .ZN(n8709) );
  INV_X1 U11079 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10050) );
  AND2_X1 U11080 ( .A1(n11542), .A2(n14367), .ZN(n10049) );
  NOR2_X1 U11081 ( .A1(n14367), .A2(n11477), .ZN(n8711) );
  NAND2_X1 U11082 ( .A1(n8713), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8714) );
  MUX2_X1 U11083 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8714), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8716) );
  NAND2_X1 U11084 ( .A1(n8716), .A2(n8715), .ZN(n10060) );
  NAND2_X1 U11085 ( .A1(n11976), .A2(n8717), .ZN(n10287) );
  NAND2_X1 U11086 ( .A1(n10295), .A2(n10287), .ZN(n12031) );
  NOR2_X1 U11087 ( .A1(n10644), .A2(n12031), .ZN(n8733) );
  NOR4_X1 U11088 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8721) );
  NOR4_X1 U11089 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8720) );
  NOR4_X1 U11090 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8719) );
  NOR4_X1 U11091 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8718) );
  NAND4_X1 U11092 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(n8727)
         );
  NOR2_X1 U11093 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n8725) );
  NOR4_X1 U11094 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n8724) );
  NOR4_X1 U11095 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8723) );
  NOR4_X1 U11096 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8722) );
  NAND4_X1 U11097 ( .A1(n8725), .A2(n8724), .A3(n8723), .A4(n8722), .ZN(n8726)
         );
  NOR2_X1 U11098 ( .A1(n8727), .A2(n8726), .ZN(n10278) );
  INV_X1 U11099 ( .A(n10278), .ZN(n8728) );
  INV_X1 U11100 ( .A(n10286), .ZN(n10294) );
  AOI21_X1 U11101 ( .B1(n10281), .B2(n8728), .A(n10294), .ZN(n8732) );
  INV_X1 U11102 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U11103 ( .A1(n10281), .A2(n10051), .ZN(n8730) );
  INV_X1 U11104 ( .A(n10279), .ZN(n8729) );
  NAND2_X1 U11105 ( .A1(n8730), .A2(n8729), .ZN(n8731) );
  AND2_X1 U11106 ( .A1(n8732), .A2(n8731), .ZN(n9363) );
  INV_X1 U11107 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8734) );
  OR2_X1 U11108 ( .A1(n14687), .A2(n8734), .ZN(n8735) );
  INV_X1 U11109 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8737) );
  INV_X1 U11110 ( .A(n8876), .ZN(n8738) );
  NAND2_X1 U11111 ( .A1(n8857), .A2(n8738), .ZN(n8741) );
  NAND2_X1 U11112 ( .A1(n8739), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11113 ( .A1(n8741), .A2(n8740), .ZN(n8889) );
  NAND2_X1 U11114 ( .A1(n9942), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11115 ( .A1(n9969), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8742) );
  AND2_X1 U11116 ( .A1(n8743), .A2(n8742), .ZN(n8888) );
  NAND2_X1 U11117 ( .A1(n8889), .A2(n8888), .ZN(n8887) );
  NAND2_X1 U11118 ( .A1(n8887), .A2(n8743), .ZN(n8903) );
  NAND2_X1 U11119 ( .A1(n9944), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11120 ( .A1(n9999), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8744) );
  AND2_X1 U11121 ( .A1(n8745), .A2(n8744), .ZN(n8902) );
  NAND2_X1 U11122 ( .A1(n8903), .A2(n8902), .ZN(n8905) );
  NAND2_X1 U11123 ( .A1(n9946), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8747) );
  INV_X1 U11124 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U11125 ( .A1(n9996), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U11126 ( .A1(n9966), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8749) );
  INV_X1 U11127 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U11128 ( .A1(n9994), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11129 ( .A1(n8750), .A2(n8749), .ZN(n8954) );
  NAND2_X1 U11130 ( .A1(n9973), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U11131 ( .A1(n8954), .A2(n8751), .ZN(n8753) );
  NAND2_X1 U11132 ( .A1(n9972), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U11133 ( .A1(n8753), .A2(n8752), .ZN(n8981) );
  NAND2_X1 U11134 ( .A1(n9991), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11135 ( .A1(n9990), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11136 ( .A1(n8755), .A2(n8754), .ZN(n8980) );
  NAND2_X1 U11137 ( .A1(n10003), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11138 ( .A1(n10006), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11139 ( .A1(n10040), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U11140 ( .A1(n10039), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11141 ( .A1(n10045), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11142 ( .A1(n10047), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U11143 ( .A1(n8762), .A2(n8760), .ZN(n9026) );
  INV_X1 U11144 ( .A(n9026), .ZN(n8761) );
  NAND2_X1 U11145 ( .A1(n10072), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U11146 ( .A1(n10070), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U11147 ( .A1(n8765), .A2(n8763), .ZN(n9052) );
  INV_X1 U11148 ( .A(n9052), .ZN(n8764) );
  NAND2_X1 U11149 ( .A1(n10092), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11150 ( .A1(n10097), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11151 ( .A1(n10447), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U11152 ( .A1(n10421), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U11153 ( .A1(n10453), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11154 ( .A1(n10452), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U11155 ( .A1(n10422), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U11156 ( .A1(n10401), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U11157 ( .A1(n10449), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11158 ( .A1(n10446), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8775) );
  INV_X1 U11159 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U11160 ( .A1(n10719), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8778) );
  INV_X1 U11161 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U11162 ( .A1(n10722), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11163 ( .A1(n10787), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U11164 ( .A1(n10789), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8779) );
  INV_X1 U11165 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U11166 ( .A1(n11237), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8785) );
  INV_X1 U11167 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11236) );
  NAND2_X1 U11168 ( .A1(n11236), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8784) );
  AND2_X1 U11169 ( .A1(n8785), .A2(n8784), .ZN(n9208) );
  INV_X1 U11170 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11253) );
  XNOR2_X1 U11171 ( .A(n11253), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11172 ( .A1(n11253), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8786) );
  XNOR2_X1 U11173 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9239) );
  INV_X1 U11174 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8787) );
  INV_X1 U11175 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U11176 ( .A1(n8788), .A2(n11441), .ZN(n8789) );
  NAND2_X1 U11177 ( .A1(n11480), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U11178 ( .A1(n11476), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8791) );
  AND2_X1 U11179 ( .A1(n14364), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U11180 ( .A1(n13689), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8794) );
  XNOR2_X1 U11181 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8795) );
  XNOR2_X1 U11182 ( .A(n9711), .B(n8795), .ZN(n12073) );
  INV_X1 U11183 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8805) );
  XNOR2_X2 U11184 ( .A(n8806), .B(n8834), .ZN(n9336) );
  XNOR2_X2 U11185 ( .A(n8809), .B(n8805), .ZN(n9885) );
  NAND2_X1 U11186 ( .A1(n12073), .A2(n12098), .ZN(n8811) );
  NAND2_X2 U11187 ( .A1(n6508), .A2(n9961), .ZN(n8984) );
  INV_X1 U11188 ( .A(SI_27_), .ZN(n12074) );
  NAND2_X1 U11189 ( .A1(n6534), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8812) );
  INV_X1 U11190 ( .A(n8813), .ZN(n8815) );
  AND2_X2 U11191 ( .A1(n8814), .A2(n8815), .ZN(n11135) );
  INV_X1 U11192 ( .A(P3_B_REG_SCAN_IN), .ZN(n9736) );
  XNOR2_X1 U11193 ( .A(n11135), .B(n9736), .ZN(n8817) );
  NAND2_X1 U11194 ( .A1(n8815), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8816) );
  INV_X1 U11195 ( .A(n9305), .ZN(n11282) );
  NAND2_X1 U11196 ( .A1(n8818), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8819) );
  INV_X1 U11197 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U11198 ( .A1(n10165), .A2(n8820), .ZN(n8822) );
  OR2_X1 U11199 ( .A1(n11135), .A2(n11346), .ZN(n8821) );
  INV_X1 U11200 ( .A(n8823), .ZN(n8824) );
  NAND2_X1 U11201 ( .A1(n8824), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U11202 ( .A1(n8827), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U11203 ( .A1(n12139), .A2(n9746), .ZN(n12132) );
  OR2_X2 U11204 ( .A1(n9318), .A2(n12132), .ZN(n8833) );
  NAND2_X1 U11205 ( .A1(n9132), .A2(n8829), .ZN(n9149) );
  NOR2_X1 U11206 ( .A1(n12139), .A2(n9746), .ZN(n8831) );
  XNOR2_X1 U11207 ( .A(n12855), .B(n8926), .ZN(n8851) );
  INV_X1 U11208 ( .A(n8836), .ZN(n8835) );
  NAND2_X1 U11209 ( .A1(n8835), .A2(n8837), .ZN(n13002) );
  NAND2_X1 U11210 ( .A1(n12083), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8850) );
  INV_X1 U11211 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12656) );
  OR2_X1 U11212 ( .A1(n12086), .A2(n12656), .ZN(n8849) );
  INV_X1 U11213 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12500) );
  NOR2_X1 U11214 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8941) );
  NAND2_X1 U11215 ( .A1(n8941), .A2(n9564), .ZN(n8960) );
  NOR2_X1 U11216 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_REG3_REG_9__SCAN_IN), 
        .ZN(n8842) );
  NAND2_X1 U11217 ( .A1(n9100), .A2(n15087), .ZN(n9120) );
  INV_X1 U11218 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9169) );
  INV_X1 U11219 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U11220 ( .A1(n12500), .A2(n9251), .ZN(n9267) );
  INV_X1 U11221 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11222 ( .A1(n9581), .A2(n9281), .ZN(n9338) );
  INV_X1 U11223 ( .A(n9281), .ZN(n8844) );
  NAND2_X1 U11224 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8844), .ZN(n8845) );
  OR2_X1 U11225 ( .A1(n9723), .A2(n12655), .ZN(n8848) );
  INV_X1 U11226 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12856) );
  OR2_X1 U11227 ( .A1(n12085), .A2(n12856), .ZN(n8847) );
  INV_X1 U11228 ( .A(n12427), .ZN(n12583) );
  NOR2_X1 U11229 ( .A1(n8851), .A2(n12583), .ZN(n12435) );
  AOI21_X1 U11230 ( .B1(n8851), .B2(n12583), .A(n12435), .ZN(n9291) );
  NAND2_X1 U11231 ( .A1(n6504), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8856) );
  INV_X1 U11232 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8852) );
  OR2_X1 U11233 ( .A1(n8913), .A2(n8852), .ZN(n8855) );
  INV_X1 U11234 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15120) );
  OR2_X1 U11235 ( .A1(n8891), .A2(n15120), .ZN(n8854) );
  INV_X1 U11236 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11107) );
  NAND4_X2 U11237 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8853), .ZN(n8879)
         );
  INV_X1 U11238 ( .A(n8879), .ZN(n8862) );
  OR2_X1 U11239 ( .A1(n8984), .A2(n9948), .ZN(n8861) );
  XNOR2_X1 U11240 ( .A(n8857), .B(n8876), .ZN(n9947) );
  NAND2_X1 U11241 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8859) );
  INV_X1 U11242 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8858) );
  XNOR2_X2 U11243 ( .A(n8859), .B(n8858), .ZN(n9830) );
  OR2_X1 U11244 ( .A1(n6502), .A2(n9830), .ZN(n8860) );
  OAI21_X1 U11245 ( .B1(n8879), .B2(n10776), .A(n9754), .ZN(n8863) );
  OR2_X1 U11246 ( .A1(n6535), .A2(n10776), .ZN(n8864) );
  NAND2_X1 U11247 ( .A1(n8863), .A2(n8864), .ZN(n8883) );
  INV_X1 U11248 ( .A(n8864), .ZN(n8865) );
  NAND2_X1 U11249 ( .A1(n8865), .A2(n8879), .ZN(n8866) );
  INV_X1 U11250 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8867) );
  OR2_X1 U11251 ( .A1(n8892), .A2(n8867), .ZN(n8870) );
  INV_X1 U11252 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9828) );
  OR2_X1 U11253 ( .A1(n8913), .A2(n9828), .ZN(n8869) );
  INV_X1 U11254 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n14993) );
  OR2_X1 U11255 ( .A1(n8891), .A2(n14993), .ZN(n8868) );
  NAND3_X1 U11256 ( .A1(n8870), .A2(n8869), .A3(n8868), .ZN(n8871) );
  AND2_X1 U11257 ( .A1(n8873), .A2(n7444), .ZN(n8878) );
  NAND2_X1 U11258 ( .A1(n8874), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8875) );
  AND2_X1 U11259 ( .A1(n8876), .A2(n8875), .ZN(n9959) );
  NAND2_X1 U11260 ( .A1(n8879), .A2(n6535), .ZN(n12140) );
  NAND2_X1 U11261 ( .A1(n9755), .A2(n10776), .ZN(n8881) );
  NAND2_X1 U11262 ( .A1(n10780), .A2(n8882), .ZN(n10779) );
  NAND2_X1 U11263 ( .A1(n10779), .A2(n8883), .ZN(n10812) );
  OR2_X1 U11264 ( .A1(n8984), .A2(SI_2_), .ZN(n8890) );
  OAI21_X1 U11265 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(n9982) );
  XNOR2_X1 U11266 ( .A(n15106), .B(n8926), .ZN(n8897) );
  NAND2_X1 U11267 ( .A1(n6503), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8896) );
  INV_X1 U11268 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15107) );
  OR2_X1 U11269 ( .A1(n8891), .A2(n15107), .ZN(n8895) );
  INV_X1 U11270 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9863) );
  XNOR2_X1 U11271 ( .A(n8897), .B(n9672), .ZN(n10811) );
  NAND2_X1 U11272 ( .A1(n10812), .A2(n10811), .ZN(n8900) );
  INV_X1 U11273 ( .A(n8897), .ZN(n8898) );
  OR2_X1 U11274 ( .A1(n9672), .A2(n8898), .ZN(n8899) );
  INV_X1 U11275 ( .A(n12409), .ZN(n8928) );
  NAND2_X1 U11276 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6572), .ZN(n8901) );
  OR2_X1 U11277 ( .A1(n8984), .A2(SI_3_), .ZN(n8907) );
  OR2_X1 U11278 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  NAND2_X1 U11279 ( .A1(n8905), .A2(n8904), .ZN(n9984) );
  OR2_X1 U11280 ( .A1(n12082), .A2(n9984), .ZN(n8906) );
  OAI211_X1 U11281 ( .C1(n11132), .C2(n6508), .A(n8907), .B(n8906), .ZN(n15140) );
  XNOR2_X1 U11282 ( .A(n15140), .B(n10776), .ZN(n8930) );
  NAND2_X1 U11283 ( .A1(n6504), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8911) );
  INV_X1 U11284 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10957) );
  OR2_X1 U11285 ( .A1(n8913), .A2(n10957), .ZN(n8909) );
  INV_X1 U11286 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9889) );
  OR2_X1 U11287 ( .A1(n12085), .A2(n9889), .ZN(n8908) );
  XNOR2_X1 U11288 ( .A(n8930), .B(n12606), .ZN(n12408) );
  NAND2_X1 U11289 ( .A1(n6504), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8919) );
  INV_X1 U11290 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n8912) );
  OR2_X1 U11291 ( .A1(n8913), .A2(n8912), .ZN(n8918) );
  AND2_X1 U11292 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8914) );
  NOR2_X1 U11293 ( .A1(n8941), .A2(n8914), .ZN(n11168) );
  INV_X1 U11294 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n8915) );
  OR2_X1 U11295 ( .A1(n12085), .A2(n8915), .ZN(n8916) );
  XNOR2_X1 U11296 ( .A(n8923), .B(n8922), .ZN(n9975) );
  OR2_X1 U11297 ( .A1(n12082), .A2(n9975), .ZN(n8925) );
  OR2_X1 U11298 ( .A1(n8984), .A2(SI_4_), .ZN(n8924) );
  OAI211_X1 U11299 ( .C1(n11084), .C2(n6508), .A(n8925), .B(n8924), .ZN(n15147) );
  XNOR2_X1 U11300 ( .A(n6467), .B(n15147), .ZN(n8929) );
  INV_X1 U11301 ( .A(n8929), .ZN(n8927) );
  NOR2_X1 U11302 ( .A1(n12605), .A2(n8927), .ZN(n8931) );
  XNOR2_X1 U11303 ( .A(n8929), .B(n12605), .ZN(n11154) );
  NAND2_X1 U11304 ( .A1(n8930), .A2(n12606), .ZN(n11150) );
  INV_X1 U11305 ( .A(n8932), .ZN(n8936) );
  NAND2_X1 U11306 ( .A1(n8933), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8934) );
  MUX2_X1 U11307 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8934), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8935) );
  NAND2_X1 U11308 ( .A1(n8936), .A2(n8935), .ZN(n9895) );
  INV_X1 U11309 ( .A(n9895), .ZN(n11057) );
  XNOR2_X1 U11310 ( .A(n8938), .B(n8937), .ZN(n9980) );
  OR2_X1 U11311 ( .A1(n12082), .A2(n9980), .ZN(n8940) );
  OR2_X1 U11312 ( .A1(n9714), .A2(SI_5_), .ZN(n8939) );
  OAI211_X1 U11313 ( .C1(n11057), .C2(n6507), .A(n8940), .B(n8939), .ZN(n15154) );
  XNOR2_X1 U11314 ( .A(n15154), .B(n8926), .ZN(n8949) );
  NAND2_X1 U11315 ( .A1(n6504), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8947) );
  INV_X2 U11316 ( .A(n9732), .ZN(n12086) );
  INV_X1 U11317 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11259) );
  OR2_X1 U11318 ( .A1(n12086), .A2(n11259), .ZN(n8946) );
  OR2_X1 U11319 ( .A1(n9564), .A2(n8941), .ZN(n8942) );
  AND2_X1 U11320 ( .A1(n8960), .A2(n8942), .ZN(n11260) );
  OR2_X1 U11321 ( .A1(n9723), .A2(n11260), .ZN(n8945) );
  INV_X1 U11322 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8943) );
  OR2_X1 U11323 ( .A1(n12085), .A2(n8943), .ZN(n8944) );
  XNOR2_X1 U11324 ( .A(n8949), .B(n12604), .ZN(n11062) );
  NAND2_X1 U11325 ( .A1(n11061), .A2(n8948), .ZN(n8952) );
  INV_X1 U11326 ( .A(n8949), .ZN(n8950) );
  OR2_X1 U11327 ( .A1(n12604), .A2(n8950), .ZN(n8951) );
  INV_X1 U11328 ( .A(SI_6_), .ZN(n9953) );
  OR2_X1 U11329 ( .A1(n8984), .A2(n9953), .ZN(n8958) );
  XNOR2_X1 U11330 ( .A(n9972), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8953) );
  XNOR2_X1 U11331 ( .A(n8954), .B(n8953), .ZN(n9954) );
  OR2_X1 U11332 ( .A1(n12082), .A2(n9954), .ZN(n8957) );
  OR2_X1 U11333 ( .A1(n8932), .A2(n8807), .ZN(n8955) );
  OR2_X1 U11334 ( .A1(n9855), .A2(n9955), .ZN(n8956) );
  XNOR2_X1 U11335 ( .A(n15158), .B(n10776), .ZN(n8967) );
  NAND2_X1 U11336 ( .A1(n6504), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8966) );
  INV_X1 U11337 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8959) );
  OR2_X1 U11338 ( .A1(n12086), .A2(n8959), .ZN(n8965) );
  NAND2_X1 U11339 ( .A1(n8960), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8961) );
  AND2_X1 U11340 ( .A1(n8969), .A2(n8961), .ZN(n11313) );
  OR2_X1 U11341 ( .A1(n9723), .A2(n11313), .ZN(n8964) );
  INV_X1 U11342 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n8962) );
  OR2_X1 U11343 ( .A1(n12085), .A2(n8962), .ZN(n8963) );
  NAND4_X1 U11344 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .ZN(n12603) );
  XNOR2_X1 U11345 ( .A(n8967), .B(n12603), .ZN(n11172) );
  NAND2_X1 U11346 ( .A1(n8967), .A2(n12603), .ZN(n8968) );
  NAND2_X1 U11347 ( .A1(n6504), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8976) );
  AND2_X1 U11348 ( .A1(n8969), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8970) );
  NOR2_X1 U11349 ( .A1(n9017), .A2(n8970), .ZN(n14971) );
  OR2_X1 U11350 ( .A1(n9723), .A2(n14971), .ZN(n8975) );
  INV_X1 U11351 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8971) );
  OR2_X1 U11352 ( .A1(n12086), .A2(n8971), .ZN(n8974) );
  INV_X1 U11353 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8972) );
  OR2_X1 U11354 ( .A1(n12085), .A2(n8972), .ZN(n8973) );
  NAND4_X1 U11355 ( .A1(n8976), .A2(n8975), .A3(n8974), .A4(n8973), .ZN(n12602) );
  INV_X1 U11356 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11357 ( .A1(n8932), .A2(n8977), .ZN(n8991) );
  NAND2_X1 U11358 ( .A1(n8991), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8979) );
  XNOR2_X1 U11359 ( .A(n8979), .B(n8978), .ZN(n11040) );
  INV_X1 U11360 ( .A(n11040), .ZN(n9977) );
  NAND2_X1 U11361 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  AND2_X1 U11362 ( .A1(n8983), .A2(n8982), .ZN(n9978) );
  OR2_X1 U11363 ( .A1(n12082), .A2(n9978), .ZN(n8986) );
  OR2_X1 U11364 ( .A1(n9714), .A2(SI_7_), .ZN(n8985) );
  OAI211_X1 U11365 ( .C1(n9977), .C2(n6502), .A(n8986), .B(n8985), .ZN(n14962)
         );
  OR2_X1 U11366 ( .A1(n12602), .A2(n14962), .ZN(n12176) );
  NAND2_X1 U11367 ( .A1(n12602), .A2(n14962), .ZN(n12177) );
  NAND2_X1 U11368 ( .A1(n12176), .A2(n12177), .ZN(n12172) );
  XNOR2_X1 U11369 ( .A(n12172), .B(n8926), .ZN(n14964) );
  NAND2_X1 U11370 ( .A1(n14965), .A2(n14964), .ZN(n14963) );
  INV_X1 U11371 ( .A(n14964), .ZN(n8987) );
  NAND2_X1 U11372 ( .A1(n8987), .A2(n12602), .ZN(n8988) );
  NAND2_X1 U11373 ( .A1(n14963), .A2(n8988), .ZN(n14977) );
  INV_X1 U11374 ( .A(SI_8_), .ZN(n9956) );
  OR2_X1 U11375 ( .A1(n9714), .A2(n9956), .ZN(n8995) );
  XNOR2_X1 U11376 ( .A(n8990), .B(n8989), .ZN(n9957) );
  OR2_X1 U11377 ( .A1(n12082), .A2(n9957), .ZN(n8994) );
  NAND2_X1 U11378 ( .A1(n9005), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8992) );
  XNOR2_X1 U11379 ( .A(n8992), .B(P3_IR_REG_8__SCAN_IN), .ZN(n9900) );
  OR2_X1 U11380 ( .A1(n6508), .A2(n10921), .ZN(n8993) );
  XNOR2_X1 U11381 ( .A(n15170), .B(n8926), .ZN(n9002) );
  NAND2_X1 U11382 ( .A1(n6503), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9001) );
  INV_X1 U11383 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n8996) );
  OR2_X1 U11384 ( .A1(n12085), .A2(n8996), .ZN(n9000) );
  XNOR2_X1 U11385 ( .A(n9017), .B(P3_REG3_REG_8__SCAN_IN), .ZN(n14984) );
  OR2_X1 U11386 ( .A1(n9723), .A2(n14984), .ZN(n8999) );
  INV_X1 U11387 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n8997) );
  OR2_X1 U11388 ( .A1(n12086), .A2(n8997), .ZN(n8998) );
  NAND4_X1 U11389 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(n12601) );
  XNOR2_X1 U11390 ( .A(n9002), .B(n12601), .ZN(n14976) );
  INV_X1 U11391 ( .A(n9002), .ZN(n9003) );
  NAND2_X1 U11392 ( .A1(n9003), .A2(n12601), .ZN(n9004) );
  NOR2_X1 U11393 ( .A1(n9005), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9008) );
  OR2_X1 U11394 ( .A1(n9008), .A2(n8807), .ZN(n9006) );
  INV_X1 U11395 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9007) );
  MUX2_X1 U11396 ( .A(n9006), .B(P3_IR_REG_31__SCAN_IN), .S(n9007), .Z(n9009)
         );
  NAND2_X1 U11397 ( .A1(n9008), .A2(n9007), .ZN(n9049) );
  NAND2_X1 U11398 ( .A1(n9009), .A2(n9049), .ZN(n9950) );
  OR2_X1 U11399 ( .A1(n9011), .A2(n9010), .ZN(n9012) );
  AND2_X1 U11400 ( .A1(n9013), .A2(n9012), .ZN(n9949) );
  OR2_X1 U11401 ( .A1(n12082), .A2(n9949), .ZN(n9015) );
  OR2_X1 U11402 ( .A1(n9714), .A2(SI_9_), .ZN(n9014) );
  OAI211_X1 U11403 ( .C1(n15003), .C2(n6508), .A(n9015), .B(n9014), .ZN(n15179) );
  XNOR2_X1 U11404 ( .A(n15179), .B(n10776), .ZN(n9041) );
  NAND2_X1 U11405 ( .A1(n12083), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9023) );
  INV_X1 U11406 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n9016) );
  OR2_X1 U11407 ( .A1(n12086), .A2(n9016), .ZN(n9022) );
  INV_X1 U11408 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n9565) );
  INV_X1 U11409 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9662) );
  AOI21_X1 U11410 ( .B1(n9017), .B2(n9565), .A(n9662), .ZN(n9018) );
  OR2_X1 U11411 ( .A1(n9032), .A2(n9018), .ZN(n11449) );
  INV_X1 U11412 ( .A(n11449), .ZN(n11428) );
  OR2_X1 U11413 ( .A1(n9723), .A2(n11428), .ZN(n9021) );
  INV_X1 U11414 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n9019) );
  OR2_X1 U11415 ( .A1(n12085), .A2(n9019), .ZN(n9020) );
  NAND4_X1 U11416 ( .A1(n9023), .A2(n9022), .A3(n9021), .A4(n9020), .ZN(n12600) );
  XNOR2_X1 U11417 ( .A(n9041), .B(n12600), .ZN(n11444) );
  NAND2_X1 U11418 ( .A1(n9049), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9025) );
  INV_X1 U11419 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9024) );
  XNOR2_X1 U11420 ( .A(n9025), .B(n9024), .ZN(n15021) );
  INV_X1 U11421 ( .A(n15021), .ZN(n9986) );
  XNOR2_X1 U11422 ( .A(n9027), .B(n9026), .ZN(n9987) );
  OR2_X1 U11423 ( .A1(n12082), .A2(n9987), .ZN(n9029) );
  OR2_X1 U11424 ( .A1(n9714), .A2(SI_10_), .ZN(n9028) );
  OAI211_X1 U11425 ( .C1(n9986), .C2(n9855), .A(n9029), .B(n9028), .ZN(n15186)
         );
  XNOR2_X1 U11426 ( .A(n15186), .B(n8926), .ZN(n9040) );
  INV_X1 U11427 ( .A(n9040), .ZN(n9039) );
  NAND2_X1 U11428 ( .A1(n12083), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9038) );
  INV_X1 U11429 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n9030) );
  OR2_X1 U11430 ( .A1(n12085), .A2(n9030), .ZN(n9037) );
  OR2_X1 U11431 ( .A1(n9032), .A2(n9031), .ZN(n9033) );
  AND2_X1 U11432 ( .A1(n9044), .A2(n9033), .ZN(n11474) );
  OR2_X1 U11433 ( .A1(n9723), .A2(n11474), .ZN(n9036) );
  INV_X1 U11434 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9034) );
  OR2_X1 U11435 ( .A1(n12086), .A2(n9034), .ZN(n9035) );
  NAND4_X1 U11436 ( .A1(n9038), .A2(n9037), .A3(n9036), .A4(n9035), .ZN(n12599) );
  AND2_X1 U11437 ( .A1(n9039), .A2(n12599), .ZN(n9042) );
  XNOR2_X1 U11438 ( .A(n9040), .B(n12599), .ZN(n11468) );
  OR2_X1 U11439 ( .A1(n12600), .A2(n9041), .ZN(n11464) );
  AND2_X1 U11440 ( .A1(n11468), .A2(n11464), .ZN(n11465) );
  NAND2_X1 U11441 ( .A1(n12083), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9048) );
  INV_X1 U11442 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9043) );
  OR2_X1 U11443 ( .A1(n12085), .A2(n9043), .ZN(n9047) );
  INV_X1 U11444 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n9594) );
  XNOR2_X1 U11445 ( .A(n9044), .B(n9594), .ZN(n12840) );
  OR2_X1 U11446 ( .A1(n9723), .A2(n12840), .ZN(n9046) );
  INV_X1 U11447 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12839) );
  OR2_X1 U11448 ( .A1(n12086), .A2(n12839), .ZN(n9045) );
  NAND4_X1 U11449 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n12598) );
  INV_X1 U11450 ( .A(n12598), .ZN(n12539) );
  OAI21_X1 U11451 ( .B1(n9049), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9051) );
  INV_X1 U11452 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9050) );
  XNOR2_X1 U11453 ( .A(n9051), .B(n9050), .ZN(n15036) );
  INV_X1 U11454 ( .A(n15036), .ZN(n9908) );
  XNOR2_X1 U11455 ( .A(n9053), .B(n9052), .ZN(n14382) );
  OR2_X1 U11456 ( .A1(n12082), .A2(n14382), .ZN(n9055) );
  OR2_X1 U11457 ( .A1(n9714), .A2(SI_11_), .ZN(n9054) );
  OAI211_X1 U11458 ( .C1(n9908), .C2(n6507), .A(n9055), .B(n9054), .ZN(n12997)
         );
  XNOR2_X1 U11459 ( .A(n12997), .B(n8926), .ZN(n12450) );
  OR2_X1 U11460 ( .A1(n9057), .A2(n9056), .ZN(n9058) );
  NAND2_X1 U11461 ( .A1(n9059), .A2(n9058), .ZN(n9968) );
  OR2_X1 U11462 ( .A1(n12082), .A2(n9968), .ZN(n9064) );
  OR2_X1 U11463 ( .A1(n9714), .A2(n9967), .ZN(n9063) );
  OR2_X1 U11464 ( .A1(n9060), .A2(n8807), .ZN(n9061) );
  XNOR2_X1 U11465 ( .A(n9061), .B(P3_IR_REG_12__SCAN_IN), .ZN(n9911) );
  INV_X1 U11466 ( .A(n9911), .ZN(n15054) );
  OR2_X1 U11467 ( .A1(n6502), .A2(n15054), .ZN(n9062) );
  XNOR2_X1 U11468 ( .A(n12993), .B(n10776), .ZN(n9071) );
  NAND2_X1 U11469 ( .A1(n12083), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9070) );
  INV_X1 U11470 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n9861) );
  OR2_X1 U11471 ( .A1(n12085), .A2(n9861), .ZN(n9069) );
  NAND2_X1 U11472 ( .A1(n9065), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9066) );
  AND2_X1 U11473 ( .A1(n9074), .A2(n9066), .ZN(n12827) );
  OR2_X1 U11474 ( .A1(n9723), .A2(n12827), .ZN(n9068) );
  INV_X1 U11475 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12826) );
  OR2_X1 U11476 ( .A1(n12086), .A2(n12826), .ZN(n9067) );
  NAND4_X1 U11477 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n12597) );
  NAND2_X1 U11478 ( .A1(n9071), .A2(n12597), .ZN(n12454) );
  OAI21_X1 U11479 ( .B1(n12539), .B2(n12450), .A(n12454), .ZN(n9073) );
  NAND3_X1 U11480 ( .A1(n12454), .A2(n12539), .A3(n12450), .ZN(n9072) );
  OR2_X1 U11481 ( .A1(n9071), .A2(n12597), .ZN(n12453) );
  NAND2_X1 U11482 ( .A1(n12083), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9081) );
  AND2_X1 U11483 ( .A1(n9074), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9075) );
  NOR2_X1 U11484 ( .A1(n9100), .A2(n9075), .ZN(n12811) );
  OR2_X1 U11485 ( .A1(n9723), .A2(n12811), .ZN(n9080) );
  INV_X1 U11486 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n9076) );
  OR2_X1 U11487 ( .A1(n12086), .A2(n9076), .ZN(n9079) );
  INV_X1 U11488 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9077) );
  OR2_X1 U11489 ( .A1(n12085), .A2(n9077), .ZN(n9078) );
  NAND4_X1 U11490 ( .A1(n9081), .A2(n9080), .A3(n9079), .A4(n9078), .ZN(n12596) );
  INV_X1 U11491 ( .A(n12596), .ZN(n12457) );
  NAND2_X1 U11492 ( .A1(n9082), .A2(n10224), .ZN(n9083) );
  NAND2_X1 U11493 ( .A1(n9084), .A2(n9083), .ZN(n10008) );
  NAND2_X1 U11494 ( .A1(n12098), .A2(n10008), .ZN(n9089) );
  NAND2_X1 U11495 ( .A1(n9085), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9086) );
  MUX2_X1 U11496 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9086), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9087) );
  NAND2_X1 U11497 ( .A1(n9087), .A2(n6516), .ZN(n15070) );
  INV_X1 U11498 ( .A(n15070), .ZN(n9914) );
  OR2_X1 U11499 ( .A1(n6508), .A2(n9914), .ZN(n9088) );
  OAI211_X1 U11500 ( .C1(n9714), .C2(SI_13_), .A(n9089), .B(n9088), .ZN(n14450) );
  XNOR2_X1 U11501 ( .A(n14450), .B(n8926), .ZN(n12512) );
  OAI21_X1 U11502 ( .B1(n12514), .B2(n12457), .A(n12512), .ZN(n9091) );
  NAND2_X1 U11503 ( .A1(n12514), .A2(n12457), .ZN(n9090) );
  NAND2_X1 U11504 ( .A1(n9091), .A2(n9090), .ZN(n12395) );
  INV_X1 U11505 ( .A(n12395), .ZN(n9107) );
  OR2_X1 U11506 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  NAND2_X1 U11507 ( .A1(n9095), .A2(n9094), .ZN(n10043) );
  NAND2_X1 U11508 ( .A1(n10043), .A2(n12098), .ZN(n9099) );
  INV_X1 U11509 ( .A(n9714), .ZN(n9182) );
  INV_X1 U11510 ( .A(n9855), .ZN(n9181) );
  NAND2_X1 U11511 ( .A1(n6516), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9097) );
  INV_X1 U11512 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9096) );
  XNOR2_X1 U11513 ( .A(n9097), .B(n9096), .ZN(n15091) );
  AOI22_X1 U11514 ( .A1(n9182), .A2(n10042), .B1(n9181), .B2(n15091), .ZN(
        n9098) );
  NAND2_X1 U11515 ( .A1(n9099), .A2(n9098), .ZN(n12389) );
  XNOR2_X1 U11516 ( .A(n12389), .B(n10776), .ZN(n9108) );
  NAND2_X1 U11517 ( .A1(n12083), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9105) );
  INV_X1 U11518 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12794) );
  OR2_X1 U11519 ( .A1(n12086), .A2(n12794), .ZN(n9104) );
  OR2_X1 U11520 ( .A1(n9100), .A2(n15087), .ZN(n9101) );
  AND2_X1 U11521 ( .A1(n9101), .A2(n9120), .ZN(n12795) );
  OR2_X1 U11522 ( .A1(n9723), .A2(n12795), .ZN(n9103) );
  INV_X1 U11523 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12900) );
  OR2_X1 U11524 ( .A1(n12085), .A2(n12900), .ZN(n9102) );
  NAND4_X1 U11525 ( .A1(n9105), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n12595) );
  XNOR2_X1 U11526 ( .A(n9108), .B(n12595), .ZN(n12396) );
  NAND2_X1 U11527 ( .A1(n9108), .A2(n12595), .ZN(n9109) );
  NAND2_X1 U11528 ( .A1(n12393), .A2(n9109), .ZN(n12571) );
  OR2_X1 U11529 ( .A1(n9111), .A2(n9110), .ZN(n9112) );
  NAND2_X1 U11530 ( .A1(n9113), .A2(n9112), .ZN(n10059) );
  OR2_X1 U11531 ( .A1(n10059), .A2(n12082), .ZN(n9119) );
  NAND2_X1 U11532 ( .A1(n9114), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9116) );
  XNOR2_X1 U11533 ( .A(n9116), .B(n9115), .ZN(n14408) );
  INV_X1 U11534 ( .A(n14408), .ZN(n9117) );
  AOI22_X1 U11535 ( .A1(n9182), .A2(SI_15_), .B1(n9181), .B2(n9117), .ZN(n9118) );
  XNOR2_X1 U11536 ( .A(n12896), .B(n8926), .ZN(n9126) );
  NAND2_X1 U11537 ( .A1(n12083), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9125) );
  INV_X1 U11538 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12897) );
  OR2_X1 U11539 ( .A1(n12085), .A2(n12897), .ZN(n9124) );
  NAND2_X1 U11540 ( .A1(n9120), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9121) );
  AND2_X1 U11541 ( .A1(n9136), .A2(n9121), .ZN(n12782) );
  OR2_X1 U11542 ( .A1(n9723), .A2(n12782), .ZN(n9123) );
  INV_X1 U11543 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14402) );
  OR2_X1 U11544 ( .A1(n12086), .A2(n14402), .ZN(n9122) );
  INV_X1 U11545 ( .A(n12477), .ZN(n12594) );
  AND2_X1 U11546 ( .A1(n9126), .A2(n12594), .ZN(n12568) );
  INV_X1 U11547 ( .A(n9126), .ZN(n9127) );
  NAND2_X1 U11548 ( .A1(n9127), .A2(n12477), .ZN(n12567) );
  OR2_X1 U11549 ( .A1(n9129), .A2(n9128), .ZN(n9130) );
  NAND2_X1 U11550 ( .A1(n9131), .A2(n9130), .ZN(n10090) );
  OR2_X1 U11551 ( .A1(n10090), .A2(n12082), .ZN(n9135) );
  OR2_X1 U11552 ( .A1(n9132), .A2(n8807), .ZN(n9133) );
  XNOR2_X1 U11553 ( .A(n9133), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U11554 ( .A1(n9182), .A2(SI_16_), .B1(n9181), .B2(n14418), .ZN(
        n9134) );
  XNOR2_X1 U11555 ( .A(n12974), .B(n10776), .ZN(n12474) );
  NAND2_X1 U11556 ( .A1(n12083), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9141) );
  INV_X1 U11557 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12892) );
  OR2_X1 U11558 ( .A1(n12085), .A2(n12892), .ZN(n9140) );
  AND2_X1 U11559 ( .A1(n9136), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9137) );
  NOR2_X1 U11560 ( .A1(n9154), .A2(n9137), .ZN(n12772) );
  OR2_X1 U11561 ( .A1(n9723), .A2(n12772), .ZN(n9139) );
  INV_X1 U11562 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12771) );
  OR2_X1 U11563 ( .A1(n12086), .A2(n12771), .ZN(n9138) );
  AND2_X1 U11564 ( .A1(n12474), .A2(n12486), .ZN(n9144) );
  INV_X1 U11565 ( .A(n12474), .ZN(n9142) );
  INV_X1 U11566 ( .A(n12486), .ZN(n12593) );
  NAND2_X1 U11567 ( .A1(n9142), .A2(n12593), .ZN(n9143) );
  OR2_X1 U11568 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  NAND2_X1 U11569 ( .A1(n9148), .A2(n9147), .ZN(n10095) );
  OR2_X1 U11570 ( .A1(n10095), .A2(n12082), .ZN(n9153) );
  NAND2_X1 U11571 ( .A1(n9149), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9150) );
  MUX2_X1 U11572 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9150), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9151) );
  AND2_X1 U11573 ( .A1(n9151), .A2(n6531), .ZN(n14433) );
  AOI22_X1 U11574 ( .A1(n9182), .A2(SI_17_), .B1(n9181), .B2(n14433), .ZN(
        n9152) );
  XNOR2_X1 U11575 ( .A(n12968), .B(n8926), .ZN(n9160) );
  NAND2_X1 U11576 ( .A1(n12083), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9159) );
  INV_X1 U11577 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12889) );
  OR2_X1 U11578 ( .A1(n12085), .A2(n12889), .ZN(n9158) );
  NOR2_X1 U11579 ( .A1(n9154), .A2(n9554), .ZN(n9155) );
  OR2_X1 U11580 ( .A1(n9170), .A2(n9155), .ZN(n12762) );
  INV_X1 U11581 ( .A(n12762), .ZN(n12489) );
  OR2_X1 U11582 ( .A1(n9723), .A2(n12489), .ZN(n9157) );
  INV_X1 U11583 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14443) );
  OR2_X1 U11584 ( .A1(n12086), .A2(n14443), .ZN(n9156) );
  XNOR2_X1 U11585 ( .A(n9160), .B(n12549), .ZN(n12484) );
  INV_X1 U11586 ( .A(n12549), .ZN(n12592) );
  NAND2_X1 U11587 ( .A1(n9160), .A2(n12592), .ZN(n9161) );
  OR2_X1 U11588 ( .A1(n9163), .A2(n9162), .ZN(n9164) );
  NAND2_X1 U11589 ( .A1(n9165), .A2(n9164), .ZN(n10246) );
  OR2_X1 U11590 ( .A1(n10246), .A2(n12082), .ZN(n9168) );
  NAND2_X1 U11591 ( .A1(n6531), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U11592 ( .A(n9166), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U11593 ( .A1(n9182), .A2(SI_18_), .B1(n9181), .B2(n12617), .ZN(
        n9167) );
  XNOR2_X1 U11594 ( .A(n12962), .B(n8926), .ZN(n9176) );
  NAND2_X1 U11595 ( .A1(n9731), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9175) );
  INV_X1 U11596 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12961) );
  OR2_X1 U11597 ( .A1(n9280), .A2(n12961), .ZN(n9174) );
  OR2_X1 U11598 ( .A1(n9170), .A2(n9169), .ZN(n9171) );
  AND2_X1 U11599 ( .A1(n9185), .A2(n9171), .ZN(n12752) );
  OR2_X1 U11600 ( .A1(n9723), .A2(n12752), .ZN(n9173) );
  INV_X1 U11601 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12751) );
  OR2_X1 U11602 ( .A1(n12086), .A2(n12751), .ZN(n9172) );
  XNOR2_X1 U11603 ( .A(n9176), .B(n12487), .ZN(n12546) );
  INV_X1 U11604 ( .A(n12487), .ZN(n12591) );
  OR2_X1 U11605 ( .A1(n9178), .A2(n9177), .ZN(n9179) );
  NAND2_X1 U11606 ( .A1(n9180), .A2(n9179), .ZN(n10329) );
  OR2_X1 U11607 ( .A1(n10329), .A2(n12082), .ZN(n9184) );
  AOI22_X1 U11608 ( .A1(n9182), .A2(SI_19_), .B1(n9181), .B2(n12614), .ZN(
        n9183) );
  XNOR2_X1 U11609 ( .A(n12956), .B(n8926), .ZN(n9191) );
  NAND2_X1 U11610 ( .A1(n12083), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9190) );
  INV_X1 U11611 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12883) );
  OR2_X1 U11612 ( .A1(n12085), .A2(n12883), .ZN(n9189) );
  NAND2_X1 U11613 ( .A1(n9185), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9186) );
  AND2_X1 U11614 ( .A1(n9199), .A2(n9186), .ZN(n12739) );
  OR2_X1 U11615 ( .A1(n9723), .A2(n12739), .ZN(n9188) );
  INV_X1 U11616 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12738) );
  OR2_X1 U11617 ( .A1(n12086), .A2(n12738), .ZN(n9187) );
  XNOR2_X1 U11618 ( .A(n9191), .B(n12551), .ZN(n12417) );
  NAND2_X1 U11619 ( .A1(n12418), .A2(n12417), .ZN(n9193) );
  INV_X1 U11620 ( .A(n12551), .ZN(n12590) );
  NAND2_X1 U11621 ( .A1(n9191), .A2(n12590), .ZN(n9192) );
  NAND2_X1 U11622 ( .A1(n9194), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11623 ( .A1(n9196), .A2(n9195), .ZN(n10577) );
  OR2_X1 U11624 ( .A1(n10577), .A2(n12082), .ZN(n9198) );
  XNOR2_X1 U11625 ( .A(n12950), .B(n10776), .ZN(n9205) );
  NAND2_X1 U11626 ( .A1(n9731), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9204) );
  INV_X1 U11627 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12949) );
  OR2_X1 U11628 ( .A1(n9280), .A2(n12949), .ZN(n9203) );
  AND2_X1 U11629 ( .A1(n9199), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9200) );
  NOR2_X1 U11630 ( .A1(n9215), .A2(n9200), .ZN(n12725) );
  OR2_X1 U11631 ( .A1(n9723), .A2(n12725), .ZN(n9202) );
  INV_X1 U11632 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12724) );
  OR2_X1 U11633 ( .A1(n12086), .A2(n12724), .ZN(n9201) );
  XNOR2_X1 U11634 ( .A(n9205), .B(n12589), .ZN(n12505) );
  INV_X1 U11635 ( .A(n9205), .ZN(n9206) );
  NAND2_X1 U11636 ( .A1(n9206), .A2(n12589), .ZN(n9207) );
  OR2_X1 U11637 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  NAND2_X1 U11638 ( .A1(n9211), .A2(n9210), .ZN(n10682) );
  OR2_X1 U11639 ( .A1(n10682), .A2(n12082), .ZN(n9213) );
  INV_X1 U11640 ( .A(SI_21_), .ZN(n10683) );
  XNOR2_X1 U11641 ( .A(n12877), .B(n10776), .ZN(n9221) );
  NAND2_X1 U11642 ( .A1(n9731), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9220) );
  INV_X1 U11643 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12945) );
  OR2_X1 U11644 ( .A1(n9280), .A2(n12945), .ZN(n9219) );
  NOR2_X1 U11645 ( .A1(n9215), .A2(n9214), .ZN(n9216) );
  OR2_X1 U11646 ( .A1(n9723), .A2(n7454), .ZN(n9218) );
  INV_X1 U11647 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12712) );
  OR2_X1 U11648 ( .A1(n12086), .A2(n12712), .ZN(n9217) );
  NAND4_X1 U11649 ( .A1(n9220), .A2(n9219), .A3(n9218), .A4(n9217), .ZN(n12588) );
  NAND2_X1 U11650 ( .A1(n9221), .A2(n12507), .ZN(n9224) );
  INV_X1 U11651 ( .A(n9221), .ZN(n9222) );
  NAND2_X1 U11652 ( .A1(n9222), .A2(n12588), .ZN(n9223) );
  NAND2_X1 U11653 ( .A1(n9224), .A2(n9223), .ZN(n12442) );
  XNOR2_X1 U11654 ( .A(n9226), .B(n9225), .ZN(n10697) );
  NAND2_X1 U11655 ( .A1(n10697), .A2(n12098), .ZN(n9228) );
  XNOR2_X1 U11656 ( .A(n12873), .B(n10776), .ZN(n9229) );
  AND2_X2 U11657 ( .A1(n9231), .A2(n9238), .ZN(n12523) );
  NAND2_X1 U11658 ( .A1(n9731), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9237) );
  INV_X1 U11659 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12941) );
  OR2_X1 U11660 ( .A1(n9280), .A2(n12941), .ZN(n9236) );
  OR2_X1 U11661 ( .A1(n9232), .A2(n12529), .ZN(n9233) );
  AND2_X1 U11662 ( .A1(n9233), .A2(n9243), .ZN(n12701) );
  OR2_X1 U11663 ( .A1(n9723), .A2(n12701), .ZN(n9235) );
  INV_X1 U11664 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12702) );
  OR2_X1 U11665 ( .A1(n12086), .A2(n12702), .ZN(n9234) );
  XNOR2_X1 U11666 ( .A(n9240), .B(n9239), .ZN(n10845) );
  NAND2_X1 U11667 ( .A1(n10845), .A2(n12098), .ZN(n9242) );
  XNOR2_X1 U11668 ( .A(n12691), .B(n10776), .ZN(n9259) );
  NAND2_X1 U11669 ( .A1(n9731), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9247) );
  INV_X1 U11670 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12937) );
  OR2_X1 U11671 ( .A1(n9280), .A2(n12937), .ZN(n9246) );
  AOI21_X1 U11672 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(n9243), .A(n9251), .ZN(
        n12688) );
  OR2_X1 U11673 ( .A1(n9723), .A2(n12688), .ZN(n9245) );
  INV_X1 U11674 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12689) );
  OR2_X1 U11675 ( .A1(n12086), .A2(n12689), .ZN(n9244) );
  NAND2_X1 U11676 ( .A1(n9259), .A2(n12526), .ZN(n9260) );
  INV_X1 U11677 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11540) );
  XNOR2_X1 U11678 ( .A(n9248), .B(n11540), .ZN(n11136) );
  NAND2_X1 U11679 ( .A1(n11136), .A2(n12098), .ZN(n9250) );
  INV_X1 U11680 ( .A(SI_24_), .ZN(n11137) );
  XNOR2_X1 U11681 ( .A(n12676), .B(n10776), .ZN(n9258) );
  NAND2_X1 U11682 ( .A1(n9731), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9257) );
  INV_X1 U11683 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12933) );
  OR2_X1 U11684 ( .A1(n9280), .A2(n12933), .ZN(n9256) );
  INV_X1 U11685 ( .A(n9251), .ZN(n9253) );
  AOI21_X1 U11686 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(n9253), .A(n9252), .ZN(
        n12673) );
  OR2_X1 U11687 ( .A1(n9723), .A2(n12673), .ZN(n9255) );
  INV_X1 U11688 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12674) );
  OR2_X1 U11689 ( .A1(n12086), .A2(n12674), .ZN(n9254) );
  NAND2_X1 U11690 ( .A1(n9258), .A2(n12403), .ZN(n9261) );
  OAI21_X1 U11691 ( .B1(n9258), .B2(n12403), .A(n9261), .ZN(n12495) );
  INV_X1 U11692 ( .A(n9259), .ZN(n12400) );
  INV_X1 U11693 ( .A(n12526), .ZN(n12587) );
  INV_X1 U11694 ( .A(n9261), .ZN(n12465) );
  XNOR2_X1 U11695 ( .A(n11480), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9262) );
  XNOR2_X1 U11696 ( .A(n9263), .B(n9262), .ZN(n11279) );
  NAND2_X1 U11697 ( .A1(n11279), .A2(n12098), .ZN(n9265) );
  XNOR2_X1 U11698 ( .A(n12858), .B(n10776), .ZN(n9272) );
  NAND2_X1 U11699 ( .A1(n9731), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9271) );
  INV_X1 U11700 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12930) );
  OR2_X1 U11701 ( .A1(n9280), .A2(n12930), .ZN(n9270) );
  INV_X1 U11702 ( .A(n9282), .ZN(n9266) );
  AOI21_X1 U11703 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n9267), .A(n9266), .ZN(
        n12470) );
  OR2_X1 U11704 ( .A1(n9723), .A2(n12470), .ZN(n9269) );
  INV_X1 U11705 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n11784) );
  OR2_X1 U11706 ( .A1(n12086), .A2(n11784), .ZN(n9268) );
  INV_X1 U11707 ( .A(n12585), .ZN(n12265) );
  NAND2_X1 U11708 ( .A1(n9272), .A2(n12265), .ZN(n9275) );
  INV_X1 U11709 ( .A(n9272), .ZN(n9273) );
  NAND2_X1 U11710 ( .A1(n9273), .A2(n12585), .ZN(n9274) );
  AND2_X1 U11711 ( .A1(n9275), .A2(n9274), .ZN(n12464) );
  NAND2_X1 U11712 ( .A1(n12462), .A2(n9275), .ZN(n12557) );
  XNOR2_X1 U11713 ( .A(n13689), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9276) );
  XNOR2_X1 U11714 ( .A(n9277), .B(n9276), .ZN(n11347) );
  NAND2_X1 U11715 ( .A1(n11347), .A2(n12098), .ZN(n9279) );
  XNOR2_X1 U11716 ( .A(n12559), .B(n6467), .ZN(n9287) );
  NAND2_X1 U11717 ( .A1(n9731), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9286) );
  INV_X1 U11718 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n11761) );
  OR2_X1 U11719 ( .A1(n9280), .A2(n11761), .ZN(n9285) );
  AOI21_X1 U11720 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n9282), .A(n9281), .ZN(
        n12563) );
  OR2_X1 U11721 ( .A1(n9723), .A2(n12563), .ZN(n9284) );
  INV_X1 U11722 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n11767) );
  OR2_X1 U11723 ( .A1(n12086), .A2(n11767), .ZN(n9283) );
  NOR2_X1 U11724 ( .A1(n9287), .A2(n12584), .ZN(n9288) );
  AOI21_X1 U11725 ( .B1(n9287), .B2(n12584), .A(n9288), .ZN(n12558) );
  NAND2_X1 U11726 ( .A1(n12557), .A2(n12558), .ZN(n12556) );
  INV_X1 U11727 ( .A(n9288), .ZN(n9289) );
  NAND2_X1 U11728 ( .A1(n12556), .A2(n9289), .ZN(n9290) );
  NAND2_X1 U11729 ( .A1(n9290), .A2(n9291), .ZN(n12434) );
  OAI21_X1 U11730 ( .B1(n9291), .B2(n9290), .A(n12434), .ZN(n9323) );
  INV_X1 U11731 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11732 ( .A1(n10165), .A2(n9292), .ZN(n9294) );
  OR2_X1 U11733 ( .A1(n11346), .A2(n9305), .ZN(n9293) );
  NOR2_X1 U11734 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9298) );
  NOR4_X1 U11735 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9297) );
  NOR4_X1 U11736 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9296) );
  NOR4_X1 U11737 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9295) );
  NAND4_X1 U11738 ( .A1(n9298), .A2(n9297), .A3(n9296), .A4(n9295), .ZN(n9304)
         );
  NOR4_X1 U11739 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9302) );
  NOR4_X1 U11740 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9301) );
  NOR4_X1 U11741 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9300) );
  NOR4_X1 U11742 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9299) );
  NAND4_X1 U11743 ( .A1(n9302), .A2(n9301), .A3(n9300), .A4(n9299), .ZN(n9303)
         );
  NAND3_X1 U11744 ( .A1(n12999), .A2(n13001), .A3(n9741), .ZN(n9327) );
  NAND2_X1 U11745 ( .A1(n6513), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9307) );
  MUX2_X1 U11746 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9307), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9308) );
  INV_X1 U11747 ( .A(n13000), .ZN(n9309) );
  INV_X1 U11748 ( .A(n12293), .ZN(n9310) );
  NOR2_X1 U11749 ( .A1(n9327), .A2(n9310), .ZN(n9808) );
  NAND2_X1 U11750 ( .A1(n9311), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9312) );
  MUX2_X1 U11751 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9312), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9313) );
  OR2_X1 U11752 ( .A1(n12614), .A2(n9797), .ZN(n9316) );
  NAND2_X1 U11753 ( .A1(n12139), .A2(n10579), .ZN(n9314) );
  XNOR2_X1 U11754 ( .A(n12297), .B(n9314), .ZN(n9315) );
  NAND2_X1 U11755 ( .A1(n9316), .A2(n9315), .ZN(n9809) );
  NAND3_X1 U11756 ( .A1(n9808), .A2(n15185), .A3(n9809), .ZN(n9322) );
  INV_X1 U11757 ( .A(n12999), .ZN(n9317) );
  NAND2_X1 U11758 ( .A1(n9332), .A2(n12293), .ZN(n9811) );
  INV_X1 U11759 ( .A(n12132), .ZN(n9319) );
  AND2_X1 U11760 ( .A1(n12297), .A2(n9319), .ZN(n9320) );
  NAND2_X1 U11761 ( .A1(n12614), .A2(n9320), .ZN(n9805) );
  OR2_X1 U11762 ( .A1(n9811), .A2(n9805), .ZN(n9321) );
  NAND2_X1 U11763 ( .A1(n9323), .A2(n14974), .ZN(n9349) );
  INV_X1 U11764 ( .A(n12855), .ZN(n12273) );
  INV_X1 U11765 ( .A(n9327), .ZN(n9324) );
  NAND2_X1 U11766 ( .A1(n9324), .A2(n9325), .ZN(n9326) );
  INV_X1 U11767 ( .A(n12655), .ZN(n9345) );
  NAND2_X1 U11768 ( .A1(n9327), .A2(n9809), .ZN(n9330) );
  INV_X2 U11769 ( .A(n12286), .ZN(n12276) );
  OAI211_X1 U11770 ( .C1(n12292), .C2(n12276), .A(n9826), .B(n9856), .ZN(n9328) );
  INV_X1 U11771 ( .A(n9328), .ZN(n9329) );
  OAI211_X1 U11772 ( .C1(n9332), .C2(n9805), .A(n9330), .B(n9329), .ZN(n9331)
         );
  NAND2_X1 U11773 ( .A1(n9331), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9335) );
  INV_X1 U11774 ( .A(n9332), .ZN(n9333) );
  NAND3_X1 U11775 ( .A1(n9333), .A2(n10678), .A3(n12293), .ZN(n9334) );
  INV_X1 U11776 ( .A(n9336), .ZN(n12294) );
  NAND2_X1 U11777 ( .A1(n12294), .A2(n9883), .ZN(n9857) );
  AND2_X1 U11778 ( .A1(n9855), .A2(n9857), .ZN(n11454) );
  NAND2_X1 U11779 ( .A1(n12083), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9343) );
  INV_X1 U11780 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12851) );
  OR2_X1 U11781 ( .A1(n12085), .A2(n12851), .ZN(n9342) );
  INV_X1 U11782 ( .A(n9338), .ZN(n9337) );
  INV_X1 U11783 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U11784 ( .A1(n9337), .A2(n9562), .ZN(n9800) );
  NAND2_X1 U11785 ( .A1(n9338), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9339) );
  OR2_X1 U11786 ( .A1(n9723), .A2(n12645), .ZN(n9341) );
  INV_X1 U11787 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12644) );
  OR2_X1 U11788 ( .A1(n12086), .A2(n12644), .ZN(n9340) );
  INV_X1 U11789 ( .A(n9738), .ZN(n12582) );
  AOI22_X1 U11790 ( .A1(n12572), .A2(n12584), .B1(n12582), .B2(n12573), .ZN(
        n12653) );
  INV_X1 U11791 ( .A(n12292), .ZN(n9745) );
  OAI22_X1 U11792 ( .A1(n12653), .A2(n12530), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9581), .ZN(n9344) );
  AOI21_X1 U11793 ( .B1(n9345), .B2(n12532), .A(n9344), .ZN(n9346) );
  INV_X1 U11794 ( .A(n9347), .ZN(n9348) );
  NAND2_X1 U11795 ( .A1(n9349), .A2(n9348), .ZN(P3_U3154) );
  NAND2_X1 U11796 ( .A1(n9377), .A2(n12382), .ZN(n9350) );
  XNOR2_X1 U11797 ( .A(n9353), .B(n9352), .ZN(n9354) );
  NAND2_X1 U11798 ( .A1(n9354), .A2(n14676), .ZN(n9358) );
  OAI22_X1 U11799 ( .A1(n9356), .A2(n14520), .B1(n9355), .B2(n14522), .ZN(
        n9357) );
  INV_X1 U11800 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9360) );
  NOR2_X1 U11801 ( .A1(n14687), .A2(n9360), .ZN(n9361) );
  INV_X1 U11802 ( .A(n12031), .ZN(n10643) );
  AND2_X1 U11803 ( .A1(n10643), .A2(n10644), .ZN(n9364) );
  NAND2_X1 U11804 ( .A1(n14695), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9366) );
  NAND2_X1 U11805 ( .A1(n9367), .A2(n9366), .ZN(P1_U3557) );
  NOR2_X1 U11806 ( .A1(n9368), .A2(n14661), .ZN(n9372) );
  NAND2_X1 U11807 ( .A1(n9368), .A2(n14676), .ZN(n9371) );
  NAND2_X1 U11808 ( .A1(n9369), .A2(n14684), .ZN(n9370) );
  AOI22_X1 U11809 ( .A1(n14498), .A2(n13871), .B1(n13869), .B2(n14642), .ZN(
        n9373) );
  OAI21_X1 U11810 ( .B1(n9374), .B2(n14672), .A(n9373), .ZN(n9375) );
  AOI21_X1 U11811 ( .B1(n6965), .B2(n14033), .A(n14644), .ZN(n9378) );
  NAND2_X1 U11812 ( .A1(n9378), .A2(n9377), .ZN(n14036) );
  NAND2_X1 U11813 ( .A1(n14039), .A2(n14036), .ZN(n9668) );
  INV_X1 U11814 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9379) );
  OR2_X1 U11815 ( .A1(n14687), .A2(n9379), .ZN(n9380) );
  INV_X1 U11816 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n9489) );
  INV_X1 U11817 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9419) );
  XOR2_X1 U11818 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9419), .Z(n9483) );
  INV_X1 U11819 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9415) );
  XNOR2_X1 U11820 ( .A(n9415), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n9479) );
  INV_X1 U11821 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10323) );
  XOR2_X1 U11822 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n13950), .Z(n9455) );
  XOR2_X1 U11823 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n9386), .Z(n9432) );
  NAND2_X1 U11824 ( .A1(n9436), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9435) );
  INV_X1 U11825 ( .A(n9435), .ZN(n9383) );
  NAND2_X1 U11826 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n9390), .ZN(n9392) );
  NAND2_X1 U11827 ( .A1(n9431), .A2(n13916), .ZN(n9391) );
  NAND2_X1 U11828 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n9394), .ZN(n9396) );
  NAND2_X1 U11829 ( .A1(n9429), .A2(n9430), .ZN(n9395) );
  NAND2_X1 U11830 ( .A1(n9396), .A2(n9395), .ZN(n9397) );
  NAND2_X1 U11831 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n9397), .ZN(n9399) );
  XOR2_X1 U11832 ( .A(n9397), .B(P3_ADDR_REG_5__SCAN_IN), .Z(n9443) );
  NAND2_X1 U11833 ( .A1(n9443), .A2(n9442), .ZN(n9398) );
  INV_X1 U11834 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11835 ( .A1(n9402), .A2(n9401), .ZN(n9404) );
  XOR2_X1 U11836 ( .A(n9402), .B(n9401), .Z(n9428) );
  NAND2_X1 U11837 ( .A1(n9428), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U11838 ( .A1(n9404), .A2(n9403), .ZN(n9456) );
  NAND2_X1 U11839 ( .A1(n9455), .A2(n9456), .ZN(n9405) );
  XNOR2_X1 U11840 ( .A(n9407), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U11841 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n9424), .ZN(n9409) );
  NOR2_X1 U11842 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n9424), .ZN(n9408) );
  XOR2_X1 U11843 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n13986), .Z(n9467) );
  NAND2_X1 U11844 ( .A1(n9468), .A2(n9467), .ZN(n9410) );
  XOR2_X1 U11845 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .Z(n9423) );
  INV_X1 U11846 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9473) );
  NOR2_X1 U11847 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n9473), .ZN(n9413) );
  INV_X1 U11848 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9412) );
  NOR2_X1 U11849 ( .A1(n9479), .A2(n9478), .ZN(n9414) );
  INV_X1 U11850 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U11851 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n9416), .ZN(n9417) );
  INV_X1 U11852 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14622) );
  AOI22_X1 U11853 ( .A1(n9421), .A2(n9417), .B1(P3_ADDR_REG_15__SCAN_IN), .B2(
        n14622), .ZN(n9482) );
  NAND2_X1 U11854 ( .A1(n9483), .A2(n9482), .ZN(n9418) );
  XNOR2_X1 U11855 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9487), .ZN(n9488) );
  XOR2_X1 U11856 ( .A(n9489), .B(n9488), .Z(n14398) );
  XNOR2_X1 U11857 ( .A(n14622), .B(P3_ADDR_REG_15__SCAN_IN), .ZN(n9420) );
  XNOR2_X1 U11858 ( .A(n9421), .B(n9420), .ZN(n14568) );
  XOR2_X1 U11859 ( .A(n9423), .B(n9422), .Z(n9469) );
  XNOR2_X1 U11860 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n9424), .ZN(n9425) );
  XNOR2_X1 U11861 ( .A(n9425), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n9465) );
  XOR2_X1 U11862 ( .A(n9427), .B(n9426), .Z(n9461) );
  XNOR2_X1 U11863 ( .A(n9428), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15215) );
  XNOR2_X1 U11864 ( .A(n9430), .B(n9429), .ZN(n9440) );
  AND2_X1 U11865 ( .A1(n9440), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9441) );
  XOR2_X1 U11866 ( .A(n9431), .B(n13916), .Z(n15218) );
  XOR2_X1 U11867 ( .A(n9433), .B(n9432), .Z(n14378) );
  NOR2_X1 U11868 ( .A1(n9437), .A2(n7038), .ZN(n9438) );
  OAI21_X1 U11869 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9436), .A(n9435), .ZN(
        n15212) );
  NAND2_X1 U11870 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15212), .ZN(n15222) );
  NOR2_X1 U11871 ( .A1(n15222), .A2(n15221), .ZN(n15220) );
  NAND2_X1 U11872 ( .A1(n14378), .A2(n14377), .ZN(n14376) );
  NAND2_X1 U11873 ( .A1(n15218), .A2(n15217), .ZN(n9439) );
  AOI21_X1 U11874 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n9439), .A(n15216), .ZN(
        n15208) );
  XNOR2_X1 U11875 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n9440), .ZN(n15207) );
  NOR2_X1 U11876 ( .A1(n15208), .A2(n15207), .ZN(n15206) );
  NAND2_X1 U11877 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  INV_X1 U11878 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15210) );
  XOR2_X1 U11879 ( .A(n9447), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n9449) );
  XOR2_X1 U11880 ( .A(n9449), .B(n9448), .Z(n14385) );
  INV_X1 U11881 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9450) );
  NOR2_X1 U11882 ( .A1(n9451), .A2(n9450), .ZN(n9452) );
  XNOR2_X1 U11883 ( .A(n9456), .B(n9455), .ZN(n9457) );
  NAND2_X1 U11884 ( .A1(n9459), .A2(n9457), .ZN(n9460) );
  XNOR2_X2 U11885 ( .A(n9459), .B(n9458), .ZN(n14389) );
  INV_X1 U11886 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14388) );
  NAND2_X1 U11887 ( .A1(n14389), .A2(n14388), .ZN(n14387) );
  NAND2_X1 U11888 ( .A1(n9460), .A2(n14387), .ZN(n9462) );
  NOR2_X1 U11889 ( .A1(n9461), .A2(n9462), .ZN(n9463) );
  XNOR2_X1 U11890 ( .A(n9462), .B(n9461), .ZN(n14392) );
  INV_X1 U11891 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14391) );
  NOR2_X1 U11892 ( .A1(n14392), .A2(n14391), .ZN(n14390) );
  INV_X1 U11893 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14394) );
  NOR2_X1 U11894 ( .A1(n9465), .A2(n9464), .ZN(n9466) );
  NOR2_X2 U11895 ( .A1(n14393), .A2(n9466), .ZN(n14551) );
  XNOR2_X1 U11896 ( .A(n9468), .B(n9467), .ZN(n14552) );
  NAND2_X1 U11897 ( .A1(n14551), .A2(n14552), .ZN(n14550) );
  NAND2_X1 U11898 ( .A1(n9469), .A2(n9471), .ZN(n9472) );
  INV_X1 U11899 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14555) );
  XOR2_X1 U11900 ( .A(n9473), .B(P3_ADDR_REG_13__SCAN_IN), .Z(n9475) );
  XOR2_X1 U11901 ( .A(n9475), .B(n9474), .Z(n9477) );
  NOR2_X2 U11902 ( .A1(n9476), .A2(n9477), .ZN(n14558) );
  INV_X1 U11903 ( .A(n14558), .ZN(n14559) );
  INV_X1 U11904 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U11905 ( .A1(n9477), .A2(n9476), .ZN(n14560) );
  NAND2_X1 U11906 ( .A1(n14561), .A2(n14560), .ZN(n14557) );
  AND2_X2 U11907 ( .A1(n14559), .A2(n14557), .ZN(n9481) );
  XOR2_X1 U11908 ( .A(n9479), .B(n9478), .Z(n9480) );
  NOR2_X2 U11909 ( .A1(n9481), .A2(n9480), .ZN(n14563) );
  INV_X1 U11910 ( .A(n14563), .ZN(n14564) );
  INV_X1 U11911 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14566) );
  NAND2_X1 U11912 ( .A1(n9481), .A2(n9480), .ZN(n14565) );
  XNOR2_X1 U11913 ( .A(n9483), .B(n9482), .ZN(n14571) );
  INV_X1 U11914 ( .A(n14396), .ZN(n9486) );
  NAND2_X1 U11915 ( .A1(n14398), .A2(n14397), .ZN(n9484) );
  NAND2_X1 U11916 ( .A1(n9484), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n9485) );
  AND2_X2 U11917 ( .A1(n9486), .A2(n9485), .ZN(n14371) );
  INV_X1 U11918 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n9497) );
  XOR2_X1 U11919 ( .A(n9497), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n9492) );
  NOR2_X1 U11920 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9487), .ZN(n9491) );
  NOR2_X1 U11921 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  NOR2_X1 U11922 ( .A1(n9491), .A2(n9490), .ZN(n9496) );
  XNOR2_X1 U11923 ( .A(n9492), .B(n9496), .ZN(n14372) );
  XNOR2_X1 U11924 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9493) );
  XNOR2_X1 U11925 ( .A(n9493), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n9494) );
  INV_X1 U11926 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14638) );
  NOR2_X1 U11927 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n14638), .ZN(n9495) );
  OAI22_X1 U11928 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9497), .B1(n9496), .B2(
        n9495), .ZN(n9664) );
  AOI22_X1 U11929 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(keyinput_f44), .ZN(n9498) );
  OAI221_X1 U11930 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P3_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n9498), .ZN(n9505) );
  AOI22_X1 U11931 ( .A1(SI_6_), .A2(keyinput_f26), .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n9499) );
  OAI221_X1 U11932 ( .B1(SI_6_), .B2(keyinput_f26), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n9499), .ZN(n9504) );
  AOI22_X1 U11933 ( .A1(SI_18_), .A2(keyinput_f14), .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n9500) );
  OAI221_X1 U11934 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n9500), .ZN(n9503) );
  AOI22_X1 U11935 ( .A1(SI_10_), .A2(keyinput_f22), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n9501) );
  OAI221_X1 U11936 ( .B1(SI_10_), .B2(keyinput_f22), .C1(SI_21_), .C2(
        keyinput_f11), .A(n9501), .ZN(n9502) );
  NOR4_X1 U11937 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n9532)
         );
  XOR2_X1 U11938 ( .A(P3_U3151), .B(keyinput_f34), .Z(n9512) );
  AOI22_X1 U11939 ( .A1(SI_16_), .A2(keyinput_f16), .B1(n14993), .B2(
        keyinput_f54), .ZN(n9506) );
  OAI221_X1 U11940 ( .B1(SI_16_), .B2(keyinput_f16), .C1(n14993), .C2(
        keyinput_f54), .A(n9506), .ZN(n9511) );
  AOI22_X1 U11941 ( .A1(SI_0_), .A2(keyinput_f32), .B1(SI_8_), .B2(
        keyinput_f24), .ZN(n9507) );
  OAI221_X1 U11942 ( .B1(SI_0_), .B2(keyinput_f32), .C1(SI_8_), .C2(
        keyinput_f24), .A(n9507), .ZN(n9510) );
  AOI22_X1 U11943 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n9508) );
  OAI221_X1 U11944 ( .B1(SI_3_), .B2(keyinput_f29), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n9508), .ZN(n9509) );
  NOR4_X1 U11945 ( .A1(n9512), .A2(n9511), .A3(n9510), .A4(n9509), .ZN(n9531)
         );
  AOI22_X1 U11946 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n9513) );
  OAI221_X1 U11947 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n9513), .ZN(n9520) );
  AOI22_X1 U11948 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n9514) );
  OAI221_X1 U11949 ( .B1(SI_23_), .B2(keyinput_f9), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n9514), .ZN(n9519) );
  AOI22_X1 U11950 ( .A1(keyinput_f33), .A2(P3_RD_REG_SCAN_IN), .B1(SI_25_), 
        .B2(keyinput_f7), .ZN(n9515) );
  OAI221_X1 U11951 ( .B1(keyinput_f33), .B2(P3_RD_REG_SCAN_IN), .C1(SI_25_), 
        .C2(keyinput_f7), .A(n9515), .ZN(n9518) );
  AOI22_X1 U11952 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(SI_28_), .B2(keyinput_f4), .ZN(n9516) );
  OAI221_X1 U11953 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        SI_28_), .C2(keyinput_f4), .A(n9516), .ZN(n9517) );
  NOR4_X1 U11954 ( .A1(n9520), .A2(n9519), .A3(n9518), .A4(n9517), .ZN(n9530)
         );
  AOI22_X1 U11955 ( .A1(SI_24_), .A2(keyinput_f8), .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n9521) );
  OAI221_X1 U11956 ( .B1(SI_24_), .B2(keyinput_f8), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n9521), .ZN(n9528) );
  AOI22_X1 U11957 ( .A1(SI_20_), .A2(keyinput_f12), .B1(SI_27_), .B2(
        keyinput_f5), .ZN(n9522) );
  OAI221_X1 U11958 ( .B1(SI_20_), .B2(keyinput_f12), .C1(SI_27_), .C2(
        keyinput_f5), .A(n9522), .ZN(n9527) );
  AOI22_X1 U11959 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n9523) );
  OAI221_X1 U11960 ( .B1(SI_2_), .B2(keyinput_f30), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n9523), .ZN(n9526) );
  AOI22_X1 U11961 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_1_), .B2(
        keyinput_f31), .ZN(n9524) );
  OAI221_X1 U11962 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_1_), .C2(
        keyinput_f31), .A(n9524), .ZN(n9525) );
  NOR4_X1 U11963 ( .A1(n9528), .A2(n9527), .A3(n9526), .A4(n9525), .ZN(n9529)
         );
  NAND4_X1 U11964 ( .A1(n9532), .A2(n9531), .A3(n9530), .A4(n9529), .ZN(n9576)
         );
  AOI22_X1 U11965 ( .A1(n10330), .A2(keyinput_f13), .B1(keyinput_f19), .B2(
        n10007), .ZN(n9533) );
  OAI221_X1 U11966 ( .B1(n10330), .B2(keyinput_f13), .C1(n10007), .C2(
        keyinput_f19), .A(n9533), .ZN(n9542) );
  XNOR2_X1 U11967 ( .A(SI_5_), .B(keyinput_f27), .ZN(n9537) );
  XNOR2_X1 U11968 ( .A(SI_4_), .B(keyinput_f28), .ZN(n9536) );
  XNOR2_X1 U11969 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_f47), .ZN(n9535)
         );
  XNOR2_X1 U11970 ( .A(SI_7_), .B(keyinput_f25), .ZN(n9534) );
  NAND4_X1 U11971 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(n9541)
         );
  INV_X1 U11972 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n9538) );
  XNOR2_X1 U11973 ( .A(keyinput_f38), .B(n9538), .ZN(n9540) );
  INV_X1 U11974 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9581) );
  XNOR2_X1 U11975 ( .A(keyinput_f36), .B(n9581), .ZN(n9539) );
  NOR4_X1 U11976 ( .A1(n9542), .A2(n9541), .A3(n9540), .A4(n9539), .ZN(n9574)
         );
  INV_X1 U11977 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9579) );
  INV_X1 U11978 ( .A(P3_WR_REG_SCAN_IN), .ZN(n9602) );
  AOI22_X1 U11979 ( .A1(n9579), .A2(keyinput_f52), .B1(keyinput_f0), .B2(n9602), .ZN(n9543) );
  OAI221_X1 U11980 ( .B1(n9579), .B2(keyinput_f52), .C1(n9602), .C2(
        keyinput_f0), .A(n9543), .ZN(n9550) );
  AOI22_X1 U11981 ( .A1(SI_31_), .A2(keyinput_f1), .B1(n15107), .B2(
        keyinput_f59), .ZN(n9544) );
  OAI221_X1 U11982 ( .B1(SI_31_), .B2(keyinput_f1), .C1(n15107), .C2(
        keyinput_f59), .A(n9544), .ZN(n9549) );
  INV_X1 U11983 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9603) );
  INV_X1 U11984 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9611) );
  AOI22_X1 U11985 ( .A1(n9603), .A2(keyinput_f55), .B1(keyinput_f41), .B2(
        n9611), .ZN(n9545) );
  OAI221_X1 U11986 ( .B1(n9603), .B2(keyinput_f55), .C1(n9611), .C2(
        keyinput_f41), .A(n9545), .ZN(n9548) );
  INV_X1 U11987 ( .A(SI_9_), .ZN(n9951) );
  AOI22_X1 U11988 ( .A1(n9967), .A2(keyinput_f20), .B1(keyinput_f23), .B2(
        n9951), .ZN(n9546) );
  OAI221_X1 U11989 ( .B1(n9967), .B2(keyinput_f20), .C1(n9951), .C2(
        keyinput_f23), .A(n9546), .ZN(n9547) );
  NOR4_X1 U11990 ( .A1(n9550), .A2(n9549), .A3(n9548), .A4(n9547), .ZN(n9573)
         );
  INV_X1 U11991 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n14961) );
  INV_X1 U11992 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15067) );
  AOI22_X1 U11993 ( .A1(n14961), .A2(keyinput_f35), .B1(n15067), .B2(
        keyinput_f56), .ZN(n9551) );
  OAI221_X1 U11994 ( .B1(n14961), .B2(keyinput_f35), .C1(n15067), .C2(
        keyinput_f56), .A(n9551), .ZN(n9559) );
  AOI22_X1 U11995 ( .A1(n10042), .A2(keyinput_f18), .B1(keyinput_f3), .B2(
        n12388), .ZN(n9552) );
  OAI221_X1 U11996 ( .B1(n10042), .B2(keyinput_f18), .C1(n12388), .C2(
        keyinput_f3), .A(n9552), .ZN(n9558) );
  INV_X1 U11997 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U11998 ( .A1(n14405), .A2(keyinput_f63), .B1(n9554), .B2(
        keyinput_f50), .ZN(n9553) );
  OAI221_X1 U11999 ( .B1(n14405), .B2(keyinput_f63), .C1(n9554), .C2(
        keyinput_f50), .A(n9553), .ZN(n9557) );
  INV_X1 U12000 ( .A(SI_17_), .ZN(n10094) );
  AOI22_X1 U12001 ( .A1(n10058), .A2(keyinput_f17), .B1(n10094), .B2(
        keyinput_f15), .ZN(n9555) );
  OAI221_X1 U12002 ( .B1(n10058), .B2(keyinput_f17), .C1(n10094), .C2(
        keyinput_f15), .A(n9555), .ZN(n9556) );
  NOR4_X1 U12003 ( .A1(n9559), .A2(n9558), .A3(n9557), .A4(n9556), .ZN(n9572)
         );
  INV_X1 U12004 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9583) );
  AOI22_X1 U12005 ( .A1(n7211), .A2(keyinput_f10), .B1(n9583), .B2(
        keyinput_f48), .ZN(n9560) );
  OAI221_X1 U12006 ( .B1(n7211), .B2(keyinput_f10), .C1(n9583), .C2(
        keyinput_f48), .A(n9560), .ZN(n9570) );
  AOI22_X1 U12007 ( .A1(n11349), .A2(keyinput_f6), .B1(n9562), .B2(
        keyinput_f42), .ZN(n9561) );
  OAI221_X1 U12008 ( .B1(n11349), .B2(keyinput_f6), .C1(n9562), .C2(
        keyinput_f42), .A(n9561), .ZN(n9569) );
  AOI22_X1 U12009 ( .A1(n9565), .A2(keyinput_f43), .B1(keyinput_f49), .B2(
        n9564), .ZN(n9563) );
  OAI221_X1 U12010 ( .B1(n9565), .B2(keyinput_f43), .C1(n9564), .C2(
        keyinput_f49), .A(n9563), .ZN(n9568) );
  AOI22_X1 U12011 ( .A1(n12529), .A2(keyinput_f57), .B1(keyinput_f45), .B2(
        n9214), .ZN(n9566) );
  OAI221_X1 U12012 ( .B1(n12529), .B2(keyinput_f57), .C1(n9214), .C2(
        keyinput_f45), .A(n9566), .ZN(n9567) );
  NOR4_X1 U12013 ( .A1(n9570), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(n9571)
         );
  NAND4_X1 U12014 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9571), .ZN(n9575)
         );
  OAI22_X1 U12015 ( .A1(n9576), .A2(n9575), .B1(keyinput_f53), .B2(
        P3_REG3_REG_9__SCAN_IN), .ZN(n9577) );
  AOI21_X1 U12016 ( .B1(keyinput_f53), .B2(P3_REG3_REG_9__SCAN_IN), .A(n9577), 
        .ZN(n9661) );
  AOI22_X1 U12017 ( .A1(n9579), .A2(keyinput_g52), .B1(n12500), .B2(
        keyinput_g51), .ZN(n9578) );
  OAI221_X1 U12018 ( .B1(n9579), .B2(keyinput_g52), .C1(n12500), .C2(
        keyinput_g51), .A(n9578), .ZN(n9589) );
  AOI22_X1 U12019 ( .A1(n9581), .A2(keyinput_g36), .B1(keyinput_g12), .B2(
        n10578), .ZN(n9580) );
  OAI221_X1 U12020 ( .B1(n9581), .B2(keyinput_g36), .C1(n10578), .C2(
        keyinput_g12), .A(n9580), .ZN(n9588) );
  AOI22_X1 U12021 ( .A1(n11137), .A2(keyinput_g8), .B1(n9583), .B2(
        keyinput_g48), .ZN(n9582) );
  OAI221_X1 U12022 ( .B1(n11137), .B2(keyinput_g8), .C1(n9583), .C2(
        keyinput_g48), .A(n9582), .ZN(n9587) );
  XNOR2_X1 U12023 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_g46), .ZN(n9585)
         );
  XNOR2_X1 U12024 ( .A(SI_4_), .B(keyinput_g28), .ZN(n9584) );
  NAND2_X1 U12025 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  NOR4_X1 U12026 ( .A1(n9589), .A2(n9588), .A3(n9587), .A4(n9586), .ZN(n9622)
         );
  AOI22_X1 U12027 ( .A1(SI_7_), .A2(keyinput_g25), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n9590) );
  OAI221_X1 U12028 ( .B1(SI_7_), .B2(keyinput_g25), .C1(SI_10_), .C2(
        keyinput_g22), .A(n9590), .ZN(n9598) );
  AOI22_X1 U12029 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n9591) );
  OAI221_X1 U12030 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n9591), .ZN(n9597) );
  AOI22_X1 U12031 ( .A1(n11349), .A2(keyinput_g6), .B1(n12529), .B2(
        keyinput_g57), .ZN(n9592) );
  OAI221_X1 U12032 ( .B1(n11349), .B2(keyinput_g6), .C1(n12529), .C2(
        keyinput_g57), .A(n9592), .ZN(n9596) );
  AOI22_X1 U12033 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(n9594), .B2(keyinput_g58), .ZN(n9593) );
  OAI221_X1 U12034 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        n9594), .C2(keyinput_g58), .A(n9593), .ZN(n9595) );
  NOR4_X1 U12035 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n9621)
         );
  AOI22_X1 U12036 ( .A1(n11281), .A2(keyinput_g7), .B1(keyinput_g44), .B2(
        n15120), .ZN(n9599) );
  OAI221_X1 U12037 ( .B1(n11281), .B2(keyinput_g7), .C1(n15120), .C2(
        keyinput_g44), .A(n9599), .ZN(n9608) );
  AOI22_X1 U12038 ( .A1(n14961), .A2(keyinput_g35), .B1(n14405), .B2(
        keyinput_g63), .ZN(n9600) );
  OAI221_X1 U12039 ( .B1(n14961), .B2(keyinput_g35), .C1(n14405), .C2(
        keyinput_g63), .A(n9600), .ZN(n9607) );
  AOI22_X1 U12040 ( .A1(n9603), .A2(keyinput_g55), .B1(keyinput_g0), .B2(n9602), .ZN(n9601) );
  OAI221_X1 U12041 ( .B1(n9603), .B2(keyinput_g55), .C1(n9602), .C2(
        keyinput_g0), .A(n9601), .ZN(n9606) );
  AOI22_X1 U12042 ( .A1(n10088), .A2(keyinput_g16), .B1(n10683), .B2(
        keyinput_g11), .ZN(n9604) );
  OAI221_X1 U12043 ( .B1(n10088), .B2(keyinput_g16), .C1(n10683), .C2(
        keyinput_g11), .A(n9604), .ZN(n9605) );
  NOR4_X1 U12044 ( .A1(n9608), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(n9620)
         );
  INV_X1 U12045 ( .A(P3_RD_REG_SCAN_IN), .ZN(n14375) );
  AOI22_X1 U12046 ( .A1(n10007), .A2(keyinput_g19), .B1(keyinput_g33), .B2(
        n14375), .ZN(n9609) );
  OAI221_X1 U12047 ( .B1(n10007), .B2(keyinput_g19), .C1(n14375), .C2(
        keyinput_g33), .A(n9609), .ZN(n9618) );
  AOI22_X1 U12048 ( .A1(n9611), .A2(keyinput_g41), .B1(keyinput_g23), .B2(
        n9951), .ZN(n9610) );
  OAI221_X1 U12049 ( .B1(n9611), .B2(keyinput_g41), .C1(n9951), .C2(
        keyinput_g23), .A(n9610), .ZN(n9617) );
  XNOR2_X1 U12050 ( .A(SI_18_), .B(keyinput_g14), .ZN(n9615) );
  XNOR2_X1 U12051 ( .A(SI_6_), .B(keyinput_g26), .ZN(n9614) );
  XNOR2_X1 U12052 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_g49), .ZN(n9613)
         );
  XNOR2_X1 U12053 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9612) );
  NAND4_X1 U12054 ( .A1(n9615), .A2(n9614), .A3(n9613), .A4(n9612), .ZN(n9616)
         );
  NOR3_X1 U12055 ( .A1(n9618), .A2(n9617), .A3(n9616), .ZN(n9619) );
  NAND4_X1 U12056 ( .A1(n9622), .A2(n9621), .A3(n9620), .A4(n9619), .ZN(n9659)
         );
  AOI22_X1 U12057 ( .A1(SI_22_), .A2(keyinput_g10), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n9623) );
  OAI221_X1 U12058 ( .B1(SI_22_), .B2(keyinput_g10), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n9623), .ZN(n9630) );
  AOI22_X1 U12059 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n9624) );
  OAI221_X1 U12060 ( .B1(SI_2_), .B2(keyinput_g30), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n9624), .ZN(n9629) );
  AOI22_X1 U12061 ( .A1(SI_14_), .A2(keyinput_g18), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n9625) );
  OAI221_X1 U12062 ( .B1(SI_14_), .B2(keyinput_g18), .C1(SI_17_), .C2(
        keyinput_g15), .A(n9625), .ZN(n9628) );
  AOI22_X1 U12063 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_g34), .ZN(n9626) );
  OAI221_X1 U12064 ( .B1(SI_30_), .B2(keyinput_g2), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_g34), .A(n9626), .ZN(n9627) );
  NOR4_X1 U12065 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(n9657)
         );
  XNOR2_X1 U12066 ( .A(n15087), .B(keyinput_g37), .ZN(n9637) );
  AOI22_X1 U12067 ( .A1(SI_15_), .A2(keyinput_g17), .B1(SI_28_), .B2(
        keyinput_g4), .ZN(n9631) );
  OAI221_X1 U12068 ( .B1(SI_15_), .B2(keyinput_g17), .C1(SI_28_), .C2(
        keyinput_g4), .A(n9631), .ZN(n9636) );
  AOI22_X1 U12069 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P3_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g43), .ZN(n9632) );
  OAI221_X1 U12070 ( .B1(SI_23_), .B2(keyinput_g9), .C1(P3_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n9632), .ZN(n9635) );
  AOI22_X1 U12071 ( .A1(SI_5_), .A2(keyinput_g27), .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n9633) );
  OAI221_X1 U12072 ( .B1(SI_5_), .B2(keyinput_g27), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n9633), .ZN(n9634) );
  NOR4_X1 U12073 ( .A1(n9637), .A2(n9636), .A3(n9635), .A4(n9634), .ZN(n9656)
         );
  AOI22_X1 U12074 ( .A1(SI_31_), .A2(keyinput_g1), .B1(SI_3_), .B2(
        keyinput_g29), .ZN(n9638) );
  OAI221_X1 U12075 ( .B1(SI_31_), .B2(keyinput_g1), .C1(SI_3_), .C2(
        keyinput_g29), .A(n9638), .ZN(n9645) );
  AOI22_X1 U12076 ( .A1(SI_12_), .A2(keyinput_g20), .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .ZN(n9639) );
  OAI221_X1 U12077 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n9639), .ZN(n9644) );
  AOI22_X1 U12078 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n9640) );
  OAI221_X1 U12079 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_27_), .C2(
        keyinput_g5), .A(n9640), .ZN(n9643) );
  AOI22_X1 U12080 ( .A1(SI_8_), .A2(keyinput_g24), .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n9641) );
  OAI221_X1 U12081 ( .B1(SI_8_), .B2(keyinput_g24), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9641), .ZN(n9642) );
  NOR4_X1 U12082 ( .A1(n9645), .A2(n9644), .A3(n9643), .A4(n9642), .ZN(n9655)
         );
  AOI22_X1 U12083 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n9646) );
  OAI221_X1 U12084 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n9646), .ZN(n9653) );
  AOI22_X1 U12085 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_19_), .B2(keyinput_g13), .ZN(n9647) );
  OAI221_X1 U12086 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        SI_19_), .C2(keyinput_g13), .A(n9647), .ZN(n9652) );
  AOI22_X1 U12087 ( .A1(SI_11_), .A2(keyinput_g21), .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n9648) );
  OAI221_X1 U12088 ( .B1(SI_11_), .B2(keyinput_g21), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n9648), .ZN(n9651) );
  AOI22_X1 U12089 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n9649) );
  OAI221_X1 U12090 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9649), .ZN(n9650) );
  NOR4_X1 U12091 ( .A1(n9653), .A2(n9652), .A3(n9651), .A4(n9650), .ZN(n9654)
         );
  NAND4_X1 U12092 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n9658)
         );
  OAI22_X1 U12093 ( .A1(keyinput_g53), .A2(n9662), .B1(n9659), .B2(n9658), 
        .ZN(n9660) );
  AOI211_X1 U12094 ( .C1(keyinput_g53), .C2(n9662), .A(n9661), .B(n9660), .ZN(
        n9663) );
  XNOR2_X1 U12095 ( .A(n9664), .B(n9663), .ZN(n9665) );
  NAND2_X1 U12096 ( .A1(n14695), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9666) );
  INV_X1 U12097 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9753) );
  INV_X1 U12098 ( .A(n6535), .ZN(n10783) );
  OR2_X1 U12099 ( .A1(n8879), .A2(n10783), .ZN(n9671) );
  NAND2_X1 U12100 ( .A1(n10775), .A2(n15116), .ZN(n9670) );
  NAND2_X1 U12101 ( .A1(n9671), .A2(n9670), .ZN(n15109) );
  OR2_X1 U12102 ( .A1(n9672), .A2(n15106), .ZN(n12148) );
  NAND2_X1 U12103 ( .A1(n9672), .A2(n15106), .ZN(n12147) );
  INV_X1 U12104 ( .A(n15106), .ZN(n9673) );
  NOR2_X1 U12105 ( .A1(n9672), .A2(n9673), .ZN(n9674) );
  OR2_X1 U12106 ( .A1(n9675), .A2(n15140), .ZN(n12152) );
  NAND2_X1 U12107 ( .A1(n9675), .A2(n15140), .ZN(n12151) );
  NAND2_X1 U12108 ( .A1(n10951), .A2(n12115), .ZN(n10955) );
  INV_X1 U12109 ( .A(n15140), .ZN(n12412) );
  NAND2_X1 U12110 ( .A1(n12606), .A2(n12412), .ZN(n9676) );
  NAND2_X1 U12111 ( .A1(n10955), .A2(n9676), .ZN(n11165) );
  NAND2_X1 U12112 ( .A1(n12605), .A2(n15147), .ZN(n12158) );
  NAND2_X1 U12113 ( .A1(n11165), .A2(n12117), .ZN(n11164) );
  INV_X1 U12114 ( .A(n15147), .ZN(n9677) );
  NAND2_X1 U12115 ( .A1(n12605), .A2(n9677), .ZN(n9678) );
  NAND2_X1 U12116 ( .A1(n11164), .A2(n9678), .ZN(n11255) );
  NAND2_X1 U12117 ( .A1(n12604), .A2(n15154), .ZN(n12166) );
  INV_X1 U12118 ( .A(n15158), .ZN(n9679) );
  AND2_X1 U12119 ( .A1(n12603), .A2(n9679), .ZN(n9680) );
  OR2_X1 U12120 ( .A1(n12604), .A2(n7435), .ZN(n11306) );
  INV_X1 U12121 ( .A(n14962), .ZN(n15168) );
  NAND2_X1 U12122 ( .A1(n12602), .A2(n15168), .ZN(n11361) );
  INV_X1 U12123 ( .A(n15170), .ZN(n9682) );
  NAND2_X1 U12124 ( .A1(n12601), .A2(n9682), .ZN(n9681) );
  AND2_X1 U12125 ( .A1(n11361), .A2(n9681), .ZN(n9683) );
  XNOR2_X1 U12126 ( .A(n12600), .B(n15179), .ZN(n12187) );
  NAND2_X1 U12127 ( .A1(n11425), .A2(n12187), .ZN(n9685) );
  INV_X1 U12128 ( .A(n15179), .ZN(n11445) );
  NAND2_X1 U12129 ( .A1(n12600), .A2(n11445), .ZN(n9684) );
  NAND2_X1 U12130 ( .A1(n9685), .A2(n9684), .ZN(n11452) );
  OR2_X1 U12131 ( .A1(n12599), .A2(n15186), .ZN(n12194) );
  NAND2_X1 U12132 ( .A1(n12599), .A2(n15186), .ZN(n12195) );
  INV_X1 U12133 ( .A(n15186), .ZN(n9686) );
  NAND2_X1 U12134 ( .A1(n12599), .A2(n9686), .ZN(n9687) );
  INV_X1 U12135 ( .A(n12997), .ZN(n9688) );
  OR2_X1 U12136 ( .A1(n12598), .A2(n9688), .ZN(n9689) );
  NAND2_X1 U12137 ( .A1(n9690), .A2(n9689), .ZN(n12820) );
  NAND2_X1 U12138 ( .A1(n12597), .A2(n12993), .ZN(n12204) );
  NAND2_X1 U12139 ( .A1(n12205), .A2(n12204), .ZN(n12113) );
  NOR2_X1 U12140 ( .A1(n12820), .A2(n12824), .ZN(n9691) );
  INV_X1 U12141 ( .A(n9691), .ZN(n12819) );
  INV_X1 U12142 ( .A(n12993), .ZN(n9692) );
  NAND2_X1 U12143 ( .A1(n12597), .A2(n9692), .ZN(n12803) );
  OR2_X1 U12144 ( .A1(n12596), .A2(n14450), .ZN(n12209) );
  NAND2_X1 U12145 ( .A1(n12209), .A2(n12210), .ZN(n12122) );
  AOI21_X2 U12146 ( .B1(n12819), .B2(n12803), .A(n12815), .ZN(n12807) );
  NOR2_X1 U12147 ( .A1(n12457), .A2(n14450), .ZN(n12789) );
  NAND2_X1 U12148 ( .A1(n12595), .A2(n12389), .ZN(n12213) );
  NAND2_X1 U12149 ( .A1(n12214), .A2(n12213), .ZN(n12788) );
  OAI21_X1 U12150 ( .B1(n12807), .B2(n12789), .A(n12788), .ZN(n12792) );
  INV_X1 U12151 ( .A(n12896), .ZN(n9695) );
  NAND2_X1 U12152 ( .A1(n9695), .A2(n12477), .ZN(n9696) );
  AOI22_X1 U12153 ( .A1(n12779), .A2(n9696), .B1(n12594), .B2(n12896), .ZN(
        n12767) );
  OR2_X1 U12154 ( .A1(n12974), .A2(n12486), .ZN(n12224) );
  NAND2_X1 U12155 ( .A1(n12974), .A2(n12486), .ZN(n12220) );
  INV_X1 U12156 ( .A(n12974), .ZN(n9697) );
  OAI22_X2 U12157 ( .A1(n12767), .A2(n12768), .B1(n12486), .B2(n9697), .ZN(
        n12759) );
  NOR2_X1 U12158 ( .A1(n12968), .A2(n12549), .ZN(n12229) );
  INV_X1 U12159 ( .A(n12229), .ZN(n9698) );
  NAND2_X1 U12160 ( .A1(n12968), .A2(n12549), .ZN(n12230) );
  NAND2_X1 U12161 ( .A1(n9698), .A2(n12230), .ZN(n12231) );
  NAND2_X1 U12162 ( .A1(n12962), .A2(n12487), .ZN(n12237) );
  NAND2_X1 U12163 ( .A1(n12956), .A2(n12590), .ZN(n12719) );
  NAND2_X1 U12164 ( .A1(n12956), .A2(n12551), .ZN(n12236) );
  NAND2_X1 U12165 ( .A1(n12239), .A2(n12236), .ZN(n12732) );
  OR2_X1 U12166 ( .A1(n12962), .A2(n12591), .ZN(n12733) );
  NAND2_X1 U12167 ( .A1(n12732), .A2(n12733), .ZN(n12717) );
  AOI21_X1 U12168 ( .B1(n12719), .B2(n12717), .A(n12720), .ZN(n9699) );
  NAND2_X1 U12169 ( .A1(n12877), .A2(n12588), .ZN(n12108) );
  OR2_X1 U12170 ( .A1(n12877), .A2(n12588), .ZN(n12109) );
  INV_X1 U12171 ( .A(n12873), .ZN(n12536) );
  INV_X1 U12172 ( .A(n12524), .ZN(n9700) );
  NAND2_X1 U12173 ( .A1(n12873), .A2(n9700), .ZN(n9701) );
  NAND2_X1 U12174 ( .A1(n12691), .A2(n12526), .ZN(n9703) );
  NAND2_X1 U12175 ( .A1(n12662), .A2(n9703), .ZN(n12256) );
  NAND2_X1 U12176 ( .A1(n12676), .A2(n12403), .ZN(n12257) );
  INV_X1 U12177 ( .A(n9705), .ZN(n11756) );
  INV_X1 U12178 ( .A(n12559), .ZN(n9706) );
  NAND2_X1 U12179 ( .A1(n12855), .A2(n12427), .ZN(n12277) );
  OR2_X1 U12180 ( .A1(n12855), .A2(n12427), .ZN(n9709) );
  INV_X1 U12181 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11656) );
  AND2_X1 U12182 ( .A1(n11656), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9710) );
  INV_X1 U12183 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14360) );
  NAND2_X1 U12184 ( .A1(n14360), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9712) );
  XNOR2_X1 U12185 ( .A(n9720), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9713) );
  XNOR2_X1 U12186 ( .A(n9719), .B(n9713), .ZN(n12319) );
  NAND2_X1 U12187 ( .A1(n12319), .A2(n12098), .ZN(n9716) );
  NAND2_X1 U12188 ( .A1(n12921), .A2(n9738), .ZN(n12278) );
  INV_X1 U12189 ( .A(n12921), .ZN(n9717) );
  AND2_X1 U12190 ( .A1(n12037), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U12191 ( .A1(n9720), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9721) );
  XNOR2_X1 U12192 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12079) );
  XNOR2_X1 U12193 ( .A(n12081), .B(n12079), .ZN(n12385) );
  NOR2_X1 U12194 ( .A1(n9714), .A2(n12388), .ZN(n9722) );
  AOI21_X1 U12195 ( .B1(n12385), .B2(n12098), .A(n9722), .ZN(n9727) );
  NAND2_X1 U12196 ( .A1(n12083), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9726) );
  OR2_X1 U12197 ( .A1(n12085), .A2(n9753), .ZN(n9725) );
  INV_X1 U12198 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9796) );
  OR2_X1 U12199 ( .A1(n12086), .A2(n9796), .ZN(n9724) );
  NAND4_X1 U12200 ( .A1(n12090), .A2(n9726), .A3(n9725), .A4(n9724), .ZN(
        n12581) );
  AND2_X1 U12201 ( .A1(n9727), .A2(n12581), .ZN(n12076) );
  INV_X1 U12202 ( .A(n9727), .ZN(n9815) );
  INV_X1 U12203 ( .A(n12581), .ZN(n9728) );
  XNOR2_X1 U12204 ( .A(n9729), .B(n12281), .ZN(n9740) );
  NAND2_X1 U12205 ( .A1(n12614), .A2(n12297), .ZN(n9730) );
  NAND2_X1 U12206 ( .A1(n9797), .A2(n9746), .ZN(n12134) );
  NAND2_X1 U12207 ( .A1(n9731), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U12208 ( .A1(n12083), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U12209 ( .A1(n9732), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9733) );
  NOR2_X1 U12210 ( .A1(n9336), .A2(n9736), .ZN(n9737) );
  OR2_X1 U12211 ( .A1(n12550), .A2(n9737), .ZN(n12631) );
  OAI22_X1 U12212 ( .A1(n12102), .A2(n12631), .B1(n9738), .B2(n12548), .ZN(
        n9739) );
  AOI21_X1 U12213 ( .B1(n9740), .B2(n12804), .A(n9739), .ZN(n9804) );
  XNOR2_X1 U12214 ( .A(n13001), .B(n12999), .ZN(n9743) );
  NAND2_X1 U12215 ( .A1(n9741), .A2(n12293), .ZN(n9742) );
  OAI22_X1 U12216 ( .A1(n15185), .A2(n9746), .B1(n12614), .B2(n12137), .ZN(
        n9744) );
  AOI21_X1 U12217 ( .B1(n9745), .B2(n9744), .A(n12286), .ZN(n9750) );
  NAND2_X1 U12218 ( .A1(n12297), .A2(n9746), .ZN(n9747) );
  NOR2_X1 U12219 ( .A1(n12614), .A2(n9747), .ZN(n9790) );
  MUX2_X1 U12220 ( .A(n9790), .B(n12292), .S(n12286), .Z(n9792) );
  INV_X1 U12221 ( .A(n9792), .ZN(n9748) );
  NAND2_X1 U12222 ( .A1(n12999), .A2(n9748), .ZN(n9749) );
  OAI21_X1 U12223 ( .B1(n12999), .B2(n9750), .A(n9749), .ZN(n9751) );
  INV_X1 U12224 ( .A(n9751), .ZN(n9752) );
  MUX2_X1 U12225 ( .A(n9753), .B(n9804), .S(n15205), .Z(n9789) );
  NAND2_X1 U12226 ( .A1(n9755), .A2(n9754), .ZN(n15105) );
  NAND2_X1 U12227 ( .A1(n15104), .A2(n15105), .ZN(n9756) );
  NAND2_X1 U12228 ( .A1(n9756), .A2(n12148), .ZN(n10950) );
  INV_X1 U12229 ( .A(n12115), .ZN(n10948) );
  NAND2_X1 U12230 ( .A1(n10949), .A2(n12152), .ZN(n11162) );
  INV_X1 U12231 ( .A(n12117), .ZN(n12154) );
  NAND2_X1 U12232 ( .A1(n11162), .A2(n12154), .ZN(n9757) );
  NAND2_X1 U12233 ( .A1(n9757), .A2(n12157), .ZN(n11254) );
  NAND2_X1 U12234 ( .A1(n11254), .A2(n12160), .ZN(n9758) );
  NAND2_X1 U12235 ( .A1(n9758), .A2(n12162), .ZN(n11303) );
  INV_X1 U12236 ( .A(n12114), .ZN(n11305) );
  NAND2_X1 U12237 ( .A1(n11304), .A2(n12163), .ZN(n11283) );
  INV_X1 U12238 ( .A(n12172), .ZN(n9759) );
  NAND2_X1 U12239 ( .A1(n11283), .A2(n9759), .ZN(n9760) );
  NAND2_X1 U12240 ( .A1(n9760), .A2(n12176), .ZN(n11360) );
  NAND2_X1 U12241 ( .A1(n12601), .A2(n15170), .ZN(n12183) );
  NAND2_X1 U12242 ( .A1(n12184), .A2(n12183), .ZN(n12180) );
  INV_X1 U12243 ( .A(n12180), .ZN(n9761) );
  NAND2_X1 U12244 ( .A1(n11360), .A2(n9761), .ZN(n9762) );
  OR2_X1 U12245 ( .A1(n12600), .A2(n15179), .ZN(n12191) );
  INV_X1 U12246 ( .A(n12191), .ZN(n9763) );
  NAND2_X1 U12247 ( .A1(n12600), .A2(n15179), .ZN(n12190) );
  INV_X1 U12248 ( .A(n12192), .ZN(n9765) );
  AOI21_X2 U12249 ( .B1(n11459), .B2(n9765), .A(n9764), .ZN(n12838) );
  OR2_X1 U12250 ( .A1(n12598), .A2(n12997), .ZN(n12201) );
  NAND2_X1 U12251 ( .A1(n12598), .A2(n12997), .ZN(n12200) );
  NAND2_X1 U12252 ( .A1(n12201), .A2(n12200), .ZN(n12833) );
  NAND2_X1 U12253 ( .A1(n12837), .A2(n12201), .ZN(n12825) );
  INV_X1 U12254 ( .A(n12816), .ZN(n9768) );
  INV_X1 U12255 ( .A(n12210), .ZN(n9767) );
  NAND2_X1 U12256 ( .A1(n12786), .A2(n12214), .ZN(n12777) );
  OR2_X1 U12257 ( .A1(n12896), .A2(n12477), .ZN(n12217) );
  NAND2_X1 U12258 ( .A1(n12896), .A2(n12477), .ZN(n12221) );
  NAND2_X1 U12259 ( .A1(n12217), .A2(n12221), .ZN(n12778) );
  INV_X1 U12260 ( .A(n12778), .ZN(n9770) );
  NAND2_X1 U12261 ( .A1(n12777), .A2(n9770), .ZN(n9771) );
  NAND2_X1 U12262 ( .A1(n9771), .A2(n12221), .ZN(n12766) );
  NAND2_X1 U12263 ( .A1(n12766), .A2(n12768), .ZN(n9772) );
  NAND2_X1 U12264 ( .A1(n9772), .A2(n12220), .ZN(n12757) );
  NAND2_X1 U12265 ( .A1(n12757), .A2(n12758), .ZN(n9773) );
  NAND2_X1 U12266 ( .A1(n9773), .A2(n12230), .ZN(n12743) );
  NAND2_X1 U12267 ( .A1(n12239), .A2(n12729), .ZN(n12228) );
  INV_X1 U12268 ( .A(n12228), .ZN(n9774) );
  NOR2_X1 U12269 ( .A1(n12950), .A2(n12443), .ZN(n12246) );
  INV_X1 U12270 ( .A(n12246), .ZN(n9775) );
  NAND2_X1 U12271 ( .A1(n12877), .A2(n12507), .ZN(n9776) );
  INV_X1 U12272 ( .A(n12662), .ZN(n9777) );
  INV_X1 U12273 ( .A(n12259), .ZN(n9780) );
  NOR2_X1 U12274 ( .A1(n11775), .A2(n11779), .ZN(n9778) );
  AND2_X1 U12275 ( .A1(n9778), .A2(n11773), .ZN(n9779) );
  NAND2_X1 U12276 ( .A1(n11774), .A2(n9779), .ZN(n9782) );
  NAND2_X1 U12277 ( .A1(n12873), .A2(n12524), .ZN(n12680) );
  NAND2_X1 U12278 ( .A1(n9782), .A2(n9781), .ZN(n11772) );
  NAND2_X1 U12279 ( .A1(n12559), .A2(n12269), .ZN(n11753) );
  INV_X1 U12280 ( .A(n9784), .ZN(n12279) );
  INV_X1 U12281 ( .A(n12281), .ZN(n12129) );
  XNOR2_X1 U12282 ( .A(n12101), .B(n12129), .ZN(n9814) );
  INV_X1 U12283 ( .A(n9790), .ZN(n9786) );
  NAND3_X1 U12284 ( .A1(n9809), .A2(n12292), .A3(n15185), .ZN(n9785) );
  NAND2_X1 U12285 ( .A1(n15205), .A2(n15190), .ZN(n12899) );
  OR2_X1 U12286 ( .A1(n9814), .A2(n12899), .ZN(n9788) );
  NAND2_X1 U12287 ( .A1(n9815), .A2(n12901), .ZN(n9787) );
  NAND2_X1 U12288 ( .A1(n9789), .A2(n7458), .ZN(P3_U3488) );
  OAI21_X1 U12289 ( .B1(n12286), .B2(n9790), .A(n12999), .ZN(n9791) );
  OAI21_X1 U12290 ( .B1(n12999), .B2(n9792), .A(n9791), .ZN(n9793) );
  INV_X1 U12291 ( .A(n9793), .ZN(n9794) );
  NAND2_X1 U12292 ( .A1(n9795), .A2(n9794), .ZN(n9799) );
  MUX2_X1 U12293 ( .A(n9796), .B(n9804), .S(n15126), .Z(n9803) );
  NAND2_X1 U12294 ( .A1(n15122), .A2(n9797), .ZN(n15119) );
  OR2_X1 U12295 ( .A1(n15128), .A2(n15164), .ZN(n9798) );
  NOR2_X1 U12296 ( .A1(n15121), .A2(n9800), .ZN(n12634) );
  AOI21_X1 U12297 ( .B1(n9815), .B2(n12798), .A(n12634), .ZN(n9801) );
  NAND2_X1 U12298 ( .A1(n9803), .A2(n7457), .ZN(P3_U3204) );
  INV_X1 U12299 ( .A(n9805), .ZN(n9806) );
  OR2_X1 U12300 ( .A1(n10678), .A2(n9806), .ZN(n9807) );
  NAND2_X1 U12301 ( .A1(n9808), .A2(n9807), .ZN(n9813) );
  INV_X1 U12302 ( .A(n9809), .ZN(n9810) );
  OR2_X1 U12303 ( .A1(n9811), .A2(n9810), .ZN(n9812) );
  NAND2_X1 U12304 ( .A1(n9815), .A2(n12985), .ZN(n9818) );
  INV_X1 U12305 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9816) );
  OR2_X1 U12306 ( .A1(n15193), .A2(n9816), .ZN(n9817) );
  AND2_X1 U12307 ( .A1(n9818), .A2(n9817), .ZN(n9819) );
  OAI21_X1 U12308 ( .B1(n9804), .B2(n15191), .A(n7456), .ZN(P3_U3456) );
  INV_X1 U12309 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U12310 ( .A1(n14698), .A2(n9822), .ZN(n9823) );
  INV_X1 U12311 ( .A(n14418), .ZN(n10089) );
  NAND2_X1 U12312 ( .A1(n15091), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U12313 ( .A1(n9828), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9829) );
  OAI21_X1 U12314 ( .B1(n9830), .B2(n9829), .A(n9831), .ZN(n11104) );
  OR2_X1 U12315 ( .A1(n11104), .A2(n8852), .ZN(n11106) );
  NAND2_X1 U12316 ( .A1(n11106), .A2(n9831), .ZN(n11016) );
  NAND2_X1 U12317 ( .A1(n6656), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9832) );
  NAND2_X1 U12318 ( .A1(n11015), .A2(n9832), .ZN(n9834) );
  AOI22_X1 U12319 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n11084), .B1(n9862), .B2(
        n8912), .ZN(n11074) );
  XNOR2_X1 U12320 ( .A(n9836), .B(n11057), .ZN(n11048) );
  AOI22_X1 U12321 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n11100), .B1(n9955), .B2(
        n8959), .ZN(n11090) );
  NOR2_X1 U12322 ( .A1(n9977), .A2(n9839), .ZN(n9840) );
  AOI22_X1 U12323 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n9900), .B1(n10921), .B2(
        n8997), .ZN(n10911) );
  NOR2_X1 U12324 ( .A1(n15003), .A2(n9841), .ZN(n9842) );
  NOR2_X1 U12325 ( .A1(n9842), .A2(n14998), .ZN(n15015) );
  AOI22_X1 U12326 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n9986), .B1(n15021), 
        .B2(n9034), .ZN(n15014) );
  NOR2_X1 U12327 ( .A1(n9908), .A2(n9843), .ZN(n9844) );
  NOR2_X1 U12328 ( .A1(n9844), .A2(n15030), .ZN(n15048) );
  AOI22_X1 U12329 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n9911), .B1(n15054), 
        .B2(n12826), .ZN(n15047) );
  NOR2_X1 U12330 ( .A1(n15048), .A2(n15047), .ZN(n15046) );
  NOR2_X1 U12331 ( .A1(n9914), .A2(n9845), .ZN(n9846) );
  OR2_X1 U12332 ( .A1(n15091), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9847) );
  NAND2_X1 U12333 ( .A1(n9917), .A2(n9847), .ZN(n15082) );
  INV_X1 U12334 ( .A(n15081), .ZN(n9848) );
  AND2_X1 U12335 ( .A1(n14408), .A2(n9849), .ZN(n9850) );
  AOI22_X1 U12336 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14418), .B1(n10089), 
        .B2(n12771), .ZN(n14427) );
  INV_X1 U12337 ( .A(n12617), .ZN(n12611) );
  NAND2_X1 U12338 ( .A1(n12611), .A2(n12751), .ZN(n9853) );
  NAND2_X1 U12339 ( .A1(n12617), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9852) );
  AND2_X1 U12340 ( .A1(n9853), .A2(n9852), .ZN(n9858) );
  NAND2_X1 U12341 ( .A1(n9856), .A2(n12286), .ZN(n9854) );
  NAND2_X1 U12342 ( .A1(n6508), .A2(n9854), .ZN(n9933) );
  NOR2_X1 U12343 ( .A1(n9856), .A2(P3_U3151), .ZN(n12290) );
  NOR2_X1 U12344 ( .A1(n12293), .A2(n12290), .ZN(n9932) );
  OR2_X1 U12345 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  INV_X1 U12346 ( .A(n15102), .ZN(n14441) );
  AOI22_X1 U12347 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n10089), .B1(n14418), 
        .B2(n12892), .ZN(n14424) );
  NAND2_X1 U12348 ( .A1(n15091), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9916) );
  OAI21_X1 U12349 ( .B1(n15091), .B2(P3_REG1_REG_14__SCAN_IN), .A(n9916), .ZN(
        n9860) );
  INV_X1 U12350 ( .A(n9860), .ZN(n15086) );
  MUX2_X1 U12351 ( .A(n9861), .B(P3_REG1_REG_12__SCAN_IN), .S(n9911), .Z(
        n15050) );
  AOI22_X1 U12352 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n15021), .B1(n9986), 
        .B2(n9030), .ZN(n15018) );
  AOI22_X1 U12353 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10921), .B1(n9900), .B2(
        n8996), .ZN(n10919) );
  AOI22_X1 U12354 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n9955), .B1(n11100), .B2(
        n8962), .ZN(n11093) );
  AOI22_X1 U12355 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n9862), .B1(n11084), .B2(
        n8915), .ZN(n11078) );
  MUX2_X1 U12356 ( .A(n9863), .B(P3_REG1_REG_2__SCAN_IN), .S(n6500), .Z(n11021) );
  AND2_X1 U12357 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n6992), .ZN(n9864) );
  OR3_X1 U12358 ( .A1(n8867), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n9865) );
  OAI21_X1 U12359 ( .B1(n9830), .B2(n9864), .A(n9865), .ZN(n11108) );
  OR2_X1 U12360 ( .A1(n11108), .A2(n11107), .ZN(n11110) );
  NAND2_X1 U12361 ( .A1(n11110), .A2(n9865), .ZN(n11020) );
  NAND2_X1 U12362 ( .A1(n11021), .A2(n11020), .ZN(n11019) );
  NAND2_X1 U12363 ( .A1(n6656), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12364 ( .A1(n11019), .A2(n9866), .ZN(n9867) );
  NAND2_X1 U12365 ( .A1(n9867), .A2(n9891), .ZN(n9868) );
  XNOR2_X1 U12366 ( .A(n9867), .B(n11132), .ZN(n11126) );
  NAND2_X1 U12367 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n11126), .ZN(n11125) );
  NAND2_X1 U12368 ( .A1(n9868), .A2(n11125), .ZN(n11077) );
  NAND2_X1 U12369 ( .A1(n11078), .A2(n11077), .ZN(n11076) );
  NAND2_X1 U12370 ( .A1(n9895), .A2(n9869), .ZN(n9870) );
  NAND2_X1 U12371 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n11050), .ZN(n11049) );
  NAND2_X1 U12372 ( .A1(n9870), .A2(n11049), .ZN(n11092) );
  NAND2_X1 U12373 ( .A1(n11093), .A2(n11092), .ZN(n11091) );
  OAI21_X1 U12374 ( .B1(n11100), .B2(n8962), .A(n11091), .ZN(n9871) );
  NAND2_X1 U12375 ( .A1(n11040), .A2(n9871), .ZN(n9872) );
  NAND2_X1 U12376 ( .A1(n9872), .A2(n11035), .ZN(n10918) );
  NAND2_X1 U12377 ( .A1(n10919), .A2(n10918), .ZN(n10917) );
  NAND2_X1 U12378 ( .A1(n9950), .A2(n9873), .ZN(n9874) );
  XNOR2_X1 U12379 ( .A(n15003), .B(n9873), .ZN(n15001) );
  NAND2_X1 U12380 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15001), .ZN(n15000) );
  NAND2_X1 U12381 ( .A1(n9874), .A2(n15000), .ZN(n15017) );
  NAND2_X1 U12382 ( .A1(n15018), .A2(n15017), .ZN(n15016) );
  NAND2_X1 U12383 ( .A1(n15036), .A2(n9875), .ZN(n9876) );
  XNOR2_X1 U12384 ( .A(n9875), .B(n9908), .ZN(n15033) );
  NAND2_X1 U12385 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15033), .ZN(n15032) );
  NAND2_X1 U12386 ( .A1(n9876), .A2(n15032), .ZN(n15051) );
  NAND2_X1 U12387 ( .A1(n15050), .A2(n15051), .ZN(n15049) );
  NAND2_X1 U12388 ( .A1(n15070), .A2(n9877), .ZN(n9878) );
  XNOR2_X1 U12389 ( .A(n9914), .B(n9877), .ZN(n15066) );
  NAND2_X1 U12390 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n15066), .ZN(n15065) );
  NAND2_X1 U12391 ( .A1(n9878), .A2(n15065), .ZN(n15085) );
  NAND2_X1 U12392 ( .A1(n15086), .A2(n15085), .ZN(n15084) );
  NAND2_X1 U12393 ( .A1(n14408), .A2(n9879), .ZN(n9880) );
  NAND2_X1 U12394 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14404), .ZN(n14403) );
  NAND2_X1 U12395 ( .A1(n9880), .A2(n14403), .ZN(n14423) );
  NAND2_X1 U12396 ( .A1(n10093), .A2(n9881), .ZN(n9882) );
  XNOR2_X1 U12397 ( .A(n14433), .B(n9881), .ZN(n14435) );
  NAND2_X1 U12398 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14435), .ZN(n14434) );
  NAND2_X1 U12399 ( .A1(n9882), .A2(n14434), .ZN(n12613) );
  XNOR2_X1 U12400 ( .A(n12617), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12612) );
  XNOR2_X1 U12401 ( .A(n12613), .B(n12612), .ZN(n9930) );
  NOR2_X2 U12402 ( .A1(n9931), .A2(n9883), .ZN(n15094) );
  MUX2_X1 U12403 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n9922), .Z(n9927) );
  MUX2_X1 U12404 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n9922), .Z(n9925) );
  MUX2_X1 U12405 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n9922), .Z(n9884) );
  MUX2_X1 U12406 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n9922), .Z(n9912) );
  INV_X1 U12407 ( .A(n9912), .ZN(n9913) );
  MUX2_X1 U12408 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n9922), .Z(n9909) );
  INV_X1 U12409 ( .A(n9909), .ZN(n9910) );
  MUX2_X1 U12410 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n9922), .Z(n9906) );
  INV_X1 U12411 ( .A(n9906), .ZN(n9907) );
  MUX2_X1 U12412 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n9922), .Z(n9904) );
  INV_X1 U12413 ( .A(n9904), .ZN(n9905) );
  MUX2_X1 U12414 ( .A(n9016), .B(n9019), .S(n9922), .Z(n9903) );
  OR2_X1 U12415 ( .A1(n9903), .A2(n15003), .ZN(n14994) );
  MUX2_X1 U12416 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n9922), .Z(n9901) );
  OR2_X1 U12417 ( .A1(n9901), .A2(n10921), .ZN(n9902) );
  MUX2_X1 U12418 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n9885), .Z(n9886) );
  XNOR2_X1 U12419 ( .A(n9886), .B(n9830), .ZN(n11103) );
  MUX2_X1 U12420 ( .A(n9828), .B(n8867), .S(n9885), .Z(n14988) );
  NAND2_X1 U12421 ( .A1(n14988), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14987) );
  OAI22_X1 U12422 ( .A1(n11103), .A2(n14987), .B1(n9886), .B2(n9830), .ZN(
        n11013) );
  MUX2_X1 U12423 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n9922), .Z(n9887) );
  XNOR2_X1 U12424 ( .A(n9887), .B(n6500), .ZN(n11014) );
  INV_X1 U12425 ( .A(n9887), .ZN(n9888) );
  AOI22_X1 U12426 ( .A1(n11013), .A2(n11014), .B1(n6500), .B2(n9888), .ZN(
        n11122) );
  MUX2_X1 U12427 ( .A(n10957), .B(n9889), .S(n9922), .Z(n9890) );
  XNOR2_X1 U12428 ( .A(n9890), .B(n11132), .ZN(n11121) );
  INV_X1 U12429 ( .A(n9890), .ZN(n9892) );
  OAI22_X1 U12430 ( .A1(n11122), .A2(n11121), .B1(n9892), .B2(n9891), .ZN(
        n11072) );
  MUX2_X1 U12431 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n9922), .Z(n9893) );
  XNOR2_X1 U12432 ( .A(n9893), .B(n11084), .ZN(n11071) );
  INV_X1 U12433 ( .A(n9893), .ZN(n9894) );
  AOI22_X1 U12434 ( .A1(n11072), .A2(n11071), .B1(n11084), .B2(n9894), .ZN(
        n11045) );
  MUX2_X1 U12435 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n9922), .Z(n9896) );
  XNOR2_X1 U12436 ( .A(n9896), .B(n9895), .ZN(n11046) );
  OAI22_X1 U12437 ( .A1(n11045), .A2(n11046), .B1(n9896), .B2(n9895), .ZN(
        n11087) );
  MUX2_X1 U12438 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n9922), .Z(n9897) );
  XNOR2_X1 U12439 ( .A(n9897), .B(n11100), .ZN(n11088) );
  INV_X1 U12440 ( .A(n9897), .ZN(n9898) );
  MUX2_X1 U12441 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n9922), .Z(n9899) );
  XNOR2_X1 U12442 ( .A(n9899), .B(n11040), .ZN(n11030) );
  OAI22_X1 U12443 ( .A1(n11031), .A2(n11030), .B1(n9899), .B2(n11040), .ZN(
        n10915) );
  XNOR2_X1 U12444 ( .A(n9901), .B(n9900), .ZN(n10914) );
  NAND2_X1 U12445 ( .A1(n10915), .A2(n10914), .ZN(n10913) );
  XNOR2_X1 U12446 ( .A(n9904), .B(n15021), .ZN(n15022) );
  XNOR2_X1 U12447 ( .A(n9906), .B(n15036), .ZN(n15040) );
  NOR2_X1 U12448 ( .A1(n15041), .A2(n15040), .ZN(n15039) );
  XNOR2_X1 U12449 ( .A(n9909), .B(n9911), .ZN(n15058) );
  XNOR2_X1 U12450 ( .A(n9912), .B(n15070), .ZN(n15075) );
  INV_X1 U12451 ( .A(n15082), .ZN(n9915) );
  MUX2_X1 U12452 ( .A(n9915), .B(n15086), .S(n9922), .Z(n15098) );
  NAND2_X1 U12453 ( .A1(n15099), .A2(n15098), .ZN(n15097) );
  MUX2_X1 U12454 ( .A(n9917), .B(n9916), .S(n9922), .Z(n9918) );
  NAND2_X1 U12455 ( .A1(n15097), .A2(n9918), .ZN(n9919) );
  MUX2_X1 U12456 ( .A(n14402), .B(n12897), .S(n9922), .Z(n14411) );
  AND2_X1 U12457 ( .A1(n14412), .A2(n14411), .ZN(n14414) );
  MUX2_X1 U12458 ( .A(n12771), .B(n12892), .S(n9922), .Z(n9924) );
  NAND2_X1 U12459 ( .A1(n9924), .A2(n14418), .ZN(n14419) );
  XNOR2_X1 U12460 ( .A(n9925), .B(n10093), .ZN(n14437) );
  XNOR2_X1 U12461 ( .A(n12618), .B(n12617), .ZN(n9926) );
  NOR2_X1 U12462 ( .A1(n9926), .A2(n9927), .ZN(n12616) );
  AOI21_X1 U12463 ( .B1(n9927), .B2(n9926), .A(n12616), .ZN(n9928) );
  NAND2_X1 U12464 ( .A1(P3_U3897), .A2(n9336), .ZN(n15076) );
  NOR2_X1 U12465 ( .A1(n9928), .A2(n15076), .ZN(n9929) );
  AOI21_X1 U12466 ( .B1(n9930), .B2(n15094), .A(n9929), .ZN(n9937) );
  NAND2_X1 U12467 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n9936) );
  MUX2_X1 U12468 ( .A(n9931), .B(n12607), .S(n12294), .Z(n15092) );
  INV_X1 U12469 ( .A(n9932), .ZN(n9934) );
  AOI22_X1 U12470 ( .A1(n15002), .A2(n12617), .B1(n15089), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n9935) );
  NAND4_X1 U12471 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(
        P3_U3200) );
  INV_X1 U12472 ( .A(n10290), .ZN(n9940) );
  NOR2_X2 U12473 ( .A1(n10274), .A2(n9940), .ZN(P1_U4016) );
  NOR2_X1 U12474 ( .A1(n6492), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13683) );
  AOI22_X1 U12475 ( .A1(n13683), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n13162), .ZN(n9941) );
  OAI21_X1 U12476 ( .B1(n9963), .B2(n13685), .A(n9941), .ZN(P2_U3326) );
  INV_X2 U12477 ( .A(n13683), .ZN(n13688) );
  INV_X1 U12478 ( .A(n10074), .ZN(n10084) );
  OAI222_X1 U12479 ( .A1(n13688), .A2(n9942), .B1(n13685), .B2(n9970), .C1(
        P2_U3088), .C2(n10084), .ZN(P2_U3325) );
  INV_X1 U12480 ( .A(n9943), .ZN(n10000) );
  INV_X1 U12481 ( .A(n14699), .ZN(n10011) );
  OAI222_X1 U12482 ( .A1(n13688), .A2(n9944), .B1(n13685), .B2(n10000), .C1(
        P2_U3088), .C2(n10011), .ZN(P2_U3324) );
  INV_X1 U12483 ( .A(n9945), .ZN(n9997) );
  INV_X1 U12484 ( .A(n14711), .ZN(n10013) );
  OAI222_X1 U12485 ( .A1(n13688), .A2(n9946), .B1(n13685), .B2(n9997), .C1(
        P2_U3088), .C2(n10013), .ZN(P2_U3323) );
  OAI222_X1 U12486 ( .A1(P3_U3151), .A2(n9830), .B1(n13004), .B2(n9948), .C1(
        n12387), .C2(n9947), .ZN(P3_U3294) );
  INV_X1 U12487 ( .A(n9949), .ZN(n9952) );
  OAI222_X1 U12488 ( .A1(n12387), .A2(n9952), .B1(n13004), .B2(n9951), .C1(
        n9950), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12489 ( .A1(n9955), .A2(P3_U3151), .B1(n12387), .B2(n9954), .C1(
        n9953), .C2(n13004), .ZN(P3_U3289) );
  OAI222_X1 U12490 ( .A1(n10921), .A2(P3_U3151), .B1(n12387), .B2(n9957), .C1(
        n9956), .C2(n13004), .ZN(P3_U3287) );
  OAI222_X1 U12491 ( .A1(n6992), .A2(P3_U3151), .B1(n12387), .B2(n9959), .C1(
        n9958), .C2(n13004), .ZN(P3_U3295) );
  INV_X1 U12492 ( .A(n13888), .ZN(n9964) );
  NAND2_X2 U12493 ( .A1(n9960), .A2(P1_U3086), .ZN(n14366) );
  OAI222_X1 U12494 ( .A1(P1_U3086), .A2(n9964), .B1(n14366), .B2(n9963), .C1(
        n9962), .C2(n14363), .ZN(P1_U3354) );
  INV_X1 U12495 ( .A(n9965), .ZN(n9995) );
  INV_X1 U12496 ( .A(n14723), .ZN(n10015) );
  OAI222_X1 U12497 ( .A1(n13688), .A2(n9966), .B1(n13685), .B2(n9995), .C1(
        P2_U3088), .C2(n10015), .ZN(P2_U3322) );
  OAI222_X1 U12498 ( .A1(n12387), .A2(n9968), .B1(n13004), .B2(n9967), .C1(
        n15054), .C2(P3_U3151), .ZN(P3_U3283) );
  OAI222_X1 U12499 ( .A1(n8316), .A2(P1_U3086), .B1(n14366), .B2(n9970), .C1(
        n9969), .C2(n14363), .ZN(P1_U3353) );
  INV_X1 U12500 ( .A(n9971), .ZN(n9974) );
  INV_X1 U12501 ( .A(n14735), .ZN(n10024) );
  OAI222_X1 U12502 ( .A1(n13688), .A2(n9972), .B1(n13685), .B2(n9974), .C1(
        P2_U3088), .C2(n10024), .ZN(P2_U3321) );
  INV_X1 U12503 ( .A(n10247), .ZN(n10259) );
  OAI222_X1 U12504 ( .A1(n10259), .A2(P1_U3086), .B1(n14366), .B2(n9974), .C1(
        n9973), .C2(n14363), .ZN(P1_U3349) );
  INV_X1 U12505 ( .A(n13004), .ZN(n14380) );
  AOI222_X1 U12506 ( .A1(n9975), .A2(n14381), .B1(SI_4_), .B2(n14380), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11084), .ZN(n9976) );
  INV_X1 U12507 ( .A(n9976), .ZN(P3_U3291) );
  AOI222_X1 U12508 ( .A1(n9978), .A2(n14381), .B1(SI_7_), .B2(n14380), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n9977), .ZN(n9979) );
  INV_X1 U12509 ( .A(n9979), .ZN(P3_U3288) );
  AOI222_X1 U12510 ( .A1(n9980), .A2(n14381), .B1(SI_5_), .B2(n14380), .C1(
        n11057), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9981) );
  INV_X1 U12511 ( .A(n9981), .ZN(P3_U3290) );
  AOI222_X1 U12512 ( .A1(n9982), .A2(n14381), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n6500), .C1(SI_2_), .C2(n14380), .ZN(n9983) );
  INV_X1 U12513 ( .A(n9983), .ZN(P3_U3293) );
  AOI222_X1 U12514 ( .A1(n9984), .A2(n14381), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11132), .C1(SI_3_), .C2(n14380), .ZN(n9985) );
  INV_X1 U12515 ( .A(n9985), .ZN(P3_U3292) );
  AOI222_X1 U12516 ( .A1(n9987), .A2(n14381), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9986), .C1(SI_10_), .C2(n14380), .ZN(n9988) );
  INV_X1 U12517 ( .A(n9988), .ZN(P3_U3285) );
  INV_X1 U12518 ( .A(n9989), .ZN(n9992) );
  INV_X1 U12519 ( .A(n13175), .ZN(n13191) );
  OAI222_X1 U12520 ( .A1(n13688), .A2(n9990), .B1(n13685), .B2(n9992), .C1(
        P2_U3088), .C2(n13191), .ZN(P2_U3320) );
  INV_X1 U12521 ( .A(n13939), .ZN(n9993) );
  OAI222_X1 U12522 ( .A1(n9993), .A2(P1_U3086), .B1(n14366), .B2(n9992), .C1(
        n9991), .C2(n14363), .ZN(P1_U3348) );
  OAI222_X1 U12523 ( .A1(n10125), .A2(P1_U3086), .B1(n14366), .B2(n9995), .C1(
        n9994), .C2(n14363), .ZN(P1_U3350) );
  INV_X1 U12524 ( .A(n14582), .ZN(n9998) );
  OAI222_X1 U12525 ( .A1(n9998), .A2(P1_U3086), .B1(n14366), .B2(n9997), .C1(
        n9996), .C2(n14363), .ZN(P1_U3351) );
  INV_X1 U12526 ( .A(n13924), .ZN(n10001) );
  OAI222_X1 U12527 ( .A1(n10001), .A2(P1_U3086), .B1(n14366), .B2(n10000), 
        .C1(n9999), .C2(n14363), .ZN(P1_U3352) );
  INV_X1 U12528 ( .A(n13955), .ZN(n10004) );
  INV_X1 U12529 ( .A(n10002), .ZN(n10005) );
  OAI222_X1 U12530 ( .A1(n10004), .A2(P1_U3086), .B1(n14366), .B2(n10005), 
        .C1(n10003), .C2(n14363), .ZN(P1_U3347) );
  INV_X1 U12531 ( .A(n14747), .ZN(n13192) );
  OAI222_X1 U12532 ( .A1(n13688), .A2(n10006), .B1(n13685), .B2(n10005), .C1(
        P2_U3088), .C2(n13192), .ZN(P2_U3319) );
  OAI222_X1 U12533 ( .A1(n12387), .A2(n10008), .B1(n13004), .B2(n10007), .C1(
        n15070), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12534 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10016) );
  INV_X1 U12535 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10014) );
  INV_X1 U12536 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10012) );
  INV_X1 U12537 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10429) );
  MUX2_X1 U12538 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10429), .S(n10074), .Z(
        n10010) );
  INV_X1 U12539 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10627) );
  MUX2_X1 U12540 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10627), .S(n13162), .Z(
        n13164) );
  AND2_X1 U12541 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n13165) );
  NAND2_X1 U12542 ( .A1(n13164), .A2(n13165), .ZN(n13163) );
  NAND2_X1 U12543 ( .A1(n13162), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U12544 ( .A1(n13163), .A2(n10009), .ZN(n10073) );
  NAND2_X1 U12545 ( .A1(n10010), .A2(n10073), .ZN(n10075) );
  OAI21_X1 U12546 ( .B1(n10429), .B2(n10084), .A(n10075), .ZN(n14702) );
  MUX2_X1 U12547 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10012), .S(n14699), .Z(
        n14701) );
  NAND2_X1 U12548 ( .A1(n14702), .A2(n14701), .ZN(n14700) );
  OAI21_X1 U12549 ( .B1(n10012), .B2(n10011), .A(n14700), .ZN(n14714) );
  MUX2_X1 U12550 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10014), .S(n14711), .Z(
        n14713) );
  NAND2_X1 U12551 ( .A1(n14714), .A2(n14713), .ZN(n14712) );
  OAI21_X1 U12552 ( .B1(n10014), .B2(n10013), .A(n14712), .ZN(n14726) );
  MUX2_X1 U12553 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10016), .S(n14723), .Z(
        n14725) );
  NAND2_X1 U12554 ( .A1(n14726), .A2(n14725), .ZN(n14724) );
  OAI21_X1 U12555 ( .B1(n10016), .B2(n10015), .A(n14724), .ZN(n14738) );
  INV_X1 U12556 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10017) );
  MUX2_X1 U12557 ( .A(n10017), .B(P2_REG2_REG_6__SCAN_IN), .S(n14735), .Z(
        n10018) );
  INV_X1 U12558 ( .A(n10018), .ZN(n14737) );
  NAND2_X1 U12559 ( .A1(n14738), .A2(n14737), .ZN(n14736) );
  NAND2_X1 U12560 ( .A1(n14735), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10021) );
  INV_X1 U12561 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10019) );
  MUX2_X1 U12562 ( .A(n10019), .B(P2_REG2_REG_7__SCAN_IN), .S(n13175), .Z(
        n10020) );
  AOI21_X1 U12563 ( .B1(n14736), .B2(n10021), .A(n10020), .ZN(n13174) );
  NOR2_X1 U12564 ( .A1(n10155), .A2(P2_U3088), .ZN(n13682) );
  AND2_X1 U12565 ( .A1(n10032), .A2(n13682), .ZN(n10029) );
  INV_X1 U12566 ( .A(n8240), .ZN(n13225) );
  AND2_X1 U12567 ( .A1(n10029), .A2(n13225), .ZN(n14851) );
  NAND3_X1 U12568 ( .A1(n14736), .A2(n10021), .A3(n10020), .ZN(n10022) );
  NAND2_X1 U12569 ( .A1(n14851), .A2(n10022), .ZN(n10037) );
  INV_X1 U12570 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10160) );
  MUX2_X1 U12571 ( .A(n10160), .B(P2_REG1_REG_1__SCAN_IN), .S(n13162), .Z(
        n13159) );
  NAND2_X1 U12572 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13160) );
  AOI21_X1 U12573 ( .B1(n13162), .B2(P2_REG1_REG_1__SCAN_IN), .A(n13158), .ZN(
        n10081) );
  INV_X1 U12574 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n14945) );
  MUX2_X1 U12575 ( .A(n14945), .B(P2_REG1_REG_2__SCAN_IN), .S(n10074), .Z(
        n10080) );
  AOI21_X1 U12576 ( .B1(n10074), .B2(P2_REG1_REG_2__SCAN_IN), .A(n10079), .ZN(
        n14705) );
  INV_X1 U12577 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10023) );
  MUX2_X1 U12578 ( .A(n10023), .B(P2_REG1_REG_3__SCAN_IN), .S(n14699), .Z(
        n14704) );
  NOR2_X1 U12579 ( .A1(n14705), .A2(n14704), .ZN(n14703) );
  AOI21_X1 U12580 ( .B1(n14699), .B2(P2_REG1_REG_3__SCAN_IN), .A(n14703), .ZN(
        n14717) );
  INV_X1 U12581 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14947) );
  MUX2_X1 U12582 ( .A(n14947), .B(P2_REG1_REG_4__SCAN_IN), .S(n14711), .Z(
        n14716) );
  AOI21_X1 U12583 ( .B1(n14711), .B2(P2_REG1_REG_4__SCAN_IN), .A(n14715), .ZN(
        n14729) );
  INV_X1 U12584 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14949) );
  MUX2_X1 U12585 ( .A(n14949), .B(P2_REG1_REG_5__SCAN_IN), .S(n14723), .Z(
        n14728) );
  NOR2_X1 U12586 ( .A1(n14729), .A2(n14728), .ZN(n14727) );
  AOI21_X1 U12587 ( .B1(n14723), .B2(P2_REG1_REG_5__SCAN_IN), .A(n14727), .ZN(
        n14741) );
  INV_X1 U12588 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14951) );
  MUX2_X1 U12589 ( .A(n14951), .B(P2_REG1_REG_6__SCAN_IN), .S(n14735), .Z(
        n14740) );
  NOR2_X1 U12590 ( .A1(n10024), .A2(n14951), .ZN(n10028) );
  INV_X1 U12591 ( .A(n10028), .ZN(n10026) );
  INV_X1 U12592 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n14953) );
  MUX2_X1 U12593 ( .A(n14953), .B(P2_REG1_REG_7__SCAN_IN), .S(n13175), .Z(
        n10025) );
  NAND2_X1 U12594 ( .A1(n10026), .A2(n10025), .ZN(n10030) );
  MUX2_X1 U12595 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n14953), .S(n13175), .Z(
        n10027) );
  OAI21_X1 U12596 ( .B1(n14739), .B2(n10028), .A(n10027), .ZN(n13190) );
  NAND2_X1 U12597 ( .A1(n10029), .A2(n8240), .ZN(n14805) );
  OAI211_X1 U12598 ( .C1(n14739), .C2(n10030), .A(n13190), .B(n14877), .ZN(
        n10036) );
  AND2_X1 U12599 ( .A1(n10155), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12600 ( .A1(n10032), .A2(n10031), .ZN(n14873) );
  NAND2_X1 U12601 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10671) );
  OAI21_X1 U12602 ( .B1(n10033), .B2(n9453), .A(n10671), .ZN(n10034) );
  AOI21_X1 U12603 ( .B1(n13175), .B2(n14823), .A(n10034), .ZN(n10035) );
  OAI211_X1 U12604 ( .C1(n13174), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        P2_U3221) );
  INV_X1 U12605 ( .A(n10038), .ZN(n10041) );
  INV_X1 U12606 ( .A(n14759), .ZN(n13194) );
  OAI222_X1 U12607 ( .A1(n13688), .A2(n10039), .B1(n13685), .B2(n10041), .C1(
        P2_U3088), .C2(n13194), .ZN(P2_U3318) );
  INV_X1 U12608 ( .A(n13972), .ZN(n13963) );
  OAI222_X1 U12609 ( .A1(n13963), .A2(P1_U3086), .B1(n14366), .B2(n10041), 
        .C1(n10040), .C2(n14363), .ZN(P1_U3346) );
  OAI222_X1 U12610 ( .A1(n12387), .A2(n10043), .B1(n13004), .B2(n10042), .C1(
        n15091), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12611 ( .A(n10317), .ZN(n10222) );
  INV_X1 U12612 ( .A(n10044), .ZN(n10046) );
  OAI222_X1 U12613 ( .A1(n10222), .A2(P1_U3086), .B1(n14366), .B2(n10046), 
        .C1(n10045), .C2(n14363), .ZN(P1_U3345) );
  INV_X1 U12614 ( .A(n14772), .ZN(n13196) );
  OAI222_X1 U12615 ( .A1(n13688), .A2(n10047), .B1(n13685), .B2(n10046), .C1(
        P2_U3088), .C2(n13196), .ZN(P2_U3317) );
  INV_X1 U12616 ( .A(n10281), .ZN(n10048) );
  AOI22_X1 U12617 ( .A1(n14639), .A2(n10050), .B1(n10290), .B2(n10049), .ZN(
        P1_U3445) );
  AOI22_X1 U12618 ( .A1(n14639), .A2(n10051), .B1(n10290), .B2(n10279), .ZN(
        P1_U3446) );
  INV_X1 U12619 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10052) );
  OAI211_X1 U12620 ( .C1(n14881), .C2(P2_REG2_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .B(n14873), .ZN(n10053) );
  AOI21_X1 U12621 ( .B1(n14877), .B2(n10052), .A(n10053), .ZN(n10057) );
  AOI21_X1 U12622 ( .B1(n14851), .B2(P2_REG2_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U12623 ( .A1(n14849), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10055) );
  NAND3_X1 U12624 ( .A1(n10053), .A2(n14877), .A3(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10054) );
  OAI211_X1 U12625 ( .C1(n10057), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        P2_U3214) );
  OAI222_X1 U12626 ( .A1(n12387), .A2(n10059), .B1(n13004), .B2(n10058), .C1(
        n14408), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12627 ( .A(n10060), .ZN(n10569) );
  NAND2_X1 U12628 ( .A1(n10569), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12034) );
  NAND2_X1 U12629 ( .A1(n10282), .A2(n12034), .ZN(n10064) );
  NAND2_X1 U12630 ( .A1(n11976), .A2(n10060), .ZN(n10061) );
  AND2_X1 U12631 ( .A1(n10061), .A2(n8304), .ZN(n10063) );
  INV_X1 U12632 ( .A(n10063), .ZN(n10062) );
  AND2_X1 U12633 ( .A1(n10064), .A2(n10063), .ZN(n10108) );
  INV_X1 U12634 ( .A(n14362), .ZN(n10065) );
  INV_X1 U12635 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10771) );
  AOI21_X1 U12636 ( .B1(n10065), .B2(n10771), .A(n8651), .ZN(n13900) );
  OAI21_X1 U12637 ( .B1(n10065), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13900), .ZN(
        n10066) );
  XNOR2_X1 U12638 ( .A(n10066), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U12639 ( .A1(n10108), .A2(n10067), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10068) );
  OAI21_X1 U12640 ( .B1(n14637), .B2(n9436), .A(n10068), .ZN(P1_U3243) );
  INV_X1 U12641 ( .A(n10069), .ZN(n10071) );
  INV_X1 U12642 ( .A(n14784), .ZN(n13197) );
  OAI222_X1 U12643 ( .A1(n13688), .A2(n10070), .B1(n13685), .B2(n10071), .C1(
        P2_U3088), .C2(n13197), .ZN(P2_U3316) );
  INV_X1 U12644 ( .A(n13988), .ZN(n10318) );
  OAI222_X1 U12645 ( .A1(n14363), .A2(n10072), .B1(n14366), .B2(n10071), .C1(
        P1_U3086), .C2(n10318), .ZN(P1_U3344) );
  INV_X1 U12646 ( .A(n10073), .ZN(n10078) );
  MUX2_X1 U12647 ( .A(n10429), .B(P2_REG2_REG_2__SCAN_IN), .S(n10074), .Z(
        n10077) );
  INV_X1 U12648 ( .A(n10075), .ZN(n10076) );
  AOI211_X1 U12649 ( .C1(n10078), .C2(n10077), .A(n10076), .B(n14881), .ZN(
        n10087) );
  AOI211_X1 U12650 ( .C1(n10081), .C2(n10080), .A(n10079), .B(n14805), .ZN(
        n10086) );
  NAND2_X1 U12651 ( .A1(n14849), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U12652 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(P2_U3088), .ZN(n10082) );
  OAI211_X1 U12653 ( .C1(n14873), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10085) );
  OR3_X1 U12654 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(P2_U3216) );
  OAI222_X1 U12655 ( .A1(n12387), .A2(n10090), .B1(n10089), .B2(P3_U3151), 
        .C1(n10088), .C2(n13004), .ZN(P3_U3279) );
  INV_X1 U12656 ( .A(n10325), .ZN(n10389) );
  INV_X1 U12657 ( .A(n10091), .ZN(n10096) );
  OAI222_X1 U12658 ( .A1(P1_U3086), .A2(n10389), .B1(n14366), .B2(n10096), 
        .C1(n10092), .C2(n14363), .ZN(P1_U3343) );
  OAI222_X1 U12659 ( .A1(n12387), .A2(n10095), .B1(n13004), .B2(n10094), .C1(
        n10093), .C2(P3_U3151), .ZN(P3_U3278) );
  OAI222_X1 U12660 ( .A1(n13688), .A2(n10097), .B1(n14796), .B2(P2_U3088), 
        .C1(n13685), .C2(n10096), .ZN(P2_U3315) );
  NAND2_X1 U12661 ( .A1(n10108), .A2(n14362), .ZN(n14626) );
  INV_X1 U12662 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10098) );
  MUX2_X1 U12663 ( .A(n10098), .B(P1_REG1_REG_5__SCAN_IN), .S(n10125), .Z(
        n10106) );
  INV_X1 U12664 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10099) );
  MUX2_X1 U12665 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10099), .S(n13907), .Z(
        n10102) );
  INV_X1 U12666 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10100) );
  MUX2_X1 U12667 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10100), .S(n13888), .Z(
        n13886) );
  AND2_X1 U12668 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13887) );
  NAND2_X1 U12669 ( .A1(n13886), .A2(n13887), .ZN(n13902) );
  NAND2_X1 U12670 ( .A1(n13888), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n13901) );
  NAND2_X1 U12671 ( .A1(n13902), .A2(n13901), .ZN(n10101) );
  NAND2_X1 U12672 ( .A1(n10102), .A2(n10101), .ZN(n13922) );
  INV_X1 U12673 ( .A(n13922), .ZN(n10104) );
  NOR2_X1 U12674 ( .A1(n8316), .A2(n10099), .ZN(n13918) );
  INV_X1 U12675 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n13919) );
  MUX2_X1 U12676 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n13919), .S(n13924), .Z(
        n10103) );
  OAI21_X1 U12677 ( .B1(n10104), .B2(n13918), .A(n10103), .ZN(n14577) );
  NAND2_X1 U12678 ( .A1(n13924), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14576) );
  INV_X1 U12679 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14689) );
  MUX2_X1 U12680 ( .A(n14689), .B(P1_REG1_REG_4__SCAN_IN), .S(n14582), .Z(
        n14575) );
  AOI21_X1 U12681 ( .B1(n14577), .B2(n14576), .A(n14575), .ZN(n14574) );
  AOI21_X1 U12682 ( .B1(n14582), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14574), .ZN(
        n10105) );
  NAND2_X1 U12683 ( .A1(n10105), .A2(n10106), .ZN(n10198) );
  OAI21_X1 U12684 ( .B1(n10106), .B2(n10105), .A(n10198), .ZN(n10122) );
  NOR2_X1 U12685 ( .A1(n8651), .A2(n14362), .ZN(n10107) );
  INV_X1 U12686 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10109) );
  MUX2_X1 U12687 ( .A(n10109), .B(P1_REG2_REG_5__SCAN_IN), .S(n10125), .Z(
        n10117) );
  INV_X1 U12688 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n13908) );
  MUX2_X1 U12689 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n13908), .S(n13907), .Z(
        n10111) );
  INV_X1 U12690 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14254) );
  MUX2_X1 U12691 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n14254), .S(n13888), .Z(
        n13889) );
  AND2_X1 U12692 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13895) );
  NAND2_X1 U12693 ( .A1(n13889), .A2(n13895), .ZN(n13910) );
  NAND2_X1 U12694 ( .A1(n13888), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U12695 ( .A1(n13910), .A2(n13909), .ZN(n10110) );
  NAND2_X1 U12696 ( .A1(n10111), .A2(n10110), .ZN(n13928) );
  NAND2_X1 U12697 ( .A1(n13907), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U12698 ( .A1(n13928), .A2(n13926), .ZN(n10113) );
  INV_X1 U12699 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n13925) );
  MUX2_X1 U12700 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n13925), .S(n13924), .Z(
        n10112) );
  NAND2_X1 U12701 ( .A1(n10113), .A2(n10112), .ZN(n14585) );
  NAND2_X1 U12702 ( .A1(n13924), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14584) );
  NAND2_X1 U12703 ( .A1(n14585), .A2(n14584), .ZN(n10115) );
  INV_X1 U12704 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10753) );
  MUX2_X1 U12705 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10753), .S(n14582), .Z(
        n10114) );
  NAND2_X1 U12706 ( .A1(n10115), .A2(n10114), .ZN(n14587) );
  NAND2_X1 U12707 ( .A1(n14582), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U12708 ( .A1(n14587), .A2(n10118), .ZN(n10116) );
  NAND2_X1 U12709 ( .A1(n10117), .A2(n10116), .ZN(n10250) );
  MUX2_X1 U12710 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10109), .S(n10125), .Z(
        n10119) );
  NAND3_X1 U12711 ( .A1(n10119), .A2(n14587), .A3(n10118), .ZN(n10120) );
  AND3_X1 U12712 ( .A1(n14628), .A2(n10250), .A3(n10120), .ZN(n10121) );
  AOI21_X1 U12713 ( .B1(n14600), .B2(n10122), .A(n10121), .ZN(n10124) );
  AND2_X1 U12714 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11239) );
  AOI21_X1 U12715 ( .B1(n14596), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n11239), .ZN(
        n10123) );
  OAI211_X1 U12716 ( .C1(n10125), .C2(n14618), .A(n10124), .B(n10123), .ZN(
        P1_U3248) );
  NAND2_X1 U12717 ( .A1(n10334), .A2(n10335), .ZN(n10345) );
  INV_X1 U12718 ( .A(n10126), .ZN(n11478) );
  XNOR2_X1 U12719 ( .A(n11440), .B(P2_B_REG_SCAN_IN), .ZN(n10127) );
  NAND2_X1 U12720 ( .A1(n11478), .A2(n10127), .ZN(n10129) );
  INV_X1 U12721 ( .A(n13690), .ZN(n10128) );
  AND2_X1 U12722 ( .A1(n10129), .A2(n10128), .ZN(n14883) );
  NOR4_X1 U12723 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n10138) );
  NOR4_X1 U12724 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n10133) );
  NOR4_X1 U12725 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n10132) );
  NOR4_X1 U12726 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n10131) );
  NOR4_X1 U12727 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n10130) );
  NAND4_X1 U12728 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10134) );
  NOR4_X1 U12729 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n10135), .A4(n10134), .ZN(n10137) );
  NOR4_X1 U12730 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n10136) );
  NAND3_X1 U12731 ( .A1(n10138), .A2(n10137), .A3(n10136), .ZN(n10139) );
  NAND2_X1 U12732 ( .A1(n14883), .A2(n10139), .ZN(n10331) );
  AND2_X1 U12733 ( .A1(n10345), .A2(n10331), .ZN(n10262) );
  INV_X1 U12734 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14890) );
  NAND2_X1 U12735 ( .A1(n14883), .A2(n14890), .ZN(n10141) );
  NAND2_X1 U12736 ( .A1(n11478), .A2(n13690), .ZN(n10140) );
  NAND2_X1 U12737 ( .A1(n10141), .A2(n10140), .ZN(n10260) );
  AND2_X1 U12738 ( .A1(n10143), .A2(n10142), .ZN(n10344) );
  AND2_X1 U12739 ( .A1(n10344), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14887) );
  AND2_X1 U12740 ( .A1(n10260), .A2(n14887), .ZN(n14888) );
  OR2_X1 U12741 ( .A1(n10265), .A2(n10348), .ZN(n10342) );
  NAND3_X1 U12742 ( .A1(n10262), .A2(n14888), .A3(n10342), .ZN(n10161) );
  INV_X1 U12743 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14885) );
  NAND2_X1 U12744 ( .A1(n14883), .A2(n14885), .ZN(n10146) );
  NAND2_X1 U12745 ( .A1(n11440), .A2(n13690), .ZN(n10145) );
  NAND2_X1 U12746 ( .A1(n10146), .A2(n10145), .ZN(n14886) );
  OR2_X1 U12747 ( .A1(n10265), .A2(n10150), .ZN(n13648) );
  XNOR2_X1 U12748 ( .A(n10227), .B(n10225), .ZN(n10630) );
  NAND2_X1 U12749 ( .A1(n10623), .A2(n10338), .ZN(n10430) );
  OAI211_X1 U12750 ( .C1(n10623), .C2(n10338), .A(n13510), .B(n10430), .ZN(
        n10149) );
  INV_X1 U12751 ( .A(n10149), .ZN(n10625) );
  NAND2_X1 U12752 ( .A1(n6469), .A2(n10150), .ZN(n10152) );
  NAND2_X2 U12753 ( .A1(n10152), .A2(n10151), .ZN(n13526) );
  NOR2_X1 U12754 ( .A1(n10338), .A2(n13157), .ZN(n10153) );
  NAND2_X1 U12755 ( .A1(n10153), .A2(n10227), .ZN(n10231) );
  OAI21_X1 U12756 ( .B1(n10153), .B2(n10227), .A(n10231), .ZN(n10156) );
  INV_X1 U12757 ( .A(n10155), .ZN(n10154) );
  NAND2_X1 U12758 ( .A1(n10335), .A2(n10155), .ZN(n13503) );
  AOI222_X1 U12759 ( .A1(n13526), .A2(n10156), .B1(n13157), .B2(n13523), .C1(
        n13155), .C2(n13521), .ZN(n10626) );
  INV_X1 U12760 ( .A(n10626), .ZN(n10157) );
  AOI211_X1 U12761 ( .C1(n14936), .C2(n13018), .A(n10625), .B(n10157), .ZN(
        n10158) );
  OAI21_X1 U12762 ( .B1(n14922), .B2(n10630), .A(n10158), .ZN(n10162) );
  NAND2_X1 U12763 ( .A1(n10162), .A2(n14960), .ZN(n10159) );
  OAI21_X1 U12764 ( .B1(n14960), .B2(n10160), .A(n10159), .ZN(P2_U3500) );
  INV_X1 U12765 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U12766 ( .A1(n10162), .A2(n14944), .ZN(n10163) );
  OAI21_X1 U12767 ( .B1(n14944), .B2(n10164), .A(n10163), .ZN(P2_U3433) );
  NOR2_X1 U12768 ( .A1(n10165), .A2(n13000), .ZN(n10167) );
  CLKBUF_X1 U12769 ( .A(n10167), .Z(n10185) );
  INV_X1 U12770 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10166) );
  NOR2_X1 U12771 ( .A1(n10185), .A2(n10166), .ZN(P3_U3261) );
  INV_X1 U12772 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10168) );
  NOR2_X1 U12773 ( .A1(n10185), .A2(n10168), .ZN(P3_U3262) );
  INV_X1 U12774 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10169) );
  NOR2_X1 U12775 ( .A1(n10167), .A2(n10169), .ZN(P3_U3260) );
  INV_X1 U12776 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10170) );
  NOR2_X1 U12777 ( .A1(n10185), .A2(n10170), .ZN(P3_U3259) );
  INV_X1 U12778 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U12779 ( .A1(n10185), .A2(n10171), .ZN(P3_U3263) );
  INV_X1 U12780 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10172) );
  NOR2_X1 U12781 ( .A1(n10185), .A2(n10172), .ZN(P3_U3257) );
  INV_X1 U12782 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10173) );
  NOR2_X1 U12783 ( .A1(n10185), .A2(n10173), .ZN(P3_U3256) );
  INV_X1 U12784 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10174) );
  NOR2_X1 U12785 ( .A1(n10185), .A2(n10174), .ZN(P3_U3255) );
  INV_X1 U12786 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U12787 ( .A1(n10185), .A2(n10175), .ZN(P3_U3254) );
  INV_X1 U12788 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10176) );
  NOR2_X1 U12789 ( .A1(n10185), .A2(n10176), .ZN(P3_U3253) );
  INV_X1 U12790 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10177) );
  NOR2_X1 U12791 ( .A1(n10167), .A2(n10177), .ZN(P3_U3258) );
  INV_X1 U12792 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U12793 ( .A1(n10185), .A2(n10178), .ZN(P3_U3251) );
  INV_X1 U12794 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10179) );
  NOR2_X1 U12795 ( .A1(n10185), .A2(n10179), .ZN(P3_U3250) );
  INV_X1 U12796 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10180) );
  NOR2_X1 U12797 ( .A1(n10185), .A2(n10180), .ZN(P3_U3249) );
  INV_X1 U12798 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10181) );
  NOR2_X1 U12799 ( .A1(n10185), .A2(n10181), .ZN(P3_U3248) );
  INV_X1 U12800 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10182) );
  NOR2_X1 U12801 ( .A1(n10185), .A2(n10182), .ZN(P3_U3247) );
  INV_X1 U12802 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10183) );
  NOR2_X1 U12803 ( .A1(n10185), .A2(n10183), .ZN(P3_U3252) );
  INV_X1 U12804 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U12805 ( .A1(n10185), .A2(n10184), .ZN(P3_U3246) );
  INV_X1 U12806 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10186) );
  NOR2_X1 U12807 ( .A1(n10167), .A2(n10186), .ZN(P3_U3245) );
  INV_X1 U12808 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10187) );
  NOR2_X1 U12809 ( .A1(n10167), .A2(n10187), .ZN(P3_U3244) );
  INV_X1 U12810 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10188) );
  NOR2_X1 U12811 ( .A1(n10167), .A2(n10188), .ZN(P3_U3243) );
  INV_X1 U12812 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10189) );
  NOR2_X1 U12813 ( .A1(n10167), .A2(n10189), .ZN(P3_U3242) );
  INV_X1 U12814 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10190) );
  NOR2_X1 U12815 ( .A1(n10167), .A2(n10190), .ZN(P3_U3241) );
  INV_X1 U12816 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10191) );
  NOR2_X1 U12817 ( .A1(n10167), .A2(n10191), .ZN(P3_U3240) );
  INV_X1 U12818 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10192) );
  NOR2_X1 U12819 ( .A1(n10167), .A2(n10192), .ZN(P3_U3239) );
  INV_X1 U12820 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10193) );
  NOR2_X1 U12821 ( .A1(n10167), .A2(n10193), .ZN(P3_U3238) );
  INV_X1 U12822 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10194) );
  NOR2_X1 U12823 ( .A1(n10167), .A2(n10194), .ZN(P3_U3237) );
  INV_X1 U12824 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U12825 ( .A1(n10185), .A2(n10195), .ZN(P3_U3236) );
  INV_X1 U12826 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U12827 ( .A1(n10185), .A2(n10196), .ZN(P3_U3235) );
  INV_X1 U12828 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10197) );
  NOR2_X1 U12829 ( .A1(n10185), .A2(n10197), .ZN(P3_U3234) );
  OAI21_X1 U12830 ( .B1(n10204), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10198), .ZN(
        n10252) );
  INV_X1 U12831 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14691) );
  MUX2_X1 U12832 ( .A(n14691), .B(P1_REG1_REG_6__SCAN_IN), .S(n10247), .Z(
        n10253) );
  OR2_X1 U12833 ( .A1(n10252), .A2(n10253), .ZN(n13936) );
  NAND2_X1 U12834 ( .A1(n10247), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n13935) );
  INV_X1 U12835 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10199) );
  MUX2_X1 U12836 ( .A(n10199), .B(P1_REG1_REG_7__SCAN_IN), .S(n13939), .Z(
        n13934) );
  AOI21_X1 U12837 ( .B1(n13936), .B2(n13935), .A(n13934), .ZN(n13933) );
  AOI21_X1 U12838 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n13939), .A(n13933), .ZN(
        n13953) );
  INV_X1 U12839 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n14693) );
  MUX2_X1 U12840 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n14693), .S(n13955), .Z(
        n13952) );
  AND2_X1 U12841 ( .A1(n13953), .A2(n13952), .ZN(n13969) );
  NOR2_X1 U12842 ( .A1(n13955), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n13967) );
  INV_X1 U12843 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10200) );
  MUX2_X1 U12844 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10200), .S(n13972), .Z(
        n13968) );
  OAI21_X1 U12845 ( .B1(n13969), .B2(n13967), .A(n13968), .ZN(n13966) );
  OAI21_X1 U12846 ( .B1(n13972), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13966), .ZN(
        n10202) );
  INV_X1 U12847 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14696) );
  MUX2_X1 U12848 ( .A(n14696), .B(P1_REG1_REG_10__SCAN_IN), .S(n10317), .Z(
        n10201) );
  NOR2_X1 U12849 ( .A1(n10202), .A2(n10201), .ZN(n10316) );
  AOI211_X1 U12850 ( .C1(n10202), .C2(n10201), .A(n14626), .B(n10316), .ZN(
        n10203) );
  INV_X1 U12851 ( .A(n10203), .ZN(n10221) );
  NAND2_X1 U12852 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11534)
         );
  NAND2_X1 U12853 ( .A1(n10204), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U12854 ( .A1(n10250), .A2(n10249), .ZN(n10206) );
  INV_X1 U12855 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10822) );
  MUX2_X1 U12856 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10822), .S(n10247), .Z(
        n10205) );
  NAND2_X1 U12857 ( .A1(n10206), .A2(n10205), .ZN(n13941) );
  NAND2_X1 U12858 ( .A1(n10247), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13940) );
  NAND2_X1 U12859 ( .A1(n13941), .A2(n13940), .ZN(n10208) );
  INV_X1 U12860 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10906) );
  MUX2_X1 U12861 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10906), .S(n13939), .Z(
        n10207) );
  NAND2_X1 U12862 ( .A1(n10208), .A2(n10207), .ZN(n13958) );
  NAND2_X1 U12863 ( .A1(n13939), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n13957) );
  NAND2_X1 U12864 ( .A1(n13958), .A2(n13957), .ZN(n10210) );
  INV_X1 U12865 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11144) );
  MUX2_X1 U12866 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11144), .S(n13955), .Z(
        n10209) );
  NAND2_X1 U12867 ( .A1(n10210), .A2(n10209), .ZN(n13975) );
  NAND2_X1 U12868 ( .A1(n13955), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n13974) );
  NAND2_X1 U12869 ( .A1(n13975), .A2(n13974), .ZN(n10213) );
  INV_X1 U12870 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10211) );
  MUX2_X1 U12871 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10211), .S(n13972), .Z(
        n10212) );
  NAND2_X1 U12872 ( .A1(n10213), .A2(n10212), .ZN(n13977) );
  NAND2_X1 U12873 ( .A1(n13972), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U12874 ( .A1(n13977), .A2(n10214), .ZN(n10217) );
  INV_X1 U12875 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10215) );
  MUX2_X1 U12876 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10215), .S(n10317), .Z(
        n10216) );
  NAND2_X1 U12877 ( .A1(n10217), .A2(n10216), .ZN(n13991) );
  OAI211_X1 U12878 ( .C1(n10217), .C2(n10216), .A(n14628), .B(n13991), .ZN(
        n10218) );
  NAND2_X1 U12879 ( .A1(n11534), .A2(n10218), .ZN(n10219) );
  AOI21_X1 U12880 ( .B1(n14596), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10219), 
        .ZN(n10220) );
  OAI211_X1 U12881 ( .C1(n14618), .C2(n10222), .A(n10221), .B(n10220), .ZN(
        P1_U3253) );
  INV_X1 U12882 ( .A(n10223), .ZN(n10244) );
  OAI222_X1 U12883 ( .A1(n13685), .A2(n10244), .B1(n13200), .B2(P2_U3088), 
        .C1(n10224), .C2(n13688), .ZN(P2_U3314) );
  INV_X1 U12884 ( .A(n13648), .ZN(n14932) );
  INV_X1 U12885 ( .A(n10438), .ZN(n10426) );
  INV_X1 U12886 ( .A(n10225), .ZN(n10340) );
  NAND2_X1 U12887 ( .A1(n8193), .A2(n10623), .ZN(n10226) );
  OAI21_X1 U12888 ( .B1(n10340), .B2(n10227), .A(n10226), .ZN(n10425) );
  NAND2_X1 U12889 ( .A1(n10426), .A2(n10425), .ZN(n10424) );
  OR2_X1 U12890 ( .A1(n10591), .A2(n13155), .ZN(n10228) );
  NAND2_X1 U12891 ( .A1(n10424), .A2(n10228), .ZN(n10229) );
  OAI21_X1 U12892 ( .B1(n10229), .B2(n10233), .A(n10470), .ZN(n10497) );
  INV_X1 U12893 ( .A(n10491), .ZN(n10377) );
  OAI211_X1 U12894 ( .C1(n10377), .C2(n10431), .A(n13510), .B(n10503), .ZN(
        n10493) );
  OAI21_X1 U12895 ( .B1(n10377), .B2(n14927), .A(n10493), .ZN(n10241) );
  INV_X1 U12896 ( .A(n10497), .ZN(n10240) );
  NAND2_X1 U12897 ( .A1(n13018), .A2(n8193), .ZN(n10230) );
  NAND2_X1 U12898 ( .A1(n10231), .A2(n10230), .ZN(n10437) );
  NAND2_X1 U12899 ( .A1(n10437), .A2(n10438), .ZN(n10436) );
  OAI21_X1 U12900 ( .B1(n10235), .B2(n10234), .A(n10509), .ZN(n10238) );
  INV_X1 U12901 ( .A(n13153), .ZN(n10478) );
  OAI22_X1 U12902 ( .A1(n10478), .A2(n13503), .B1(n10236), .B2(n13505), .ZN(
        n10237) );
  AOI21_X1 U12903 ( .B1(n10238), .B2(n13526), .A(n10237), .ZN(n10239) );
  OAI21_X1 U12904 ( .B1(n10240), .B2(n10353), .A(n10239), .ZN(n10494) );
  AOI211_X1 U12905 ( .C1(n14932), .C2(n10497), .A(n10241), .B(n10494), .ZN(
        n10299) );
  NAND2_X1 U12906 ( .A1(n14957), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10242) );
  OAI21_X1 U12907 ( .B1(n10299), .B2(n14957), .A(n10242), .ZN(P2_U3502) );
  INV_X1 U12908 ( .A(n10385), .ZN(n14598) );
  OAI222_X1 U12909 ( .A1(P1_U3086), .A2(n14598), .B1(n14366), .B2(n10244), 
        .C1(n10243), .C2(n14363), .ZN(P1_U3342) );
  INV_X1 U12910 ( .A(SI_18_), .ZN(n10245) );
  OAI222_X1 U12911 ( .A1(n12387), .A2(n10246), .B1(n13004), .B2(n10245), .C1(
        n12611), .C2(P3_U3151), .ZN(P3_U3277) );
  MUX2_X1 U12912 ( .A(n10822), .B(P1_REG2_REG_6__SCAN_IN), .S(n10247), .Z(
        n10248) );
  NAND3_X1 U12913 ( .A1(n10250), .A2(n10249), .A3(n10248), .ZN(n10251) );
  NAND3_X1 U12914 ( .A1(n14628), .A2(n13941), .A3(n10251), .ZN(n10258) );
  NAND2_X1 U12915 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11208) );
  NAND2_X1 U12916 ( .A1(n10253), .A2(n10252), .ZN(n10254) );
  NAND3_X1 U12917 ( .A1(n14600), .A2(n13936), .A3(n10254), .ZN(n10255) );
  NAND2_X1 U12918 ( .A1(n11208), .A2(n10255), .ZN(n10256) );
  AOI21_X1 U12919 ( .B1(n14596), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10256), .ZN(
        n10257) );
  OAI211_X1 U12920 ( .C1(n14618), .C2(n10259), .A(n10258), .B(n10257), .ZN(
        P1_U3249) );
  INV_X1 U12921 ( .A(n10260), .ZN(n10332) );
  AND3_X1 U12922 ( .A1(n10332), .A2(n14887), .A3(n14886), .ZN(n10261) );
  NAND2_X1 U12923 ( .A1(n10262), .A2(n10261), .ZN(n10264) );
  NAND2_X1 U12924 ( .A1(n14887), .A2(n10267), .ZN(n10263) );
  OR2_X1 U12925 ( .A1(n10265), .A2(n11235), .ZN(n10499) );
  INV_X1 U12926 ( .A(n10499), .ZN(n10266) );
  AND2_X1 U12927 ( .A1(n13527), .A2(n10266), .ZN(n10741) );
  INV_X1 U12928 ( .A(n10741), .ZN(n10767) );
  NAND2_X1 U12929 ( .A1(n10354), .A2(n10267), .ZN(n13645) );
  INV_X1 U12930 ( .A(n13526), .ZN(n13500) );
  AOI21_X1 U12931 ( .B1(n13500), .B2(n10353), .A(n13647), .ZN(n10268) );
  AOI21_X1 U12932 ( .B1(n13521), .B2(n13156), .A(n10268), .ZN(n13646) );
  OAI21_X1 U12933 ( .B1(n10269), .B2(n13645), .A(n13646), .ZN(n10270) );
  AOI22_X1 U12934 ( .A1(n10270), .A2(n13527), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13529), .ZN(n10272) );
  INV_X2 U12935 ( .A(n13527), .ZN(n13512) );
  NAND2_X1 U12936 ( .A1(n13512), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10271) );
  OAI211_X1 U12937 ( .C1(n10767), .C2(n13647), .A(n10272), .B(n10271), .ZN(
        P2_U3265) );
  INV_X1 U12938 ( .A(n14240), .ZN(n10302) );
  NAND2_X1 U12939 ( .A1(n10303), .A2(n11584), .ZN(n10276) );
  INV_X1 U12940 ( .A(n10274), .ZN(n10277) );
  NAND2_X1 U12941 ( .A1(n10277), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10275) );
  OAI211_X1 U12942 ( .C1(n11638), .C2(n10302), .A(n10276), .B(n10275), .ZN(
        n10458) );
  AOI222_X1 U12943 ( .A1(n10303), .A2(n12372), .B1(n14240), .B2(n11584), .C1(
        n10277), .C2(P1_IR_REG_0__SCAN_IN), .ZN(n10459) );
  XOR2_X1 U12944 ( .A(n10458), .B(n10459), .Z(n13894) );
  NAND2_X1 U12945 ( .A1(n10278), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10280) );
  AOI21_X1 U12946 ( .B1(n10281), .B2(n10280), .A(n10279), .ZN(n10642) );
  NAND2_X1 U12947 ( .A1(n10644), .A2(n10642), .ZN(n10292) );
  OR2_X1 U12948 ( .A1(n10292), .A2(n10282), .ZN(n10296) );
  INV_X1 U12949 ( .A(n10296), .ZN(n10285) );
  AND2_X1 U12950 ( .A1(n10283), .A2(n14680), .ZN(n10284) );
  NAND2_X1 U12951 ( .A1(n10292), .A2(n10286), .ZN(n10289) );
  AND2_X1 U12952 ( .A1(n10274), .A2(n10287), .ZN(n10288) );
  NAND2_X1 U12953 ( .A1(n10289), .A2(n10288), .ZN(n10570) );
  INV_X1 U12954 ( .A(n10570), .ZN(n10291) );
  NAND2_X1 U12955 ( .A1(n10291), .A2(n10290), .ZN(n13738) );
  AOI22_X1 U12956 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n13738), .B1(n13825), 
        .B2(n14248), .ZN(n10298) );
  AND2_X1 U12957 ( .A1(n11794), .A2(n11795), .ZN(n11982) );
  NAND2_X1 U12958 ( .A1(n11791), .A2(n11982), .ZN(n10650) );
  NAND2_X1 U12959 ( .A1(n13817), .A2(n14240), .ZN(n10297) );
  OAI211_X1 U12960 ( .C1(n13894), .C2(n13864), .A(n10298), .B(n10297), .ZN(
        P1_U3232) );
  NOR2_X1 U12961 ( .A1(n14596), .A2(n13881), .ZN(P1_U3085) );
  INV_X1 U12962 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10301) );
  OR2_X1 U12963 ( .A1(n10299), .A2(n14942), .ZN(n10300) );
  OAI21_X1 U12964 ( .B1(n14944), .B2(n10301), .A(n10300), .ZN(P2_U3439) );
  INV_X1 U12965 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U12966 ( .A1(n10303), .A2(n10302), .ZN(n11789) );
  NAND2_X1 U12967 ( .A1(n11796), .A2(n11789), .ZN(n11988) );
  NAND2_X1 U12968 ( .A1(n14672), .A2(n14661), .ZN(n10304) );
  AOI22_X1 U12969 ( .A1(n11988), .A2(n10304), .B1(n14642), .B2(n14248), .ZN(
        n10774) );
  NAND3_X1 U12970 ( .A1(n14240), .A2(n11794), .A3(n11791), .ZN(n10305) );
  NAND2_X1 U12971 ( .A1(n10774), .A2(n10305), .ZN(n14325) );
  NAND2_X1 U12972 ( .A1(n14325), .A2(n14687), .ZN(n10306) );
  OAI21_X1 U12973 ( .B1(n14687), .B2(n10307), .A(n10306), .ZN(P1_U3459) );
  NAND2_X1 U12974 ( .A1(n10317), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n13990) );
  NAND2_X1 U12975 ( .A1(n13991), .A2(n13990), .ZN(n10310) );
  INV_X1 U12976 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10308) );
  MUX2_X1 U12977 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10308), .S(n13988), .Z(
        n10309) );
  NAND2_X1 U12978 ( .A1(n10310), .A2(n10309), .ZN(n13993) );
  NAND2_X1 U12979 ( .A1(n13988), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10311) );
  AND2_X1 U12980 ( .A1(n13993), .A2(n10311), .ZN(n10313) );
  INV_X1 U12981 ( .A(n10313), .ZN(n10315) );
  INV_X1 U12982 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10390) );
  MUX2_X1 U12983 ( .A(n10390), .B(P1_REG2_REG_12__SCAN_IN), .S(n10325), .Z(
        n10314) );
  MUX2_X1 U12984 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10390), .S(n10325), .Z(
        n10312) );
  AND2_X1 U12985 ( .A1(n10313), .A2(n10312), .ZN(n10388) );
  AOI21_X1 U12986 ( .B1(n10315), .B2(n10314), .A(n10388), .ZN(n10328) );
  INV_X1 U12987 ( .A(n14628), .ZN(n14616) );
  AOI21_X1 U12988 ( .B1(n10317), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10316), 
        .ZN(n13982) );
  INV_X1 U12989 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14535) );
  MUX2_X1 U12990 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14535), .S(n13988), .Z(
        n13983) );
  NAND2_X1 U12991 ( .A1(n13982), .A2(n13983), .ZN(n13981) );
  NAND2_X1 U12992 ( .A1(n10318), .A2(n14535), .ZN(n10320) );
  INV_X1 U12993 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10319) );
  MUX2_X1 U12994 ( .A(n10319), .B(P1_REG1_REG_12__SCAN_IN), .S(n10325), .Z(
        n10321) );
  AOI21_X1 U12995 ( .B1(n13981), .B2(n10320), .A(n10321), .ZN(n10380) );
  AND3_X1 U12996 ( .A1(n13981), .A2(n10321), .A3(n10320), .ZN(n10322) );
  OAI21_X1 U12997 ( .B1(n10380), .B2(n10322), .A(n14600), .ZN(n10327) );
  INV_X1 U12998 ( .A(n14618), .ZN(n14634) );
  NAND2_X1 U12999 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n13755)
         );
  OAI21_X1 U13000 ( .B1(n14637), .B2(n10323), .A(n13755), .ZN(n10324) );
  AOI21_X1 U13001 ( .B1(n10325), .B2(n14634), .A(n10324), .ZN(n10326) );
  OAI211_X1 U13002 ( .C1(n10328), .C2(n14616), .A(n10327), .B(n10326), .ZN(
        P1_U3255) );
  OAI222_X1 U13003 ( .A1(P3_U3151), .A2(n12105), .B1(n13004), .B2(n10330), 
        .C1(n12387), .C2(n10329), .ZN(P3_U3276) );
  NAND3_X1 U13004 ( .A1(n10333), .A2(n10332), .A3(n10331), .ZN(n10343) );
  INV_X1 U13005 ( .A(n14887), .ZN(n14889) );
  AND2_X1 U13006 ( .A1(n13122), .A2(n13521), .ZN(n13136) );
  INV_X1 U13007 ( .A(n13157), .ZN(n10339) );
  INV_X1 U13008 ( .A(n10335), .ZN(n10336) );
  NAND2_X1 U13009 ( .A1(n14927), .A2(n10336), .ZN(n10337) );
  OAI22_X1 U13010 ( .A1(n10339), .A2(n13132), .B1(n14462), .B2(n10338), .ZN(
        n10341) );
  NAND2_X1 U13011 ( .A1(n10340), .A2(n10602), .ZN(n10355) );
  NAND2_X1 U13012 ( .A1(n10341), .A2(n10355), .ZN(n10351) );
  NAND2_X1 U13013 ( .A1(n10343), .A2(n10342), .ZN(n10347) );
  AND2_X1 U13014 ( .A1(n10345), .A2(n10344), .ZN(n10346) );
  NAND2_X1 U13015 ( .A1(n10347), .A2(n10346), .ZN(n10374) );
  NOR2_X1 U13016 ( .A1(n10374), .A2(P2_U3088), .ZN(n10583) );
  INV_X1 U13017 ( .A(n10583), .ZN(n13019) );
  OR2_X1 U13018 ( .A1(n10348), .A2(n11012), .ZN(n10427) );
  OAI21_X2 U13019 ( .B1(n10349), .B2(n10427), .A(n13466), .ZN(n14467) );
  AOI22_X1 U13020 ( .A1(n13019), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n10354), 
        .B2(n14467), .ZN(n10350) );
  OAI211_X1 U13021 ( .C1(n8193), .C2(n14458), .A(n10351), .B(n10350), .ZN(
        P2_U3204) );
  INV_X1 U13022 ( .A(n11730), .ZN(n11742) );
  NOR2_X1 U13023 ( .A1(n8193), .A2(n13510), .ZN(n10358) );
  OR2_X1 U13024 ( .A1(n11708), .A2(n10354), .ZN(n10356) );
  AND2_X1 U13025 ( .A1(n10356), .A2(n10355), .ZN(n13021) );
  NAND2_X1 U13026 ( .A1(n13020), .A2(n13021), .ZN(n10585) );
  INV_X1 U13027 ( .A(n10358), .ZN(n10359) );
  NAND2_X1 U13028 ( .A1(n6468), .A2(n10359), .ZN(n10360) );
  NAND2_X1 U13029 ( .A1(n10585), .A2(n10360), .ZN(n10361) );
  INV_X2 U13030 ( .A(n11730), .ZN(n10851) );
  XNOR2_X1 U13031 ( .A(n10851), .B(n10591), .ZN(n10364) );
  NAND2_X1 U13032 ( .A1(n13470), .A2(n13155), .ZN(n10362) );
  XNOR2_X1 U13033 ( .A(n10364), .B(n10362), .ZN(n10586) );
  NAND2_X1 U13034 ( .A1(n10361), .A2(n10586), .ZN(n10593) );
  INV_X1 U13035 ( .A(n10362), .ZN(n10363) );
  OR2_X1 U13036 ( .A1(n10364), .A2(n10363), .ZN(n10365) );
  XNOR2_X1 U13037 ( .A(n10491), .B(n10851), .ZN(n10366) );
  BUF_X1 U13038 ( .A(n10602), .Z(n10857) );
  AND2_X1 U13039 ( .A1(n10857), .A2(n13154), .ZN(n10367) );
  NAND2_X1 U13040 ( .A1(n10366), .A2(n10367), .ZN(n10402) );
  INV_X1 U13041 ( .A(n10366), .ZN(n13077) );
  INV_X1 U13042 ( .A(n10367), .ZN(n10368) );
  NAND2_X1 U13043 ( .A1(n13077), .A2(n10368), .ZN(n10369) );
  NAND2_X1 U13044 ( .A1(n10402), .A2(n10369), .ZN(n10372) );
  INV_X1 U13045 ( .A(n13071), .ZN(n10371) );
  AOI211_X1 U13046 ( .C1(n10373), .C2(n10372), .A(n14462), .B(n10371), .ZN(
        n10379) );
  AND2_X1 U13047 ( .A1(n13122), .A2(n13523), .ZN(n13135) );
  AOI22_X1 U13048 ( .A1(n13136), .A2(n13153), .B1(n13135), .B2(n13155), .ZN(
        n10376) );
  INV_X1 U13049 ( .A(n14470), .ZN(n13098) );
  AOI22_X1 U13050 ( .A1(n13098), .A2(n10490), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10375) );
  OAI211_X1 U13051 ( .C1(n10377), .C2(n13139), .A(n10376), .B(n10375), .ZN(
        n10378) );
  OR2_X1 U13052 ( .A1(n10379), .A2(n10378), .ZN(P2_U3190) );
  MUX2_X1 U13053 ( .A(n14519), .B(P1_REG1_REG_14__SCAN_IN), .S(n10383), .Z(
        n10382) );
  INV_X1 U13054 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14529) );
  AOI21_X1 U13055 ( .B1(n10319), .B2(n10389), .A(n10380), .ZN(n14603) );
  MUX2_X1 U13056 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14529), .S(n10385), .Z(
        n14602) );
  NAND2_X1 U13057 ( .A1(n14603), .A2(n14602), .ZN(n14601) );
  OAI21_X1 U13058 ( .B1(n14529), .B2(n14598), .A(n14601), .ZN(n10381) );
  NOR2_X1 U13059 ( .A1(n10381), .A2(n10382), .ZN(n10967) );
  AOI21_X1 U13060 ( .B1(n10382), .B2(n10381), .A(n10967), .ZN(n10399) );
  INV_X1 U13061 ( .A(n10383), .ZN(n10968) );
  INV_X1 U13062 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10384) );
  MUX2_X1 U13063 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10384), .S(n10383), .Z(
        n10393) );
  NAND2_X1 U13064 ( .A1(n10385), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10391) );
  INV_X1 U13065 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10386) );
  MUX2_X1 U13066 ( .A(n10386), .B(P1_REG2_REG_13__SCAN_IN), .S(n10385), .Z(
        n10387) );
  INV_X1 U13067 ( .A(n10387), .ZN(n14606) );
  AOI21_X1 U13068 ( .B1(n10390), .B2(n10389), .A(n10388), .ZN(n14605) );
  NAND2_X1 U13069 ( .A1(n14606), .A2(n14605), .ZN(n14604) );
  NAND2_X1 U13070 ( .A1(n10391), .A2(n14604), .ZN(n10392) );
  NAND2_X1 U13071 ( .A1(n10393), .A2(n10392), .ZN(n10961) );
  OAI211_X1 U13072 ( .C1(n10393), .C2(n10392), .A(n14628), .B(n10961), .ZN(
        n10396) );
  NAND2_X1 U13073 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13706)
         );
  INV_X1 U13074 ( .A(n13706), .ZN(n10394) );
  AOI21_X1 U13075 ( .B1(n14596), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n10394), 
        .ZN(n10395) );
  OAI211_X1 U13076 ( .C1(n14618), .C2(n10968), .A(n10396), .B(n10395), .ZN(
        n10397) );
  INV_X1 U13077 ( .A(n10397), .ZN(n10398) );
  OAI21_X1 U13078 ( .B1(n10399), .B2(n14626), .A(n10398), .ZN(P1_U3257) );
  INV_X1 U13079 ( .A(n10400), .ZN(n10423) );
  INV_X1 U13080 ( .A(n13172), .ZN(n14856) );
  OAI222_X1 U13081 ( .A1(n13685), .A2(n10423), .B1(n14856), .B2(P2_U3088), 
        .C1(n10401), .C2(n13688), .ZN(P2_U3311) );
  NAND2_X1 U13082 ( .A1(n13470), .A2(n13153), .ZN(n10403) );
  INV_X1 U13083 ( .A(n10408), .ZN(n10404) );
  NAND2_X1 U13084 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  XNOR2_X1 U13085 ( .A(n14904), .B(n10851), .ZN(n10530) );
  NAND2_X1 U13086 ( .A1(n13470), .A2(n13524), .ZN(n10531) );
  XNOR2_X1 U13087 ( .A(n10530), .B(n10531), .ZN(n10407) );
  INV_X1 U13088 ( .A(n10407), .ZN(n10411) );
  NAND2_X1 U13089 ( .A1(n10408), .A2(n13126), .ZN(n10409) );
  OAI21_X1 U13090 ( .B1(n13132), .B2(n10478), .A(n10409), .ZN(n10410) );
  NAND3_X1 U13091 ( .A1(n13070), .A2(n10411), .A3(n10410), .ZN(n10418) );
  INV_X1 U13092 ( .A(n10474), .ZN(n10413) );
  OAI22_X1 U13093 ( .A1(n14470), .A2(n10413), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10412), .ZN(n10414) );
  INV_X1 U13094 ( .A(n10414), .ZN(n10417) );
  AOI22_X1 U13095 ( .A1(n13136), .A2(n13152), .B1(n13135), .B2(n13153), .ZN(
        n10416) );
  NAND2_X1 U13096 ( .A1(n14467), .A2(n14904), .ZN(n10415) );
  AND4_X1 U13097 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10419) );
  OAI21_X1 U13098 ( .B1(n10534), .B2(n14462), .A(n10419), .ZN(P2_U3199) );
  INV_X1 U13099 ( .A(n10420), .ZN(n10448) );
  INV_X1 U13100 ( .A(n14822), .ZN(n13202) );
  OAI222_X1 U13101 ( .A1(n13685), .A2(n10448), .B1(n13202), .B2(P2_U3088), 
        .C1(n10421), .C2(n13688), .ZN(P2_U3313) );
  INV_X1 U13102 ( .A(n10973), .ZN(n11227) );
  OAI222_X1 U13103 ( .A1(P1_U3086), .A2(n11227), .B1(n14366), .B2(n10423), 
        .C1(n10422), .C2(n14363), .ZN(P1_U3339) );
  OAI21_X1 U13104 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(n14897) );
  INV_X1 U13105 ( .A(n14897), .ZN(n10444) );
  INV_X1 U13106 ( .A(n10427), .ZN(n10428) );
  INV_X1 U13107 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10582) );
  OAI22_X1 U13108 ( .A1(n13527), .A2(n10429), .B1(n10582), .B2(n13466), .ZN(
        n10435) );
  INV_X1 U13109 ( .A(n10430), .ZN(n10433) );
  INV_X1 U13110 ( .A(n10431), .ZN(n10432) );
  OAI211_X1 U13111 ( .C1(n8191), .C2(n10433), .A(n10432), .B(n13510), .ZN(
        n14894) );
  NOR2_X1 U13112 ( .A1(n13515), .A2(n14894), .ZN(n10434) );
  AOI211_X1 U13113 ( .C1(n13530), .C2(n10591), .A(n10435), .B(n10434), .ZN(
        n10443) );
  OAI21_X1 U13114 ( .B1(n10438), .B2(n10437), .A(n10436), .ZN(n10440) );
  OAI22_X1 U13115 ( .A1(n10476), .A2(n13503), .B1(n8193), .B2(n13505), .ZN(
        n10439) );
  AOI21_X1 U13116 ( .B1(n10440), .B2(n13526), .A(n10439), .ZN(n10441) );
  OAI21_X1 U13117 ( .B1(n10444), .B2(n10353), .A(n10441), .ZN(n14895) );
  NAND2_X1 U13118 ( .A1(n14895), .A2(n13527), .ZN(n10442) );
  OAI211_X1 U13119 ( .C1(n10444), .C2(n10767), .A(n10443), .B(n10442), .ZN(
        P2_U3263) );
  INV_X1 U13120 ( .A(n10445), .ZN(n10450) );
  OAI222_X1 U13121 ( .A1(n13685), .A2(n10450), .B1(n14865), .B2(P2_U3088), 
        .C1(n10446), .C2(n13688), .ZN(P2_U3310) );
  OAI222_X1 U13122 ( .A1(P1_U3086), .A2(n10968), .B1(n14366), .B2(n10448), 
        .C1(n10447), .C2(n14363), .ZN(P1_U3341) );
  OAI222_X1 U13123 ( .A1(P1_U3086), .A2(n13998), .B1(n14366), .B2(n10450), 
        .C1(n10449), .C2(n14363), .ZN(P1_U3338) );
  INV_X1 U13124 ( .A(n10451), .ZN(n10454) );
  INV_X1 U13125 ( .A(n13203), .ZN(n14834) );
  OAI222_X1 U13126 ( .A1(n13685), .A2(n10454), .B1(n14834), .B2(P2_U3088), 
        .C1(n10452), .C2(n13688), .ZN(P2_U3312) );
  INV_X1 U13127 ( .A(n10969), .ZN(n14617) );
  OAI222_X1 U13128 ( .A1(P1_U3086), .A2(n14617), .B1(n14366), .B2(n10454), 
        .C1(n10453), .C2(n14363), .ZN(P1_U3340) );
  AOI22_X1 U13129 ( .A1(n12372), .A2(n8319), .B1(n11584), .B2(n11809), .ZN(
        n10562) );
  AOI22_X1 U13130 ( .A1(n8319), .A2(n11584), .B1(n12360), .B2(n11809), .ZN(
        n10455) );
  XNOR2_X1 U13131 ( .A(n10455), .B(n12370), .ZN(n10563) );
  XOR2_X1 U13132 ( .A(n10562), .B(n10563), .Z(n10564) );
  AOI22_X1 U13133 ( .A1(n14248), .A2(n11584), .B1(n12360), .B2(n14641), .ZN(
        n10456) );
  XNOR2_X1 U13134 ( .A(n10456), .B(n12370), .ZN(n10461) );
  XNOR2_X1 U13135 ( .A(n10461), .B(n10457), .ZN(n13736) );
  MUX2_X1 U13136 ( .A(n12370), .B(n10459), .S(n10458), .Z(n13735) );
  NAND2_X1 U13137 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  NAND2_X1 U13138 ( .A1(n13734), .A2(n10462), .ZN(n10565) );
  XOR2_X1 U13139 ( .A(n10564), .B(n10565), .Z(n10468) );
  NOR2_X1 U13140 ( .A1(n13858), .A2(n10653), .ZN(n10466) );
  NOR2_X2 U13141 ( .A1(n13847), .A2(n14520), .ZN(n13855) );
  INV_X1 U13142 ( .A(n13855), .ZN(n13828) );
  OAI22_X1 U13143 ( .A1(n10464), .A2(n13857), .B1(n13828), .B2(n10463), .ZN(
        n10465) );
  AOI211_X1 U13144 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n13738), .A(n10466), .B(
        n10465), .ZN(n10467) );
  OAI21_X1 U13145 ( .B1(n10468), .B2(n13864), .A(n10467), .ZN(P1_U3237) );
  OR2_X1 U13146 ( .A1(n10491), .A2(n13154), .ZN(n10469) );
  NAND2_X1 U13147 ( .A1(n10470), .A2(n10469), .ZN(n10502) );
  NAND2_X1 U13148 ( .A1(n10502), .A2(n10508), .ZN(n10501) );
  NAND2_X1 U13149 ( .A1(n10501), .A2(n10471), .ZN(n10595) );
  XNOR2_X1 U13150 ( .A(n10595), .B(n10479), .ZN(n10486) );
  INV_X1 U13151 ( .A(n10486), .ZN(n14909) );
  NAND2_X1 U13152 ( .A1(n14904), .A2(n10504), .ZN(n10472) );
  NAND2_X1 U13153 ( .A1(n10472), .A2(n13510), .ZN(n10473) );
  OR2_X1 U13154 ( .A1(n13535), .A2(n10473), .ZN(n14905) );
  AOI22_X1 U13155 ( .A1(n13530), .A2(n14904), .B1(n10474), .B2(n13529), .ZN(
        n10475) );
  OAI21_X1 U13156 ( .B1(n14905), .B2(n13515), .A(n10475), .ZN(n10488) );
  AOI22_X1 U13157 ( .A1(n13521), .A2(n13152), .B1(n13153), .B2(n13523), .ZN(
        n10485) );
  NAND2_X1 U13158 ( .A1(n10491), .A2(n10476), .ZN(n10507) );
  INV_X1 U13159 ( .A(n10508), .ZN(n10477) );
  NAND2_X1 U13160 ( .A1(n13076), .A2(n10478), .ZN(n10480) );
  INV_X1 U13161 ( .A(n10605), .ZN(n10483) );
  AND3_X1 U13162 ( .A1(n10511), .A2(n10481), .A3(n10480), .ZN(n10482) );
  OAI21_X1 U13163 ( .B1(n10483), .B2(n10482), .A(n13526), .ZN(n10484) );
  OAI211_X1 U13164 ( .C1(n10486), .C2(n10353), .A(n10485), .B(n10484), .ZN(
        n14907) );
  MUX2_X1 U13165 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n14907), .S(n13527), .Z(
        n10487) );
  AOI211_X1 U13166 ( .C1(n10741), .C2(n14909), .A(n10488), .B(n10487), .ZN(
        n10489) );
  INV_X1 U13167 ( .A(n10489), .ZN(P2_U3260) );
  AOI22_X1 U13168 ( .A1(n13530), .A2(n10491), .B1(n13529), .B2(n10490), .ZN(
        n10492) );
  OAI21_X1 U13169 ( .B1(n13515), .B2(n10493), .A(n10492), .ZN(n10496) );
  MUX2_X1 U13170 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10494), .S(n13527), .Z(
        n10495) );
  AOI211_X1 U13171 ( .C1(n10741), .C2(n10497), .A(n10496), .B(n10495), .ZN(
        n10498) );
  INV_X1 U13172 ( .A(n10498), .ZN(P2_U3262) );
  NAND2_X1 U13173 ( .A1(n10499), .A2(n10353), .ZN(n10500) );
  OAI21_X1 U13174 ( .B1(n10502), .B2(n10508), .A(n10501), .ZN(n14902) );
  OAI211_X1 U13175 ( .C1(n6980), .C2(n6979), .A(n13510), .B(n10504), .ZN(
        n14899) );
  AOI22_X1 U13176 ( .A1(n13530), .A2(n13076), .B1(n13529), .B2(n10505), .ZN(
        n10506) );
  OAI21_X1 U13177 ( .B1(n14899), .B2(n13515), .A(n10506), .ZN(n10516) );
  NAND3_X1 U13178 ( .A1(n10509), .A2(n10508), .A3(n10507), .ZN(n10510) );
  NAND2_X1 U13179 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  NAND2_X1 U13180 ( .A1(n10512), .A2(n13526), .ZN(n10514) );
  AOI22_X1 U13181 ( .A1(n13521), .A2(n13524), .B1(n13154), .B2(n13523), .ZN(
        n10513) );
  NAND2_X1 U13182 ( .A1(n10514), .A2(n10513), .ZN(n14900) );
  MUX2_X1 U13183 ( .A(n14900), .B(P2_REG2_REG_4__SCAN_IN), .S(n13512), .Z(
        n10515) );
  AOI211_X1 U13184 ( .C1(n13534), .C2(n14902), .A(n10516), .B(n10515), .ZN(
        n10517) );
  INV_X1 U13185 ( .A(n10517), .ZN(P2_U3261) );
  XNOR2_X1 U13186 ( .A(n11801), .B(n10518), .ZN(n10523) );
  XNOR2_X1 U13187 ( .A(n11990), .B(n10519), .ZN(n10520) );
  NAND2_X1 U13188 ( .A1(n10520), .A2(n14684), .ZN(n10522) );
  AOI22_X1 U13189 ( .A1(n14498), .A2(n14248), .B1(n13885), .B2(n14642), .ZN(
        n10521) );
  OAI211_X1 U13190 ( .C1(n14661), .C2(n10523), .A(n10522), .B(n10521), .ZN(
        n10648) );
  OAI211_X1 U13191 ( .C1(n14242), .C2(n10653), .A(n14302), .B(n10553), .ZN(
        n10657) );
  INV_X1 U13192 ( .A(n10657), .ZN(n10524) );
  NOR2_X1 U13193 ( .A1(n10648), .A2(n10524), .ZN(n10529) );
  INV_X1 U13194 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10525) );
  OAI22_X1 U13195 ( .A1(n14348), .A2(n10653), .B1(n14687), .B2(n10525), .ZN(
        n10526) );
  INV_X1 U13196 ( .A(n10526), .ZN(n10527) );
  OAI21_X1 U13197 ( .B1(n10529), .B2(n14685), .A(n10527), .ZN(P1_U3465) );
  AOI22_X1 U13198 ( .A1(n9824), .A2(n11809), .B1(n14695), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n10528) );
  OAI21_X1 U13199 ( .B1(n10529), .B2(n14695), .A(n10528), .ZN(P1_U3530) );
  INV_X1 U13200 ( .A(n14912), .ZN(n13536) );
  INV_X1 U13201 ( .A(n10530), .ZN(n10532) );
  NAND2_X1 U13202 ( .A1(n10532), .A2(n10531), .ZN(n10533) );
  XNOR2_X1 U13203 ( .A(n14912), .B(n10851), .ZN(n10535) );
  AND2_X1 U13204 ( .A1(n10857), .A2(n13152), .ZN(n10536) );
  NAND2_X1 U13205 ( .A1(n10535), .A2(n10536), .ZN(n10665) );
  INV_X1 U13206 ( .A(n10535), .ZN(n10664) );
  INV_X1 U13207 ( .A(n10536), .ZN(n10537) );
  NAND2_X1 U13208 ( .A1(n10664), .A2(n10537), .ZN(n10538) );
  NAND2_X1 U13209 ( .A1(n10665), .A2(n10538), .ZN(n10540) );
  AOI21_X1 U13210 ( .B1(n10539), .B2(n10540), .A(n14462), .ZN(n10542) );
  NAND2_X1 U13211 ( .A1(n10542), .A2(n10666), .ZN(n10547) );
  NAND2_X1 U13212 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14745) );
  INV_X1 U13213 ( .A(n14745), .ZN(n10545) );
  INV_X1 U13214 ( .A(n13522), .ZN(n12062) );
  INV_X1 U13215 ( .A(n13135), .ZN(n14457) );
  OAI22_X1 U13216 ( .A1(n12062), .A2(n14458), .B1(n14457), .B2(n10543), .ZN(
        n10544) );
  AOI211_X1 U13217 ( .C1(n13528), .C2(n13098), .A(n10545), .B(n10544), .ZN(
        n10546) );
  OAI211_X1 U13218 ( .C1(n13536), .C2(n13139), .A(n10547), .B(n10546), .ZN(
        P2_U3211) );
  XNOR2_X1 U13219 ( .A(n10548), .B(n11989), .ZN(n10549) );
  NAND2_X1 U13220 ( .A1(n10549), .A2(n14684), .ZN(n10551) );
  AOI22_X1 U13221 ( .A1(n14498), .A2(n8319), .B1(n13884), .B2(n14642), .ZN(
        n10550) );
  OAI211_X1 U13222 ( .C1(n14661), .C2(n10552), .A(n10551), .B(n10550), .ZN(
        n10712) );
  AOI21_X1 U13223 ( .B1(n10553), .B2(n10714), .A(n14644), .ZN(n10554) );
  NAND2_X1 U13224 ( .A1(n10554), .A2(n10745), .ZN(n10717) );
  INV_X1 U13225 ( .A(n10717), .ZN(n10555) );
  NOR2_X1 U13226 ( .A1(n10712), .A2(n10555), .ZN(n10561) );
  AOI22_X1 U13227 ( .A1(n9824), .A2(n10714), .B1(n14695), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n10556) );
  OAI21_X1 U13228 ( .B1(n10561), .B2(n14695), .A(n10556), .ZN(P1_U3531) );
  INV_X1 U13229 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10557) );
  OAI22_X1 U13230 ( .A1(n14348), .A2(n10558), .B1(n14687), .B2(n10557), .ZN(
        n10559) );
  INV_X1 U13231 ( .A(n10559), .ZN(n10560) );
  OAI21_X1 U13232 ( .B1(n10561), .B2(n14685), .A(n10560), .ZN(P1_U3468) );
  AOI22_X1 U13233 ( .A1(n10565), .A2(n10564), .B1(n10563), .B2(n10562), .ZN(
        n10568) );
  AOI22_X1 U13234 ( .A1(n12364), .A2(n13885), .B1(n11584), .B2(n10714), .ZN(
        n10933) );
  AOI22_X1 U13235 ( .A1(n13885), .A2(n11584), .B1(n12360), .B2(n10714), .ZN(
        n10566) );
  XNOR2_X1 U13236 ( .A(n10566), .B(n12370), .ZN(n10932) );
  XOR2_X1 U13237 ( .A(n10933), .B(n10932), .Z(n10567) );
  NAND2_X1 U13238 ( .A1(n10568), .A2(n10567), .ZN(n10937) );
  OAI211_X1 U13239 ( .C1(n10568), .C2(n10567), .A(n10937), .B(n13844), .ZN(
        n10576) );
  OR2_X1 U13240 ( .A1(n10570), .A2(n10569), .ZN(n10571) );
  NAND2_X1 U13241 ( .A1(n10571), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13786) );
  INV_X1 U13242 ( .A(n13786), .ZN(n13862) );
  MUX2_X1 U13243 ( .A(n13862), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10574) );
  OAI22_X1 U13244 ( .A1(n10572), .A2(n13857), .B1(n13828), .B2(n11808), .ZN(
        n10573) );
  AOI211_X1 U13245 ( .C1(n10714), .C2(n13817), .A(n10574), .B(n10573), .ZN(
        n10575) );
  NAND2_X1 U13246 ( .A1(n10576), .A2(n10575), .ZN(P1_U3218) );
  OAI222_X1 U13247 ( .A1(P3_U3151), .A2(n10579), .B1(n13004), .B2(n10578), 
        .C1(n12387), .C2(n10577), .ZN(P3_U3275) );
  NAND2_X1 U13248 ( .A1(n13136), .A2(n13154), .ZN(n10581) );
  NAND2_X1 U13249 ( .A1(n13135), .A2(n13156), .ZN(n10580) );
  OAI211_X1 U13250 ( .C1(n10583), .C2(n10582), .A(n10581), .B(n10580), .ZN(
        n10590) );
  INV_X1 U13251 ( .A(n13132), .ZN(n13097) );
  INV_X1 U13252 ( .A(n6468), .ZN(n10584) );
  AOI22_X1 U13253 ( .A1(n13097), .A2(n13156), .B1(n13126), .B2(n10584), .ZN(
        n10588) );
  INV_X1 U13254 ( .A(n10585), .ZN(n10587) );
  NOR3_X1 U13255 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(n10589) );
  AOI211_X1 U13256 ( .C1(n10591), .C2(n14467), .A(n10590), .B(n10589), .ZN(
        n10592) );
  OAI21_X1 U13257 ( .B1(n14462), .B2(n10593), .A(n10592), .ZN(P2_U3209) );
  INV_X1 U13258 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10615) );
  NAND2_X1 U13259 ( .A1(n14904), .A2(n13524), .ZN(n10594) );
  OR2_X1 U13260 ( .A1(n14904), .A2(n13524), .ZN(n10596) );
  NAND2_X1 U13261 ( .A1(n14912), .A2(n13152), .ZN(n10598) );
  NAND2_X1 U13262 ( .A1(n13531), .A2(n10598), .ZN(n10631) );
  OR2_X1 U13263 ( .A1(n14919), .A2(n13522), .ZN(n10599) );
  NAND2_X1 U13264 ( .A1(n10631), .A2(n10599), .ZN(n10601) );
  NAND2_X1 U13265 ( .A1(n14919), .A2(n13522), .ZN(n10600) );
  NAND2_X1 U13266 ( .A1(n10601), .A2(n10600), .ZN(n10724) );
  INV_X1 U13267 ( .A(n10729), .ZN(n10723) );
  XNOR2_X1 U13268 ( .A(n10724), .B(n10723), .ZN(n10691) );
  NAND2_X1 U13269 ( .A1(n13536), .A2(n13535), .ZN(n10637) );
  INV_X1 U13270 ( .A(n10764), .ZN(n10603) );
  AOI211_X1 U13271 ( .C1(n12070), .C2(n10636), .A(n10602), .B(n10603), .ZN(
        n10694) );
  AOI21_X1 U13272 ( .B1(n14936), .B2(n12070), .A(n10694), .ZN(n10613) );
  NAND2_X1 U13273 ( .A1(n10605), .A2(n10604), .ZN(n13520) );
  NAND2_X1 U13274 ( .A1(n13520), .A2(n13533), .ZN(n13519) );
  INV_X1 U13275 ( .A(n13152), .ZN(n10663) );
  NAND2_X1 U13276 ( .A1(n14912), .A2(n10663), .ZN(n10606) );
  OR2_X1 U13277 ( .A1(n14919), .A2(n12062), .ZN(n10607) );
  NAND2_X1 U13278 ( .A1(n10633), .A2(n10607), .ZN(n10609) );
  NAND2_X1 U13279 ( .A1(n14919), .A2(n12062), .ZN(n10608) );
  NAND2_X1 U13280 ( .A1(n10609), .A2(n10608), .ZN(n10730) );
  XNOR2_X1 U13281 ( .A(n10730), .B(n10729), .ZN(n10612) );
  NAND2_X1 U13282 ( .A1(n13149), .A2(n13521), .ZN(n10611) );
  NAND2_X1 U13283 ( .A1(n13522), .A2(n13523), .ZN(n10610) );
  NAND2_X1 U13284 ( .A1(n10611), .A2(n10610), .ZN(n12058) );
  AOI21_X1 U13285 ( .B1(n10612), .B2(n13526), .A(n12058), .ZN(n10696) );
  OAI211_X1 U13286 ( .C1(n14922), .C2(n10691), .A(n10613), .B(n10696), .ZN(
        n10616) );
  NAND2_X1 U13287 ( .A1(n10616), .A2(n14944), .ZN(n10614) );
  OAI21_X1 U13288 ( .B1(n14944), .B2(n10615), .A(n10614), .ZN(P2_U3454) );
  INV_X1 U13289 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n13193) );
  NAND2_X1 U13290 ( .A1(n10616), .A2(n14960), .ZN(n10617) );
  OAI21_X1 U13291 ( .B1(n14960), .B2(n13193), .A(n10617), .ZN(P2_U3507) );
  NAND2_X1 U13292 ( .A1(n14985), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10814) );
  INV_X1 U13293 ( .A(n10814), .ZN(n10786) );
  AND2_X1 U13294 ( .A1(n8879), .A2(n12573), .ZN(n10679) );
  AOI22_X1 U13295 ( .A1(n10679), .A2(n14982), .B1(n10618), .B2(n12577), .ZN(
        n10621) );
  NOR2_X1 U13296 ( .A1(n12608), .A2(n10618), .ZN(n12136) );
  INV_X1 U13297 ( .A(n12136), .ZN(n10619) );
  NAND2_X1 U13298 ( .A1(n10777), .A2(n10619), .ZN(n12111) );
  NAND2_X1 U13299 ( .A1(n12111), .A2(n14974), .ZN(n10620) );
  OAI211_X1 U13300 ( .C1(n10786), .C2(n14993), .A(n10621), .B(n10620), .ZN(
        P3_U3172) );
  INV_X1 U13301 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10622) );
  OAI22_X1 U13302 ( .A1(n13489), .A2(n10623), .B1(n10622), .B2(n13466), .ZN(
        n10624) );
  AOI21_X1 U13303 ( .B1(n13538), .B2(n10625), .A(n10624), .ZN(n10629) );
  MUX2_X1 U13304 ( .A(n10627), .B(n10626), .S(n13527), .Z(n10628) );
  OAI211_X1 U13305 ( .C1(n13475), .C2(n10630), .A(n10629), .B(n10628), .ZN(
        P2_U3264) );
  XOR2_X1 U13306 ( .A(n10632), .B(n10631), .Z(n14923) );
  XNOR2_X1 U13307 ( .A(n10633), .B(n10632), .ZN(n10635) );
  AOI22_X1 U13308 ( .A1(n13521), .A2(n13151), .B1(n13152), .B2(n13523), .ZN(
        n10672) );
  INV_X1 U13309 ( .A(n10672), .ZN(n10634) );
  AOI21_X1 U13310 ( .B1(n10635), .B2(n13526), .A(n10634), .ZN(n14921) );
  MUX2_X1 U13311 ( .A(n10019), .B(n14921), .S(n13527), .Z(n10641) );
  AOI211_X1 U13312 ( .C1(n14919), .C2(n10637), .A(n10602), .B(n6984), .ZN(
        n14918) );
  INV_X1 U13313 ( .A(n14919), .ZN(n10677) );
  INV_X1 U13314 ( .A(n10674), .ZN(n10638) );
  OAI22_X1 U13315 ( .A1(n10677), .A2(n13489), .B1(n10638), .B2(n13466), .ZN(
        n10639) );
  AOI21_X1 U13316 ( .B1(n14918), .B2(n13538), .A(n10639), .ZN(n10640) );
  OAI211_X1 U13317 ( .C1(n14923), .C2(n13475), .A(n10641), .B(n10640), .ZN(
        P2_U3258) );
  AND2_X1 U13318 ( .A1(n10643), .A2(n10642), .ZN(n10646) );
  INV_X1 U13319 ( .A(n10644), .ZN(n10645) );
  INV_X1 U13320 ( .A(n10647), .ZN(n12311) );
  MUX2_X1 U13321 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10648), .S(n14253), .Z(
        n10649) );
  INV_X1 U13322 ( .A(n10649), .ZN(n10656) );
  INV_X1 U13323 ( .A(n10650), .ZN(n10651) );
  INV_X1 U13324 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10652) );
  OAI22_X1 U13325 ( .A1(n14196), .A2(n10653), .B1(n14206), .B2(n10652), .ZN(
        n10654) );
  INV_X1 U13326 ( .A(n10654), .ZN(n10655) );
  OAI211_X1 U13327 ( .C1(n14239), .C2(n10657), .A(n10656), .B(n10655), .ZN(
        P1_U3291) );
  XNOR2_X1 U13328 ( .A(n14919), .B(n10851), .ZN(n10658) );
  AND2_X1 U13329 ( .A1(n10857), .A2(n13522), .ZN(n10659) );
  NAND2_X1 U13330 ( .A1(n10658), .A2(n10659), .ZN(n10848) );
  INV_X1 U13331 ( .A(n10658), .ZN(n12063) );
  INV_X1 U13332 ( .A(n10659), .ZN(n10660) );
  NAND2_X1 U13333 ( .A1(n12063), .A2(n10660), .ZN(n10661) );
  AND2_X1 U13334 ( .A1(n10848), .A2(n10661), .ZN(n10667) );
  INV_X1 U13335 ( .A(n10667), .ZN(n10662) );
  AOI21_X1 U13336 ( .B1(n10666), .B2(n10662), .A(n14462), .ZN(n10670) );
  NOR3_X1 U13337 ( .A1(n10664), .A2(n10663), .A3(n13132), .ZN(n10669) );
  NAND2_X1 U13338 ( .A1(n10666), .A2(n10665), .ZN(n10668) );
  NAND2_X2 U13339 ( .A1(n10668), .A2(n10667), .ZN(n12061) );
  OAI21_X1 U13340 ( .B1(n10670), .B2(n10669), .A(n12061), .ZN(n10676) );
  INV_X1 U13341 ( .A(n13122), .ZN(n13101) );
  OAI21_X1 U13342 ( .B1(n13101), .B2(n10672), .A(n10671), .ZN(n10673) );
  AOI21_X1 U13343 ( .B1(n10674), .B2(n13098), .A(n10673), .ZN(n10675) );
  OAI211_X1 U13344 ( .C1(n10677), .C2(n13139), .A(n10676), .B(n10675), .ZN(
        P2_U3185) );
  NOR2_X1 U13345 ( .A1(n10678), .A2(n15167), .ZN(n10680) );
  AOI21_X1 U13346 ( .B1(n12111), .B2(n10680), .A(n10679), .ZN(n10944) );
  AOI22_X1 U13347 ( .A1(n12901), .A2(n10618), .B1(n15203), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n10681) );
  OAI21_X1 U13348 ( .B1(n10944), .B2(n15203), .A(n10681), .ZN(P3_U3459) );
  OAI222_X1 U13349 ( .A1(n12139), .A2(P3_U3151), .B1(n13004), .B2(n10683), 
        .C1(n12387), .C2(n10682), .ZN(P3_U3274) );
  INV_X1 U13350 ( .A(n12985), .ZN(n12998) );
  INV_X1 U13351 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10684) );
  OAI22_X1 U13352 ( .A1(n12998), .A2(n10685), .B1(n10684), .B2(n15193), .ZN(
        n10686) );
  INV_X1 U13353 ( .A(n10686), .ZN(n10687) );
  OAI21_X1 U13354 ( .B1(n15191), .B2(n10944), .A(n10687), .ZN(P3_U3390) );
  NAND2_X1 U13355 ( .A1(n12607), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10688) );
  OAI21_X1 U13356 ( .B1(n12102), .B2(n12607), .A(n10688), .ZN(P3_U3521) );
  AOI22_X1 U13357 ( .A1(n13512), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10689), 
        .B2(n13529), .ZN(n10690) );
  OAI21_X1 U13358 ( .B1(n6983), .B2(n13489), .A(n10690), .ZN(n10693) );
  NOR2_X1 U13359 ( .A1(n10691), .A2(n13475), .ZN(n10692) );
  AOI211_X1 U13360 ( .C1(n10694), .C2(n13538), .A(n10693), .B(n10692), .ZN(
        n10695) );
  OAI21_X1 U13361 ( .B1(n13512), .B2(n10696), .A(n10695), .ZN(P2_U3257) );
  INV_X1 U13362 ( .A(n10697), .ZN(n10699) );
  OAI22_X1 U13363 ( .A1(n12297), .A2(P3_U3151), .B1(SI_22_), .B2(n13004), .ZN(
        n10698) );
  AOI21_X1 U13364 ( .B1(n10699), .B2(n14381), .A(n10698), .ZN(P3_U3273) );
  XNOR2_X1 U13365 ( .A(n10700), .B(n10701), .ZN(n10705) );
  NAND2_X1 U13366 ( .A1(n10702), .A2(n14684), .ZN(n10704) );
  AOI22_X1 U13367 ( .A1(n14498), .A2(n13884), .B1(n13882), .B2(n14642), .ZN(
        n10703) );
  OAI211_X1 U13368 ( .C1(n14661), .C2(n10705), .A(n10704), .B(n10703), .ZN(
        n10892) );
  OAI21_X1 U13369 ( .B1(n10744), .B2(n10891), .A(n14302), .ZN(n10706) );
  NOR2_X1 U13370 ( .A1(n10706), .A2(n10825), .ZN(n10895) );
  NOR2_X1 U13371 ( .A1(n10892), .A2(n10895), .ZN(n10711) );
  AOI22_X1 U13372 ( .A1(n9824), .A2(n11829), .B1(n14695), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n10707) );
  OAI21_X1 U13373 ( .B1(n10711), .B2(n14695), .A(n10707), .ZN(P1_U3533) );
  INV_X1 U13374 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10708) );
  OAI22_X1 U13375 ( .A1(n14348), .A2(n10891), .B1(n14687), .B2(n10708), .ZN(
        n10709) );
  INV_X1 U13376 ( .A(n10709), .ZN(n10710) );
  OAI21_X1 U13377 ( .B1(n10711), .B2(n14685), .A(n10710), .ZN(P1_U3474) );
  INV_X2 U13378 ( .A(n14253), .ZN(n14147) );
  MUX2_X1 U13379 ( .A(n10712), .B(P1_REG2_REG_3__SCAN_IN), .S(n14147), .Z(
        n10713) );
  INV_X1 U13380 ( .A(n10713), .ZN(n10716) );
  AOI22_X1 U13381 ( .A1(n14246), .A2(n10714), .B1(n8322), .B2(n14243), .ZN(
        n10715) );
  OAI211_X1 U13382 ( .C1(n14239), .C2(n10717), .A(n10716), .B(n10715), .ZN(
        P1_U3290) );
  INV_X1 U13383 ( .A(n14633), .ZN(n10720) );
  INV_X1 U13384 ( .A(n10718), .ZN(n10721) );
  OAI222_X1 U13385 ( .A1(n10720), .A2(P1_U3086), .B1(n14366), .B2(n10721), 
        .C1(n10719), .C2(n14363), .ZN(P1_U3337) );
  INV_X1 U13386 ( .A(n13209), .ZN(n14872) );
  OAI222_X1 U13387 ( .A1(n13688), .A2(n10722), .B1(n13685), .B2(n10721), .C1(
        P2_U3088), .C2(n14872), .ZN(P2_U3309) );
  NAND2_X1 U13388 ( .A1(n10724), .A2(n10723), .ZN(n10726) );
  NAND2_X1 U13389 ( .A1(n12070), .A2(n13151), .ZN(n10725) );
  NAND2_X1 U13390 ( .A1(n10726), .A2(n10725), .ZN(n10759) );
  NAND2_X1 U13391 ( .A1(n10759), .A2(n10758), .ZN(n10728) );
  NAND2_X1 U13392 ( .A1(n11703), .A2(n13149), .ZN(n10727) );
  NAND2_X1 U13393 ( .A1(n10728), .A2(n10727), .ZN(n10790) );
  XNOR2_X1 U13394 ( .A(n10790), .B(n10794), .ZN(n10737) );
  NAND2_X1 U13395 ( .A1(n10730), .A2(n10729), .ZN(n10732) );
  INV_X1 U13396 ( .A(n13151), .ZN(n10757) );
  NAND2_X1 U13397 ( .A1(n12070), .A2(n10757), .ZN(n10731) );
  NAND2_X1 U13398 ( .A1(n10732), .A2(n10731), .ZN(n10756) );
  OR2_X1 U13399 ( .A1(n11703), .A2(n10868), .ZN(n10733) );
  XNOR2_X1 U13400 ( .A(n10796), .B(n10794), .ZN(n10735) );
  OAI22_X1 U13401 ( .A1(n11005), .A2(n13503), .B1(n10868), .B2(n13505), .ZN(
        n10734) );
  AOI21_X1 U13402 ( .B1(n10735), .B2(n13526), .A(n10734), .ZN(n10736) );
  OAI21_X1 U13403 ( .B1(n10737), .B2(n10353), .A(n10736), .ZN(n14929) );
  INV_X1 U13404 ( .A(n14929), .ZN(n10743) );
  INV_X1 U13405 ( .A(n10737), .ZN(n14931) );
  OAI211_X1 U13406 ( .C1(n14928), .C2(n10763), .A(n13510), .B(n10802), .ZN(
        n14926) );
  AOI22_X1 U13407 ( .A1(n13512), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10871), 
        .B2(n13529), .ZN(n10739) );
  NAND2_X1 U13408 ( .A1(n10856), .A2(n13530), .ZN(n10738) );
  OAI211_X1 U13409 ( .C1(n14926), .C2(n13515), .A(n10739), .B(n10738), .ZN(
        n10740) );
  AOI21_X1 U13410 ( .B1(n14931), .B2(n10741), .A(n10740), .ZN(n10742) );
  OAI21_X1 U13411 ( .B1(n10743), .B2(n13512), .A(n10742), .ZN(P2_U3255) );
  AOI211_X1 U13412 ( .C1(n14652), .C2(n10745), .A(n14644), .B(n10744), .ZN(
        n14651) );
  XNOR2_X1 U13413 ( .A(n10746), .B(n11991), .ZN(n10747) );
  NAND2_X1 U13414 ( .A1(n10747), .A2(n14676), .ZN(n10751) );
  NAND2_X1 U13415 ( .A1(n13883), .A2(n14642), .ZN(n10749) );
  NAND2_X1 U13416 ( .A1(n13885), .A2(n14498), .ZN(n10748) );
  NAND2_X1 U13417 ( .A1(n10749), .A2(n10748), .ZN(n10928) );
  INV_X1 U13418 ( .A(n10928), .ZN(n10750) );
  NAND2_X1 U13419 ( .A1(n10751), .A2(n10750), .ZN(n14655) );
  AOI21_X1 U13420 ( .B1(n14651), .B2(n6857), .A(n14655), .ZN(n10752) );
  MUX2_X1 U13421 ( .A(n10753), .B(n10752), .S(n14253), .Z(n10755) );
  AOI22_X1 U13422 ( .A1(n14246), .A2(n14652), .B1(n10927), .B2(n14243), .ZN(
        n10754) );
  OAI211_X1 U13423 ( .C1(n14219), .C2(n14654), .A(n10755), .B(n10754), .ZN(
        P1_U3289) );
  XOR2_X1 U13424 ( .A(n10758), .B(n10756), .Z(n10762) );
  OAI22_X1 U13425 ( .A1(n14456), .A2(n13503), .B1(n10757), .B2(n13505), .ZN(
        n10761) );
  XNOR2_X1 U13426 ( .A(n10759), .B(n10758), .ZN(n10900) );
  NOR2_X1 U13427 ( .A1(n10900), .A2(n10353), .ZN(n10760) );
  AOI211_X1 U13428 ( .C1(n13526), .C2(n10762), .A(n10761), .B(n10760), .ZN(
        n10899) );
  AOI211_X1 U13429 ( .C1(n11703), .C2(n10764), .A(n10602), .B(n10763), .ZN(
        n10897) );
  INV_X1 U13430 ( .A(n11703), .ZN(n10766) );
  AOI22_X1 U13431 ( .A1(n13512), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11694), 
        .B2(n13529), .ZN(n10765) );
  OAI21_X1 U13432 ( .B1(n10766), .B2(n13489), .A(n10765), .ZN(n10769) );
  NOR2_X1 U13433 ( .A1(n10900), .A2(n10767), .ZN(n10768) );
  AOI211_X1 U13434 ( .C1(n10897), .C2(n13538), .A(n10769), .B(n10768), .ZN(
        n10770) );
  OAI21_X1 U13435 ( .B1(n10899), .B2(n13512), .A(n10770), .ZN(P2_U3256) );
  NOR2_X1 U13436 ( .A1(n14239), .A2(n14644), .ZN(n14244) );
  OAI21_X1 U13437 ( .B1(n14244), .B2(n14246), .A(n14240), .ZN(n10773) );
  AOI22_X1 U13438 ( .A1(n14147), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14243), .ZN(n10772) );
  OAI211_X1 U13439 ( .C1(n14147), .C2(n10774), .A(n10773), .B(n10772), .ZN(
        P1_U3293) );
  NAND3_X1 U13440 ( .A1(n10775), .A2(n10777), .A3(n10776), .ZN(n10778) );
  OAI211_X1 U13441 ( .C1(n10780), .C2(n15116), .A(n10779), .B(n10778), .ZN(
        n10781) );
  NAND2_X1 U13442 ( .A1(n10781), .A2(n14974), .ZN(n10785) );
  INV_X1 U13443 ( .A(n9672), .ZN(n10782) );
  OAI22_X1 U13444 ( .A1(n10782), .A2(n12550), .B1(n12608), .B2(n12548), .ZN(
        n15131) );
  AOI22_X1 U13445 ( .A1(n15131), .A2(n14982), .B1(n10783), .B2(n12577), .ZN(
        n10784) );
  OAI211_X1 U13446 ( .C1(n10786), .C2(n15120), .A(n10785), .B(n10784), .ZN(
        P3_U3162) );
  OAI222_X1 U13447 ( .A1(P1_U3086), .A2(n6857), .B1(n14366), .B2(n10788), .C1(
        n10787), .C2(n14363), .ZN(P1_U3336) );
  OAI222_X1 U13448 ( .A1(n13688), .A2(n10789), .B1(n13685), .B2(n10788), .C1(
        n13216), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U13449 ( .A1(n10856), .A2(n13148), .ZN(n10791) );
  XNOR2_X1 U13450 ( .A(n10880), .B(n10798), .ZN(n14935) );
  INV_X1 U13451 ( .A(n14935), .ZN(n10810) );
  NOR2_X1 U13452 ( .A1(n10856), .A2(n14456), .ZN(n10795) );
  OAI21_X1 U13453 ( .B1(n10798), .B2(n10797), .A(n10875), .ZN(n10799) );
  NAND2_X1 U13454 ( .A1(n10799), .A2(n13526), .ZN(n10801) );
  AOI22_X1 U13455 ( .A1(n13521), .A2(n13146), .B1(n13148), .B2(n13523), .ZN(
        n10800) );
  NAND2_X1 U13456 ( .A1(n10801), .A2(n10800), .ZN(n14941) );
  INV_X1 U13457 ( .A(n14937), .ZN(n10807) );
  AOI21_X1 U13458 ( .B1(n10802), .B2(n14937), .A(n10602), .ZN(n10803) );
  OR2_X1 U13459 ( .A1(n10802), .A2(n14937), .ZN(n10883) );
  AND2_X1 U13460 ( .A1(n10803), .A2(n10883), .ZN(n14939) );
  NAND2_X1 U13461 ( .A1(n14939), .A2(n13538), .ZN(n10806) );
  AOI22_X1 U13462 ( .A1(n13512), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10804), 
        .B2(n13529), .ZN(n10805) );
  OAI211_X1 U13463 ( .C1(n10807), .C2(n13489), .A(n10806), .B(n10805), .ZN(
        n10808) );
  AOI21_X1 U13464 ( .B1(n14941), .B2(n13527), .A(n10808), .ZN(n10809) );
  OAI21_X1 U13465 ( .B1(n13475), .B2(n10810), .A(n10809), .ZN(P2_U3254) );
  XOR2_X1 U13466 ( .A(n10811), .B(n10812), .Z(n10816) );
  AOI22_X1 U13467 ( .A1(n12572), .A2(n8879), .B1(n12606), .B2(n12573), .ZN(
        n15110) );
  OAI22_X1 U13468 ( .A1(n15110), .A2(n12530), .B1(n14973), .B2(n15106), .ZN(
        n10813) );
  AOI21_X1 U13469 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10814), .A(n10813), .ZN(
        n10815) );
  OAI21_X1 U13470 ( .B1(n10816), .B2(n12579), .A(n10815), .ZN(P3_U3177) );
  XNOR2_X1 U13471 ( .A(n10817), .B(n10819), .ZN(n14662) );
  NOR2_X1 U13472 ( .A1(n14147), .A2(n14661), .ZN(n14180) );
  INV_X1 U13473 ( .A(n14180), .ZN(n14131) );
  XNOR2_X1 U13474 ( .A(n10818), .B(n10819), .ZN(n14665) );
  INV_X1 U13475 ( .A(n14219), .ZN(n14256) );
  NAND2_X1 U13476 ( .A1(n14665), .A2(n14256), .ZN(n10829) );
  INV_X1 U13477 ( .A(n11207), .ZN(n10824) );
  NAND2_X1 U13478 ( .A1(n13880), .A2(n14642), .ZN(n10821) );
  NAND2_X1 U13479 ( .A1(n13883), .A2(n14498), .ZN(n10820) );
  AND2_X1 U13480 ( .A1(n10821), .A2(n10820), .ZN(n14658) );
  MUX2_X1 U13481 ( .A(n10822), .B(n14658), .S(n14253), .Z(n10823) );
  OAI21_X1 U13482 ( .B1(n14206), .B2(n10824), .A(n10823), .ZN(n10827) );
  OAI211_X1 U13483 ( .C1(n10825), .C2(n14660), .A(n14302), .B(n10837), .ZN(
        n14659) );
  NOR2_X1 U13484 ( .A1(n14659), .A2(n14239), .ZN(n10826) );
  AOI211_X1 U13485 ( .C1(n14246), .C2(n11836), .A(n10827), .B(n10826), .ZN(
        n10828) );
  OAI211_X1 U13486 ( .C1(n14662), .C2(n14131), .A(n10829), .B(n10828), .ZN(
        P1_U3287) );
  XNOR2_X1 U13487 ( .A(n10830), .B(n11997), .ZN(n10831) );
  NAND2_X1 U13488 ( .A1(n10831), .A2(n14676), .ZN(n10836) );
  XNOR2_X1 U13489 ( .A(n10832), .B(n11997), .ZN(n10833) );
  NAND2_X1 U13490 ( .A1(n10833), .A2(n14684), .ZN(n10835) );
  AOI22_X1 U13491 ( .A1(n14498), .A2(n13882), .B1(n13879), .B2(n14642), .ZN(
        n10834) );
  AOI21_X1 U13492 ( .B1(n10837), .B2(n11839), .A(n14644), .ZN(n10838) );
  NAND2_X1 U13493 ( .A1(n10838), .A2(n11145), .ZN(n10909) );
  AND2_X1 U13494 ( .A1(n10905), .A2(n10909), .ZN(n10844) );
  INV_X1 U13495 ( .A(n11839), .ZN(n10840) );
  INV_X1 U13496 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10839) );
  OAI22_X1 U13497 ( .A1(n14348), .A2(n10840), .B1(n14687), .B2(n10839), .ZN(
        n10841) );
  INV_X1 U13498 ( .A(n10841), .ZN(n10842) );
  OAI21_X1 U13499 ( .B1(n10844), .B2(n14685), .A(n10842), .ZN(P1_U3480) );
  AOI22_X1 U13500 ( .A1(n9824), .A2(n11839), .B1(n14695), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n10843) );
  OAI21_X1 U13501 ( .B1(n10844), .B2(n14695), .A(n10843), .ZN(P1_U3535) );
  NAND2_X1 U13502 ( .A1(n10845), .A2(n14381), .ZN(n10846) );
  INV_X1 U13503 ( .A(n12290), .ZN(n12296) );
  OAI211_X1 U13504 ( .C1(n10847), .C2(n13004), .A(n10846), .B(n12296), .ZN(
        P3_U3272) );
  XNOR2_X1 U13505 ( .A(n12070), .B(n10851), .ZN(n11697) );
  NAND2_X1 U13506 ( .A1(n13470), .A2(n13151), .ZN(n10849) );
  XNOR2_X1 U13507 ( .A(n11697), .B(n10849), .ZN(n12066) );
  INV_X1 U13508 ( .A(n11697), .ZN(n10850) );
  XNOR2_X1 U13509 ( .A(n11703), .B(n10851), .ZN(n10852) );
  NAND2_X1 U13510 ( .A1(n13470), .A2(n13149), .ZN(n10853) );
  XNOR2_X1 U13511 ( .A(n10852), .B(n10853), .ZN(n11698) );
  INV_X1 U13512 ( .A(n10852), .ZN(n10854) );
  NAND2_X1 U13513 ( .A1(n10854), .A2(n10853), .ZN(n10855) );
  XNOR2_X1 U13514 ( .A(n10856), .B(n11708), .ZN(n10858) );
  AND2_X1 U13515 ( .A1(n10857), .A2(n13148), .ZN(n10859) );
  NAND2_X1 U13516 ( .A1(n10858), .A2(n10859), .ZN(n10994) );
  INV_X1 U13517 ( .A(n10858), .ZN(n10861) );
  INV_X1 U13518 ( .A(n10859), .ZN(n10860) );
  NAND2_X1 U13519 ( .A1(n10861), .A2(n10860), .ZN(n10862) );
  NAND2_X1 U13520 ( .A1(n10994), .A2(n10862), .ZN(n10864) );
  AOI21_X1 U13521 ( .B1(n10863), .B2(n10864), .A(n14462), .ZN(n10867) );
  INV_X1 U13522 ( .A(n10863), .ZN(n10866) );
  NAND2_X1 U13523 ( .A1(n10867), .A2(n10995), .ZN(n10873) );
  NAND2_X1 U13524 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14782)
         );
  INV_X1 U13525 ( .A(n14782), .ZN(n10870) );
  OAI22_X1 U13526 ( .A1(n11005), .A2(n14458), .B1(n14457), .B2(n10868), .ZN(
        n10869) );
  AOI211_X1 U13527 ( .C1(n10871), .C2(n13098), .A(n10870), .B(n10869), .ZN(
        n10872) );
  OAI211_X1 U13528 ( .C1(n14928), .C2(n13139), .A(n10873), .B(n10872), .ZN(
        P2_U3189) );
  NAND2_X1 U13529 ( .A1(n10875), .A2(n10874), .ZN(n10981) );
  XNOR2_X1 U13530 ( .A(n10981), .B(n10881), .ZN(n10876) );
  NAND2_X1 U13531 ( .A1(n10876), .A2(n13526), .ZN(n10878) );
  AOI22_X1 U13532 ( .A1(n13145), .A2(n13521), .B1(n13523), .B2(n13147), .ZN(
        n10877) );
  NAND2_X1 U13533 ( .A1(n10878), .A2(n10877), .ZN(n14475) );
  INV_X1 U13534 ( .A(n14475), .ZN(n10889) );
  AND2_X1 U13535 ( .A1(n14937), .A2(n13147), .ZN(n10879) );
  INV_X1 U13536 ( .A(n10881), .ZN(n10882) );
  XNOR2_X1 U13537 ( .A(n10990), .B(n10882), .ZN(n14471) );
  AOI21_X1 U13538 ( .B1(n11003), .B2(n10883), .A(n10602), .ZN(n10884) );
  NAND2_X1 U13539 ( .A1(n10884), .A2(n10986), .ZN(n14472) );
  OAI22_X1 U13540 ( .A1(n13527), .A2(n13180), .B1(n11000), .B2(n13466), .ZN(
        n10885) );
  AOI21_X1 U13541 ( .B1(n11003), .B2(n13530), .A(n10885), .ZN(n10886) );
  OAI21_X1 U13542 ( .B1(n14472), .B2(n13515), .A(n10886), .ZN(n10887) );
  AOI21_X1 U13543 ( .B1(n14471), .B2(n13534), .A(n10887), .ZN(n10888) );
  OAI21_X1 U13544 ( .B1(n10889), .B2(n13512), .A(n10888), .ZN(P2_U3253) );
  INV_X1 U13545 ( .A(n10890), .ZN(n11242) );
  OAI22_X1 U13546 ( .A1(n14196), .A2(n10891), .B1(n14206), .B2(n11242), .ZN(
        n10894) );
  MUX2_X1 U13547 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10892), .S(n14253), .Z(
        n10893) );
  AOI211_X1 U13548 ( .C1(n14124), .C2(n10895), .A(n10894), .B(n10893), .ZN(
        n10896) );
  INV_X1 U13549 ( .A(n10896), .ZN(P1_U3288) );
  INV_X1 U13550 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10902) );
  AOI21_X1 U13551 ( .B1(n14936), .B2(n11703), .A(n10897), .ZN(n10898) );
  OAI211_X1 U13552 ( .C1(n10900), .C2(n13648), .A(n10899), .B(n10898), .ZN(
        n10903) );
  NAND2_X1 U13553 ( .A1(n10903), .A2(n14944), .ZN(n10901) );
  OAI21_X1 U13554 ( .B1(n14944), .B2(n10902), .A(n10901), .ZN(P2_U3457) );
  INV_X1 U13555 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n13195) );
  NAND2_X1 U13556 ( .A1(n10903), .A2(n14960), .ZN(n10904) );
  OAI21_X1 U13557 ( .B1(n14960), .B2(n13195), .A(n10904), .ZN(P2_U3508) );
  MUX2_X1 U13558 ( .A(n10906), .B(n10905), .S(n14253), .Z(n10908) );
  AOI22_X1 U13559 ( .A1(n14246), .A2(n11839), .B1(n14243), .B2(n11396), .ZN(
        n10907) );
  OAI211_X1 U13560 ( .C1(n14239), .C2(n10909), .A(n10908), .B(n10907), .ZN(
        P1_U3286) );
  AOI21_X1 U13561 ( .B1(n10912), .B2(n10911), .A(n10910), .ZN(n10926) );
  OAI21_X1 U13562 ( .B1(n10915), .B2(n10914), .A(n10913), .ZN(n10916) );
  INV_X1 U13563 ( .A(n15076), .ZN(n15096) );
  NAND2_X1 U13564 ( .A1(n10916), .A2(n15096), .ZN(n10925) );
  OAI21_X1 U13565 ( .B1(n10919), .B2(n10918), .A(n10917), .ZN(n10923) );
  NAND2_X1 U13566 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n14972) );
  NAND2_X1 U13567 ( .A1(n15089), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10920) );
  OAI211_X1 U13568 ( .C1(n15092), .C2(n10921), .A(n14972), .B(n10920), .ZN(
        n10922) );
  AOI21_X1 U13569 ( .B1(n15094), .B2(n10923), .A(n10922), .ZN(n10924) );
  OAI211_X1 U13570 ( .C1(n10926), .C2(n15102), .A(n10925), .B(n10924), .ZN(
        P3_U3190) );
  INV_X1 U13571 ( .A(n10927), .ZN(n10930) );
  INV_X1 U13572 ( .A(n13847), .ZN(n13805) );
  AOI22_X1 U13573 ( .A1(n13805), .A2(n10928), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10929) );
  OAI21_X1 U13574 ( .B1(n13786), .B2(n10930), .A(n10929), .ZN(n10942) );
  AOI22_X1 U13575 ( .A1(n13884), .A2(n11584), .B1(n12360), .B2(n14652), .ZN(
        n10931) );
  XNOR2_X1 U13576 ( .A(n10931), .B(n12370), .ZN(n10940) );
  INV_X1 U13577 ( .A(n10932), .ZN(n10935) );
  INV_X1 U13578 ( .A(n10933), .ZN(n10934) );
  AOI22_X1 U13579 ( .A1(n12364), .A2(n13884), .B1(n11584), .B2(n14652), .ZN(
        n11196) );
  AOI211_X1 U13580 ( .C1(n10940), .C2(n10939), .A(n13864), .B(n11195), .ZN(
        n10941) );
  AOI211_X1 U13581 ( .C1(n14652), .C2(n13817), .A(n10942), .B(n10941), .ZN(
        n10943) );
  INV_X1 U13582 ( .A(n10943), .ZN(P1_U3230) );
  INV_X1 U13583 ( .A(n10944), .ZN(n10945) );
  NAND2_X1 U13584 ( .A1(n10945), .A2(n15126), .ZN(n10947) );
  INV_X1 U13585 ( .A(n15121), .ZN(n12797) );
  AOI22_X1 U13586 ( .A1(n12813), .A2(n10618), .B1(n12797), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10946) );
  OAI211_X1 U13587 ( .C1(n9828), .C2(n15126), .A(n10947), .B(n10946), .ZN(
        P3_U3233) );
  OAI21_X1 U13588 ( .B1(n10950), .B2(n10948), .A(n10949), .ZN(n15145) );
  INV_X1 U13589 ( .A(n15145), .ZN(n15141) );
  INV_X1 U13590 ( .A(n10951), .ZN(n10952) );
  AOI21_X1 U13591 ( .B1(n10952), .B2(n10948), .A(n15117), .ZN(n10956) );
  NAND2_X1 U13592 ( .A1(n12605), .A2(n12573), .ZN(n10954) );
  NAND2_X1 U13593 ( .A1(n9672), .A2(n12572), .ZN(n10953) );
  NAND2_X1 U13594 ( .A1(n10954), .A2(n10953), .ZN(n12413) );
  AOI21_X1 U13595 ( .B1(n10956), .B2(n10955), .A(n12413), .ZN(n15142) );
  MUX2_X1 U13596 ( .A(n10957), .B(n15142), .S(n15126), .Z(n10960) );
  INV_X1 U13597 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13598 ( .A1(n12813), .A2(n12412), .B1(n12797), .B2(n10958), .ZN(
        n10959) );
  OAI211_X1 U13599 ( .C1(n12802), .C2(n15141), .A(n10960), .B(n10959), .ZN(
        P3_U3230) );
  OAI21_X1 U13600 ( .B1(n10384), .B2(n10968), .A(n10961), .ZN(n10962) );
  NOR2_X1 U13601 ( .A1(n10962), .A2(n10969), .ZN(n10964) );
  AOI21_X1 U13602 ( .B1(n10969), .B2(n10962), .A(n10964), .ZN(n10963) );
  INV_X1 U13603 ( .A(n10963), .ZN(n14611) );
  NOR2_X1 U13604 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14611), .ZN(n14610) );
  NOR2_X1 U13605 ( .A1(n10964), .A2(n14610), .ZN(n10966) );
  INV_X1 U13606 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U13607 ( .A1(n10973), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11221), 
        .B2(n11227), .ZN(n10965) );
  NAND2_X1 U13608 ( .A1(n10965), .A2(n10966), .ZN(n11220) );
  OAI211_X1 U13609 ( .C1(n10966), .C2(n10965), .A(n14628), .B(n11220), .ZN(
        n10979) );
  NAND2_X1 U13610 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13776)
         );
  INV_X1 U13611 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14519) );
  AOI21_X1 U13612 ( .B1(n14519), .B2(n10968), .A(n10967), .ZN(n10970) );
  INV_X1 U13613 ( .A(n10970), .ZN(n10971) );
  XNOR2_X1 U13614 ( .A(n10970), .B(n10969), .ZN(n14613) );
  NOR2_X1 U13615 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14613), .ZN(n14612) );
  AOI21_X1 U13616 ( .B1(n14617), .B2(n10971), .A(n14612), .ZN(n10975) );
  NOR2_X1 U13617 ( .A1(n10973), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10972) );
  AOI21_X1 U13618 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n10973), .A(n10972), 
        .ZN(n10974) );
  NAND2_X1 U13619 ( .A1(n10974), .A2(n10975), .ZN(n11226) );
  OAI211_X1 U13620 ( .C1(n10975), .C2(n10974), .A(n14600), .B(n11226), .ZN(
        n10976) );
  NAND2_X1 U13621 ( .A1(n13776), .A2(n10976), .ZN(n10977) );
  AOI21_X1 U13622 ( .B1(n14596), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10977), 
        .ZN(n10978) );
  OAI211_X1 U13623 ( .C1(n14618), .C2(n11227), .A(n10979), .B(n10978), .ZN(
        P1_U3259) );
  INV_X1 U13624 ( .A(n13146), .ZN(n14459) );
  INV_X1 U13625 ( .A(n11003), .ZN(n14473) );
  XNOR2_X1 U13626 ( .A(n11266), .B(n10991), .ZN(n10984) );
  NAND2_X1 U13627 ( .A1(n13257), .A2(n13521), .ZN(n10983) );
  NAND2_X1 U13628 ( .A1(n13146), .A2(n13523), .ZN(n10982) );
  NAND2_X1 U13629 ( .A1(n10983), .A2(n10982), .ZN(n11406) );
  AOI21_X1 U13630 ( .B1(n10984), .B2(n13526), .A(n11406), .ZN(n13642) );
  INV_X1 U13631 ( .A(n11271), .ZN(n10985) );
  AOI211_X1 U13632 ( .C1(n13641), .C2(n10986), .A(n10602), .B(n10985), .ZN(
        n13640) );
  NOR2_X1 U13633 ( .A1(n6981), .A2(n13489), .ZN(n10988) );
  INV_X1 U13634 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13173) );
  OAI22_X1 U13635 ( .A1(n13527), .A2(n13173), .B1(n11408), .B2(n13466), .ZN(
        n10987) );
  AOI211_X1 U13636 ( .C1(n13640), .C2(n13538), .A(n10988), .B(n10987), .ZN(
        n10993) );
  NOR2_X1 U13637 ( .A1(n11003), .A2(n13146), .ZN(n10989) );
  INV_X1 U13638 ( .A(n10991), .ZN(n11265) );
  XNOR2_X1 U13639 ( .A(n11268), .B(n11265), .ZN(n13644) );
  OR2_X1 U13640 ( .A1(n13644), .A2(n13475), .ZN(n10992) );
  OAI211_X1 U13641 ( .C1(n13642), .C2(n13512), .A(n10993), .B(n10992), .ZN(
        P2_U3252) );
  XNOR2_X1 U13642 ( .A(n14937), .B(n11730), .ZN(n11006) );
  NAND2_X1 U13643 ( .A1(n13470), .A2(n13147), .ZN(n10997) );
  XNOR2_X1 U13644 ( .A(n11006), .B(n10997), .ZN(n14460) );
  INV_X1 U13645 ( .A(n14460), .ZN(n10996) );
  NAND2_X1 U13646 ( .A1(n11006), .A2(n10997), .ZN(n10998) );
  XNOR2_X1 U13647 ( .A(n11003), .B(n11708), .ZN(n11413) );
  NAND2_X1 U13648 ( .A1(n13470), .A2(n13146), .ZN(n11414) );
  XNOR2_X1 U13649 ( .A(n11413), .B(n11414), .ZN(n11004) );
  OAI22_X1 U13650 ( .A1(n14470), .A2(n11000), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10999), .ZN(n11002) );
  OAI22_X1 U13651 ( .A1(n12049), .A2(n14458), .B1(n14457), .B2(n11005), .ZN(
        n11001) );
  AOI211_X1 U13652 ( .C1(n11003), .C2(n14467), .A(n11002), .B(n11001), .ZN(
        n11009) );
  OAI22_X1 U13653 ( .A1(n11006), .A2(n14462), .B1(n11005), .B2(n13132), .ZN(
        n11007) );
  NAND3_X1 U13654 ( .A1(n14464), .A2(n6796), .A3(n11007), .ZN(n11008) );
  OAI211_X1 U13655 ( .C1(n11417), .C2(n14462), .A(n11009), .B(n11008), .ZN(
        P2_U3196) );
  INV_X1 U13656 ( .A(n11010), .ZN(n11119) );
  INV_X1 U13657 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11011) );
  OAI222_X1 U13658 ( .A1(n13685), .A2(n11119), .B1(P2_U3088), .B2(n11012), 
        .C1(n11011), .C2(n13688), .ZN(P2_U3307) );
  XOR2_X1 U13659 ( .A(n11014), .B(n11013), .Z(n11029) );
  OAI21_X1 U13660 ( .B1(n11017), .B2(n11016), .A(n11015), .ZN(n11018) );
  NAND2_X1 U13661 ( .A1(n14441), .A2(n11018), .ZN(n11025) );
  AOI22_X1 U13662 ( .A1(n15089), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11024) );
  OAI21_X1 U13663 ( .B1(n11021), .B2(n11020), .A(n11019), .ZN(n11022) );
  NAND2_X1 U13664 ( .A1(n15094), .A2(n11022), .ZN(n11023) );
  NAND3_X1 U13665 ( .A1(n11025), .A2(n11024), .A3(n11023), .ZN(n11026) );
  AOI21_X1 U13666 ( .B1(n6500), .B2(n15002), .A(n11026), .ZN(n11028) );
  OAI21_X1 U13667 ( .B1(n11029), .B2(n15076), .A(n11028), .ZN(P3_U3184) );
  XNOR2_X1 U13668 ( .A(n11031), .B(n11030), .ZN(n11043) );
  AOI21_X1 U13669 ( .B1(n11033), .B2(n8971), .A(n11032), .ZN(n11034) );
  NOR2_X1 U13670 ( .A1(n11034), .A2(n15102), .ZN(n11042) );
  AOI22_X1 U13671 ( .A1(n15089), .A2(P3_ADDR_REG_7__SCAN_IN), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(P3_U3151), .ZN(n11039) );
  OAI21_X1 U13672 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n11036), .A(n11035), .ZN(
        n11037) );
  NAND2_X1 U13673 ( .A1(n15094), .A2(n11037), .ZN(n11038) );
  OAI211_X1 U13674 ( .C1(n15092), .C2(n11040), .A(n11039), .B(n11038), .ZN(
        n11041) );
  AOI211_X1 U13675 ( .C1(n11043), .C2(n15096), .A(n11042), .B(n11041), .ZN(
        n11044) );
  INV_X1 U13676 ( .A(n11044), .ZN(P3_U3189) );
  XOR2_X1 U13677 ( .A(n11046), .B(n11045), .Z(n11059) );
  AOI21_X1 U13678 ( .B1(n11048), .B2(n11259), .A(n11047), .ZN(n11055) );
  OAI21_X1 U13679 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n11050), .A(n11049), .ZN(
        n11053) );
  INV_X1 U13680 ( .A(n15089), .ZN(n15011) );
  INV_X1 U13681 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n11051) );
  NAND2_X1 U13682 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11067) );
  OAI21_X1 U13683 ( .B1(n15011), .B2(n11051), .A(n11067), .ZN(n11052) );
  AOI21_X1 U13684 ( .B1(n15094), .B2(n11053), .A(n11052), .ZN(n11054) );
  OAI21_X1 U13685 ( .B1(n11055), .B2(n15102), .A(n11054), .ZN(n11056) );
  AOI21_X1 U13686 ( .B1(n11057), .B2(n15002), .A(n11056), .ZN(n11058) );
  OAI21_X1 U13687 ( .B1(n11059), .B2(n15076), .A(n11058), .ZN(P3_U3187) );
  AND2_X1 U13688 ( .A1(n11061), .A2(n11060), .ZN(n11063) );
  XNOR2_X1 U13689 ( .A(n11063), .B(n11062), .ZN(n11064) );
  NAND2_X1 U13690 ( .A1(n11064), .A2(n14974), .ZN(n11070) );
  NAND2_X1 U13691 ( .A1(n12603), .A2(n12573), .ZN(n11066) );
  NAND2_X1 U13692 ( .A1(n12605), .A2(n12572), .ZN(n11065) );
  NAND2_X1 U13693 ( .A1(n11066), .A2(n11065), .ZN(n11257) );
  OAI21_X1 U13694 ( .B1(n14973), .B2(n15154), .A(n11067), .ZN(n11068) );
  AOI21_X1 U13695 ( .B1(n11257), .B2(n14982), .A(n11068), .ZN(n11069) );
  OAI211_X1 U13696 ( .C1(n11260), .C2(n14985), .A(n11070), .B(n11069), .ZN(
        P3_U3167) );
  XOR2_X1 U13697 ( .A(n11072), .B(n11071), .Z(n11086) );
  AOI21_X1 U13698 ( .B1(n11075), .B2(n11074), .A(n11073), .ZN(n11082) );
  OAI21_X1 U13699 ( .B1(n11078), .B2(n11077), .A(n11076), .ZN(n11080) );
  NAND2_X1 U13700 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11158) );
  OAI21_X1 U13701 ( .B1(n15011), .B2(n9393), .A(n11158), .ZN(n11079) );
  AOI21_X1 U13702 ( .B1(n15094), .B2(n11080), .A(n11079), .ZN(n11081) );
  OAI21_X1 U13703 ( .B1(n11082), .B2(n15102), .A(n11081), .ZN(n11083) );
  AOI21_X1 U13704 ( .B1(n11084), .B2(n15002), .A(n11083), .ZN(n11085) );
  OAI21_X1 U13705 ( .B1(n11086), .B2(n15076), .A(n11085), .ZN(P3_U3186) );
  XOR2_X1 U13706 ( .A(n11088), .B(n11087), .Z(n11102) );
  AOI21_X1 U13707 ( .B1(n6648), .B2(n11090), .A(n11089), .ZN(n11098) );
  OAI21_X1 U13708 ( .B1(n11093), .B2(n11092), .A(n11091), .ZN(n11096) );
  INV_X1 U13709 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U13710 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11178) );
  OAI21_X1 U13711 ( .B1(n15011), .B2(n11094), .A(n11178), .ZN(n11095) );
  AOI21_X1 U13712 ( .B1(n15094), .B2(n11096), .A(n11095), .ZN(n11097) );
  OAI21_X1 U13713 ( .B1(n11098), .B2(n15102), .A(n11097), .ZN(n11099) );
  AOI21_X1 U13714 ( .B1(n11100), .B2(n15002), .A(n11099), .ZN(n11101) );
  OAI21_X1 U13715 ( .B1(n11102), .B2(n15076), .A(n11101), .ZN(P3_U3188) );
  XOR2_X1 U13716 ( .A(n14987), .B(n11103), .Z(n11118) );
  INV_X1 U13717 ( .A(n9830), .ZN(n11116) );
  NAND2_X1 U13718 ( .A1(n11104), .A2(n8852), .ZN(n11105) );
  AND2_X1 U13719 ( .A1(n11106), .A2(n11105), .ZN(n11114) );
  AOI22_X1 U13720 ( .A1(n15089), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11113) );
  NAND2_X1 U13721 ( .A1(n11108), .A2(n11107), .ZN(n11109) );
  NAND2_X1 U13722 ( .A1(n11110), .A2(n11109), .ZN(n11111) );
  NAND2_X1 U13723 ( .A1(n15094), .A2(n11111), .ZN(n11112) );
  OAI211_X1 U13724 ( .C1(n11114), .C2(n15102), .A(n11113), .B(n11112), .ZN(
        n11115) );
  AOI21_X1 U13725 ( .B1(n11116), .B2(n15002), .A(n11115), .ZN(n11117) );
  OAI21_X1 U13726 ( .B1(n15076), .B2(n11118), .A(n11117), .ZN(P3_U3183) );
  OAI222_X1 U13727 ( .A1(n11120), .A2(P1_U3086), .B1(n14366), .B2(n11119), 
        .C1(n6887), .C2(n14363), .ZN(P1_U3335) );
  XOR2_X1 U13728 ( .A(n11122), .B(n11121), .Z(n11134) );
  AOI21_X1 U13729 ( .B1(n11124), .B2(n10957), .A(n11123), .ZN(n11130) );
  AOI22_X1 U13730 ( .A1(n15089), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11129) );
  OAI21_X1 U13731 ( .B1(n11126), .B2(P3_REG1_REG_3__SCAN_IN), .A(n11125), .ZN(
        n11127) );
  NAND2_X1 U13732 ( .A1(n15094), .A2(n11127), .ZN(n11128) );
  OAI211_X1 U13733 ( .C1(n11130), .C2(n15102), .A(n11129), .B(n11128), .ZN(
        n11131) );
  AOI21_X1 U13734 ( .B1(n11132), .B2(n15002), .A(n11131), .ZN(n11133) );
  OAI21_X1 U13735 ( .B1(n11134), .B2(n15076), .A(n11133), .ZN(P3_U3185) );
  INV_X1 U13736 ( .A(n11135), .ZN(n11139) );
  INV_X1 U13737 ( .A(n11136), .ZN(n11138) );
  OAI222_X1 U13738 ( .A1(P3_U3151), .A2(n11139), .B1(n12387), .B2(n11138), 
        .C1(n11137), .C2(n13004), .ZN(P3_U3271) );
  XOR2_X1 U13739 ( .A(n11140), .B(n11996), .Z(n14673) );
  XOR2_X1 U13740 ( .A(n11996), .B(n11141), .Z(n11143) );
  OAI22_X1 U13741 ( .A1(n11142), .A2(n14520), .B1(n11535), .B2(n14522), .ZN(
        n11340) );
  AOI21_X1 U13742 ( .B1(n11143), .B2(n14676), .A(n11340), .ZN(n14671) );
  MUX2_X1 U13743 ( .A(n11144), .B(n14671), .S(n14253), .Z(n11149) );
  AOI211_X1 U13744 ( .C1(n14668), .C2(n11145), .A(n14644), .B(n6966), .ZN(
        n14667) );
  INV_X1 U13745 ( .A(n14668), .ZN(n11146) );
  OAI22_X1 U13746 ( .A1(n11146), .A2(n14196), .B1(n11342), .B2(n14206), .ZN(
        n11147) );
  AOI21_X1 U13747 ( .B1(n14667), .B2(n14124), .A(n11147), .ZN(n11148) );
  OAI211_X1 U13748 ( .C1(n14219), .C2(n14673), .A(n11149), .B(n11148), .ZN(
        P1_U3285) );
  OR2_X1 U13749 ( .A1(n12409), .A2(n12408), .ZN(n12410) );
  AND2_X1 U13750 ( .A1(n12410), .A2(n11150), .ZN(n11153) );
  NAND2_X1 U13751 ( .A1(n12410), .A2(n11151), .ZN(n11152) );
  OAI21_X1 U13752 ( .B1(n11154), .B2(n11153), .A(n11152), .ZN(n11155) );
  NAND2_X1 U13753 ( .A1(n11155), .A2(n14974), .ZN(n11161) );
  NAND2_X1 U13754 ( .A1(n12604), .A2(n12573), .ZN(n11157) );
  NAND2_X1 U13755 ( .A1(n12606), .A2(n12572), .ZN(n11156) );
  NAND2_X1 U13756 ( .A1(n11157), .A2(n11156), .ZN(n11163) );
  OAI21_X1 U13757 ( .B1(n14973), .B2(n15147), .A(n11158), .ZN(n11159) );
  AOI21_X1 U13758 ( .B1(n11163), .B2(n14982), .A(n11159), .ZN(n11160) );
  OAI211_X1 U13759 ( .C1(n11168), .C2(n14985), .A(n11161), .B(n11160), .ZN(
        P3_U3170) );
  XNOR2_X1 U13760 ( .A(n11162), .B(n12117), .ZN(n15148) );
  INV_X1 U13761 ( .A(n11163), .ZN(n11167) );
  OAI211_X1 U13762 ( .C1(n11165), .C2(n12117), .A(n11164), .B(n12804), .ZN(
        n11166) );
  OAI211_X1 U13763 ( .C1(n15148), .C2(n15164), .A(n11167), .B(n11166), .ZN(
        n15150) );
  NAND2_X1 U13764 ( .A1(n15150), .A2(n15126), .ZN(n11171) );
  INV_X1 U13765 ( .A(n12798), .ZN(n12841) );
  OAI22_X1 U13766 ( .A1(n12841), .A2(n15147), .B1(n11168), .B2(n15121), .ZN(
        n11169) );
  AOI21_X1 U13767 ( .B1(n15128), .B2(P3_REG2_REG_4__SCAN_IN), .A(n11169), .ZN(
        n11170) );
  OAI211_X1 U13768 ( .C1(n15148), .C2(n12694), .A(n11171), .B(n11170), .ZN(
        P3_U3229) );
  AOI21_X1 U13769 ( .B1(n11173), .B2(n11172), .A(n12579), .ZN(n11175) );
  NAND2_X1 U13770 ( .A1(n11175), .A2(n11174), .ZN(n11182) );
  NAND2_X1 U13771 ( .A1(n12602), .A2(n12573), .ZN(n11177) );
  NAND2_X1 U13772 ( .A1(n12604), .A2(n12572), .ZN(n11176) );
  AND2_X1 U13773 ( .A1(n11177), .A2(n11176), .ZN(n11312) );
  INV_X1 U13774 ( .A(n11312), .ZN(n11180) );
  OAI21_X1 U13775 ( .B1(n14973), .B2(n15158), .A(n11178), .ZN(n11179) );
  AOI21_X1 U13776 ( .B1(n11180), .B2(n14982), .A(n11179), .ZN(n11181) );
  OAI211_X1 U13777 ( .C1(n11313), .C2(n14985), .A(n11182), .B(n11181), .ZN(
        P3_U3179) );
  XNOR2_X1 U13778 ( .A(n11183), .B(n11999), .ZN(n11189) );
  OAI21_X1 U13779 ( .B1(n6640), .B2(n11999), .A(n11184), .ZN(n11187) );
  OAI22_X1 U13780 ( .A1(n11185), .A2(n14520), .B1(n13827), .B2(n14522), .ZN(
        n11186) );
  AOI21_X1 U13781 ( .B1(n11187), .B2(n14676), .A(n11186), .ZN(n11188) );
  OAI21_X1 U13782 ( .B1(n14672), .B2(n11189), .A(n11188), .ZN(n11214) );
  INV_X1 U13783 ( .A(n11214), .ZN(n11194) );
  AOI211_X1 U13784 ( .C1(n11849), .C2(n11190), .A(n14644), .B(n11296), .ZN(
        n11213) );
  AOI22_X1 U13785 ( .A1(n14147), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11504), 
        .B2(n14243), .ZN(n11191) );
  OAI21_X1 U13786 ( .B1(n6970), .B2(n14196), .A(n11191), .ZN(n11192) );
  AOI21_X1 U13787 ( .B1(n11213), .B2(n14124), .A(n11192), .ZN(n11193) );
  OAI21_X1 U13788 ( .B1(n11194), .B2(n14147), .A(n11193), .ZN(P1_U3284) );
  INV_X1 U13789 ( .A(n11195), .ZN(n11199) );
  NAND2_X1 U13790 ( .A1(n11197), .A2(n10938), .ZN(n11198) );
  NAND2_X1 U13791 ( .A1(n12364), .A2(n13883), .ZN(n11201) );
  NAND2_X1 U13792 ( .A1(n11829), .A2(n11633), .ZN(n11200) );
  NAND2_X1 U13793 ( .A1(n11201), .A2(n11200), .ZN(n11243) );
  INV_X1 U13794 ( .A(n11243), .ZN(n11203) );
  AOI22_X1 U13795 ( .A1(n11829), .A2(n12360), .B1(n13883), .B2(n11584), .ZN(
        n11202) );
  XOR2_X1 U13796 ( .A(n12370), .B(n11202), .Z(n11244) );
  NAND2_X1 U13797 ( .A1(n11836), .A2(n12360), .ZN(n11205) );
  NAND2_X1 U13798 ( .A1(n13882), .A2(n11584), .ZN(n11204) );
  NAND2_X1 U13799 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  XNOR2_X1 U13800 ( .A(n11206), .B(n12370), .ZN(n11324) );
  AOI22_X1 U13801 ( .A1(n11836), .A2(n11633), .B1(n12364), .B2(n13882), .ZN(
        n11323) );
  XNOR2_X1 U13802 ( .A(n11324), .B(n11323), .ZN(n11326) );
  XNOR2_X1 U13803 ( .A(n11327), .B(n11326), .ZN(n11212) );
  NAND2_X1 U13804 ( .A1(n13862), .A2(n11207), .ZN(n11209) );
  OAI211_X1 U13805 ( .C1(n14658), .C2(n13847), .A(n11209), .B(n11208), .ZN(
        n11210) );
  AOI21_X1 U13806 ( .B1(n11836), .B2(n13817), .A(n11210), .ZN(n11211) );
  OAI21_X1 U13807 ( .B1(n11212), .B2(n13864), .A(n11211), .ZN(P1_U3239) );
  NOR2_X1 U13808 ( .A1(n11214), .A2(n11213), .ZN(n11219) );
  INV_X1 U13809 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11215) );
  OAI22_X1 U13810 ( .A1(n6970), .A2(n14348), .B1(n14687), .B2(n11215), .ZN(
        n11216) );
  INV_X1 U13811 ( .A(n11216), .ZN(n11217) );
  OAI21_X1 U13812 ( .B1(n11219), .B2(n14685), .A(n11217), .ZN(P1_U3486) );
  AOI22_X1 U13813 ( .A1(n11849), .A2(n9824), .B1(n14695), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11218) );
  OAI21_X1 U13814 ( .B1(n11219), .B2(n14695), .A(n11218), .ZN(P1_U3537) );
  OAI21_X1 U13815 ( .B1(n11221), .B2(n11227), .A(n11220), .ZN(n11223) );
  INV_X1 U13816 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14208) );
  AOI22_X1 U13817 ( .A1(n14003), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14208), 
        .B2(n13998), .ZN(n11222) );
  NAND2_X1 U13818 ( .A1(n11222), .A2(n11223), .ZN(n14004) );
  OAI211_X1 U13819 ( .C1(n11223), .C2(n11222), .A(n14628), .B(n14004), .ZN(
        n11233) );
  NAND2_X1 U13820 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13787)
         );
  NOR2_X1 U13821 ( .A1(n13998), .A2(n11224), .ZN(n11225) );
  AOI21_X1 U13822 ( .B1(n11224), .B2(n13998), .A(n11225), .ZN(n11229) );
  INV_X1 U13823 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14497) );
  OAI21_X1 U13824 ( .B1(n14497), .B2(n11227), .A(n11226), .ZN(n11228) );
  NAND2_X1 U13825 ( .A1(n11229), .A2(n11228), .ZN(n13997) );
  OAI211_X1 U13826 ( .C1(n11229), .C2(n11228), .A(n13997), .B(n14600), .ZN(
        n11230) );
  NAND2_X1 U13827 ( .A1(n13787), .A2(n11230), .ZN(n11231) );
  AOI21_X1 U13828 ( .B1(n14596), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11231), 
        .ZN(n11232) );
  OAI211_X1 U13829 ( .C1(n14618), .C2(n13998), .A(n11233), .B(n11232), .ZN(
        P1_U3260) );
  INV_X1 U13830 ( .A(n11234), .ZN(n11238) );
  OAI222_X1 U13831 ( .A1(n13688), .A2(n11236), .B1(n13685), .B2(n11238), .C1(
        P2_U3088), .C2(n11235), .ZN(P2_U3306) );
  OAI222_X1 U13832 ( .A1(P1_U3086), .A2(n11794), .B1(n14366), .B2(n11238), 
        .C1(n11237), .C2(n14363), .ZN(P1_U3334) );
  AOI21_X1 U13833 ( .B1(n13825), .B2(n13882), .A(n11239), .ZN(n11241) );
  NAND2_X1 U13834 ( .A1(n13855), .A2(n13884), .ZN(n11240) );
  OAI211_X1 U13835 ( .C1(n13786), .C2(n11242), .A(n11241), .B(n11240), .ZN(
        n11249) );
  XNOR2_X1 U13836 ( .A(n11244), .B(n11243), .ZN(n11245) );
  XNOR2_X1 U13837 ( .A(n11246), .B(n11245), .ZN(n11247) );
  NOR2_X1 U13838 ( .A1(n11247), .A2(n13864), .ZN(n11248) );
  AOI211_X1 U13839 ( .C1(n11829), .C2(n13817), .A(n11249), .B(n11248), .ZN(
        n11250) );
  INV_X1 U13840 ( .A(n11250), .ZN(P1_U3227) );
  INV_X1 U13841 ( .A(n11251), .ZN(n11252) );
  OAI222_X1 U13842 ( .A1(n13688), .A2(n11253), .B1(n13685), .B2(n11252), .C1(
        P2_U3088), .C2(n10144), .ZN(P2_U3305) );
  XNOR2_X1 U13843 ( .A(n11254), .B(n12112), .ZN(n15152) );
  OR2_X1 U13844 ( .A1(n11255), .A2(n12160), .ZN(n11308) );
  OAI21_X1 U13845 ( .B1(n11256), .B2(n12112), .A(n11308), .ZN(n11258) );
  AOI21_X1 U13846 ( .B1(n11258), .B2(n12804), .A(n11257), .ZN(n15153) );
  MUX2_X1 U13847 ( .A(n11259), .B(n15153), .S(n15126), .Z(n11263) );
  INV_X1 U13848 ( .A(n11260), .ZN(n11261) );
  AOI22_X1 U13849 ( .A1(n12813), .A2(n7435), .B1(n12797), .B2(n11261), .ZN(
        n11262) );
  OAI211_X1 U13850 ( .C1(n12802), .C2(n15152), .A(n11263), .B(n11262), .ZN(
        P3_U3228) );
  XNOR2_X1 U13851 ( .A(n13237), .B(n11269), .ZN(n11267) );
  OAI22_X1 U13852 ( .A1(n13261), .A2(n13503), .B1(n12049), .B2(n13505), .ZN(
        n12046) );
  AOI21_X1 U13853 ( .B1(n11267), .B2(n13526), .A(n12046), .ZN(n13638) );
  NAND2_X1 U13854 ( .A1(n11270), .A2(n11269), .ZN(n13259) );
  OAI21_X1 U13855 ( .B1(n11270), .B2(n11269), .A(n13259), .ZN(n13639) );
  INV_X1 U13856 ( .A(n13639), .ZN(n11277) );
  AND2_X1 U13857 ( .A1(n13636), .A2(n11271), .ZN(n11272) );
  OR3_X1 U13858 ( .A1(n13511), .A2(n11272), .A3(n10602), .ZN(n13634) );
  INV_X1 U13859 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11273) );
  OAI22_X1 U13860 ( .A1(n13527), .A2(n11273), .B1(n12048), .B2(n13466), .ZN(
        n11274) );
  AOI21_X1 U13861 ( .B1(n13636), .B2(n13530), .A(n11274), .ZN(n11275) );
  OAI21_X1 U13862 ( .B1(n13634), .B2(n13515), .A(n11275), .ZN(n11276) );
  AOI21_X1 U13863 ( .B1(n11277), .B2(n13534), .A(n11276), .ZN(n11278) );
  OAI21_X1 U13864 ( .B1(n13638), .B2(n13512), .A(n11278), .ZN(P2_U3251) );
  INV_X1 U13865 ( .A(n11279), .ZN(n11280) );
  OAI222_X1 U13866 ( .A1(n11282), .A2(P3_U3151), .B1(n13004), .B2(n11281), 
        .C1(n12387), .C2(n11280), .ZN(P3_U3270) );
  XNOR2_X1 U13867 ( .A(n11283), .B(n12172), .ZN(n15163) );
  OAI211_X1 U13868 ( .C1(n11284), .C2(n12172), .A(n11362), .B(n12804), .ZN(
        n11288) );
  NAND2_X1 U13869 ( .A1(n12601), .A2(n12573), .ZN(n11286) );
  NAND2_X1 U13870 ( .A1(n12603), .A2(n12572), .ZN(n11285) );
  NAND2_X1 U13871 ( .A1(n11286), .A2(n11285), .ZN(n14969) );
  INV_X1 U13872 ( .A(n14969), .ZN(n11287) );
  NAND2_X1 U13873 ( .A1(n11288), .A2(n11287), .ZN(n15166) );
  NAND2_X1 U13874 ( .A1(n15166), .A2(n15126), .ZN(n11291) );
  OAI22_X1 U13875 ( .A1(n12841), .A2(n14962), .B1(n14971), .B2(n15121), .ZN(
        n11289) );
  AOI21_X1 U13876 ( .B1(n15128), .B2(P3_REG2_REG_7__SCAN_IN), .A(n11289), .ZN(
        n11290) );
  OAI211_X1 U13877 ( .C1(n12802), .C2(n15163), .A(n11291), .B(n11290), .ZN(
        P3_U3226) );
  XNOR2_X1 U13878 ( .A(n11292), .B(n11998), .ZN(n14683) );
  INV_X1 U13879 ( .A(n14683), .ZN(n11302) );
  INV_X1 U13880 ( .A(n11293), .ZN(n11294) );
  AOI21_X1 U13881 ( .B1(n11998), .B2(n11295), .A(n11294), .ZN(n14677) );
  XNOR2_X1 U13882 ( .A(n11296), .B(n11854), .ZN(n11297) );
  AOI222_X1 U13883 ( .A1(n13878), .A2(n14498), .B1(n14302), .B2(n11297), .C1(
        n13876), .C2(n14642), .ZN(n14678) );
  NAND2_X1 U13884 ( .A1(n14253), .A2(n6857), .ZN(n14178) );
  AOI22_X1 U13885 ( .A1(n14147), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11537), 
        .B2(n14243), .ZN(n11299) );
  NAND2_X1 U13886 ( .A1(n11854), .A2(n14246), .ZN(n11298) );
  OAI211_X1 U13887 ( .C1(n14678), .C2(n14178), .A(n11299), .B(n11298), .ZN(
        n11300) );
  AOI21_X1 U13888 ( .B1(n14677), .B2(n14180), .A(n11300), .ZN(n11301) );
  OAI21_X1 U13889 ( .B1(n11302), .B2(n14219), .A(n11301), .ZN(P1_U3283) );
  OAI21_X1 U13890 ( .B1(n11303), .B2(n11305), .A(n11304), .ZN(n15161) );
  INV_X1 U13891 ( .A(n15161), .ZN(n11317) );
  AND2_X1 U13892 ( .A1(n11308), .A2(n11306), .ZN(n11310) );
  NAND2_X1 U13893 ( .A1(n11308), .A2(n11307), .ZN(n11309) );
  OAI211_X1 U13894 ( .C1(n11310), .C2(n12114), .A(n12804), .B(n11309), .ZN(
        n11311) );
  OAI211_X1 U13895 ( .C1(n11317), .C2(n15164), .A(n11312), .B(n11311), .ZN(
        n15159) );
  NAND2_X1 U13896 ( .A1(n15159), .A2(n15126), .ZN(n11316) );
  OAI22_X1 U13897 ( .A1(n12841), .A2(n15158), .B1(n11313), .B2(n15121), .ZN(
        n11314) );
  AOI21_X1 U13898 ( .B1(n15128), .B2(P3_REG2_REG_6__SCAN_IN), .A(n11314), .ZN(
        n11315) );
  OAI211_X1 U13899 ( .C1(n11317), .C2(n12694), .A(n11316), .B(n11315), .ZN(
        P3_U3227) );
  INV_X1 U13900 ( .A(n11318), .ZN(n11322) );
  INV_X1 U13901 ( .A(n14363), .ZN(n14354) );
  NAND2_X1 U13902 ( .A1(n14354), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11319) );
  OAI211_X1 U13903 ( .C1(n11322), .C2(n14366), .A(n11319), .B(n12034), .ZN(
        P1_U3332) );
  NAND2_X1 U13904 ( .A1(n13683), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11320) );
  OAI211_X1 U13905 ( .C1(n11322), .C2(n13685), .A(n11321), .B(n11320), .ZN(
        P2_U3304) );
  INV_X1 U13906 ( .A(n11323), .ZN(n11325) );
  AOI22_X1 U13907 ( .A1(n11839), .A2(n12360), .B1(n11633), .B2(n13880), .ZN(
        n11328) );
  XNOR2_X1 U13908 ( .A(n11328), .B(n12370), .ZN(n11330) );
  AND2_X1 U13909 ( .A1(n12364), .A2(n13880), .ZN(n11329) );
  AOI21_X1 U13910 ( .B1(n11839), .B2(n11633), .A(n11329), .ZN(n11331) );
  XNOR2_X1 U13911 ( .A(n11330), .B(n11331), .ZN(n11400) );
  NAND2_X1 U13912 ( .A1(n14668), .A2(n12360), .ZN(n11333) );
  NAND2_X1 U13913 ( .A1(n13879), .A2(n11633), .ZN(n11332) );
  NAND2_X1 U13914 ( .A1(n11333), .A2(n11332), .ZN(n11334) );
  XNOR2_X1 U13915 ( .A(n11334), .B(n12343), .ZN(n11337) );
  AND2_X1 U13916 ( .A1(n12364), .A2(n13879), .ZN(n11335) );
  AOI21_X1 U13917 ( .B1(n14668), .B2(n11633), .A(n11335), .ZN(n11336) );
  NAND2_X1 U13918 ( .A1(n11337), .A2(n11336), .ZN(n11496) );
  OAI21_X1 U13919 ( .B1(n11337), .B2(n11336), .A(n11496), .ZN(n11338) );
  AOI21_X1 U13920 ( .B1(n11339), .B2(n11338), .A(n6644), .ZN(n11345) );
  NAND2_X1 U13921 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n13949) );
  NAND2_X1 U13922 ( .A1(n13805), .A2(n11340), .ZN(n11341) );
  OAI211_X1 U13923 ( .C1(n13786), .C2(n11342), .A(n13949), .B(n11341), .ZN(
        n11343) );
  AOI21_X1 U13924 ( .B1(n14668), .B2(n13817), .A(n11343), .ZN(n11344) );
  OAI21_X1 U13925 ( .B1(n11345), .B2(n13864), .A(n11344), .ZN(P1_U3221) );
  INV_X1 U13926 ( .A(n11347), .ZN(n11348) );
  OAI222_X1 U13927 ( .A1(n6664), .A2(P3_U3151), .B1(n13004), .B2(n11349), .C1(
        n12387), .C2(n11348), .ZN(P3_U3269) );
  XNOR2_X1 U13928 ( .A(n11857), .B(n13876), .ZN(n12000) );
  XNOR2_X1 U13929 ( .A(n11350), .B(n12000), .ZN(n11351) );
  OAI222_X1 U13930 ( .A1(n14522), .A2(n14521), .B1(n11351), .B2(n14661), .C1(
        n14520), .C2(n13827), .ZN(n14532) );
  INV_X1 U13931 ( .A(n14532), .ZN(n11359) );
  XOR2_X1 U13932 ( .A(n11352), .B(n12000), .Z(n14534) );
  INV_X1 U13933 ( .A(n11380), .ZN(n11353) );
  OAI211_X1 U13934 ( .C1(n14531), .C2(n11354), .A(n11353), .B(n14302), .ZN(
        n14530) );
  AOI22_X1 U13935 ( .A1(n14147), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n13830), 
        .B2(n14243), .ZN(n11356) );
  NAND2_X1 U13936 ( .A1(n11857), .A2(n14246), .ZN(n11355) );
  OAI211_X1 U13937 ( .C1(n14530), .C2(n14239), .A(n11356), .B(n11355), .ZN(
        n11357) );
  AOI21_X1 U13938 ( .B1(n14534), .B2(n14256), .A(n11357), .ZN(n11358) );
  OAI21_X1 U13939 ( .B1(n11359), .B2(n14147), .A(n11358), .ZN(P1_U3282) );
  XNOR2_X1 U13940 ( .A(n11360), .B(n12180), .ZN(n15172) );
  NAND2_X1 U13941 ( .A1(n11362), .A2(n11361), .ZN(n11363) );
  XNOR2_X1 U13942 ( .A(n11363), .B(n12180), .ZN(n11367) );
  NAND2_X1 U13943 ( .A1(n12600), .A2(n12573), .ZN(n11365) );
  NAND2_X1 U13944 ( .A1(n12602), .A2(n12572), .ZN(n11364) );
  NAND2_X1 U13945 ( .A1(n11365), .A2(n11364), .ZN(n14981) );
  INV_X1 U13946 ( .A(n14981), .ZN(n11366) );
  OAI21_X1 U13947 ( .B1(n11367), .B2(n15117), .A(n11366), .ZN(n15173) );
  NAND2_X1 U13948 ( .A1(n15173), .A2(n15126), .ZN(n11370) );
  OAI22_X1 U13949 ( .A1(n12841), .A2(n15170), .B1(n14984), .B2(n15121), .ZN(
        n11368) );
  AOI21_X1 U13950 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15128), .A(n11368), .ZN(
        n11369) );
  OAI211_X1 U13951 ( .C1(n12802), .C2(n15172), .A(n11370), .B(n11369), .ZN(
        P3_U3225) );
  XOR2_X1 U13952 ( .A(n11371), .B(n12002), .Z(n11378) );
  OAI22_X1 U13953 ( .A1(n14510), .A2(n14522), .B1(n11372), .B2(n14520), .ZN(
        n11377) );
  NAND2_X1 U13954 ( .A1(n11373), .A2(n12002), .ZN(n11374) );
  AOI21_X1 U13955 ( .B1(n11375), .B2(n11374), .A(n14672), .ZN(n11376) );
  AOI211_X1 U13956 ( .C1(n11378), .C2(n14676), .A(n11377), .B(n11376), .ZN(
        n11433) );
  INV_X1 U13957 ( .A(n13757), .ZN(n11379) );
  OAI22_X1 U13958 ( .A1(n14253), .A2(n10390), .B1(n11379), .B2(n14206), .ZN(
        n11382) );
  OAI211_X1 U13959 ( .C1(n11380), .C2(n13760), .A(n14302), .B(n11391), .ZN(
        n11432) );
  NOR2_X1 U13960 ( .A1(n11432), .A2(n14239), .ZN(n11381) );
  AOI211_X1 U13961 ( .C1(n14246), .C2(n11866), .A(n11382), .B(n11381), .ZN(
        n11383) );
  OAI21_X1 U13962 ( .B1(n11433), .B2(n14147), .A(n11383), .ZN(P1_U3281) );
  XNOR2_X1 U13963 ( .A(n11384), .B(n12004), .ZN(n11388) );
  OAI21_X1 U13964 ( .B1(n12004), .B2(n11386), .A(n11385), .ZN(n11387) );
  AOI22_X1 U13965 ( .A1(n11388), .A2(n14676), .B1(n11387), .B2(n14684), .ZN(
        n14528) );
  NAND2_X1 U13966 ( .A1(n14253), .A2(n14498), .ZN(n14210) );
  AOI22_X1 U13967 ( .A1(n14147), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n13816), 
        .B2(n14243), .ZN(n11390) );
  AND2_X1 U13968 ( .A1(n14253), .A2(n14642), .ZN(n14245) );
  NAND2_X1 U13969 ( .A1(n14245), .A2(n14499), .ZN(n11389) );
  OAI211_X1 U13970 ( .C1(n14521), .C2(n14210), .A(n11390), .B(n11389), .ZN(
        n11394) );
  AOI21_X1 U13971 ( .B1(n11391), .B2(n14525), .A(n14644), .ZN(n11392) );
  NAND2_X1 U13972 ( .A1(n11392), .A2(n11508), .ZN(n14526) );
  NOR2_X1 U13973 ( .A1(n14526), .A2(n14239), .ZN(n11393) );
  AOI211_X1 U13974 ( .C1(n14246), .C2(n14525), .A(n11394), .B(n11393), .ZN(
        n11395) );
  OAI21_X1 U13975 ( .B1(n14528), .B2(n14147), .A(n11395), .ZN(P1_U3280) );
  INV_X1 U13976 ( .A(n11396), .ZN(n11399) );
  AND2_X1 U13977 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13944) );
  AOI21_X1 U13978 ( .B1(n13855), .B2(n13882), .A(n13944), .ZN(n11398) );
  NAND2_X1 U13979 ( .A1(n13825), .A2(n13879), .ZN(n11397) );
  OAI211_X1 U13980 ( .C1(n13786), .C2(n11399), .A(n11398), .B(n11397), .ZN(
        n11404) );
  XNOR2_X1 U13981 ( .A(n11401), .B(n11400), .ZN(n11402) );
  NOR2_X1 U13982 ( .A1(n11402), .A2(n13864), .ZN(n11403) );
  AOI211_X1 U13983 ( .C1(n11839), .C2(n13817), .A(n11404), .B(n11403), .ZN(
        n11405) );
  INV_X1 U13984 ( .A(n11405), .ZN(P1_U3213) );
  AOI22_X1 U13985 ( .A1(n13122), .A2(n11406), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11407) );
  OAI21_X1 U13986 ( .B1(n11408), .B2(n14470), .A(n11407), .ZN(n11422) );
  XNOR2_X1 U13987 ( .A(n13641), .B(n11708), .ZN(n11409) );
  AND2_X1 U13988 ( .A1(n13470), .A2(n13145), .ZN(n11410) );
  NAND2_X1 U13989 ( .A1(n11409), .A2(n11410), .ZN(n11657) );
  INV_X1 U13990 ( .A(n11409), .ZN(n12050) );
  INV_X1 U13991 ( .A(n11410), .ZN(n11411) );
  NAND2_X1 U13992 ( .A1(n12050), .A2(n11411), .ZN(n11412) );
  NAND2_X1 U13993 ( .A1(n11657), .A2(n11412), .ZN(n11420) );
  INV_X1 U13994 ( .A(n11413), .ZN(n11415) );
  NAND2_X1 U13995 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  AOI211_X1 U13996 ( .C1(n11420), .C2(n11419), .A(n14462), .B(n11418), .ZN(
        n11421) );
  AOI211_X1 U13997 ( .C1(n13641), .C2(n14467), .A(n11422), .B(n11421), .ZN(
        n11423) );
  INV_X1 U13998 ( .A(n11423), .ZN(P2_U3206) );
  XNOR2_X1 U13999 ( .A(n11424), .B(n12187), .ZN(n15178) );
  INV_X1 U14000 ( .A(n12187), .ZN(n12119) );
  XNOR2_X1 U14001 ( .A(n11425), .B(n12119), .ZN(n11426) );
  NAND2_X1 U14002 ( .A1(n11426), .A2(n12804), .ZN(n11427) );
  AOI22_X1 U14003 ( .A1(n12572), .A2(n12601), .B1(n12599), .B2(n12573), .ZN(
        n11447) );
  OAI211_X1 U14004 ( .C1(n15164), .C2(n15178), .A(n11427), .B(n11447), .ZN(
        n15180) );
  NAND2_X1 U14005 ( .A1(n15180), .A2(n15126), .ZN(n11431) );
  OAI22_X1 U14006 ( .A1(n12841), .A2(n15179), .B1(n11428), .B2(n15121), .ZN(
        n11429) );
  AOI21_X1 U14007 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15128), .A(n11429), .ZN(
        n11430) );
  OAI211_X1 U14008 ( .C1(n15178), .C2(n12694), .A(n11431), .B(n11430), .ZN(
        P3_U3224) );
  AND2_X1 U14009 ( .A1(n11433), .A2(n11432), .ZN(n11438) );
  AOI22_X1 U14010 ( .A1(n11866), .A2(n9824), .B1(n14695), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11434) );
  OAI21_X1 U14011 ( .B1(n11438), .B2(n14695), .A(n11434), .ZN(P1_U3540) );
  INV_X1 U14012 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11435) );
  OAI22_X1 U14013 ( .A1(n13760), .A2(n14348), .B1(n14687), .B2(n11435), .ZN(
        n11436) );
  INV_X1 U14014 ( .A(n11436), .ZN(n11437) );
  OAI21_X1 U14015 ( .B1(n11438), .B2(n14685), .A(n11437), .ZN(P1_U3495) );
  INV_X1 U14016 ( .A(n11439), .ZN(n11541) );
  OAI222_X1 U14017 ( .A1(n13688), .A2(n11441), .B1(n13685), .B2(n11541), .C1(
        P2_U3088), .C2(n11440), .ZN(P2_U3303) );
  OR2_X1 U14018 ( .A1(n11442), .A2(n11444), .ZN(n11466) );
  INV_X1 U14019 ( .A(n11466), .ZN(n11443) );
  AOI21_X1 U14020 ( .B1(n11444), .B2(n11442), .A(n11443), .ZN(n11451) );
  NAND2_X1 U14021 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15009) );
  NAND2_X1 U14022 ( .A1(n12577), .A2(n11445), .ZN(n11446) );
  OAI211_X1 U14023 ( .C1(n11447), .C2(n12530), .A(n15009), .B(n11446), .ZN(
        n11448) );
  AOI21_X1 U14024 ( .B1(n11449), .B2(n12532), .A(n11448), .ZN(n11450) );
  OAI21_X1 U14025 ( .B1(n11451), .B2(n12579), .A(n11450), .ZN(P3_U3171) );
  XNOR2_X1 U14026 ( .A(n11452), .B(n12192), .ZN(n11458) );
  INV_X1 U14027 ( .A(n11454), .ZN(n11453) );
  OR2_X1 U14028 ( .A1(n12600), .A2(n11453), .ZN(n11456) );
  OR2_X1 U14029 ( .A1(n12598), .A2(n11454), .ZN(n11455) );
  AND3_X1 U14030 ( .A1(n11456), .A2(n11455), .A3(n12286), .ZN(n11471) );
  INV_X1 U14031 ( .A(n11471), .ZN(n11457) );
  OAI21_X1 U14032 ( .B1(n11458), .B2(n15117), .A(n11457), .ZN(n15187) );
  INV_X1 U14033 ( .A(n15187), .ZN(n11463) );
  XNOR2_X1 U14034 ( .A(n11459), .B(n12192), .ZN(n15189) );
  INV_X1 U14035 ( .A(n12802), .ZN(n12844) );
  NOR2_X1 U14036 ( .A1(n15126), .A2(n9034), .ZN(n11461) );
  OAI22_X1 U14037 ( .A1(n12841), .A2(n15186), .B1(n11474), .B2(n15121), .ZN(
        n11460) );
  AOI211_X1 U14038 ( .C1(n15189), .C2(n12844), .A(n11461), .B(n11460), .ZN(
        n11462) );
  OAI21_X1 U14039 ( .B1(n11463), .B2(n15128), .A(n11462), .ZN(P3_U3223) );
  AND2_X1 U14040 ( .A1(n11466), .A2(n11464), .ZN(n11469) );
  NAND2_X1 U14041 ( .A1(n11466), .A2(n11465), .ZN(n11467) );
  OAI211_X1 U14042 ( .C1(n11469), .C2(n11468), .A(n11467), .B(n14974), .ZN(
        n11473) );
  NAND2_X1 U14043 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n15020)
         );
  OAI21_X1 U14044 ( .B1(n14973), .B2(n15186), .A(n15020), .ZN(n11470) );
  AOI21_X1 U14045 ( .B1(n11471), .B2(n14982), .A(n11470), .ZN(n11472) );
  OAI211_X1 U14046 ( .C1(n11474), .C2(n14985), .A(n11473), .B(n11472), .ZN(
        P3_U3157) );
  INV_X1 U14047 ( .A(n11475), .ZN(n11479) );
  OAI222_X1 U14048 ( .A1(P1_U3086), .A2(n11477), .B1(n14366), .B2(n11479), 
        .C1(n11476), .C2(n14363), .ZN(P1_U3330) );
  OAI222_X1 U14049 ( .A1(n13688), .A2(n11480), .B1(n13685), .B2(n11479), .C1(
        P2_U3088), .C2(n11478), .ZN(P2_U3302) );
  OR2_X1 U14050 ( .A1(n11516), .A2(n12007), .ZN(n11515) );
  AND2_X1 U14051 ( .A1(n11515), .A2(n11481), .ZN(n11484) );
  NAND2_X1 U14052 ( .A1(n11515), .A2(n11482), .ZN(n11483) );
  OAI21_X1 U14053 ( .B1(n11484), .B2(n11986), .A(n11483), .ZN(n14508) );
  INV_X1 U14054 ( .A(n14508), .ZN(n11494) );
  AOI22_X1 U14055 ( .A1(n14147), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13861), 
        .B2(n14243), .ZN(n11486) );
  NAND2_X1 U14056 ( .A1(n14245), .A2(n14500), .ZN(n11485) );
  OAI211_X1 U14057 ( .C1(n14523), .C2(n14210), .A(n11486), .B(n11485), .ZN(
        n11490) );
  INV_X1 U14058 ( .A(n11487), .ZN(n11509) );
  AOI21_X1 U14059 ( .B1(n6670), .B2(n11509), .A(n14644), .ZN(n11488) );
  NAND2_X1 U14060 ( .A1(n11488), .A2(n14220), .ZN(n14502) );
  NOR2_X1 U14061 ( .A1(n14502), .A2(n14239), .ZN(n11489) );
  AOI211_X1 U14062 ( .C1(n14246), .C2(n6670), .A(n11490), .B(n11489), .ZN(
        n11493) );
  NAND2_X1 U14063 ( .A1(n11491), .A2(n11986), .ZN(n14504) );
  NAND3_X1 U14064 ( .A1(n14505), .A2(n14504), .A3(n14180), .ZN(n11492) );
  OAI211_X1 U14065 ( .C1(n11494), .C2(n14219), .A(n11493), .B(n11492), .ZN(
        P1_U3278) );
  AOI22_X1 U14066 ( .A1(n11849), .A2(n12360), .B1(n11633), .B2(n13878), .ZN(
        n11495) );
  XNOR2_X1 U14067 ( .A(n11495), .B(n12370), .ZN(n11499) );
  AND2_X1 U14068 ( .A1(n12364), .A2(n13878), .ZN(n11497) );
  AOI21_X1 U14069 ( .B1(n11849), .B2(n11633), .A(n11497), .ZN(n11521) );
  XNOR2_X1 U14070 ( .A(n11520), .B(n11521), .ZN(n11498) );
  NAND2_X1 U14071 ( .A1(n11498), .A2(n11499), .ZN(n11530) );
  OAI21_X1 U14072 ( .B1(n11499), .B2(n11498), .A(n11530), .ZN(n11500) );
  NAND2_X1 U14073 ( .A1(n11500), .A2(n13844), .ZN(n11506) );
  NOR2_X1 U14074 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11501), .ZN(n13965) );
  AOI21_X1 U14075 ( .B1(n13855), .B2(n13879), .A(n13965), .ZN(n11502) );
  OAI21_X1 U14076 ( .B1(n13857), .B2(n13827), .A(n11502), .ZN(n11503) );
  AOI21_X1 U14077 ( .B1(n11504), .B2(n13862), .A(n11503), .ZN(n11505) );
  OAI211_X1 U14078 ( .C1(n6970), .C2(n13858), .A(n11506), .B(n11505), .ZN(
        P1_U3231) );
  XNOR2_X1 U14079 ( .A(n11507), .B(n11870), .ZN(n14518) );
  AOI21_X1 U14080 ( .B1(n14513), .B2(n11508), .A(n14644), .ZN(n11510) );
  NAND2_X1 U14081 ( .A1(n11510), .A2(n11509), .ZN(n14514) );
  AOI22_X1 U14082 ( .A1(n14147), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n13708), 
        .B2(n14243), .ZN(n11512) );
  NAND2_X1 U14083 ( .A1(n14245), .A2(n13873), .ZN(n11511) );
  OAI211_X1 U14084 ( .C1(n14510), .C2(n14210), .A(n11512), .B(n11511), .ZN(
        n11513) );
  AOI21_X1 U14085 ( .B1(n14513), .B2(n14246), .A(n11513), .ZN(n11514) );
  OAI21_X1 U14086 ( .B1(n14514), .B2(n14239), .A(n11514), .ZN(n11518) );
  OAI21_X1 U14087 ( .B1(n6491), .B2(n11870), .A(n11515), .ZN(n14516) );
  NOR2_X1 U14088 ( .A1(n14516), .A2(n14219), .ZN(n11517) );
  AOI211_X1 U14089 ( .C1(n14180), .C2(n14518), .A(n11518), .B(n11517), .ZN(
        n11519) );
  INV_X1 U14090 ( .A(n11519), .ZN(P1_U3279) );
  NAND2_X1 U14091 ( .A1(n6739), .A2(n11521), .ZN(n11526) );
  AND2_X1 U14092 ( .A1(n11530), .A2(n11526), .ZN(n11532) );
  NAND2_X1 U14093 ( .A1(n11854), .A2(n12360), .ZN(n11523) );
  NAND2_X1 U14094 ( .A1(n13877), .A2(n11633), .ZN(n11522) );
  NAND2_X1 U14095 ( .A1(n11523), .A2(n11522), .ZN(n11524) );
  XNOR2_X1 U14096 ( .A(n11524), .B(n12370), .ZN(n11549) );
  AND2_X1 U14097 ( .A1(n12364), .A2(n13877), .ZN(n11525) );
  AOI21_X1 U14098 ( .B1(n11854), .B2(n11633), .A(n11525), .ZN(n11547) );
  XNOR2_X1 U14099 ( .A(n11549), .B(n11547), .ZN(n11531) );
  INV_X1 U14100 ( .A(n11531), .ZN(n11527) );
  OAI211_X1 U14101 ( .C1(n11532), .C2(n11531), .A(n13844), .B(n11551), .ZN(
        n11539) );
  NAND2_X1 U14102 ( .A1(n13825), .A2(n13876), .ZN(n11533) );
  OAI211_X1 U14103 ( .C1(n13828), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        n11536) );
  AOI21_X1 U14104 ( .B1(n11537), .B2(n13862), .A(n11536), .ZN(n11538) );
  OAI211_X1 U14105 ( .C1(n14681), .C2(n13858), .A(n11539), .B(n11538), .ZN(
        P1_U3217) );
  OAI222_X1 U14106 ( .A1(P1_U3086), .A2(n11542), .B1(n14366), .B2(n11541), 
        .C1(n11540), .C2(n14363), .ZN(P1_U3331) );
  NAND2_X1 U14107 ( .A1(n11857), .A2(n12360), .ZN(n11544) );
  NAND2_X1 U14108 ( .A1(n13876), .A2(n11633), .ZN(n11543) );
  NAND2_X1 U14109 ( .A1(n11544), .A2(n11543), .ZN(n11545) );
  XNOR2_X1 U14110 ( .A(n11545), .B(n12370), .ZN(n11556) );
  AND2_X1 U14111 ( .A1(n12364), .A2(n13876), .ZN(n11546) );
  AOI21_X1 U14112 ( .B1(n11857), .B2(n11633), .A(n11546), .ZN(n11557) );
  XNOR2_X1 U14113 ( .A(n11556), .B(n11557), .ZN(n13821) );
  INV_X1 U14114 ( .A(n11547), .ZN(n11548) );
  NAND2_X1 U14115 ( .A1(n11549), .A2(n11548), .ZN(n13822) );
  AND2_X1 U14116 ( .A1(n13821), .A2(n13822), .ZN(n11550) );
  NAND2_X1 U14117 ( .A1(n11866), .A2(n12360), .ZN(n11553) );
  NAND2_X1 U14118 ( .A1(n13875), .A2(n11633), .ZN(n11552) );
  NAND2_X1 U14119 ( .A1(n11553), .A2(n11552), .ZN(n11554) );
  XNOR2_X1 U14120 ( .A(n11554), .B(n12370), .ZN(n11560) );
  AND2_X1 U14121 ( .A1(n12364), .A2(n13875), .ZN(n11555) );
  AOI21_X1 U14122 ( .B1(n11866), .B2(n11633), .A(n11555), .ZN(n11561) );
  XNOR2_X1 U14123 ( .A(n11560), .B(n11561), .ZN(n13752) );
  INV_X1 U14124 ( .A(n11556), .ZN(n11558) );
  NAND2_X1 U14125 ( .A1(n11558), .A2(n11557), .ZN(n13750) );
  INV_X1 U14126 ( .A(n11560), .ZN(n11562) );
  AND2_X1 U14127 ( .A1(n12364), .A2(n13874), .ZN(n11563) );
  AOI21_X1 U14128 ( .B1(n14525), .B2(n11633), .A(n11563), .ZN(n11566) );
  AOI22_X1 U14129 ( .A1(n14525), .A2(n12360), .B1(n11633), .B2(n13874), .ZN(
        n11564) );
  XNOR2_X1 U14130 ( .A(n11564), .B(n12370), .ZN(n11565) );
  XOR2_X1 U14131 ( .A(n11566), .B(n11565), .Z(n13813) );
  INV_X1 U14132 ( .A(n11565), .ZN(n11568) );
  INV_X1 U14133 ( .A(n11566), .ZN(n11567) );
  NAND2_X1 U14134 ( .A1(n14513), .A2(n12360), .ZN(n11570) );
  NAND2_X1 U14135 ( .A1(n14499), .A2(n11633), .ZN(n11569) );
  NAND2_X1 U14136 ( .A1(n11570), .A2(n11569), .ZN(n11571) );
  XNOR2_X1 U14137 ( .A(n11571), .B(n12343), .ZN(n11574) );
  AND2_X1 U14138 ( .A1(n12364), .A2(n14499), .ZN(n11572) );
  AOI21_X1 U14139 ( .B1(n14513), .B2(n11633), .A(n11572), .ZN(n11573) );
  NAND2_X1 U14140 ( .A1(n11574), .A2(n11573), .ZN(n11577) );
  OAI21_X1 U14141 ( .B1(n11574), .B2(n11573), .A(n11577), .ZN(n13704) );
  NAND2_X1 U14142 ( .A1(n13701), .A2(n11577), .ZN(n11582) );
  AOI22_X1 U14143 ( .A1(n6670), .A2(n12360), .B1(n11633), .B2(n13873), .ZN(
        n11575) );
  XNOR2_X1 U14144 ( .A(n11575), .B(n12370), .ZN(n11581) );
  INV_X1 U14145 ( .A(n11581), .ZN(n11578) );
  OR2_X1 U14146 ( .A1(n13704), .A2(n11578), .ZN(n11576) );
  OR2_X1 U14147 ( .A1(n11578), .A2(n11577), .ZN(n11579) );
  OAI21_X1 U14148 ( .B1(n11582), .B2(n11581), .A(n11586), .ZN(n13853) );
  INV_X1 U14149 ( .A(n6670), .ZN(n14503) );
  INV_X1 U14150 ( .A(n11584), .ZN(n11636) );
  OAI22_X1 U14151 ( .A1(n14503), .A2(n11636), .B1(n14511), .B2(n11585), .ZN(
        n13854) );
  NAND2_X1 U14152 ( .A1(n14236), .A2(n12360), .ZN(n11588) );
  NAND2_X1 U14153 ( .A1(n14500), .A2(n11633), .ZN(n11587) );
  NAND2_X1 U14154 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  XNOR2_X1 U14155 ( .A(n11589), .B(n12370), .ZN(n11593) );
  NAND2_X1 U14156 ( .A1(n14236), .A2(n11633), .ZN(n11591) );
  NAND2_X1 U14157 ( .A1(n12364), .A2(n14500), .ZN(n11590) );
  NAND2_X1 U14158 ( .A1(n11591), .A2(n11590), .ZN(n11592) );
  NOR2_X1 U14159 ( .A1(n11593), .A2(n11592), .ZN(n13781) );
  AOI21_X1 U14160 ( .B1(n11593), .B2(n11592), .A(n13781), .ZN(n13774) );
  INV_X1 U14161 ( .A(n13781), .ZN(n11594) );
  NAND2_X1 U14162 ( .A1(n14213), .A2(n12360), .ZN(n11596) );
  NAND2_X1 U14163 ( .A1(n13872), .A2(n11633), .ZN(n11595) );
  NAND2_X1 U14164 ( .A1(n11596), .A2(n11595), .ZN(n11597) );
  XNOR2_X1 U14165 ( .A(n11597), .B(n12343), .ZN(n11599) );
  AND2_X1 U14166 ( .A1(n12364), .A2(n13872), .ZN(n11598) );
  AOI21_X1 U14167 ( .B1(n14213), .B2(n11633), .A(n11598), .ZN(n11600) );
  NAND2_X1 U14168 ( .A1(n11599), .A2(n11600), .ZN(n13724) );
  INV_X1 U14169 ( .A(n11599), .ZN(n11602) );
  INV_X1 U14170 ( .A(n11600), .ZN(n11601) );
  NAND2_X1 U14171 ( .A1(n11602), .A2(n11601), .ZN(n11603) );
  AOI22_X1 U14172 ( .A1(n8544), .A2(n12360), .B1(n11633), .B2(n14199), .ZN(
        n11604) );
  XNOR2_X1 U14173 ( .A(n11604), .B(n12370), .ZN(n11617) );
  AND2_X1 U14174 ( .A1(n14199), .A2(n12364), .ZN(n11605) );
  AOI21_X1 U14175 ( .B1(n8544), .B2(n11633), .A(n11605), .ZN(n11618) );
  XNOR2_X1 U14176 ( .A(n11617), .B(n11618), .ZN(n13725) );
  NAND2_X1 U14177 ( .A1(n14182), .A2(n12360), .ZN(n11607) );
  NAND2_X1 U14178 ( .A1(n14485), .A2(n11633), .ZN(n11606) );
  NAND2_X1 U14179 ( .A1(n11607), .A2(n11606), .ZN(n11608) );
  XNOR2_X1 U14180 ( .A(n11608), .B(n12370), .ZN(n11611) );
  AOI22_X1 U14181 ( .A1(n14182), .A2(n11633), .B1(n12364), .B2(n14485), .ZN(
        n11610) );
  INV_X1 U14182 ( .A(n11610), .ZN(n11609) );
  NOR2_X1 U14183 ( .A1(n11611), .A2(n11609), .ZN(n13726) );
  NOR2_X1 U14184 ( .A1(n13725), .A2(n13726), .ZN(n11614) );
  INV_X1 U14185 ( .A(n11614), .ZN(n11612) );
  XNOR2_X1 U14186 ( .A(n11611), .B(n11610), .ZN(n13835) );
  OR2_X1 U14187 ( .A1(n11612), .A2(n13835), .ZN(n11613) );
  INV_X1 U14188 ( .A(n11613), .ZN(n11616) );
  AND2_X1 U14189 ( .A1(n13724), .A2(n11614), .ZN(n11615) );
  INV_X1 U14190 ( .A(n11617), .ZN(n11620) );
  INV_X1 U14191 ( .A(n11618), .ZN(n11619) );
  NAND2_X1 U14192 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U14193 ( .A1(n13728), .A2(n11621), .ZN(n13802) );
  NAND2_X1 U14194 ( .A1(n14160), .A2(n12360), .ZN(n11623) );
  NAND2_X1 U14195 ( .A1(n14317), .A2(n11633), .ZN(n11622) );
  NAND2_X1 U14196 ( .A1(n11623), .A2(n11622), .ZN(n11624) );
  XNOR2_X1 U14197 ( .A(n11624), .B(n12370), .ZN(n11627) );
  AOI22_X1 U14198 ( .A1(n14160), .A2(n11633), .B1(n12364), .B2(n14317), .ZN(
        n11625) );
  XNOR2_X1 U14199 ( .A(n11627), .B(n11625), .ZN(n13801) );
  INV_X1 U14200 ( .A(n11625), .ZN(n11626) );
  NAND2_X1 U14201 ( .A1(n11627), .A2(n11626), .ZN(n11628) );
  NAND2_X1 U14202 ( .A1(n14301), .A2(n12360), .ZN(n11630) );
  NAND2_X1 U14203 ( .A1(n14152), .A2(n11633), .ZN(n11629) );
  NAND2_X1 U14204 ( .A1(n11630), .A2(n11629), .ZN(n11631) );
  XNOR2_X1 U14205 ( .A(n11631), .B(n12343), .ZN(n11635) );
  AND2_X1 U14206 ( .A1(n14152), .A2(n12364), .ZN(n11632) );
  AOI21_X1 U14207 ( .B1(n14301), .B2(n11633), .A(n11632), .ZN(n11634) );
  NAND2_X1 U14208 ( .A1(n11635), .A2(n11634), .ZN(n11646) );
  OAI21_X1 U14209 ( .B1(n11635), .B2(n11634), .A(n11646), .ZN(n13742) );
  OAI22_X1 U14210 ( .A1(n14295), .A2(n11638), .B1(n11637), .B2(n11636), .ZN(
        n11639) );
  XNOR2_X1 U14211 ( .A(n11639), .B(n12343), .ZN(n11641) );
  AND2_X1 U14212 ( .A1(n14134), .A2(n12364), .ZN(n11640) );
  AOI21_X1 U14213 ( .B1(n14123), .B2(n11633), .A(n11640), .ZN(n11642) );
  NAND2_X1 U14214 ( .A1(n11641), .A2(n11642), .ZN(n13712) );
  INV_X1 U14215 ( .A(n11641), .ZN(n11644) );
  INV_X1 U14216 ( .A(n11642), .ZN(n11643) );
  NAND2_X1 U14217 ( .A1(n11644), .A2(n11643), .ZN(n11645) );
  NOR3_X1 U14218 ( .A1(n6532), .A2(n7331), .A3(n11647), .ZN(n11649) );
  INV_X1 U14219 ( .A(n12322), .ZN(n13715) );
  OAI21_X1 U14220 ( .B1(n11649), .B2(n13715), .A(n13844), .ZN(n11654) );
  AOI22_X1 U14221 ( .A1(n14152), .A2(n14498), .B1(n14642), .B2(n14079), .ZN(
        n14294) );
  INV_X1 U14222 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n11650) );
  OAI22_X1 U14223 ( .A1(n14294), .A2(n13847), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11650), .ZN(n11651) );
  AOI21_X1 U14224 ( .B1(n11652), .B2(n13862), .A(n11651), .ZN(n11653) );
  OAI211_X1 U14225 ( .C1(n13858), .C2(n14295), .A(n11654), .B(n11653), .ZN(
        P1_U3235) );
  INV_X1 U14226 ( .A(n11655), .ZN(n14361) );
  OAI222_X1 U14227 ( .A1(n13685), .A2(n14361), .B1(n8240), .B2(P2_U3088), .C1(
        n11656), .C2(n13688), .ZN(P2_U3300) );
  XNOR2_X1 U14228 ( .A(n13636), .B(n11708), .ZN(n11660) );
  NAND2_X1 U14229 ( .A1(n13257), .A2(n10857), .ZN(n11661) );
  XNOR2_X1 U14230 ( .A(n11660), .B(n11661), .ZN(n12052) );
  INV_X1 U14231 ( .A(n11660), .ZN(n11662) );
  NAND2_X1 U14232 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  XNOR2_X1 U14233 ( .A(n13629), .B(n11730), .ZN(n11666) );
  NOR2_X1 U14234 ( .A1(n13261), .A2(n13510), .ZN(n11664) );
  INV_X1 U14235 ( .A(n11665), .ZN(n11667) );
  NAND2_X1 U14236 ( .A1(n11667), .A2(n11666), .ZN(n11668) );
  XNOR2_X1 U14237 ( .A(n13485), .B(n11730), .ZN(n13054) );
  NAND2_X1 U14238 ( .A1(n13264), .A2(n10857), .ZN(n11669) );
  XNOR2_X1 U14239 ( .A(n13054), .B(n11669), .ZN(n13044) );
  NAND2_X1 U14240 ( .A1(n13054), .A2(n11669), .ZN(n11670) );
  NAND2_X1 U14241 ( .A1(n13057), .A2(n11670), .ZN(n11671) );
  XNOR2_X1 U14242 ( .A(n13618), .B(n11708), .ZN(n11672) );
  NAND2_X1 U14243 ( .A1(n13481), .A2(n10857), .ZN(n11673) );
  XNOR2_X1 U14244 ( .A(n11672), .B(n11673), .ZN(n13053) );
  NAND2_X1 U14245 ( .A1(n11671), .A2(n13053), .ZN(n13060) );
  INV_X1 U14246 ( .A(n11672), .ZN(n11674) );
  NAND2_X1 U14247 ( .A1(n11674), .A2(n11673), .ZN(n11675) );
  NAND2_X1 U14248 ( .A1(n13060), .A2(n11675), .ZN(n13112) );
  XNOR2_X1 U14249 ( .A(n13612), .B(n10851), .ZN(n11683) );
  AND2_X1 U14250 ( .A1(n13267), .A2(n13470), .ZN(n11676) );
  NAND2_X1 U14251 ( .A1(n11683), .A2(n11676), .ZN(n11681) );
  INV_X1 U14252 ( .A(n11683), .ZN(n11678) );
  INV_X1 U14253 ( .A(n11676), .ZN(n11677) );
  NAND2_X1 U14254 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  NAND2_X1 U14255 ( .A1(n11681), .A2(n11679), .ZN(n13111) );
  XNOR2_X1 U14256 ( .A(n13608), .B(n10851), .ZN(n11706) );
  NAND2_X1 U14257 ( .A1(n13270), .A2(n10857), .ZN(n11707) );
  XNOR2_X1 U14258 ( .A(n11706), .B(n11707), .ZN(n11685) );
  AND2_X1 U14259 ( .A1(n11685), .A2(n11681), .ZN(n11682) );
  NAND3_X1 U14260 ( .A1(n11683), .A2(n13097), .A3(n13267), .ZN(n11684) );
  OAI21_X1 U14261 ( .B1(n13109), .B2(n14462), .A(n11684), .ZN(n11687) );
  INV_X1 U14262 ( .A(n11685), .ZN(n11686) );
  NAND2_X1 U14263 ( .A1(n11687), .A2(n11686), .ZN(n11693) );
  NOR2_X1 U14264 ( .A1(n14470), .A2(n13439), .ZN(n11691) );
  AND2_X1 U14265 ( .A1(n13267), .A2(n13523), .ZN(n11688) );
  AOI21_X1 U14266 ( .B1(n13271), .B2(n13521), .A(n11688), .ZN(n13435) );
  OAI22_X1 U14267 ( .A1(n13435), .A2(n13101), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11689), .ZN(n11690) );
  AOI211_X1 U14268 ( .C1(n13608), .C2(n14467), .A(n11691), .B(n11690), .ZN(
        n11692) );
  OAI211_X1 U14269 ( .C1(n13090), .C2(n14462), .A(n11693), .B(n11692), .ZN(
        P2_U3191) );
  INV_X1 U14270 ( .A(n11694), .ZN(n11696) );
  AOI22_X1 U14271 ( .A1(n13136), .A2(n13148), .B1(n13135), .B2(n13151), .ZN(
        n11695) );
  NAND2_X1 U14272 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14770) );
  OAI211_X1 U14273 ( .C1(n11696), .C2(n14470), .A(n11695), .B(n14770), .ZN(
        n11702) );
  INV_X1 U14274 ( .A(n12072), .ZN(n11700) );
  AOI22_X1 U14275 ( .A1(n11697), .A2(n13126), .B1(n13097), .B2(n13151), .ZN(
        n11699) );
  NOR3_X1 U14276 ( .A1(n11700), .A2(n11699), .A3(n11698), .ZN(n11701) );
  AOI211_X1 U14277 ( .C1(n11703), .C2(n14467), .A(n11702), .B(n11701), .ZN(
        n11704) );
  OAI21_X1 U14278 ( .B1(n14462), .B2(n11705), .A(n11704), .ZN(P2_U3203) );
  NAND2_X1 U14279 ( .A1(n13347), .A2(n10602), .ZN(n11726) );
  INV_X1 U14280 ( .A(n11726), .ZN(n11728) );
  XNOR2_X1 U14281 ( .A(n13578), .B(n11708), .ZN(n11727) );
  INV_X1 U14282 ( .A(n11706), .ZN(n13087) );
  XNOR2_X1 U14283 ( .A(n13602), .B(n11708), .ZN(n11710) );
  NAND2_X1 U14284 ( .A1(n13271), .A2(n13470), .ZN(n11711) );
  XNOR2_X1 U14285 ( .A(n11710), .B(n11711), .ZN(n13086) );
  INV_X1 U14286 ( .A(n11710), .ZN(n11712) );
  NAND2_X1 U14287 ( .A1(n11712), .A2(n11711), .ZN(n11713) );
  XNOR2_X1 U14288 ( .A(n13597), .B(n10851), .ZN(n11714) );
  AND2_X1 U14289 ( .A1(n13274), .A2(n13470), .ZN(n11715) );
  NAND2_X1 U14290 ( .A1(n11714), .A2(n11715), .ZN(n11720) );
  INV_X1 U14291 ( .A(n11714), .ZN(n11717) );
  INV_X1 U14292 ( .A(n11715), .ZN(n11716) );
  NAND2_X1 U14293 ( .A1(n11717), .A2(n11716), .ZN(n11718) );
  NAND2_X1 U14294 ( .A1(n11720), .A2(n11718), .ZN(n13026) );
  NAND2_X1 U14295 ( .A1(n13028), .A2(n11720), .ZN(n11721) );
  XNOR2_X1 U14296 ( .A(n13591), .B(n10851), .ZN(n11722) );
  NAND2_X1 U14297 ( .A1(n11721), .A2(n11722), .ZN(n13094) );
  NAND2_X1 U14298 ( .A1(n13278), .A2(n10602), .ZN(n13096) );
  NAND2_X1 U14299 ( .A1(n13094), .A2(n13096), .ZN(n11725) );
  INV_X1 U14300 ( .A(n11721), .ZN(n11724) );
  INV_X1 U14301 ( .A(n11722), .ZN(n11723) );
  NAND2_X1 U14302 ( .A1(n11724), .A2(n11723), .ZN(n13095) );
  XNOR2_X1 U14303 ( .A(n11727), .B(n11726), .ZN(n13062) );
  NAND2_X1 U14304 ( .A1(n13063), .A2(n13062), .ZN(n13061) );
  XNOR2_X1 U14305 ( .A(n13572), .B(n11708), .ZN(n13117) );
  AND2_X1 U14306 ( .A1(n13470), .A2(n13282), .ZN(n11729) );
  NAND2_X1 U14307 ( .A1(n13117), .A2(n11729), .ZN(n11731) );
  OAI21_X1 U14308 ( .B1(n13117), .B2(n11729), .A(n11731), .ZN(n13037) );
  XNOR2_X1 U14309 ( .A(n13566), .B(n11730), .ZN(n11735) );
  NAND2_X1 U14310 ( .A1(n13470), .A2(n13346), .ZN(n11734) );
  XNOR2_X1 U14311 ( .A(n11735), .B(n11734), .ZN(n13120) );
  INV_X1 U14312 ( .A(n11731), .ZN(n11732) );
  XNOR2_X1 U14313 ( .A(n13319), .B(n10851), .ZN(n11737) );
  NAND2_X1 U14314 ( .A1(n13249), .A2(n10602), .ZN(n11736) );
  NOR2_X1 U14315 ( .A1(n11737), .A2(n11736), .ZN(n11744) );
  AOI21_X1 U14316 ( .B1(n11737), .B2(n11736), .A(n11744), .ZN(n13011) );
  INV_X1 U14317 ( .A(n13010), .ZN(n11739) );
  NOR3_X1 U14318 ( .A1(n11737), .A2(n13284), .A3(n13132), .ZN(n11738) );
  AOI21_X1 U14319 ( .B1(n11739), .B2(n13126), .A(n11738), .ZN(n11752) );
  NOR2_X1 U14320 ( .A1(n11740), .A2(n13510), .ZN(n11741) );
  XNOR2_X1 U14321 ( .A(n11742), .B(n11741), .ZN(n11743) );
  XNOR2_X1 U14322 ( .A(n13308), .B(n11743), .ZN(n11751) );
  INV_X1 U14323 ( .A(n11744), .ZN(n11745) );
  NAND4_X1 U14324 ( .A1(n13010), .A2(n13126), .A3(n11745), .A4(n11751), .ZN(
        n11750) );
  OAI22_X1 U14325 ( .A1(n13284), .A2(n13505), .B1(n11746), .B2(n13503), .ZN(
        n13300) );
  AOI22_X1 U14326 ( .A1(n13122), .A2(n13300), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11747) );
  OAI21_X1 U14327 ( .B1(n13303), .B2(n14470), .A(n11747), .ZN(n11748) );
  AOI21_X1 U14328 ( .B1(n13555), .B2(n14467), .A(n11748), .ZN(n11749) );
  OAI211_X1 U14329 ( .C1(n11752), .C2(n11751), .A(n11750), .B(n11749), .ZN(
        P2_U3192) );
  NAND2_X1 U14330 ( .A1(n11754), .A2(n11753), .ZN(n12260) );
  XOR2_X1 U14331 ( .A(n12260), .B(n11755), .Z(n11771) );
  XOR2_X1 U14332 ( .A(n12260), .B(n9705), .Z(n11760) );
  OR2_X1 U14333 ( .A1(n12427), .A2(n12550), .ZN(n11758) );
  NAND2_X1 U14334 ( .A1(n12585), .A2(n12572), .ZN(n11757) );
  NAND2_X1 U14335 ( .A1(n11758), .A2(n11757), .ZN(n12560) );
  INV_X1 U14336 ( .A(n12560), .ZN(n11759) );
  OAI21_X1 U14337 ( .B1(n11760), .B2(n15117), .A(n11759), .ZN(n11766) );
  AOI21_X1 U14338 ( .B1(n15167), .B2(n12559), .A(n11766), .ZN(n11763) );
  MUX2_X1 U14339 ( .A(n11761), .B(n11763), .S(n15193), .Z(n11762) );
  OAI21_X1 U14340 ( .B1(n11771), .B2(n12981), .A(n11762), .ZN(P3_U3453) );
  INV_X1 U14341 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n11764) );
  MUX2_X1 U14342 ( .A(n11764), .B(n11763), .S(n15205), .Z(n11765) );
  OAI21_X1 U14343 ( .B1(n12899), .B2(n11771), .A(n11765), .ZN(P3_U3485) );
  NAND2_X1 U14344 ( .A1(n11766), .A2(n15126), .ZN(n11770) );
  OAI22_X1 U14345 ( .A1(n15126), .A2(n11767), .B1(n12563), .B2(n15121), .ZN(
        n11768) );
  AOI21_X1 U14346 ( .B1(n12559), .B2(n12813), .A(n11768), .ZN(n11769) );
  OAI211_X1 U14347 ( .C1(n12802), .C2(n11771), .A(n11770), .B(n11769), .ZN(
        P3_U3207) );
  NAND2_X1 U14348 ( .A1(n12666), .A2(n11776), .ZN(n11777) );
  INV_X1 U14349 ( .A(n12860), .ZN(n11788) );
  OR2_X1 U14350 ( .A1(n12403), .A2(n12548), .ZN(n11782) );
  OR2_X1 U14351 ( .A1(n12269), .A2(n12550), .ZN(n11781) );
  NAND2_X1 U14352 ( .A1(n11782), .A2(n11781), .ZN(n12468) );
  NAND2_X1 U14353 ( .A1(n12859), .A2(n15126), .ZN(n11787) );
  OAI22_X1 U14354 ( .A1(n15126), .A2(n11784), .B1(n12470), .B2(n15121), .ZN(
        n11785) );
  AOI21_X1 U14355 ( .B1(n12858), .B2(n12813), .A(n11785), .ZN(n11786) );
  OAI211_X1 U14356 ( .C1(n11788), .C2(n12694), .A(n11787), .B(n11786), .ZN(
        P3_U3208) );
  NAND2_X1 U14357 ( .A1(n11789), .A2(n11977), .ZN(n11790) );
  NAND2_X1 U14358 ( .A1(n11796), .A2(n11790), .ZN(n11797) );
  NAND2_X1 U14359 ( .A1(n11791), .A2(n14106), .ZN(n11792) );
  MUX2_X1 U14360 ( .A(n11797), .B(n11796), .S(n11952), .Z(n11799) );
  MUX2_X1 U14361 ( .A(n11802), .B(n11800), .S(n11835), .Z(n11798) );
  NAND2_X1 U14362 ( .A1(n11799), .A2(n11798), .ZN(n11807) );
  OAI21_X1 U14363 ( .B1(n11802), .B2(n11952), .A(n11801), .ZN(n11803) );
  INV_X1 U14364 ( .A(n11803), .ZN(n11804) );
  NAND2_X1 U14365 ( .A1(n11807), .A2(n11806), .ZN(n11814) );
  NAND2_X1 U14366 ( .A1(n8319), .A2(n11835), .ZN(n11811) );
  NAND2_X1 U14367 ( .A1(n11808), .A2(n11952), .ZN(n11810) );
  MUX2_X1 U14368 ( .A(n11811), .B(n11810), .S(n11809), .Z(n11813) );
  NAND3_X1 U14369 ( .A1(n11814), .A2(n11813), .A3(n11812), .ZN(n11821) );
  NAND2_X1 U14370 ( .A1(n11822), .A2(n13884), .ZN(n11815) );
  NAND3_X1 U14371 ( .A1(n11821), .A2(n11820), .A3(n11819), .ZN(n11827) );
  OAI21_X1 U14372 ( .B1(n13884), .B2(n11961), .A(n14652), .ZN(n11825) );
  NAND2_X1 U14373 ( .A1(n13884), .A2(n11961), .ZN(n11823) );
  NAND2_X1 U14374 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  NAND2_X1 U14375 ( .A1(n11825), .A2(n11824), .ZN(n11826) );
  INV_X1 U14376 ( .A(n11828), .ZN(n11831) );
  MUX2_X1 U14377 ( .A(n13883), .B(n11829), .S(n11952), .Z(n11830) );
  OAI21_X1 U14378 ( .B1(n11832), .B2(n11831), .A(n11830), .ZN(n11834) );
  NAND2_X1 U14379 ( .A1(n11832), .A2(n11831), .ZN(n11833) );
  NAND2_X1 U14380 ( .A1(n11834), .A2(n11833), .ZN(n11838) );
  MUX2_X1 U14381 ( .A(n13882), .B(n11836), .S(n11835), .Z(n11837) );
  MUX2_X1 U14382 ( .A(n13880), .B(n11839), .S(n11961), .Z(n11842) );
  MUX2_X1 U14383 ( .A(n13880), .B(n11839), .S(n11952), .Z(n11840) );
  NAND2_X1 U14384 ( .A1(n11841), .A2(n11840), .ZN(n11845) );
  INV_X1 U14385 ( .A(n11842), .ZN(n11843) );
  NAND2_X1 U14386 ( .A1(n6582), .A2(n11843), .ZN(n11844) );
  MUX2_X1 U14387 ( .A(n13879), .B(n14668), .S(n11952), .Z(n11847) );
  MUX2_X1 U14388 ( .A(n13879), .B(n14668), .S(n11835), .Z(n11846) );
  INV_X1 U14389 ( .A(n11847), .ZN(n11848) );
  MUX2_X1 U14390 ( .A(n13878), .B(n11849), .S(n11835), .Z(n11852) );
  MUX2_X1 U14391 ( .A(n13878), .B(n11849), .S(n11952), .Z(n11850) );
  INV_X1 U14392 ( .A(n11852), .ZN(n11853) );
  MUX2_X1 U14393 ( .A(n13877), .B(n11854), .S(n11952), .Z(n11856) );
  MUX2_X1 U14395 ( .A(n13877), .B(n11854), .S(n11961), .Z(n11855) );
  MUX2_X1 U14396 ( .A(n13876), .B(n11857), .S(n11961), .Z(n11861) );
  NAND2_X1 U14397 ( .A1(n11860), .A2(n11861), .ZN(n11859) );
  MUX2_X1 U14398 ( .A(n13876), .B(n11857), .S(n11952), .Z(n11858) );
  NAND2_X1 U14399 ( .A1(n11859), .A2(n11858), .ZN(n11865) );
  INV_X1 U14400 ( .A(n11860), .ZN(n11863) );
  INV_X1 U14401 ( .A(n11861), .ZN(n11862) );
  NAND2_X1 U14402 ( .A1(n11863), .A2(n11862), .ZN(n11864) );
  MUX2_X1 U14403 ( .A(n13875), .B(n11866), .S(n11952), .Z(n11869) );
  MUX2_X1 U14404 ( .A(n13875), .B(n11866), .S(n11961), .Z(n11867) );
  MUX2_X1 U14405 ( .A(n13874), .B(n14525), .S(n11961), .Z(n11875) );
  OR2_X1 U14406 ( .A1(n11870), .A2(n11875), .ZN(n11873) );
  AND2_X1 U14407 ( .A1(n11886), .A2(n11871), .ZN(n11872) );
  NAND2_X1 U14408 ( .A1(n11874), .A2(n11881), .ZN(n11885) );
  NAND2_X1 U14409 ( .A1(n11876), .A2(n11875), .ZN(n11879) );
  AND2_X1 U14410 ( .A1(n11881), .A2(n13874), .ZN(n11877) );
  MUX2_X1 U14411 ( .A(n14525), .B(n11877), .S(n11961), .Z(n11878) );
  NAND3_X1 U14412 ( .A1(n11879), .A2(n12007), .A3(n11878), .ZN(n11884) );
  NAND2_X1 U14413 ( .A1(n11881), .A2(n11880), .ZN(n11882) );
  NAND2_X1 U14414 ( .A1(n11882), .A2(n11952), .ZN(n11883) );
  MUX2_X1 U14415 ( .A(n14500), .B(n14236), .S(n11961), .Z(n11902) );
  NOR2_X1 U14416 ( .A1(n14500), .A2(n11952), .ZN(n11894) );
  AOI21_X1 U14417 ( .B1(n11902), .B2(n13872), .A(n11894), .ZN(n11892) );
  NAND2_X1 U14418 ( .A1(n13872), .A2(n11952), .ZN(n11899) );
  OR2_X1 U14419 ( .A1(n14236), .A2(n11899), .ZN(n11888) );
  NOR2_X1 U14420 ( .A1(n13872), .A2(n11952), .ZN(n11895) );
  INV_X1 U14421 ( .A(n14500), .ZN(n14209) );
  NAND2_X1 U14422 ( .A1(n11895), .A2(n14209), .ZN(n11887) );
  AND2_X1 U14423 ( .A1(n11888), .A2(n11887), .ZN(n11903) );
  NAND2_X1 U14424 ( .A1(n11902), .A2(n14233), .ZN(n11889) );
  OR2_X1 U14425 ( .A1(n14236), .A2(n11961), .ZN(n11898) );
  NAND2_X1 U14426 ( .A1(n11889), .A2(n11898), .ZN(n11890) );
  NAND2_X1 U14427 ( .A1(n11890), .A2(n14488), .ZN(n11891) );
  OAI211_X1 U14428 ( .C1(n11892), .C2(n14488), .A(n11903), .B(n11891), .ZN(
        n11893) );
  NAND2_X1 U14429 ( .A1(n11902), .A2(n11894), .ZN(n11897) );
  INV_X1 U14430 ( .A(n11895), .ZN(n11896) );
  AOI21_X1 U14431 ( .B1(n11897), .B2(n11896), .A(n14488), .ZN(n11907) );
  INV_X1 U14432 ( .A(n11898), .ZN(n11901) );
  INV_X1 U14433 ( .A(n11899), .ZN(n11900) );
  AOI21_X1 U14434 ( .B1(n11902), .B2(n11901), .A(n11900), .ZN(n11905) );
  INV_X1 U14435 ( .A(n11902), .ZN(n11904) );
  OAI22_X1 U14436 ( .A1(n11905), .A2(n14213), .B1(n11904), .B2(n11903), .ZN(
        n11906) );
  MUX2_X1 U14437 ( .A(n11909), .B(n11908), .S(n11961), .Z(n11910) );
  OR3_X1 U14438 ( .A1(n14182), .A2(n11952), .A3(n14175), .ZN(n11912) );
  NAND3_X1 U14439 ( .A1(n14182), .A2(n11952), .A3(n14175), .ZN(n11911) );
  AND2_X1 U14440 ( .A1(n11912), .A2(n11911), .ZN(n11913) );
  NOR2_X1 U14441 ( .A1(n14168), .A2(n11913), .ZN(n11914) );
  INV_X1 U14442 ( .A(n14160), .ZN(n14349) );
  MUX2_X1 U14443 ( .A(n11917), .B(n14349), .S(n11961), .Z(n11919) );
  MUX2_X1 U14444 ( .A(n14317), .B(n14160), .S(n11952), .Z(n11918) );
  NAND2_X1 U14445 ( .A1(n11922), .A2(n11921), .ZN(n11924) );
  MUX2_X1 U14446 ( .A(n14152), .B(n14301), .S(n11952), .Z(n11925) );
  MUX2_X1 U14447 ( .A(n14152), .B(n14301), .S(n11961), .Z(n11923) );
  INV_X1 U14448 ( .A(n11925), .ZN(n11926) );
  MUX2_X1 U14449 ( .A(n14134), .B(n14123), .S(n11961), .Z(n11928) );
  MUX2_X1 U14450 ( .A(n14134), .B(n14123), .S(n11952), .Z(n11927) );
  MUX2_X1 U14451 ( .A(n14079), .B(n14289), .S(n11952), .Z(n11931) );
  MUX2_X1 U14452 ( .A(n14079), .B(n14289), .S(n11961), .Z(n11929) );
  MUX2_X1 U14453 ( .A(n14112), .B(n14087), .S(n11835), .Z(n11935) );
  MUX2_X1 U14454 ( .A(n14112), .B(n14087), .S(n11952), .Z(n11932) );
  NAND2_X1 U14455 ( .A1(n11933), .A2(n11932), .ZN(n11939) );
  INV_X1 U14456 ( .A(n11934), .ZN(n11937) );
  INV_X1 U14457 ( .A(n11935), .ZN(n11936) );
  NAND2_X1 U14458 ( .A1(n11937), .A2(n11936), .ZN(n11938) );
  MUX2_X1 U14459 ( .A(n14078), .B(n14058), .S(n11952), .Z(n11941) );
  MUX2_X1 U14460 ( .A(n14078), .B(n14058), .S(n11835), .Z(n11940) );
  INV_X1 U14461 ( .A(n11941), .ZN(n11942) );
  MUX2_X1 U14462 ( .A(n13871), .B(n14046), .S(n11835), .Z(n11944) );
  MUX2_X1 U14463 ( .A(n13871), .B(n14046), .S(n11952), .Z(n11943) );
  INV_X1 U14464 ( .A(n11944), .ZN(n11945) );
  MUX2_X1 U14465 ( .A(n13870), .B(n14033), .S(n11952), .Z(n11948) );
  MUX2_X1 U14466 ( .A(n13870), .B(n14033), .S(n11835), .Z(n11946) );
  INV_X1 U14467 ( .A(n11948), .ZN(n11949) );
  MUX2_X1 U14468 ( .A(n13869), .B(n12382), .S(n11835), .Z(n11950) );
  MUX2_X1 U14469 ( .A(n13868), .B(n12308), .S(n11952), .Z(n11953) );
  MUX2_X1 U14470 ( .A(n13868), .B(n12308), .S(n11961), .Z(n11954) );
  NAND2_X1 U14471 ( .A1(n11972), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U14472 ( .A1(n6470), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U14473 ( .A1(n8647), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U14474 ( .A1(n8570), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11957) );
  AND3_X1 U14475 ( .A1(n11959), .A2(n11958), .A3(n11957), .ZN(n14023) );
  OAI22_X1 U14476 ( .A1(n14023), .A2(n11961), .B1(n11960), .B2(n6650), .ZN(
        n11962) );
  AOI22_X1 U14477 ( .A1(n11985), .A2(n11835), .B1(n13867), .B2(n11962), .ZN(
        n11966) );
  NAND2_X1 U14478 ( .A1(n11965), .A2(n11966), .ZN(n11970) );
  INV_X1 U14479 ( .A(n14023), .ZN(n13866) );
  OAI21_X1 U14480 ( .B1(n13866), .B2(n11963), .A(n13867), .ZN(n11964) );
  MUX2_X1 U14481 ( .A(n14333), .B(n11964), .S(n11835), .Z(n11969) );
  INV_X1 U14482 ( .A(n11965), .ZN(n11968) );
  INV_X1 U14483 ( .A(n11966), .ZN(n11967) );
  NAND2_X1 U14484 ( .A1(n13670), .A2(n11971), .ZN(n11974) );
  NAND2_X1 U14485 ( .A1(n11972), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11973) );
  XNOR2_X1 U14486 ( .A(n14019), .B(n14023), .ZN(n12021) );
  OR2_X1 U14487 ( .A1(n11976), .A2(n11975), .ZN(n11979) );
  NAND2_X1 U14488 ( .A1(n11977), .A2(n14106), .ZN(n11978) );
  NAND2_X1 U14489 ( .A1(n11979), .A2(n11978), .ZN(n12024) );
  NOR3_X1 U14490 ( .A1(n11984), .A2(n12021), .A3(n12024), .ZN(n12030) );
  NOR2_X1 U14491 ( .A1(n14019), .A2(n14023), .ZN(n11981) );
  AND2_X1 U14492 ( .A1(n14019), .A2(n14023), .ZN(n11980) );
  MUX2_X1 U14493 ( .A(n11981), .B(n11980), .S(n11952), .Z(n12022) );
  INV_X1 U14494 ( .A(n12022), .ZN(n11983) );
  INV_X1 U14495 ( .A(n11982), .ZN(n12026) );
  XOR2_X1 U14496 ( .A(n13867), .B(n11985), .Z(n12019) );
  NOR4_X1 U14497 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11994) );
  NAND4_X1 U14498 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n11995) );
  NOR4_X1 U14499 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n12001) );
  NAND4_X1 U14500 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12003) );
  NOR3_X1 U14501 ( .A1(n14204), .A2(n12004), .A3(n12003), .ZN(n12006) );
  NAND4_X1 U14502 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12009) );
  NOR4_X1 U14503 ( .A1(n14161), .A2(n14186), .A3(n14168), .A4(n12009), .ZN(
        n12010) );
  NAND4_X1 U14504 ( .A1(n14099), .A2(n12011), .A3(n12010), .A4(n14144), .ZN(
        n12012) );
  NOR3_X1 U14505 ( .A1(n14060), .A2(n12013), .A3(n12012), .ZN(n12015) );
  NAND4_X1 U14506 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n14043), .ZN(
        n12017) );
  NOR4_X1 U14507 ( .A1(n12021), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(
        n12020) );
  XNOR2_X1 U14508 ( .A(n12020), .B(n14106), .ZN(n12027) );
  NAND2_X1 U14509 ( .A1(n12021), .A2(n7451), .ZN(n12023) );
  MUX2_X1 U14510 ( .A(n12024), .B(n12023), .S(n11983), .Z(n12025) );
  OAI21_X1 U14511 ( .B1(n12027), .B2(n12026), .A(n12025), .ZN(n12028) );
  NOR3_X1 U14512 ( .A1(n12031), .A2(n14362), .A3(n14520), .ZN(n12033) );
  OAI21_X1 U14513 ( .B1(n12034), .B2(n6858), .A(P1_B_REG_SCAN_IN), .ZN(n12032)
         );
  OAI22_X1 U14514 ( .A1(n12035), .A2(n12034), .B1(n12033), .B2(n12032), .ZN(
        P1_U3242) );
  INV_X1 U14515 ( .A(n12036), .ZN(n13686) );
  INV_X1 U14516 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U14517 ( .A1(n6559), .A2(n13126), .B1(n13097), .B2(n13280), .ZN(
        n12045) );
  AND2_X1 U14518 ( .A1(n13278), .A2(n13523), .ZN(n12040) );
  AOI21_X1 U14519 ( .B1(n13347), .B2(n13521), .A(n12040), .ZN(n13583) );
  INV_X1 U14520 ( .A(n12041), .ZN(n13379) );
  AOI22_X1 U14521 ( .A1(n13379), .A2(n13098), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12042) );
  OAI21_X1 U14522 ( .B1(n13583), .B2(n13101), .A(n12042), .ZN(n12043) );
  AOI21_X1 U14523 ( .B1(n13383), .B2(n14467), .A(n12043), .ZN(n12044) );
  OAI21_X1 U14524 ( .B1(n12039), .B2(n12045), .A(n12044), .ZN(P2_U3188) );
  AOI22_X1 U14525 ( .A1(n13122), .A2(n12046), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12047) );
  OAI21_X1 U14526 ( .B1(n12048), .B2(n14470), .A(n12047), .ZN(n12055) );
  NOR3_X1 U14527 ( .A1(n12050), .A2(n12049), .A3(n13132), .ZN(n12051) );
  AOI21_X1 U14528 ( .B1(n11418), .B2(n13126), .A(n12051), .ZN(n12053) );
  NOR2_X1 U14529 ( .A1(n12053), .A2(n12052), .ZN(n12054) );
  AOI211_X1 U14530 ( .C1(n13636), .C2(n14467), .A(n12055), .B(n12054), .ZN(
        n12056) );
  OAI21_X1 U14531 ( .B1(n14462), .B2(n12057), .A(n12056), .ZN(P2_U3187) );
  AOI22_X1 U14532 ( .A1(n13122), .A2(n12058), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12059) );
  OAI21_X1 U14533 ( .B1(n12060), .B2(n14470), .A(n12059), .ZN(n12069) );
  INV_X1 U14534 ( .A(n12061), .ZN(n12065) );
  NOR3_X1 U14535 ( .A1(n12063), .A2(n12062), .A3(n13132), .ZN(n12064) );
  AOI21_X1 U14536 ( .B1(n12065), .B2(n13126), .A(n12064), .ZN(n12067) );
  NOR2_X1 U14537 ( .A1(n12067), .A2(n12066), .ZN(n12068) );
  AOI211_X1 U14538 ( .C1(n12070), .C2(n14467), .A(n12069), .B(n12068), .ZN(
        n12071) );
  OAI21_X1 U14539 ( .B1(n14462), .B2(n12072), .A(n12071), .ZN(P2_U3193) );
  INV_X1 U14540 ( .A(n12073), .ZN(n12075) );
  OAI222_X1 U14541 ( .A1(P3_U3151), .A2(n9922), .B1(n12387), .B2(n12075), .C1(
        n12074), .C2(n13004), .ZN(P3_U3268) );
  INV_X1 U14542 ( .A(n12076), .ZN(n12284) );
  INV_X1 U14543 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U14544 ( .A1(n13675), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U14545 ( .A1(n12077), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12078) );
  NAND2_X1 U14546 ( .A1(n12093), .A2(n12078), .ZN(n12091) );
  INV_X1 U14547 ( .A(n12079), .ZN(n12080) );
  INV_X1 U14548 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13679) );
  INV_X1 U14549 ( .A(SI_30_), .ZN(n12306) );
  INV_X1 U14550 ( .A(n12915), .ZN(n12850) );
  NAND2_X1 U14551 ( .A1(n12083), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12089) );
  INV_X1 U14552 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12084) );
  OR2_X1 U14553 ( .A1(n12085), .A2(n12084), .ZN(n12088) );
  INV_X1 U14554 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12636) );
  OR2_X1 U14555 ( .A1(n12086), .A2(n12636), .ZN(n12087) );
  NAND4_X1 U14556 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n12087), .ZN(
        n12633) );
  NAND2_X1 U14557 ( .A1(n12094), .A2(n12093), .ZN(n12096) );
  XNOR2_X1 U14558 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12095) );
  INV_X1 U14559 ( .A(SI_31_), .ZN(n13005) );
  NOR2_X1 U14560 ( .A1(n9714), .A2(n13005), .ZN(n12097) );
  INV_X1 U14561 ( .A(n12099), .ZN(n12285) );
  OAI211_X1 U14562 ( .C1(n12850), .C2(n12633), .A(n12107), .B(n12285), .ZN(
        n12100) );
  AOI21_X1 U14563 ( .B1(n12101), .B2(n12284), .A(n12100), .ZN(n12104) );
  OAI22_X1 U14564 ( .A1(n12915), .A2(n12102), .B1(n12914), .B2(n12633), .ZN(
        n12287) );
  INV_X1 U14565 ( .A(n12914), .ZN(n12630) );
  NOR2_X1 U14566 ( .A1(n12104), .A2(n12103), .ZN(n12106) );
  INV_X1 U14567 ( .A(n12107), .ZN(n12130) );
  NAND2_X1 U14568 ( .A1(n12110), .A2(n12680), .ZN(n12697) );
  INV_X1 U14569 ( .A(n12697), .ZN(n12695) );
  OR4_X1 U14570 ( .A1(n10775), .A2(n12112), .A3(n12180), .A4(n12111), .ZN(
        n12116) );
  NOR4_X1 U14571 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12120) );
  NOR4_X1 U14572 ( .A1(n12143), .A2(n12192), .A3(n12117), .A4(n12172), .ZN(
        n12118) );
  NAND4_X1 U14573 ( .A1(n12120), .A2(n12119), .A3(n9766), .A4(n12118), .ZN(
        n12121) );
  NOR4_X1 U14574 ( .A1(n12122), .A2(n12788), .A3(n12121), .A4(n12778), .ZN(
        n12123) );
  NAND2_X1 U14575 ( .A1(n12123), .A2(n12768), .ZN(n12124) );
  NOR4_X1 U14576 ( .A1(n12124), .A2(n12231), .A3(n12747), .A4(n12732), .ZN(
        n12125) );
  NAND4_X1 U14577 ( .A1(n12707), .A2(n12695), .A3(n12125), .A4(n12720), .ZN(
        n12126) );
  NOR4_X1 U14578 ( .A1(n12260), .A2(n12663), .A3(n12256), .A4(n12126), .ZN(
        n12127) );
  NAND4_X1 U14579 ( .A1(n12640), .A2(n12651), .A3(n12127), .A4(n12261), .ZN(
        n12128) );
  XNOR2_X1 U14580 ( .A(n12131), .B(n12614), .ZN(n12133) );
  INV_X1 U14581 ( .A(n12680), .ZN(n12135) );
  MUX2_X1 U14582 ( .A(n12660), .B(n12135), .S(n12276), .Z(n12255) );
  INV_X1 U14583 ( .A(n9754), .ZN(n12142) );
  NAND2_X1 U14584 ( .A1(n12138), .A2(n12139), .ZN(n12145) );
  INV_X1 U14585 ( .A(n12140), .ZN(n12141) );
  MUX2_X1 U14586 ( .A(n12142), .B(n12141), .S(n12276), .Z(n12144) );
  AOI211_X1 U14587 ( .C1(n12146), .C2(n12145), .A(n12144), .B(n12143), .ZN(
        n12156) );
  NAND2_X1 U14588 ( .A1(n12151), .A2(n12147), .ZN(n12150) );
  NAND2_X1 U14589 ( .A1(n12152), .A2(n12148), .ZN(n12149) );
  MUX2_X1 U14590 ( .A(n12150), .B(n12149), .S(n12276), .Z(n12155) );
  MUX2_X1 U14591 ( .A(n12152), .B(n12151), .S(n12276), .Z(n12153) );
  OAI211_X1 U14592 ( .C1(n12156), .C2(n12155), .A(n12154), .B(n12153), .ZN(
        n12161) );
  MUX2_X1 U14593 ( .A(n12158), .B(n12157), .S(n12276), .Z(n12159) );
  NAND3_X1 U14594 ( .A1(n12161), .A2(n12160), .A3(n12159), .ZN(n12175) );
  INV_X1 U14595 ( .A(n12162), .ZN(n12164) );
  INV_X1 U14596 ( .A(n12163), .ZN(n12170) );
  NOR2_X1 U14597 ( .A1(n12164), .A2(n12170), .ZN(n12169) );
  INV_X1 U14598 ( .A(n12166), .ZN(n12167) );
  NOR2_X1 U14599 ( .A1(n12171), .A2(n12167), .ZN(n12168) );
  MUX2_X1 U14600 ( .A(n12169), .B(n12168), .S(n12276), .Z(n12174) );
  MUX2_X1 U14601 ( .A(n12171), .B(n12170), .S(n12276), .Z(n12173) );
  AOI211_X1 U14602 ( .C1(n12175), .C2(n12174), .A(n12173), .B(n12172), .ZN(
        n12182) );
  INV_X1 U14603 ( .A(n12176), .ZN(n12179) );
  INV_X1 U14604 ( .A(n12177), .ZN(n12178) );
  MUX2_X1 U14605 ( .A(n12179), .B(n12178), .S(n12276), .Z(n12181) );
  NOR3_X1 U14606 ( .A1(n12182), .A2(n12181), .A3(n12180), .ZN(n12189) );
  INV_X1 U14607 ( .A(n12183), .ZN(n12186) );
  INV_X1 U14608 ( .A(n12184), .ZN(n12185) );
  MUX2_X1 U14609 ( .A(n12186), .B(n12185), .S(n12276), .Z(n12188) );
  MUX2_X1 U14610 ( .A(n12191), .B(n12190), .S(n12276), .Z(n12193) );
  NOR2_X1 U14611 ( .A1(n12193), .A2(n12192), .ZN(n12198) );
  INV_X1 U14612 ( .A(n12194), .ZN(n12196) );
  MUX2_X1 U14613 ( .A(n12196), .B(n9764), .S(n12276), .Z(n12197) );
  NOR4_X1 U14614 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12833), .ZN(
        n12208) );
  NAND2_X1 U14615 ( .A1(n12204), .A2(n12200), .ZN(n12203) );
  NAND2_X1 U14616 ( .A1(n12205), .A2(n12201), .ZN(n12202) );
  MUX2_X1 U14617 ( .A(n12203), .B(n12202), .S(n12276), .Z(n12207) );
  MUX2_X1 U14618 ( .A(n12205), .B(n12204), .S(n12276), .Z(n12206) );
  OAI211_X1 U14619 ( .C1(n12208), .C2(n12207), .A(n12815), .B(n12206), .ZN(
        n12212) );
  MUX2_X1 U14620 ( .A(n12210), .B(n12209), .S(n12276), .Z(n12211) );
  NAND3_X1 U14621 ( .A1(n12212), .A2(n9769), .A3(n12211), .ZN(n12216) );
  MUX2_X1 U14622 ( .A(n12214), .B(n12213), .S(n12276), .Z(n12215) );
  AOI21_X1 U14623 ( .B1(n12216), .B2(n12215), .A(n12778), .ZN(n12219) );
  AOI21_X1 U14624 ( .B1(n12224), .B2(n12217), .A(n12286), .ZN(n12218) );
  OAI21_X1 U14625 ( .B1(n12219), .B2(n12218), .A(n12220), .ZN(n12227) );
  INV_X1 U14626 ( .A(n12220), .ZN(n12223) );
  INV_X1 U14627 ( .A(n12221), .ZN(n12222) );
  OAI21_X1 U14628 ( .B1(n12223), .B2(n12222), .A(n12286), .ZN(n12226) );
  INV_X1 U14629 ( .A(n12224), .ZN(n12225) );
  AOI22_X1 U14630 ( .A1(n12227), .A2(n12226), .B1(n12286), .B2(n12225), .ZN(
        n12232) );
  AOI211_X1 U14631 ( .C1(n12229), .C2(n12237), .A(n12276), .B(n12228), .ZN(
        n12233) );
  OAI22_X1 U14632 ( .A1(n12232), .A2(n12231), .B1(n12233), .B2(n12230), .ZN(
        n12235) );
  INV_X1 U14633 ( .A(n12233), .ZN(n12238) );
  NAND3_X1 U14634 ( .A1(n12236), .A2(n12276), .A3(n12237), .ZN(n12234) );
  AOI22_X1 U14635 ( .A1(n12235), .A2(n12729), .B1(n12238), .B2(n12234), .ZN(
        n12243) );
  OAI21_X1 U14636 ( .B1(n12238), .B2(n12237), .A(n12236), .ZN(n12241) );
  INV_X1 U14637 ( .A(n12239), .ZN(n12240) );
  MUX2_X1 U14638 ( .A(n12241), .B(n12240), .S(n12276), .Z(n12242) );
  NOR2_X1 U14639 ( .A1(n12243), .A2(n12242), .ZN(n12249) );
  INV_X1 U14640 ( .A(n12950), .ZN(n12244) );
  NOR2_X1 U14641 ( .A1(n12244), .A2(n12589), .ZN(n12245) );
  MUX2_X1 U14642 ( .A(n12246), .B(n12245), .S(n12276), .Z(n12247) );
  NOR2_X1 U14643 ( .A1(n12507), .A2(n12286), .ZN(n12251) );
  NOR2_X1 U14644 ( .A1(n12588), .A2(n12276), .ZN(n12250) );
  MUX2_X1 U14645 ( .A(n12251), .B(n12250), .S(n12877), .Z(n12252) );
  NOR3_X1 U14646 ( .A1(n12253), .A2(n12252), .A3(n12697), .ZN(n12254) );
  XOR2_X1 U14647 ( .A(n12276), .B(n12257), .Z(n12258) );
  NOR2_X1 U14648 ( .A1(n12259), .A2(n12258), .ZN(n12262) );
  AOI21_X1 U14649 ( .B1(n12262), .B2(n12261), .A(n12260), .ZN(n12263) );
  AOI22_X1 U14650 ( .A1(n12264), .A2(n12263), .B1(n12286), .B2(n12266), .ZN(
        n12272) );
  NOR2_X1 U14651 ( .A1(n12265), .A2(n12286), .ZN(n12268) );
  NOR3_X1 U14652 ( .A1(n12266), .A2(n12585), .A3(n12276), .ZN(n12267) );
  MUX2_X1 U14653 ( .A(n12268), .B(n12267), .S(n12858), .Z(n12271) );
  NAND3_X1 U14654 ( .A1(n12559), .A2(n12269), .A3(n12276), .ZN(n12270) );
  OAI211_X1 U14655 ( .C1(n12272), .C2(n12271), .A(n12651), .B(n12270), .ZN(
        n12275) );
  NAND3_X1 U14656 ( .A1(n12273), .A2(n12276), .A3(n12583), .ZN(n12274) );
  AOI21_X1 U14657 ( .B1(n12275), .B2(n12274), .A(n12425), .ZN(n12283) );
  AOI21_X1 U14658 ( .B1(n12278), .B2(n12277), .A(n12276), .ZN(n12280) );
  MUX2_X1 U14659 ( .A(n12280), .B(n12276), .S(n12279), .Z(n12282) );
  NAND4_X1 U14660 ( .A1(n12572), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12295) );
  OAI211_X1 U14661 ( .C1(n12297), .C2(n12296), .A(n12295), .B(P3_B_REG_SCAN_IN), .ZN(n12298) );
  AOI22_X1 U14662 ( .A1(n14147), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n12377), 
        .B2(n14243), .ZN(n12300) );
  OAI21_X1 U14663 ( .B1(n12301), .B2(n14196), .A(n12300), .ZN(n12302) );
  AOI21_X1 U14664 ( .B1(n12303), .B2(n14244), .A(n12302), .ZN(n12304) );
  OAI21_X1 U14665 ( .B1(n12305), .B2(n14147), .A(n12304), .ZN(P1_U3265) );
  OAI222_X1 U14666 ( .A1(n8839), .A2(P3_U3151), .B1(n12387), .B2(n12307), .C1(
        n12306), .C2(n13004), .ZN(P3_U3265) );
  INV_X1 U14667 ( .A(n12308), .ZN(n12314) );
  AOI22_X1 U14668 ( .A1(n12311), .A2(n12310), .B1(n12309), .B2(n14243), .ZN(
        n12313) );
  NAND2_X1 U14669 ( .A1(n14147), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12312) );
  OAI211_X1 U14670 ( .C1(n12314), .C2(n14196), .A(n12313), .B(n12312), .ZN(
        n12316) );
  OAI21_X1 U14671 ( .B1(n12318), .B2(n14147), .A(n6608), .ZN(P1_U3356) );
  INV_X1 U14672 ( .A(n12319), .ZN(n12320) );
  NAND2_X1 U14673 ( .A1(n14289), .A2(n12360), .ZN(n12324) );
  NAND2_X1 U14674 ( .A1(n14079), .A2(n11633), .ZN(n12323) );
  NAND2_X1 U14675 ( .A1(n12324), .A2(n12323), .ZN(n12325) );
  XNOR2_X1 U14676 ( .A(n12325), .B(n12343), .ZN(n12327) );
  AND2_X1 U14677 ( .A1(n12364), .A2(n14079), .ZN(n12326) );
  AOI21_X1 U14678 ( .B1(n14289), .B2(n11633), .A(n12326), .ZN(n12328) );
  NAND2_X1 U14679 ( .A1(n12327), .A2(n12328), .ZN(n13792) );
  INV_X1 U14680 ( .A(n12327), .ZN(n12330) );
  INV_X1 U14681 ( .A(n12328), .ZN(n12329) );
  NAND2_X1 U14682 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  NAND2_X1 U14683 ( .A1(n14087), .A2(n12360), .ZN(n12333) );
  NAND2_X1 U14684 ( .A1(n14112), .A2(n11633), .ZN(n12332) );
  NAND2_X1 U14685 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  XNOR2_X1 U14686 ( .A(n12334), .B(n12343), .ZN(n12336) );
  AND2_X1 U14687 ( .A1(n12364), .A2(n14112), .ZN(n12335) );
  AOI21_X1 U14688 ( .B1(n14087), .B2(n11633), .A(n12335), .ZN(n12337) );
  NAND2_X1 U14689 ( .A1(n12336), .A2(n12337), .ZN(n13761) );
  INV_X1 U14690 ( .A(n12336), .ZN(n12339) );
  INV_X1 U14691 ( .A(n12337), .ZN(n12338) );
  NAND2_X1 U14692 ( .A1(n12339), .A2(n12338), .ZN(n12340) );
  NAND2_X1 U14693 ( .A1(n14058), .A2(n12360), .ZN(n12342) );
  NAND2_X1 U14694 ( .A1(n14078), .A2(n11584), .ZN(n12341) );
  NAND2_X1 U14695 ( .A1(n12342), .A2(n12341), .ZN(n12344) );
  XNOR2_X1 U14696 ( .A(n12344), .B(n12343), .ZN(n12346) );
  AND2_X1 U14697 ( .A1(n12364), .A2(n14078), .ZN(n12345) );
  AOI21_X1 U14698 ( .B1(n14058), .B2(n11584), .A(n12345), .ZN(n12347) );
  NAND2_X1 U14699 ( .A1(n12346), .A2(n12347), .ZN(n12351) );
  INV_X1 U14700 ( .A(n12346), .ZN(n12349) );
  INV_X1 U14701 ( .A(n12347), .ZN(n12348) );
  NAND2_X1 U14702 ( .A1(n12349), .A2(n12348), .ZN(n12350) );
  NAND2_X1 U14703 ( .A1(n14046), .A2(n12360), .ZN(n12353) );
  NAND2_X1 U14704 ( .A1(n13871), .A2(n11633), .ZN(n12352) );
  NAND2_X1 U14705 ( .A1(n12353), .A2(n12352), .ZN(n12354) );
  XNOR2_X1 U14706 ( .A(n12354), .B(n12370), .ZN(n12358) );
  NAND2_X1 U14707 ( .A1(n14046), .A2(n11584), .ZN(n12356) );
  NAND2_X1 U14708 ( .A1(n12364), .A2(n13871), .ZN(n12355) );
  NAND2_X1 U14709 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  NOR2_X1 U14710 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  AOI21_X1 U14711 ( .B1(n12358), .B2(n12357), .A(n12359), .ZN(n13843) );
  NAND2_X1 U14712 ( .A1(n14033), .A2(n12360), .ZN(n12362) );
  NAND2_X1 U14713 ( .A1(n13870), .A2(n11584), .ZN(n12361) );
  NAND2_X1 U14714 ( .A1(n12362), .A2(n12361), .ZN(n12363) );
  XNOR2_X1 U14715 ( .A(n12363), .B(n12370), .ZN(n12368) );
  NAND2_X1 U14716 ( .A1(n14033), .A2(n11584), .ZN(n12366) );
  NAND2_X1 U14717 ( .A1(n12364), .A2(n13870), .ZN(n12365) );
  NAND2_X1 U14718 ( .A1(n12366), .A2(n12365), .ZN(n12367) );
  NOR2_X1 U14719 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  AOI21_X1 U14720 ( .B1(n12368), .B2(n12367), .A(n12369), .ZN(n13693) );
  AOI22_X1 U14721 ( .A1(n12382), .A2(n12360), .B1(n11584), .B2(n13869), .ZN(
        n12371) );
  XNOR2_X1 U14722 ( .A(n12371), .B(n12370), .ZN(n12374) );
  AOI22_X1 U14723 ( .A1(n12382), .A2(n11584), .B1(n12372), .B2(n13869), .ZN(
        n12373) );
  XNOR2_X1 U14724 ( .A(n12374), .B(n12373), .ZN(n12375) );
  XNOR2_X1 U14725 ( .A(n12376), .B(n12375), .ZN(n12384) );
  INV_X1 U14726 ( .A(n12377), .ZN(n12380) );
  AOI22_X1 U14727 ( .A1(n13825), .A2(n13868), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12379) );
  NAND2_X1 U14728 ( .A1(n13855), .A2(n13870), .ZN(n12378) );
  OAI211_X1 U14729 ( .C1(n13786), .C2(n12380), .A(n12379), .B(n12378), .ZN(
        n12381) );
  AOI21_X1 U14730 ( .B1(n12382), .B2(n13817), .A(n12381), .ZN(n12383) );
  OAI21_X1 U14731 ( .B1(n12384), .B2(n13864), .A(n12383), .ZN(P1_U3220) );
  INV_X1 U14732 ( .A(n12385), .ZN(n12386) );
  OAI222_X1 U14733 ( .A1(n13004), .A2(n12388), .B1(n12387), .B2(n12386), .C1(
        P3_U3151), .C2(n8840), .ZN(P3_U3266) );
  OR2_X1 U14734 ( .A1(n12477), .A2(n12550), .ZN(n12391) );
  NAND2_X1 U14735 ( .A1(n12596), .A2(n12572), .ZN(n12390) );
  NAND2_X1 U14736 ( .A1(n12391), .A2(n12390), .ZN(n12791) );
  AOI22_X1 U14737 ( .A1(n12791), .A2(n14982), .B1(P3_REG3_REG_14__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12392) );
  OAI21_X1 U14738 ( .B1(n12795), .B2(n14985), .A(n12392), .ZN(n12398) );
  INV_X1 U14739 ( .A(n12393), .ZN(n12394) );
  AOI211_X1 U14740 ( .C1(n12396), .C2(n12395), .A(n12579), .B(n12394), .ZN(
        n12397) );
  AOI211_X1 U14741 ( .C1(n9693), .C2(n12577), .A(n12398), .B(n12397), .ZN(
        n12399) );
  INV_X1 U14742 ( .A(n12399), .ZN(P3_U3155) );
  NOR2_X1 U14743 ( .A1(n7440), .A2(n12400), .ZN(n12493) );
  NAND2_X1 U14744 ( .A1(n12401), .A2(n12526), .ZN(n12496) );
  OAI21_X1 U14745 ( .B1(n12526), .B2(n12401), .A(n12496), .ZN(n12402) );
  NAND2_X1 U14746 ( .A1(n12402), .A2(n14974), .ZN(n12407) );
  INV_X1 U14747 ( .A(n12688), .ZN(n12405) );
  INV_X1 U14748 ( .A(n12403), .ZN(n12586) );
  AOI22_X1 U14749 ( .A1(n12572), .A2(n9700), .B1(n12586), .B2(n12573), .ZN(
        n12686) );
  OAI22_X1 U14750 ( .A1(n12686), .A2(n12530), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9538), .ZN(n12404) );
  AOI21_X1 U14751 ( .B1(n12405), .B2(n12532), .A(n12404), .ZN(n12406) );
  OAI211_X1 U14752 ( .C1(n12939), .C2(n14973), .A(n12407), .B(n12406), .ZN(
        P3_U3156) );
  AOI21_X1 U14753 ( .B1(n12409), .B2(n12408), .A(n12579), .ZN(n12411) );
  NAND2_X1 U14754 ( .A1(n12411), .A2(n12410), .ZN(n12416) );
  AOI22_X1 U14755 ( .A1(n12413), .A2(n14982), .B1(n12412), .B2(n12577), .ZN(
        n12415) );
  MUX2_X1 U14756 ( .A(n14985), .B(P3_STATE_REG_SCAN_IN), .S(
        P3_REG3_REG_3__SCAN_IN), .Z(n12414) );
  NAND3_X1 U14757 ( .A1(n12416), .A2(n12415), .A3(n12414), .ZN(P3_U3158) );
  XNOR2_X1 U14758 ( .A(n12418), .B(n12417), .ZN(n12424) );
  OR2_X1 U14759 ( .A1(n12487), .A2(n12548), .ZN(n12420) );
  OR2_X1 U14760 ( .A1(n12443), .A2(n12550), .ZN(n12419) );
  NAND2_X1 U14761 ( .A1(n12420), .A2(n12419), .ZN(n12736) );
  AOI22_X1 U14762 ( .A1(n12736), .A2(n14982), .B1(P3_REG3_REG_19__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12421) );
  OAI21_X1 U14763 ( .B1(n12739), .B2(n14985), .A(n12421), .ZN(n12422) );
  AOI21_X1 U14764 ( .B1(n12956), .B2(n12577), .A(n12422), .ZN(n12423) );
  OAI21_X1 U14765 ( .B1(n12424), .B2(n12579), .A(n12423), .ZN(P3_U3159) );
  INV_X1 U14766 ( .A(n12434), .ZN(n12426) );
  XNOR2_X1 U14767 ( .A(n12425), .B(n6467), .ZN(n12436) );
  NAND3_X1 U14768 ( .A1(n12426), .A2(n12436), .A3(n14974), .ZN(n12440) );
  OR2_X1 U14769 ( .A1(n12427), .A2(n12548), .ZN(n12429) );
  NAND2_X1 U14770 ( .A1(n12581), .A2(n12573), .ZN(n12428) );
  NAND2_X1 U14771 ( .A1(n12429), .A2(n12428), .ZN(n12642) );
  AOI22_X1 U14772 ( .A1(n12642), .A2(n14982), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12430) );
  OAI21_X1 U14773 ( .B1(n12645), .B2(n14985), .A(n12430), .ZN(n12431) );
  AOI21_X1 U14774 ( .B1(n12921), .B2(n12577), .A(n12431), .ZN(n12439) );
  INV_X1 U14775 ( .A(n12435), .ZN(n12433) );
  INV_X1 U14776 ( .A(n12436), .ZN(n12432) );
  NAND4_X1 U14777 ( .A1(n12434), .A2(n12433), .A3(n14974), .A4(n12432), .ZN(
        n12438) );
  NAND3_X1 U14778 ( .A1(n12436), .A2(n12435), .A3(n14974), .ZN(n12437) );
  NAND4_X1 U14779 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        P3_U3160) );
  AOI21_X1 U14780 ( .B1(n12442), .B2(n12441), .A(n6576), .ZN(n12449) );
  OR2_X1 U14781 ( .A1(n12524), .A2(n12550), .ZN(n12445) );
  OR2_X1 U14782 ( .A1(n12443), .A2(n12548), .ZN(n12444) );
  NAND2_X1 U14783 ( .A1(n12445), .A2(n12444), .ZN(n12709) );
  AOI22_X1 U14784 ( .A1(n12709), .A2(n14982), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12446) );
  OAI21_X1 U14785 ( .B1(n7454), .B2(n14985), .A(n12446), .ZN(n12447) );
  AOI21_X1 U14786 ( .B1(n12877), .B2(n12577), .A(n12447), .ZN(n12448) );
  OAI21_X1 U14787 ( .B1(n12449), .B2(n12579), .A(n12448), .ZN(P3_U3163) );
  INV_X1 U14788 ( .A(n12450), .ZN(n12451) );
  XOR2_X1 U14789 ( .A(n12450), .B(n12452), .Z(n12538) );
  NOR2_X1 U14790 ( .A1(n12538), .A2(n12539), .ZN(n12537) );
  AOI21_X1 U14791 ( .B1(n12452), .B2(n12451), .A(n12537), .ZN(n12456) );
  NAND2_X1 U14792 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  XNOR2_X1 U14793 ( .A(n12456), .B(n12455), .ZN(n12461) );
  OAI22_X1 U14794 ( .A1(n12539), .A2(n12548), .B1(n12457), .B2(n12550), .ZN(
        n12821) );
  NAND2_X1 U14795 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n15053)
         );
  OAI21_X1 U14796 ( .B1(n14973), .B2(n12993), .A(n15053), .ZN(n12459) );
  NOR2_X1 U14797 ( .A1(n14985), .A2(n12827), .ZN(n12458) );
  AOI211_X1 U14798 ( .C1(n12821), .C2(n14982), .A(n12459), .B(n12458), .ZN(
        n12460) );
  OAI21_X1 U14799 ( .B1(n12461), .B2(n12579), .A(n12460), .ZN(P3_U3164) );
  INV_X1 U14800 ( .A(n12462), .ZN(n12467) );
  NOR3_X1 U14801 ( .A1(n12463), .A2(n12465), .A3(n12464), .ZN(n12466) );
  OAI21_X1 U14802 ( .B1(n12467), .B2(n12466), .A(n14974), .ZN(n12473) );
  AOI22_X1 U14803 ( .A1(n12468), .A2(n14982), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12469) );
  OAI21_X1 U14804 ( .B1(n12470), .B2(n14985), .A(n12469), .ZN(n12471) );
  AOI21_X1 U14805 ( .B1(n12858), .B2(n12577), .A(n12471), .ZN(n12472) );
  NAND2_X1 U14806 ( .A1(n12473), .A2(n12472), .ZN(P3_U3165) );
  XNOR2_X1 U14807 ( .A(n12474), .B(n12486), .ZN(n12475) );
  XNOR2_X1 U14808 ( .A(n12476), .B(n12475), .ZN(n12483) );
  OR2_X1 U14809 ( .A1(n12477), .A2(n12548), .ZN(n12479) );
  OR2_X1 U14810 ( .A1(n12549), .A2(n12550), .ZN(n12478) );
  NAND2_X1 U14811 ( .A1(n12479), .A2(n12478), .ZN(n12769) );
  AOI22_X1 U14812 ( .A1(n12769), .A2(n14982), .B1(P3_REG3_REG_16__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12480) );
  OAI21_X1 U14813 ( .B1(n12772), .B2(n14985), .A(n12480), .ZN(n12481) );
  AOI21_X1 U14814 ( .B1(n12974), .B2(n12577), .A(n12481), .ZN(n12482) );
  OAI21_X1 U14815 ( .B1(n12483), .B2(n12579), .A(n12482), .ZN(P3_U3166) );
  XNOR2_X1 U14816 ( .A(n12485), .B(n12484), .ZN(n12492) );
  OAI22_X1 U14817 ( .A1(n12487), .A2(n12550), .B1(n12486), .B2(n12548), .ZN(
        n12760) );
  AOI22_X1 U14818 ( .A1(n12760), .A2(n14982), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12488) );
  OAI21_X1 U14819 ( .B1(n12489), .B2(n14985), .A(n12488), .ZN(n12490) );
  AOI21_X1 U14820 ( .B1(n12968), .B2(n12577), .A(n12490), .ZN(n12491) );
  OAI21_X1 U14821 ( .B1(n12492), .B2(n12579), .A(n12491), .ZN(P3_U3168) );
  INV_X1 U14822 ( .A(n12493), .ZN(n12494) );
  AND3_X1 U14823 ( .A1(n12496), .A2(n12495), .A3(n12494), .ZN(n12497) );
  OAI21_X1 U14824 ( .B1(n12497), .B2(n12463), .A(n14974), .ZN(n12504) );
  INV_X1 U14825 ( .A(n12673), .ZN(n12502) );
  OR2_X1 U14826 ( .A1(n12526), .A2(n12548), .ZN(n12499) );
  NAND2_X1 U14827 ( .A1(n12585), .A2(n12573), .ZN(n12498) );
  AND2_X1 U14828 ( .A1(n12499), .A2(n12498), .ZN(n12671) );
  OAI22_X1 U14829 ( .A1(n12671), .A2(n12530), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12500), .ZN(n12501) );
  AOI21_X1 U14830 ( .B1(n12502), .B2(n12532), .A(n12501), .ZN(n12503) );
  OAI211_X1 U14831 ( .C1(n12935), .C2(n14973), .A(n12504), .B(n12503), .ZN(
        P3_U3169) );
  XNOR2_X1 U14832 ( .A(n12506), .B(n12505), .ZN(n12511) );
  OAI22_X1 U14833 ( .A1(n12507), .A2(n12550), .B1(n12551), .B2(n12548), .ZN(
        n12722) );
  AOI22_X1 U14834 ( .A1(n12722), .A2(n14982), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12508) );
  OAI21_X1 U14835 ( .B1(n12725), .B2(n14985), .A(n12508), .ZN(n12509) );
  AOI21_X1 U14836 ( .B1(n12950), .B2(n12577), .A(n12509), .ZN(n12510) );
  OAI21_X1 U14837 ( .B1(n12511), .B2(n12579), .A(n12510), .ZN(P3_U3173) );
  XNOR2_X1 U14838 ( .A(n12512), .B(n12596), .ZN(n12513) );
  XNOR2_X1 U14839 ( .A(n12514), .B(n12513), .ZN(n12515) );
  NAND2_X1 U14840 ( .A1(n12515), .A2(n14974), .ZN(n12521) );
  NAND2_X1 U14841 ( .A1(n12595), .A2(n12573), .ZN(n12517) );
  NAND2_X1 U14842 ( .A1(n12597), .A2(n12572), .ZN(n12516) );
  NAND2_X1 U14843 ( .A1(n12517), .A2(n12516), .ZN(n12808) );
  AOI22_X1 U14844 ( .A1(n12808), .A2(n14982), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12520) );
  OR2_X1 U14845 ( .A1(n14973), .A2(n14450), .ZN(n12519) );
  OR2_X1 U14846 ( .A1(n14985), .A2(n12811), .ZN(n12518) );
  NAND4_X1 U14847 ( .A1(n12521), .A2(n12520), .A3(n12519), .A4(n12518), .ZN(
        P3_U3174) );
  OAI21_X1 U14848 ( .B1(n12524), .B2(n12523), .A(n12522), .ZN(n12525) );
  NAND2_X1 U14849 ( .A1(n12525), .A2(n14974), .ZN(n12535) );
  INV_X1 U14850 ( .A(n12701), .ZN(n12533) );
  OR2_X1 U14851 ( .A1(n12526), .A2(n12550), .ZN(n12528) );
  NAND2_X1 U14852 ( .A1(n12588), .A2(n12572), .ZN(n12527) );
  AND2_X1 U14853 ( .A1(n12528), .A2(n12527), .ZN(n12699) );
  OAI22_X1 U14854 ( .A1(n12699), .A2(n12530), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12529), .ZN(n12531) );
  AOI21_X1 U14855 ( .B1(n12533), .B2(n12532), .A(n12531), .ZN(n12534) );
  OAI211_X1 U14856 ( .C1(n12536), .C2(n14973), .A(n12535), .B(n12534), .ZN(
        P3_U3175) );
  AOI211_X1 U14857 ( .C1(n12539), .C2(n12538), .A(n12579), .B(n12537), .ZN(
        n12540) );
  INV_X1 U14858 ( .A(n12540), .ZN(n12545) );
  NAND2_X1 U14859 ( .A1(n12597), .A2(n12573), .ZN(n12542) );
  NAND2_X1 U14860 ( .A1(n12599), .A2(n12572), .ZN(n12541) );
  NAND2_X1 U14861 ( .A1(n12542), .A2(n12541), .ZN(n12834) );
  NAND2_X1 U14862 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n15035)
         );
  OAI21_X1 U14863 ( .B1(n14973), .B2(n12997), .A(n15035), .ZN(n12543) );
  AOI21_X1 U14864 ( .B1(n12834), .B2(n14982), .A(n12543), .ZN(n12544) );
  OAI211_X1 U14865 ( .C1(n14985), .C2(n12840), .A(n12545), .B(n12544), .ZN(
        P3_U3176) );
  XNOR2_X1 U14866 ( .A(n12547), .B(n12546), .ZN(n12555) );
  OAI22_X1 U14867 ( .A1(n12551), .A2(n12550), .B1(n12549), .B2(n12548), .ZN(
        n12749) );
  AOI22_X1 U14868 ( .A1(n12749), .A2(n14982), .B1(P3_REG3_REG_18__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12552) );
  OAI21_X1 U14869 ( .B1(n12752), .B2(n14985), .A(n12552), .ZN(n12553) );
  AOI21_X1 U14870 ( .B1(n12962), .B2(n12577), .A(n12553), .ZN(n12554) );
  OAI21_X1 U14871 ( .B1(n12555), .B2(n12579), .A(n12554), .ZN(P3_U3178) );
  OAI21_X1 U14872 ( .B1(n12558), .B2(n12557), .A(n12556), .ZN(n12565) );
  NAND2_X1 U14873 ( .A1(n12559), .A2(n12577), .ZN(n12562) );
  AOI22_X1 U14874 ( .A1(n12560), .A2(n14982), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12561) );
  OAI211_X1 U14875 ( .C1(n12563), .C2(n14985), .A(n12562), .B(n12561), .ZN(
        n12564) );
  AOI21_X1 U14876 ( .B1(n12565), .B2(n14974), .A(n12564), .ZN(n12566) );
  INV_X1 U14877 ( .A(n12566), .ZN(P3_U3180) );
  INV_X1 U14878 ( .A(n12567), .ZN(n12569) );
  NOR2_X1 U14879 ( .A1(n12569), .A2(n12568), .ZN(n12570) );
  XNOR2_X1 U14880 ( .A(n12571), .B(n12570), .ZN(n12580) );
  AOI22_X1 U14881 ( .A1(n12593), .A2(n12573), .B1(n12572), .B2(n12595), .ZN(
        n12780) );
  INV_X1 U14882 ( .A(n12780), .ZN(n12574) );
  AOI22_X1 U14883 ( .A1(n12574), .A2(n14982), .B1(P3_REG3_REG_15__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12575) );
  OAI21_X1 U14884 ( .B1(n12782), .B2(n14985), .A(n12575), .ZN(n12576) );
  AOI21_X1 U14885 ( .B1(n12896), .B2(n12577), .A(n12576), .ZN(n12578) );
  OAI21_X1 U14886 ( .B1(n12580), .B2(n12579), .A(n12578), .ZN(P3_U3181) );
  MUX2_X1 U14887 ( .A(n12633), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12607), .Z(
        P3_U3522) );
  MUX2_X1 U14888 ( .A(n12581), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12607), .Z(
        P3_U3520) );
  MUX2_X1 U14889 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12582), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14890 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12583), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14891 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12584), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14892 ( .A(n12585), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12607), .Z(
        P3_U3516) );
  MUX2_X1 U14893 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12586), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14894 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12587), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14895 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n9700), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14896 ( .A(n12588), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12607), .Z(
        P3_U3512) );
  MUX2_X1 U14897 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12589), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14898 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12590), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14899 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12591), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14900 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12592), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12593), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14902 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12594), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14903 ( .A(n12595), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12607), .Z(
        P3_U3505) );
  MUX2_X1 U14904 ( .A(n12596), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12607), .Z(
        P3_U3504) );
  MUX2_X1 U14905 ( .A(n12597), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12607), .Z(
        P3_U3503) );
  MUX2_X1 U14906 ( .A(n12598), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12607), .Z(
        P3_U3502) );
  MUX2_X1 U14907 ( .A(n12599), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12607), .Z(
        P3_U3501) );
  MUX2_X1 U14908 ( .A(n12600), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12607), .Z(
        P3_U3500) );
  MUX2_X1 U14909 ( .A(n12601), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12607), .Z(
        P3_U3499) );
  MUX2_X1 U14910 ( .A(n12602), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12607), .Z(
        P3_U3498) );
  MUX2_X1 U14911 ( .A(n12603), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12607), .Z(
        P3_U3497) );
  MUX2_X1 U14912 ( .A(n12604), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12607), .Z(
        P3_U3496) );
  MUX2_X1 U14913 ( .A(n12605), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12607), .Z(
        P3_U3495) );
  MUX2_X1 U14914 ( .A(n12606), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12607), .Z(
        P3_U3494) );
  MUX2_X1 U14915 ( .A(n9672), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12607), .Z(
        P3_U3493) );
  MUX2_X1 U14916 ( .A(n8879), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12607), .Z(
        P3_U3492) );
  INV_X1 U14917 ( .A(n12608), .ZN(n12609) );
  MUX2_X1 U14918 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n12609), .S(P3_U3897), .Z(
        P3_U3491) );
  XNOR2_X1 U14919 ( .A(n12614), .B(n12738), .ZN(n12619) );
  AOI22_X1 U14920 ( .A1(n12613), .A2(n12612), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12611), .ZN(n12615) );
  XNOR2_X1 U14921 ( .A(n12614), .B(n12883), .ZN(n12620) );
  XNOR2_X1 U14922 ( .A(n12615), .B(n12620), .ZN(n12628) );
  AOI21_X1 U14923 ( .B1(n12618), .B2(n12617), .A(n12616), .ZN(n12624) );
  INV_X1 U14924 ( .A(n12619), .ZN(n12622) );
  INV_X1 U14925 ( .A(n12620), .ZN(n12621) );
  MUX2_X1 U14926 ( .A(n12622), .B(n12621), .S(n9922), .Z(n12623) );
  NAND2_X1 U14927 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n12626)
         );
  NAND2_X1 U14928 ( .A1(n15089), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12625) );
  OAI211_X1 U14929 ( .C1(n15092), .C2(n12105), .A(n12626), .B(n12625), .ZN(
        n12627) );
  NAND2_X1 U14930 ( .A1(n12630), .A2(n12813), .ZN(n12635) );
  INV_X1 U14931 ( .A(n12631), .ZN(n12632) );
  OAI21_X1 U14932 ( .B1(n12912), .B2(n12634), .A(n15126), .ZN(n12637) );
  OAI211_X1 U14933 ( .C1(n15126), .C2(n12636), .A(n12635), .B(n12637), .ZN(
        P3_U3202) );
  NAND2_X1 U14934 ( .A1(n15128), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12638) );
  OAI211_X1 U14935 ( .C1(n12850), .C2(n12841), .A(n12638), .B(n12637), .ZN(
        P3_U3203) );
  XNOR2_X1 U14936 ( .A(n12639), .B(n12640), .ZN(n12924) );
  AOI21_X1 U14937 ( .B1(n7414), .B2(n12640), .A(n15117), .ZN(n12643) );
  AOI21_X1 U14938 ( .B1(n12643), .B2(n12641), .A(n12642), .ZN(n12919) );
  MUX2_X1 U14939 ( .A(n12644), .B(n12919), .S(n15126), .Z(n12648) );
  INV_X1 U14940 ( .A(n12645), .ZN(n12646) );
  AOI22_X1 U14941 ( .A1(n12921), .A2(n12813), .B1(n12797), .B2(n12646), .ZN(
        n12647) );
  OAI211_X1 U14942 ( .C1(n12802), .C2(n12924), .A(n12648), .B(n12647), .ZN(
        P3_U3205) );
  XNOR2_X1 U14943 ( .A(n12650), .B(n12649), .ZN(n12928) );
  XNOR2_X1 U14944 ( .A(n12652), .B(n12651), .ZN(n12654) );
  OAI21_X1 U14945 ( .B1(n12654), .B2(n15117), .A(n12653), .ZN(n12854) );
  NAND2_X1 U14946 ( .A1(n12854), .A2(n15126), .ZN(n12659) );
  OAI22_X1 U14947 ( .A1(n15126), .A2(n12656), .B1(n12655), .B2(n15121), .ZN(
        n12657) );
  AOI21_X1 U14948 ( .B1(n12855), .B2(n12813), .A(n12657), .ZN(n12658) );
  OAI211_X1 U14949 ( .C1(n12802), .C2(n12928), .A(n12659), .B(n12658), .ZN(
        P3_U3206) );
  OR2_X2 U14950 ( .A1(n12696), .A2(n12660), .ZN(n12681) );
  NAND2_X1 U14951 ( .A1(n12681), .A2(n12661), .ZN(n12682) );
  NAND2_X1 U14952 ( .A1(n12682), .A2(n12662), .ZN(n12664) );
  NAND2_X1 U14953 ( .A1(n12664), .A2(n12663), .ZN(n12668) );
  INV_X1 U14954 ( .A(n12864), .ZN(n12679) );
  XNOR2_X1 U14955 ( .A(n12670), .B(n12669), .ZN(n12672) );
  NAND2_X1 U14956 ( .A1(n12863), .A2(n15126), .ZN(n12678) );
  OAI22_X1 U14957 ( .A1(n15126), .A2(n12674), .B1(n12673), .B2(n15121), .ZN(
        n12675) );
  AOI21_X1 U14958 ( .B1(n12676), .B2(n12813), .A(n12675), .ZN(n12677) );
  OAI211_X1 U14959 ( .C1(n12679), .C2(n12694), .A(n12678), .B(n12677), .ZN(
        P3_U3209) );
  AND2_X1 U14960 ( .A1(n12681), .A2(n12680), .ZN(n12683) );
  OAI21_X2 U14961 ( .B1(n12683), .B2(n7407), .A(n12682), .ZN(n12867) );
  XNOR2_X1 U14962 ( .A(n12684), .B(n7407), .ZN(n12685) );
  NAND2_X1 U14963 ( .A1(n12685), .A2(n12804), .ZN(n12687) );
  OAI211_X1 U14964 ( .C1(n15164), .C2(n12867), .A(n12687), .B(n12686), .ZN(
        n12868) );
  NAND2_X1 U14965 ( .A1(n12868), .A2(n15126), .ZN(n12693) );
  OAI22_X1 U14966 ( .A1(n15126), .A2(n12689), .B1(n12688), .B2(n15121), .ZN(
        n12690) );
  AOI21_X1 U14967 ( .B1(n12691), .B2(n12813), .A(n12690), .ZN(n12692) );
  OAI211_X1 U14968 ( .C1(n12867), .C2(n12694), .A(n12693), .B(n12692), .ZN(
        P3_U3210) );
  XNOR2_X1 U14969 ( .A(n12696), .B(n12695), .ZN(n12943) );
  XNOR2_X1 U14970 ( .A(n12698), .B(n12697), .ZN(n12700) );
  OAI21_X1 U14971 ( .B1(n12700), .B2(n15117), .A(n12699), .ZN(n12872) );
  NAND2_X1 U14972 ( .A1(n12872), .A2(n15126), .ZN(n12705) );
  OAI22_X1 U14973 ( .A1(n15126), .A2(n12702), .B1(n12701), .B2(n15121), .ZN(
        n12703) );
  AOI21_X1 U14974 ( .B1(n12873), .B2(n12798), .A(n12703), .ZN(n12704) );
  OAI211_X1 U14975 ( .C1(n12802), .C2(n12943), .A(n12705), .B(n12704), .ZN(
        P3_U3211) );
  XNOR2_X1 U14976 ( .A(n12706), .B(n12707), .ZN(n12947) );
  XNOR2_X1 U14977 ( .A(n12708), .B(n12707), .ZN(n12711) );
  INV_X1 U14978 ( .A(n12709), .ZN(n12710) );
  OAI21_X1 U14979 ( .B1(n12711), .B2(n15117), .A(n12710), .ZN(n12876) );
  NAND2_X1 U14980 ( .A1(n12876), .A2(n15126), .ZN(n12715) );
  OAI22_X1 U14981 ( .A1(n15126), .A2(n12712), .B1(n7454), .B2(n15121), .ZN(
        n12713) );
  AOI21_X1 U14982 ( .B1(n12877), .B2(n12813), .A(n12713), .ZN(n12714) );
  OAI211_X1 U14983 ( .C1(n12802), .C2(n12947), .A(n12715), .B(n12714), .ZN(
        P3_U3212) );
  OAI21_X1 U14984 ( .B1(n7439), .B2(n12720), .A(n12716), .ZN(n12953) );
  NAND2_X1 U14985 ( .A1(n12748), .A2(n12747), .ZN(n12746) );
  INV_X1 U14986 ( .A(n12717), .ZN(n12718) );
  NAND2_X1 U14987 ( .A1(n12746), .A2(n12718), .ZN(n12731) );
  NAND2_X1 U14988 ( .A1(n12731), .A2(n12719), .ZN(n12721) );
  XNOR2_X1 U14989 ( .A(n12721), .B(n12720), .ZN(n12723) );
  AOI21_X1 U14990 ( .B1(n12723), .B2(n12804), .A(n12722), .ZN(n12948) );
  MUX2_X1 U14991 ( .A(n12724), .B(n12948), .S(n15126), .Z(n12728) );
  INV_X1 U14992 ( .A(n12725), .ZN(n12726) );
  AOI22_X1 U14993 ( .A1(n12950), .A2(n12813), .B1(n12797), .B2(n12726), .ZN(
        n12727) );
  OAI211_X1 U14994 ( .C1(n12802), .C2(n12953), .A(n12728), .B(n12727), .ZN(
        P3_U3213) );
  NAND2_X1 U14995 ( .A1(n12744), .A2(n12729), .ZN(n12730) );
  XOR2_X1 U14996 ( .A(n12732), .B(n12730), .Z(n12959) );
  INV_X1 U14997 ( .A(n12731), .ZN(n12735) );
  AOI21_X1 U14998 ( .B1(n12746), .B2(n12733), .A(n12732), .ZN(n12734) );
  NOR3_X1 U14999 ( .A1(n12735), .A2(n12734), .A3(n15117), .ZN(n12737) );
  NOR2_X1 U15000 ( .A1(n12737), .A2(n12736), .ZN(n12954) );
  MUX2_X1 U15001 ( .A(n12738), .B(n12954), .S(n15126), .Z(n12742) );
  INV_X1 U15002 ( .A(n12739), .ZN(n12740) );
  AOI22_X1 U15003 ( .A1(n12956), .A2(n12813), .B1(n12797), .B2(n12740), .ZN(
        n12741) );
  OAI211_X1 U15004 ( .C1(n12802), .C2(n12959), .A(n12742), .B(n12741), .ZN(
        P3_U3214) );
  INV_X1 U15005 ( .A(n12744), .ZN(n12745) );
  AOI21_X1 U15006 ( .B1(n12743), .B2(n12747), .A(n12745), .ZN(n12963) );
  INV_X1 U15007 ( .A(n12963), .ZN(n12756) );
  OAI21_X1 U15008 ( .B1(n12748), .B2(n12747), .A(n12746), .ZN(n12750) );
  AOI21_X1 U15009 ( .B1(n12750), .B2(n12804), .A(n12749), .ZN(n12960) );
  MUX2_X1 U15010 ( .A(n12751), .B(n12960), .S(n15126), .Z(n12755) );
  INV_X1 U15011 ( .A(n12752), .ZN(n12753) );
  AOI22_X1 U15012 ( .A1(n12962), .A2(n12813), .B1(n12797), .B2(n12753), .ZN(
        n12754) );
  OAI211_X1 U15013 ( .C1(n12802), .C2(n12756), .A(n12755), .B(n12754), .ZN(
        P3_U3215) );
  XNOR2_X1 U15014 ( .A(n12757), .B(n12758), .ZN(n12969) );
  INV_X1 U15015 ( .A(n12969), .ZN(n12765) );
  XNOR2_X1 U15016 ( .A(n12759), .B(n12758), .ZN(n12761) );
  AOI21_X1 U15017 ( .B1(n12761), .B2(n12804), .A(n12760), .ZN(n12966) );
  MUX2_X1 U15018 ( .A(n14443), .B(n12966), .S(n15126), .Z(n12764) );
  AOI22_X1 U15019 ( .A1(n12968), .A2(n12798), .B1(n12797), .B2(n12762), .ZN(
        n12763) );
  OAI211_X1 U15020 ( .C1(n12802), .C2(n12765), .A(n12764), .B(n12763), .ZN(
        P3_U3216) );
  XNOR2_X1 U15021 ( .A(n12766), .B(n12768), .ZN(n12975) );
  INV_X1 U15022 ( .A(n12975), .ZN(n12776) );
  XOR2_X1 U15023 ( .A(n12768), .B(n12767), .Z(n12770) );
  AOI21_X1 U15024 ( .B1(n12770), .B2(n12804), .A(n12769), .ZN(n12972) );
  MUX2_X1 U15025 ( .A(n12771), .B(n12972), .S(n15126), .Z(n12775) );
  INV_X1 U15026 ( .A(n12772), .ZN(n12773) );
  AOI22_X1 U15027 ( .A1(n12798), .A2(n12974), .B1(n12797), .B2(n12773), .ZN(
        n12774) );
  OAI211_X1 U15028 ( .C1(n12802), .C2(n12776), .A(n12775), .B(n12774), .ZN(
        P3_U3217) );
  XNOR2_X1 U15029 ( .A(n12777), .B(n12778), .ZN(n12982) );
  XNOR2_X1 U15030 ( .A(n12779), .B(n12778), .ZN(n12781) );
  OAI21_X1 U15031 ( .B1(n12781), .B2(n15117), .A(n12780), .ZN(n12895) );
  NAND2_X1 U15032 ( .A1(n12895), .A2(n15126), .ZN(n12785) );
  OAI22_X1 U15033 ( .A1(n15126), .A2(n14402), .B1(n12782), .B2(n15121), .ZN(
        n12783) );
  AOI21_X1 U15034 ( .B1(n12813), .B2(n12896), .A(n12783), .ZN(n12784) );
  OAI211_X1 U15035 ( .C1(n12802), .C2(n12982), .A(n12785), .B(n12784), .ZN(
        P3_U3218) );
  OAI21_X1 U15036 ( .B1(n12787), .B2(n9769), .A(n12786), .ZN(n12987) );
  INV_X1 U15037 ( .A(n12987), .ZN(n12801) );
  NOR3_X1 U15038 ( .A1(n12807), .A2(n12789), .A3(n12788), .ZN(n12790) );
  NOR2_X1 U15039 ( .A1(n12790), .A2(n15117), .ZN(n12793) );
  AOI21_X1 U15040 ( .B1(n12793), .B2(n12792), .A(n12791), .ZN(n12983) );
  MUX2_X1 U15041 ( .A(n12794), .B(n12983), .S(n15126), .Z(n12800) );
  INV_X1 U15042 ( .A(n12795), .ZN(n12796) );
  AOI22_X1 U15043 ( .A1(n12798), .A2(n9693), .B1(n12797), .B2(n12796), .ZN(
        n12799) );
  OAI211_X1 U15044 ( .C1(n12802), .C2(n12801), .A(n12800), .B(n12799), .ZN(
        P3_U3219) );
  NAND3_X1 U15045 ( .A1(n12819), .A2(n12815), .A3(n12803), .ZN(n12805) );
  NAND2_X1 U15046 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  OR2_X1 U15047 ( .A1(n12807), .A2(n12806), .ZN(n12810) );
  INV_X1 U15048 ( .A(n12808), .ZN(n12809) );
  INV_X1 U15049 ( .A(n14450), .ZN(n12814) );
  OAI22_X1 U15050 ( .A1(n15126), .A2(n9076), .B1(n12811), .B2(n15121), .ZN(
        n12812) );
  AOI21_X1 U15051 ( .B1(n12814), .B2(n12813), .A(n12812), .ZN(n12818) );
  XNOR2_X1 U15052 ( .A(n12816), .B(n12815), .ZN(n14449) );
  NAND2_X1 U15053 ( .A1(n14449), .A2(n12844), .ZN(n12817) );
  OAI211_X1 U15054 ( .C1(n14453), .C2(n15128), .A(n12818), .B(n12817), .ZN(
        P3_U3220) );
  AOI211_X1 U15055 ( .C1(n12824), .C2(n12820), .A(n15117), .B(n9691), .ZN(
        n12822) );
  OR2_X1 U15056 ( .A1(n12822), .A2(n12821), .ZN(n12905) );
  INV_X1 U15057 ( .A(n12905), .ZN(n12831) );
  OAI21_X1 U15058 ( .B1(n12825), .B2(n12824), .A(n12823), .ZN(n12906) );
  NOR2_X1 U15059 ( .A1(n15126), .A2(n12826), .ZN(n12829) );
  OAI22_X1 U15060 ( .A1(n12841), .A2(n12993), .B1(n12827), .B2(n15121), .ZN(
        n12828) );
  AOI211_X1 U15061 ( .C1(n12906), .C2(n12844), .A(n12829), .B(n12828), .ZN(
        n12830) );
  OAI21_X1 U15062 ( .B1(n12831), .B2(n15128), .A(n12830), .ZN(P3_U3221) );
  XNOR2_X1 U15063 ( .A(n12832), .B(n12833), .ZN(n12836) );
  INV_X1 U15064 ( .A(n12834), .ZN(n12835) );
  OAI21_X1 U15065 ( .B1(n12836), .B2(n15117), .A(n12835), .ZN(n12908) );
  INV_X1 U15066 ( .A(n12908), .ZN(n12846) );
  OAI21_X1 U15067 ( .B1(n12838), .B2(n9766), .A(n12837), .ZN(n12909) );
  NOR2_X1 U15068 ( .A1(n15126), .A2(n12839), .ZN(n12843) );
  OAI22_X1 U15069 ( .A1(n12841), .A2(n12997), .B1(n12840), .B2(n15121), .ZN(
        n12842) );
  AOI211_X1 U15070 ( .C1(n12909), .C2(n12844), .A(n12843), .B(n12842), .ZN(
        n12845) );
  OAI21_X1 U15071 ( .B1(n12846), .B2(n15128), .A(n12845), .ZN(P3_U3222) );
  NAND2_X1 U15072 ( .A1(n12912), .A2(n15205), .ZN(n12848) );
  NAND2_X1 U15073 ( .A1(n15203), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12847) );
  OAI211_X1 U15074 ( .C1(n12914), .C2(n12911), .A(n12848), .B(n12847), .ZN(
        P3_U3490) );
  NAND2_X1 U15075 ( .A1(n15203), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12849) );
  OAI211_X1 U15076 ( .C1(n12850), .C2(n12911), .A(n12849), .B(n12848), .ZN(
        P3_U3489) );
  MUX2_X1 U15077 ( .A(n12851), .B(n12919), .S(n15205), .Z(n12853) );
  NAND2_X1 U15078 ( .A1(n12921), .A2(n12901), .ZN(n12852) );
  OAI211_X1 U15079 ( .C1(n12899), .C2(n12924), .A(n12853), .B(n12852), .ZN(
        P3_U3487) );
  AOI21_X1 U15080 ( .B1(n15167), .B2(n12855), .A(n12854), .ZN(n12925) );
  MUX2_X1 U15081 ( .A(n12856), .B(n12925), .S(n15205), .Z(n12857) );
  OAI21_X1 U15082 ( .B1(n12899), .B2(n12928), .A(n12857), .ZN(P3_U3486) );
  INV_X1 U15083 ( .A(n12858), .ZN(n12931) );
  INV_X1 U15084 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12861) );
  INV_X1 U15085 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12865) );
  AOI21_X1 U15086 ( .B1(n15182), .B2(n12864), .A(n12863), .ZN(n12932) );
  MUX2_X1 U15087 ( .A(n12865), .B(n12932), .S(n15205), .Z(n12866) );
  INV_X1 U15088 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12870) );
  INV_X1 U15089 ( .A(n12867), .ZN(n12869) );
  AOI21_X1 U15090 ( .B1(n15182), .B2(n12869), .A(n12868), .ZN(n12936) );
  MUX2_X1 U15091 ( .A(n12870), .B(n12936), .S(n15205), .Z(n12871) );
  OAI21_X1 U15092 ( .B1(n12939), .B2(n12911), .A(n12871), .ZN(P3_U3482) );
  INV_X1 U15093 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12874) );
  AOI21_X1 U15094 ( .B1(n15167), .B2(n12873), .A(n12872), .ZN(n12940) );
  MUX2_X1 U15095 ( .A(n12874), .B(n12940), .S(n15205), .Z(n12875) );
  OAI21_X1 U15096 ( .B1(n12943), .B2(n12899), .A(n12875), .ZN(P3_U3481) );
  INV_X1 U15097 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12878) );
  AOI21_X1 U15098 ( .B1(n15167), .B2(n12877), .A(n12876), .ZN(n12944) );
  MUX2_X1 U15099 ( .A(n12878), .B(n12944), .S(n15205), .Z(n12879) );
  OAI21_X1 U15100 ( .B1(n12899), .B2(n12947), .A(n12879), .ZN(P3_U3480) );
  INV_X1 U15101 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12880) );
  MUX2_X1 U15102 ( .A(n12880), .B(n12948), .S(n15205), .Z(n12882) );
  NAND2_X1 U15103 ( .A1(n12950), .A2(n12901), .ZN(n12881) );
  OAI211_X1 U15104 ( .C1(n12899), .C2(n12953), .A(n12882), .B(n12881), .ZN(
        P3_U3479) );
  MUX2_X1 U15105 ( .A(n12883), .B(n12954), .S(n15205), .Z(n12885) );
  NAND2_X1 U15106 ( .A1(n12956), .A2(n12901), .ZN(n12884) );
  OAI211_X1 U15107 ( .C1(n12959), .C2(n12899), .A(n12885), .B(n12884), .ZN(
        P3_U3478) );
  INV_X1 U15108 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12886) );
  MUX2_X1 U15109 ( .A(n12886), .B(n12960), .S(n15205), .Z(n12888) );
  INV_X1 U15110 ( .A(n12899), .ZN(n12902) );
  AOI22_X1 U15111 ( .A1(n12963), .A2(n12902), .B1(n12901), .B2(n12962), .ZN(
        n12887) );
  NAND2_X1 U15112 ( .A1(n12888), .A2(n12887), .ZN(P3_U3477) );
  MUX2_X1 U15113 ( .A(n12889), .B(n12966), .S(n15205), .Z(n12891) );
  AOI22_X1 U15114 ( .A1(n12969), .A2(n12902), .B1(n12901), .B2(n12968), .ZN(
        n12890) );
  NAND2_X1 U15115 ( .A1(n12891), .A2(n12890), .ZN(P3_U3476) );
  MUX2_X1 U15116 ( .A(n12892), .B(n12972), .S(n15205), .Z(n12894) );
  AOI22_X1 U15117 ( .A1(n12975), .A2(n12902), .B1(n12901), .B2(n12974), .ZN(
        n12893) );
  NAND2_X1 U15118 ( .A1(n12894), .A2(n12893), .ZN(P3_U3475) );
  AOI21_X1 U15119 ( .B1(n15167), .B2(n12896), .A(n12895), .ZN(n12978) );
  MUX2_X1 U15120 ( .A(n12897), .B(n12978), .S(n15205), .Z(n12898) );
  OAI21_X1 U15121 ( .B1(n12899), .B2(n12982), .A(n12898), .ZN(P3_U3474) );
  MUX2_X1 U15122 ( .A(n12900), .B(n12983), .S(n15205), .Z(n12904) );
  AOI22_X1 U15123 ( .A1(n12987), .A2(n12902), .B1(n9693), .B2(n12901), .ZN(
        n12903) );
  NAND2_X1 U15124 ( .A1(n12904), .A2(n12903), .ZN(P3_U3473) );
  AOI21_X1 U15125 ( .B1(n15190), .B2(n12906), .A(n12905), .ZN(n12990) );
  MUX2_X1 U15126 ( .A(n9861), .B(n12990), .S(n15205), .Z(n12907) );
  OAI21_X1 U15127 ( .B1(n12993), .B2(n12911), .A(n12907), .ZN(P3_U3471) );
  AOI21_X1 U15128 ( .B1(n15190), .B2(n12909), .A(n12908), .ZN(n12994) );
  MUX2_X1 U15129 ( .A(n9043), .B(n12994), .S(n15205), .Z(n12910) );
  OAI21_X1 U15130 ( .B1(n12911), .B2(n12997), .A(n12910), .ZN(P3_U3470) );
  NAND2_X1 U15131 ( .A1(n15193), .A2(n12912), .ZN(n12916) );
  NAND2_X1 U15132 ( .A1(n15191), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12913) );
  OAI211_X1 U15133 ( .C1(n12914), .C2(n12998), .A(n12916), .B(n12913), .ZN(
        P3_U3458) );
  INV_X1 U15134 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12918) );
  NAND2_X1 U15135 ( .A1(n12915), .A2(n12985), .ZN(n12917) );
  OAI211_X1 U15136 ( .C1(n12918), .C2(n15193), .A(n12917), .B(n12916), .ZN(
        P3_U3457) );
  INV_X1 U15137 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12920) );
  MUX2_X1 U15138 ( .A(n12920), .B(n12919), .S(n15193), .Z(n12923) );
  NAND2_X1 U15139 ( .A1(n12921), .A2(n12985), .ZN(n12922) );
  OAI211_X1 U15140 ( .C1(n12924), .C2(n12981), .A(n12923), .B(n12922), .ZN(
        P3_U3455) );
  INV_X1 U15141 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12926) );
  MUX2_X1 U15142 ( .A(n12926), .B(n12925), .S(n15193), .Z(n12927) );
  OAI21_X1 U15143 ( .B1(n12928), .B2(n12981), .A(n12927), .ZN(P3_U3454) );
  MUX2_X1 U15144 ( .A(n12933), .B(n12932), .S(n15193), .Z(n12934) );
  MUX2_X1 U15145 ( .A(n12937), .B(n12936), .S(n15193), .Z(n12938) );
  OAI21_X1 U15146 ( .B1(n12939), .B2(n12998), .A(n12938), .ZN(P3_U3450) );
  MUX2_X1 U15147 ( .A(n12941), .B(n12940), .S(n15193), .Z(n12942) );
  OAI21_X1 U15148 ( .B1(n12943), .B2(n12981), .A(n12942), .ZN(P3_U3449) );
  MUX2_X1 U15149 ( .A(n12945), .B(n12944), .S(n15193), .Z(n12946) );
  OAI21_X1 U15150 ( .B1(n12947), .B2(n12981), .A(n12946), .ZN(P3_U3448) );
  MUX2_X1 U15151 ( .A(n12949), .B(n12948), .S(n15193), .Z(n12952) );
  NAND2_X1 U15152 ( .A1(n12950), .A2(n12985), .ZN(n12951) );
  OAI211_X1 U15153 ( .C1(n12953), .C2(n12981), .A(n12952), .B(n12951), .ZN(
        P3_U3447) );
  INV_X1 U15154 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12955) );
  MUX2_X1 U15155 ( .A(n12955), .B(n12954), .S(n15193), .Z(n12958) );
  NAND2_X1 U15156 ( .A1(n12956), .A2(n12985), .ZN(n12957) );
  OAI211_X1 U15157 ( .C1(n12959), .C2(n12981), .A(n12958), .B(n12957), .ZN(
        P3_U3446) );
  MUX2_X1 U15158 ( .A(n12961), .B(n12960), .S(n15193), .Z(n12965) );
  INV_X1 U15159 ( .A(n12981), .ZN(n12986) );
  AOI22_X1 U15160 ( .A1(n12963), .A2(n12986), .B1(n12985), .B2(n12962), .ZN(
        n12964) );
  NAND2_X1 U15161 ( .A1(n12965), .A2(n12964), .ZN(P3_U3444) );
  INV_X1 U15162 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12967) );
  MUX2_X1 U15163 ( .A(n12967), .B(n12966), .S(n15193), .Z(n12971) );
  AOI22_X1 U15164 ( .A1(n12969), .A2(n12986), .B1(n12985), .B2(n12968), .ZN(
        n12970) );
  NAND2_X1 U15165 ( .A1(n12971), .A2(n12970), .ZN(P3_U3441) );
  INV_X1 U15166 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12973) );
  MUX2_X1 U15167 ( .A(n12973), .B(n12972), .S(n15193), .Z(n12977) );
  AOI22_X1 U15168 ( .A1(n12975), .A2(n12986), .B1(n12985), .B2(n12974), .ZN(
        n12976) );
  NAND2_X1 U15169 ( .A1(n12977), .A2(n12976), .ZN(P3_U3438) );
  INV_X1 U15170 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12979) );
  MUX2_X1 U15171 ( .A(n12979), .B(n12978), .S(n15193), .Z(n12980) );
  OAI21_X1 U15172 ( .B1(n12982), .B2(n12981), .A(n12980), .ZN(P3_U3435) );
  INV_X1 U15173 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12984) );
  MUX2_X1 U15174 ( .A(n12984), .B(n12983), .S(n15193), .Z(n12989) );
  AOI22_X1 U15175 ( .A1(n12987), .A2(n12986), .B1(n9693), .B2(n12985), .ZN(
        n12988) );
  NAND2_X1 U15176 ( .A1(n12989), .A2(n12988), .ZN(P3_U3432) );
  INV_X1 U15177 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12991) );
  MUX2_X1 U15178 ( .A(n12991), .B(n12990), .S(n15193), .Z(n12992) );
  OAI21_X1 U15179 ( .B1(n12993), .B2(n12998), .A(n12992), .ZN(P3_U3426) );
  INV_X1 U15180 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12995) );
  MUX2_X1 U15181 ( .A(n12995), .B(n12994), .S(n15193), .Z(n12996) );
  OAI21_X1 U15182 ( .B1(n12998), .B2(n12997), .A(n12996), .ZN(P3_U3423) );
  MUX2_X1 U15183 ( .A(n12999), .B(P3_D_REG_1__SCAN_IN), .S(n13000), .Z(
        P3_U3377) );
  MUX2_X1 U15184 ( .A(n13001), .B(P3_D_REG_0__SCAN_IN), .S(n13000), .Z(
        P3_U3376) );
  NAND3_X1 U15185 ( .A1(n13003), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13006) );
  OAI22_X1 U15186 ( .A1(n13002), .A2(n13006), .B1(n13005), .B2(n13004), .ZN(
        n13007) );
  AOI21_X1 U15187 ( .B1(n13008), .B2(n14381), .A(n13007), .ZN(n13009) );
  INV_X1 U15188 ( .A(n13009), .ZN(P3_U3264) );
  OAI211_X1 U15189 ( .C1(n13012), .C2(n13011), .A(n13010), .B(n13126), .ZN(
        n13017) );
  INV_X1 U15190 ( .A(n13322), .ZN(n13015) );
  AOI22_X1 U15191 ( .A1(n13285), .A2(n13521), .B1(n13523), .B2(n13346), .ZN(
        n13314) );
  OAI22_X1 U15192 ( .A1(n13101), .A2(n13314), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13013), .ZN(n13014) );
  AOI21_X1 U15193 ( .B1(n13015), .B2(n13098), .A(n13014), .ZN(n13016) );
  OAI211_X1 U15194 ( .C1(n13319), .C2(n13139), .A(n13017), .B(n13016), .ZN(
        P2_U3186) );
  AOI22_X1 U15195 ( .A1(n13136), .A2(n13155), .B1(n13135), .B2(n13157), .ZN(
        n13025) );
  AOI22_X1 U15196 ( .A1(n13019), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n13018), 
        .B2(n14467), .ZN(n13024) );
  OAI21_X1 U15197 ( .B1(n13021), .B2(n13020), .A(n10585), .ZN(n13022) );
  NAND2_X1 U15198 ( .A1(n13022), .A2(n13126), .ZN(n13023) );
  NAND3_X1 U15199 ( .A1(n13025), .A2(n13024), .A3(n13023), .ZN(P2_U3194) );
  AOI21_X1 U15200 ( .B1(n13027), .B2(n13026), .A(n14462), .ZN(n13029) );
  NAND2_X1 U15201 ( .A1(n13029), .A2(n13028), .ZN(n13035) );
  INV_X1 U15202 ( .A(n13271), .ZN(n13240) );
  OAI22_X1 U15203 ( .A1(n13030), .A2(n13503), .B1(n13240), .B2(n13505), .ZN(
        n13406) );
  INV_X1 U15204 ( .A(n13413), .ZN(n13032) );
  OAI22_X1 U15205 ( .A1(n13032), .A2(n14470), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13031), .ZN(n13033) );
  AOI21_X1 U15206 ( .B1(n13406), .B2(n13122), .A(n13033), .ZN(n13034) );
  OAI211_X1 U15207 ( .C1(n13222), .C2(n13139), .A(n13035), .B(n13034), .ZN(
        P2_U3195) );
  AOI211_X1 U15208 ( .C1(n13037), .C2(n13036), .A(n14462), .B(n13119), .ZN(
        n13041) );
  AOI22_X1 U15209 ( .A1(n13098), .A2(n13354), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13039) );
  AOI22_X1 U15210 ( .A1(n13347), .A2(n13135), .B1(n13136), .B2(n13346), .ZN(
        n13038) );
  OAI211_X1 U15211 ( .C1(n13223), .C2(n13139), .A(n13039), .B(n13038), .ZN(
        n13040) );
  OR2_X1 U15212 ( .A1(n13041), .A2(n13040), .ZN(P2_U3197) );
  INV_X1 U15213 ( .A(n13057), .ZN(n13042) );
  AOI21_X1 U15214 ( .B1(n13044), .B2(n13043), .A(n13042), .ZN(n13049) );
  INV_X1 U15215 ( .A(n13484), .ZN(n13046) );
  AOI22_X1 U15216 ( .A1(n13136), .A2(n13481), .B1(n13135), .B2(n13480), .ZN(
        n13045) );
  NAND2_X1 U15217 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14847)
         );
  OAI211_X1 U15218 ( .C1(n14470), .C2(n13046), .A(n13045), .B(n14847), .ZN(
        n13047) );
  AOI21_X1 U15219 ( .B1(n13485), .B2(n14467), .A(n13047), .ZN(n13048) );
  OAI21_X1 U15220 ( .B1(n13049), .B2(n14462), .A(n13048), .ZN(P2_U3198) );
  INV_X1 U15221 ( .A(n13050), .ZN(n13467) );
  AOI22_X1 U15222 ( .A1(n13136), .A2(n13267), .B1(n13135), .B2(n13264), .ZN(
        n13051) );
  NAND2_X1 U15223 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14863)
         );
  OAI211_X1 U15224 ( .C1(n14470), .C2(n13467), .A(n13051), .B(n14863), .ZN(
        n13052) );
  AOI21_X1 U15225 ( .B1(n13618), .B2(n14467), .A(n13052), .ZN(n13059) );
  INV_X1 U15226 ( .A(n13053), .ZN(n13056) );
  INV_X1 U15227 ( .A(n13264), .ZN(n13502) );
  OAI22_X1 U15228 ( .A1(n13054), .A2(n14462), .B1(n13502), .B2(n13132), .ZN(
        n13055) );
  NAND3_X1 U15229 ( .A1(n13057), .A2(n13056), .A3(n13055), .ZN(n13058) );
  OAI211_X1 U15230 ( .C1(n13060), .C2(n14462), .A(n13059), .B(n13058), .ZN(
        P2_U3200) );
  INV_X1 U15231 ( .A(n13578), .ZN(n13245) );
  OAI21_X1 U15232 ( .B1(n13063), .B2(n13062), .A(n13061), .ZN(n13064) );
  NAND2_X1 U15233 ( .A1(n13064), .A2(n13126), .ZN(n13069) );
  INV_X1 U15234 ( .A(n13282), .ZN(n13116) );
  OAI22_X1 U15235 ( .A1(n13065), .A2(n13505), .B1(n13116), .B2(n13503), .ZN(
        n13361) );
  INV_X1 U15236 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13066) );
  OAI22_X1 U15237 ( .A1(n13366), .A2(n14470), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13066), .ZN(n13067) );
  AOI21_X1 U15238 ( .B1(n13361), .B2(n13122), .A(n13067), .ZN(n13068) );
  OAI211_X1 U15239 ( .C1(n13245), .C2(n13139), .A(n13069), .B(n13068), .ZN(
        P2_U3201) );
  OAI21_X1 U15240 ( .B1(n13071), .B2(n13078), .A(n13070), .ZN(n13072) );
  NAND2_X1 U15241 ( .A1(n13072), .A2(n13126), .ZN(n13082) );
  NAND2_X1 U15242 ( .A1(n13136), .A2(n13524), .ZN(n13073) );
  NAND2_X1 U15243 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14721) );
  OAI211_X1 U15244 ( .C1(n14470), .C2(n13074), .A(n13073), .B(n14721), .ZN(
        n13075) );
  AOI21_X1 U15245 ( .B1(n13076), .B2(n14467), .A(n13075), .ZN(n13081) );
  NOR3_X1 U15246 ( .A1(n13078), .A2(n13077), .A3(n13132), .ZN(n13079) );
  OAI21_X1 U15247 ( .B1(n13079), .B2(n13135), .A(n13154), .ZN(n13080) );
  NAND3_X1 U15248 ( .A1(n13082), .A2(n13081), .A3(n13080), .ZN(P2_U3202) );
  INV_X1 U15249 ( .A(n13270), .ZN(n13107) );
  OAI22_X1 U15250 ( .A1(n13242), .A2(n13503), .B1(n13107), .B2(n13505), .ZN(
        n13420) );
  OAI22_X1 U15251 ( .A1(n14470), .A2(n13423), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13083), .ZN(n13085) );
  INV_X1 U15252 ( .A(n13602), .ZN(n13426) );
  NOR2_X1 U15253 ( .A1(n13426), .A2(n13139), .ZN(n13084) );
  AOI211_X1 U15254 ( .C1(n13122), .C2(n13420), .A(n13085), .B(n13084), .ZN(
        n13092) );
  INV_X1 U15255 ( .A(n13086), .ZN(n13089) );
  OAI22_X1 U15256 ( .A1(n13087), .A2(n14462), .B1(n13107), .B2(n13132), .ZN(
        n13088) );
  NAND3_X1 U15257 ( .A1(n13090), .A2(n13089), .A3(n13088), .ZN(n13091) );
  OAI211_X1 U15258 ( .C1(n13093), .C2(n14462), .A(n13092), .B(n13091), .ZN(
        P2_U3205) );
  NAND2_X1 U15259 ( .A1(n13095), .A2(n13094), .ZN(n13106) );
  NAND2_X1 U15260 ( .A1(n13096), .A2(n13126), .ZN(n13105) );
  NAND3_X1 U15261 ( .A1(n13106), .A2(n13097), .A3(n13278), .ZN(n13104) );
  AOI22_X1 U15262 ( .A1(n13280), .A2(n13521), .B1(n13523), .B2(n13274), .ZN(
        n13390) );
  INV_X1 U15263 ( .A(n13400), .ZN(n13099) );
  AOI22_X1 U15264 ( .A1(n13099), .A2(n13098), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13100) );
  OAI21_X1 U15265 ( .B1(n13390), .B2(n13101), .A(n13100), .ZN(n13102) );
  AOI21_X1 U15266 ( .B1(n13591), .B2(n14467), .A(n13102), .ZN(n13103) );
  OAI211_X1 U15267 ( .C1(n13106), .C2(n13105), .A(n13104), .B(n13103), .ZN(
        P2_U3207) );
  OAI22_X1 U15268 ( .A1(n13107), .A2(n13503), .B1(n13238), .B2(n13505), .ZN(
        n13445) );
  AOI22_X1 U15269 ( .A1(n13445), .A2(n13122), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13108) );
  OAI21_X1 U15270 ( .B1(n13448), .B2(n14470), .A(n13108), .ZN(n13114) );
  INV_X1 U15271 ( .A(n13109), .ZN(n13110) );
  AOI211_X1 U15272 ( .C1(n13112), .C2(n13111), .A(n14462), .B(n13110), .ZN(
        n13113) );
  AOI211_X1 U15273 ( .C1(n13612), .C2(n14467), .A(n13114), .B(n13113), .ZN(
        n13115) );
  INV_X1 U15274 ( .A(n13115), .ZN(P2_U3210) );
  NOR2_X1 U15275 ( .A1(n13132), .A2(n13116), .ZN(n13118) );
  AOI22_X1 U15276 ( .A1(n13119), .A2(n13126), .B1(n13118), .B2(n13117), .ZN(
        n13130) );
  INV_X1 U15277 ( .A(n13120), .ZN(n13129) );
  NAND2_X1 U15278 ( .A1(n13566), .A2(n14467), .ZN(n13124) );
  NAND2_X1 U15279 ( .A1(n13282), .A2(n13523), .ZN(n13121) );
  OAI21_X1 U15280 ( .B1(n13284), .B2(n13503), .A(n13121), .ZN(n13330) );
  AOI22_X1 U15281 ( .A1(n13122), .A2(n13330), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13123) );
  OAI211_X1 U15282 ( .C1(n14470), .C2(n13335), .A(n13124), .B(n13123), .ZN(
        n13125) );
  AOI21_X1 U15283 ( .B1(n13127), .B2(n13126), .A(n13125), .ZN(n13128) );
  OAI21_X1 U15284 ( .B1(n13130), .B2(n13129), .A(n13128), .ZN(P2_U3212) );
  INV_X1 U15285 ( .A(n13131), .ZN(n13133) );
  OAI22_X1 U15286 ( .A1(n13133), .A2(n14462), .B1(n13261), .B2(n13132), .ZN(
        n13142) );
  NAND2_X1 U15287 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n14833)
         );
  OAI21_X1 U15288 ( .B1(n14470), .B2(n13498), .A(n14833), .ZN(n13134) );
  INV_X1 U15289 ( .A(n13134), .ZN(n13138) );
  AOI22_X1 U15290 ( .A1(n13136), .A2(n13264), .B1(n13135), .B2(n13257), .ZN(
        n13137) );
  OAI211_X1 U15291 ( .C1(n13629), .C2(n13139), .A(n13138), .B(n13137), .ZN(
        n13140) );
  AOI21_X1 U15292 ( .B1(n13142), .B2(n13141), .A(n13140), .ZN(n13143) );
  INV_X1 U15293 ( .A(n13143), .ZN(P2_U3213) );
  INV_X2 U15294 ( .A(P2_U3947), .ZN(n13150) );
  MUX2_X1 U15295 ( .A(n13226), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13150), .Z(
        P2_U3562) );
  MUX2_X1 U15296 ( .A(n13254), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13150), .Z(
        P2_U3561) );
  MUX2_X1 U15297 ( .A(n13144), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13150), .Z(
        P2_U3560) );
  MUX2_X1 U15298 ( .A(n13285), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13150), .Z(
        P2_U3559) );
  MUX2_X1 U15299 ( .A(n13249), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13150), .Z(
        P2_U3558) );
  MUX2_X1 U15300 ( .A(n13346), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13150), .Z(
        P2_U3557) );
  MUX2_X1 U15301 ( .A(n13282), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13150), .Z(
        P2_U3556) );
  MUX2_X1 U15302 ( .A(n13347), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13150), .Z(
        P2_U3555) );
  MUX2_X1 U15303 ( .A(n13280), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13150), .Z(
        P2_U3554) );
  MUX2_X1 U15304 ( .A(n13278), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13150), .Z(
        P2_U3553) );
  MUX2_X1 U15305 ( .A(n13274), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13150), .Z(
        P2_U3552) );
  MUX2_X1 U15306 ( .A(n13271), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13150), .Z(
        P2_U3551) );
  MUX2_X1 U15307 ( .A(n13270), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13150), .Z(
        P2_U3550) );
  MUX2_X1 U15308 ( .A(n13267), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13150), .Z(
        P2_U3549) );
  MUX2_X1 U15309 ( .A(n13481), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13150), .Z(
        P2_U3548) );
  MUX2_X1 U15310 ( .A(n13264), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13150), .Z(
        P2_U3547) );
  MUX2_X1 U15311 ( .A(n13480), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13150), .Z(
        P2_U3546) );
  MUX2_X1 U15312 ( .A(n13257), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13150), .Z(
        P2_U3545) );
  MUX2_X1 U15313 ( .A(n13145), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13150), .Z(
        P2_U3544) );
  MUX2_X1 U15314 ( .A(n13146), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13150), .Z(
        P2_U3543) );
  MUX2_X1 U15315 ( .A(n13147), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13150), .Z(
        P2_U3542) );
  MUX2_X1 U15316 ( .A(n13148), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13150), .Z(
        P2_U3541) );
  MUX2_X1 U15317 ( .A(n13149), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13150), .Z(
        P2_U3540) );
  MUX2_X1 U15318 ( .A(n13151), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13150), .Z(
        P2_U3539) );
  MUX2_X1 U15319 ( .A(n13522), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13150), .Z(
        P2_U3538) );
  MUX2_X1 U15320 ( .A(n13152), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13150), .Z(
        P2_U3537) );
  MUX2_X1 U15321 ( .A(n13524), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13150), .Z(
        P2_U3536) );
  MUX2_X1 U15322 ( .A(n13153), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13150), .Z(
        P2_U3535) );
  MUX2_X1 U15323 ( .A(n13154), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13150), .Z(
        P2_U3534) );
  MUX2_X1 U15324 ( .A(n13155), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13150), .Z(
        P2_U3533) );
  MUX2_X1 U15325 ( .A(n13156), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13150), .Z(
        P2_U3532) );
  MUX2_X1 U15326 ( .A(n13157), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13150), .Z(
        P2_U3531) );
  AOI211_X1 U15327 ( .C1(n13160), .C2(n13159), .A(n13158), .B(n14805), .ZN(
        n13161) );
  INV_X1 U15328 ( .A(n13161), .ZN(n13169) );
  AOI22_X1 U15329 ( .A1(n14849), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n13168) );
  NAND2_X1 U15330 ( .A1(n14823), .A2(n13162), .ZN(n13167) );
  OAI211_X1 U15331 ( .C1(n13165), .C2(n13164), .A(n14851), .B(n13163), .ZN(
        n13166) );
  NAND4_X1 U15332 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        P2_U3215) );
  INV_X1 U15333 ( .A(n14865), .ZN(n13171) );
  NAND2_X1 U15334 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n13171), .ZN(n13186) );
  INV_X1 U15335 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U15336 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n13171), .B1(n14865), 
        .B2(n13170), .ZN(n14859) );
  AOI22_X1 U15337 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n13172), .B1(n14856), 
        .B2(n13488), .ZN(n14853) );
  NAND2_X1 U15338 ( .A1(n14817), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U15339 ( .A1(n14817), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13173), 
        .B2(n13200), .ZN(n14813) );
  INV_X1 U15340 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13179) );
  INV_X1 U15341 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n13178) );
  AOI21_X1 U15342 ( .B1(n13175), .B2(P2_REG2_REG_7__SCAN_IN), .A(n13174), .ZN(
        n14750) );
  INV_X1 U15343 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n13176) );
  MUX2_X1 U15344 ( .A(n13176), .B(P2_REG2_REG_8__SCAN_IN), .S(n14747), .Z(
        n14749) );
  NOR2_X1 U15345 ( .A1(n14750), .A2(n14749), .ZN(n14748) );
  AOI21_X1 U15346 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n14747), .A(n14748), .ZN(
        n14761) );
  INV_X1 U15347 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13177) );
  MUX2_X1 U15348 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n13177), .S(n14759), .Z(
        n14762) );
  NAND2_X1 U15349 ( .A1(n14761), .A2(n14762), .ZN(n14760) );
  OAI21_X1 U15350 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n14759), .A(n14760), .ZN(
        n14777) );
  MUX2_X1 U15351 ( .A(n13178), .B(P2_REG2_REG_10__SCAN_IN), .S(n14772), .Z(
        n14776) );
  OR2_X1 U15352 ( .A1(n14777), .A2(n14776), .ZN(n14778) );
  OAI21_X1 U15353 ( .B1(n13178), .B2(n13196), .A(n14778), .ZN(n14786) );
  MUX2_X1 U15354 ( .A(n13179), .B(P2_REG2_REG_11__SCAN_IN), .S(n14784), .Z(
        n14787) );
  NOR2_X1 U15355 ( .A1(n14786), .A2(n14787), .ZN(n14785) );
  AOI21_X1 U15356 ( .B1(n13179), .B2(n13197), .A(n14785), .ZN(n14800) );
  MUX2_X1 U15357 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n13180), .S(n14796), .Z(
        n14799) );
  NOR2_X1 U15358 ( .A1(n14800), .A2(n14799), .ZN(n14798) );
  AOI21_X1 U15359 ( .B1(n13180), .B2(n14796), .A(n14798), .ZN(n14812) );
  NAND2_X1 U15360 ( .A1(n14813), .A2(n14812), .ZN(n14811) );
  NAND2_X1 U15361 ( .A1(n13181), .A2(n14811), .ZN(n13182) );
  NAND2_X1 U15362 ( .A1(n14822), .A2(n13182), .ZN(n13183) );
  XNOR2_X1 U15363 ( .A(n13182), .B(n13202), .ZN(n14825) );
  NAND2_X1 U15364 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14825), .ZN(n14824) );
  NAND2_X1 U15365 ( .A1(n13183), .A2(n14824), .ZN(n13184) );
  NAND2_X1 U15366 ( .A1(n13203), .A2(n13184), .ZN(n13185) );
  XNOR2_X1 U15367 ( .A(n13184), .B(n14834), .ZN(n14839) );
  NAND2_X1 U15368 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14839), .ZN(n14838) );
  NAND2_X1 U15369 ( .A1(n13185), .A2(n14838), .ZN(n14852) );
  NAND2_X1 U15370 ( .A1(n14853), .A2(n14852), .ZN(n14850) );
  OAI21_X1 U15371 ( .B1(n14856), .B2(n13488), .A(n14850), .ZN(n14858) );
  NAND2_X1 U15372 ( .A1(n14859), .A2(n14858), .ZN(n14857) );
  NAND2_X1 U15373 ( .A1(n13186), .A2(n14857), .ZN(n13187) );
  NOR2_X1 U15374 ( .A1(n13209), .A2(n13187), .ZN(n13188) );
  XNOR2_X1 U15375 ( .A(n13209), .B(n13187), .ZN(n14870) );
  NOR2_X1 U15376 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14870), .ZN(n14869) );
  NOR2_X1 U15377 ( .A1(n13188), .A2(n14869), .ZN(n13189) );
  XOR2_X1 U15378 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13189), .Z(n13215) );
  INV_X1 U15379 ( .A(n13215), .ZN(n13213) );
  XNOR2_X1 U15380 ( .A(n14865), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14862) );
  INV_X1 U15381 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13206) );
  XNOR2_X1 U15382 ( .A(n14856), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14844) );
  INV_X1 U15383 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13201) );
  XNOR2_X1 U15384 ( .A(n13202), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14828) );
  INV_X1 U15385 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n13199) );
  INV_X1 U15386 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14958) );
  INV_X1 U15387 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14955) );
  MUX2_X1 U15388 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n13193), .S(n14747), .Z(
        n14753) );
  OAI21_X1 U15389 ( .B1(n13193), .B2(n13192), .A(n14752), .ZN(n14765) );
  MUX2_X1 U15390 ( .A(n13195), .B(P2_REG1_REG_9__SCAN_IN), .S(n14759), .Z(
        n14766) );
  NOR2_X1 U15391 ( .A1(n14765), .A2(n14766), .ZN(n14764) );
  MUX2_X1 U15392 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14955), .S(n14772), .Z(
        n14774) );
  NAND2_X1 U15393 ( .A1(n14775), .A2(n14774), .ZN(n14773) );
  OAI21_X1 U15394 ( .B1(n14955), .B2(n13196), .A(n14773), .ZN(n14791) );
  MUX2_X1 U15395 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14958), .S(n14784), .Z(
        n14790) );
  MUX2_X1 U15396 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13198), .S(n14796), .Z(
        n14804) );
  NOR2_X1 U15397 ( .A1(n14803), .A2(n14804), .ZN(n14802) );
  XNOR2_X1 U15398 ( .A(n13200), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14815) );
  NAND2_X1 U15399 ( .A1(n14816), .A2(n14815), .ZN(n14814) );
  OAI21_X1 U15400 ( .B1(n13200), .B2(n13199), .A(n14814), .ZN(n14827) );
  NAND2_X1 U15401 ( .A1(n14828), .A2(n14827), .ZN(n14826) );
  NAND2_X1 U15402 ( .A1(n13203), .A2(n13204), .ZN(n13205) );
  XNOR2_X1 U15403 ( .A(n14834), .B(n13204), .ZN(n14837) );
  NAND2_X1 U15404 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14837), .ZN(n14836) );
  NAND2_X1 U15405 ( .A1(n13205), .A2(n14836), .ZN(n14845) );
  NAND2_X1 U15406 ( .A1(n14862), .A2(n14861), .ZN(n14860) );
  XNOR2_X1 U15407 ( .A(n14872), .B(n13208), .ZN(n14878) );
  NAND2_X1 U15408 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14878), .ZN(n14876) );
  NAND2_X1 U15409 ( .A1(n13209), .A2(n13208), .ZN(n13210) );
  NAND2_X1 U15410 ( .A1(n14876), .A2(n13210), .ZN(n13211) );
  XOR2_X1 U15411 ( .A(n13211), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13214) );
  OAI21_X1 U15412 ( .B1(n13214), .B2(n14805), .A(n14873), .ZN(n13212) );
  AOI21_X1 U15413 ( .B1(n13213), .B2(n14851), .A(n13212), .ZN(n13218) );
  AOI22_X1 U15414 ( .A1(n13215), .A2(n14851), .B1(n14877), .B2(n13214), .ZN(
        n13217) );
  MUX2_X1 U15415 ( .A(n13218), .B(n13217), .S(n13216), .Z(n13220) );
  NAND2_X1 U15416 ( .A1(n14849), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n13219) );
  OAI211_X1 U15417 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n11689), .A(n13220), .B(
        n13219), .ZN(P2_U3233) );
  NOR2_X2 U15418 ( .A1(n13509), .A2(n13485), .ZN(n13469) );
  AND2_X2 U15419 ( .A1(n13334), .A2(n13319), .ZN(n13321) );
  XNOR2_X1 U15420 ( .A(n13230), .B(n13543), .ZN(n13224) );
  NAND2_X1 U15421 ( .A1(n13224), .A2(n13510), .ZN(n13544) );
  AOI21_X1 U15422 ( .B1(n13225), .B2(P2_B_REG_SCAN_IN), .A(n13503), .ZN(n13253) );
  NAND2_X1 U15423 ( .A1(n13253), .A2(n13226), .ZN(n13546) );
  NOR2_X1 U15424 ( .A1(n13512), .A2(n13546), .ZN(n13234) );
  AOI21_X1 U15425 ( .B1(n13512), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13234), 
        .ZN(n13228) );
  NAND2_X1 U15426 ( .A1(n13543), .A2(n13530), .ZN(n13227) );
  OAI211_X1 U15427 ( .C1(n13544), .C2(n13515), .A(n13228), .B(n13227), .ZN(
        P2_U3234) );
  INV_X1 U15428 ( .A(n13289), .ZN(n13232) );
  OAI211_X1 U15429 ( .C1(n13548), .C2(n13232), .A(n13231), .B(n13510), .ZN(
        n13547) );
  NOR2_X1 U15430 ( .A1(n13548), .A2(n13489), .ZN(n13233) );
  AOI211_X1 U15431 ( .C1(n13512), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13234), 
        .B(n13233), .ZN(n13235) );
  OAI21_X1 U15432 ( .B1(n13515), .B2(n13547), .A(n13235), .ZN(P2_U3235) );
  INV_X1 U15433 ( .A(n13267), .ZN(n13462) );
  INV_X1 U15434 ( .A(n13612), .ZN(n13451) );
  NAND2_X1 U15435 ( .A1(n13636), .A2(n13504), .ZN(n13236) );
  INV_X1 U15436 ( .A(n13508), .ZN(n13260) );
  AOI22_X1 U15437 ( .A1(n13499), .A2(n13260), .B1(n13261), .B2(n13513), .ZN(
        n13479) );
  NAND2_X1 U15438 ( .A1(n13479), .A2(n13494), .ZN(n13478) );
  OAI21_X1 U15439 ( .B1(n13502), .B2(n13485), .A(n13478), .ZN(n13460) );
  INV_X1 U15440 ( .A(n13433), .ZN(n13239) );
  OAI21_X1 U15441 ( .B1(n13222), .B2(n13274), .A(n13405), .ZN(n13241) );
  INV_X1 U15442 ( .A(n13591), .ZN(n13243) );
  INV_X1 U15443 ( .A(n13381), .ZN(n13375) );
  NAND2_X1 U15444 ( .A1(n13374), .A2(n13375), .ZN(n13373) );
  NAND2_X1 U15445 ( .A1(n13373), .A2(n13244), .ZN(n13360) );
  NAND2_X1 U15446 ( .A1(n13360), .A2(n13363), .ZN(n13359) );
  OAI21_X1 U15447 ( .B1(n13245), .B2(n13347), .A(n13359), .ZN(n13345) );
  NAND2_X1 U15448 ( .A1(n13345), .A2(n13344), .ZN(n13343) );
  INV_X1 U15449 ( .A(n13246), .ZN(n13247) );
  XNOR2_X1 U15450 ( .A(n13251), .B(n13287), .ZN(n13252) );
  AND2_X1 U15451 ( .A1(n13254), .A2(n13253), .ZN(n13255) );
  NAND2_X1 U15452 ( .A1(n13636), .A2(n13257), .ZN(n13258) );
  NAND2_X1 U15453 ( .A1(n13629), .A2(n13261), .ZN(n13262) );
  INV_X1 U15454 ( .A(n13494), .ZN(n13263) );
  NAND2_X1 U15455 ( .A1(n13485), .A2(n13264), .ZN(n13265) );
  NAND2_X1 U15456 ( .A1(n13492), .A2(n13265), .ZN(n13465) );
  OR2_X1 U15457 ( .A1(n13612), .A2(n13267), .ZN(n13268) );
  NOR2_X1 U15458 ( .A1(n13608), .A2(n13270), .ZN(n13269) );
  AND2_X1 U15459 ( .A1(n13602), .A2(n13271), .ZN(n13273) );
  NAND2_X1 U15460 ( .A1(n13409), .A2(n13408), .ZN(n13276) );
  OR2_X1 U15461 ( .A1(n13597), .A2(n13274), .ZN(n13275) );
  NAND2_X1 U15462 ( .A1(n13276), .A2(n13275), .ZN(n13395) );
  INV_X1 U15463 ( .A(n13395), .ZN(n13277) );
  NAND2_X1 U15464 ( .A1(n13591), .A2(n13278), .ZN(n13279) );
  INV_X1 U15465 ( .A(n13344), .ZN(n13350) );
  INV_X1 U15466 ( .A(n13312), .ZN(n13317) );
  XNOR2_X1 U15467 ( .A(n13288), .B(n13287), .ZN(n13552) );
  INV_X1 U15468 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13291) );
  OAI22_X1 U15469 ( .A1(n13527), .A2(n13291), .B1(n13290), .B2(n13466), .ZN(
        n13292) );
  AOI21_X1 U15470 ( .B1(n13293), .B2(n13530), .A(n13292), .ZN(n13294) );
  OAI21_X1 U15471 ( .B1(n13549), .B2(n13515), .A(n13294), .ZN(n13295) );
  AOI21_X1 U15472 ( .B1(n13552), .B2(n13534), .A(n13295), .ZN(n13296) );
  OAI21_X1 U15473 ( .B1(n13553), .B2(n13512), .A(n13296), .ZN(P2_U3236) );
  XNOR2_X1 U15474 ( .A(n13297), .B(n13298), .ZN(n13558) );
  AOI21_X1 U15475 ( .B1(n13299), .B2(n13298), .A(n13500), .ZN(n13302) );
  OAI21_X1 U15476 ( .B1(n13303), .B2(n13466), .A(n13557), .ZN(n13304) );
  NAND2_X1 U15477 ( .A1(n13304), .A2(n13527), .ZN(n13311) );
  NOR2_X1 U15478 ( .A1(n13308), .A2(n13321), .ZN(n13305) );
  INV_X1 U15479 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13307) );
  OAI22_X1 U15480 ( .A1(n13308), .A2(n13489), .B1(n13527), .B2(n13307), .ZN(
        n13309) );
  AOI21_X1 U15481 ( .B1(n7460), .B2(n13538), .A(n13309), .ZN(n13310) );
  OAI211_X1 U15482 ( .C1(n13475), .C2(n13558), .A(n13311), .B(n13310), .ZN(
        P2_U3237) );
  XNOR2_X1 U15483 ( .A(n13313), .B(n13312), .ZN(n13316) );
  INV_X1 U15484 ( .A(n13314), .ZN(n13315) );
  AOI21_X1 U15485 ( .B1(n13316), .B2(n13526), .A(n13315), .ZN(n13563) );
  XNOR2_X1 U15486 ( .A(n13318), .B(n13317), .ZN(n13564) );
  INV_X1 U15487 ( .A(n13564), .ZN(n13327) );
  NOR2_X1 U15488 ( .A1(n13319), .A2(n13334), .ZN(n13320) );
  INV_X1 U15489 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13323) );
  OAI22_X1 U15490 ( .A1(n13527), .A2(n13323), .B1(n13322), .B2(n13466), .ZN(
        n13324) );
  AOI21_X1 U15491 ( .B1(n13561), .B2(n13530), .A(n13324), .ZN(n13325) );
  OAI21_X1 U15492 ( .B1(n13559), .B2(n13515), .A(n13325), .ZN(n13326) );
  AOI21_X1 U15493 ( .B1(n13327), .B2(n13534), .A(n13326), .ZN(n13328) );
  OAI21_X1 U15494 ( .B1(n13563), .B2(n13512), .A(n13328), .ZN(P2_U3238) );
  XNOR2_X1 U15495 ( .A(n13329), .B(n13338), .ZN(n13331) );
  AOI21_X1 U15496 ( .B1(n13331), .B2(n13526), .A(n13330), .ZN(n13568) );
  NAND2_X1 U15497 ( .A1(n13566), .A2(n13352), .ZN(n13332) );
  NAND2_X1 U15498 ( .A1(n13332), .A2(n13510), .ZN(n13333) );
  NOR2_X1 U15499 ( .A1(n13334), .A2(n13333), .ZN(n13565) );
  INV_X1 U15500 ( .A(n13335), .ZN(n13336) );
  AOI22_X1 U15501 ( .A1(n13512), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13336), 
        .B2(n13529), .ZN(n13337) );
  OAI21_X1 U15502 ( .B1(n6973), .B2(n13489), .A(n13337), .ZN(n13341) );
  XNOR2_X1 U15503 ( .A(n13339), .B(n13338), .ZN(n13569) );
  NOR2_X1 U15504 ( .A1(n13569), .A2(n13475), .ZN(n13340) );
  AOI211_X1 U15505 ( .C1(n13565), .C2(n13538), .A(n13341), .B(n13340), .ZN(
        n13342) );
  OAI21_X1 U15506 ( .B1(n13568), .B2(n13512), .A(n13342), .ZN(P2_U3239) );
  OAI21_X1 U15507 ( .B1(n13345), .B2(n13344), .A(n13343), .ZN(n13348) );
  AOI222_X1 U15508 ( .A1(n13526), .A2(n13348), .B1(n13347), .B2(n13523), .C1(
        n13346), .C2(n13521), .ZN(n13574) );
  OAI21_X1 U15509 ( .B1(n13351), .B2(n13350), .A(n13349), .ZN(n13570) );
  AOI21_X1 U15510 ( .B1(n13572), .B2(n6545), .A(n10602), .ZN(n13353) );
  AND2_X1 U15511 ( .A1(n13353), .A2(n13352), .ZN(n13571) );
  NAND2_X1 U15512 ( .A1(n13571), .A2(n13538), .ZN(n13356) );
  AOI22_X1 U15513 ( .A1(n13512), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13354), 
        .B2(n13529), .ZN(n13355) );
  OAI211_X1 U15514 ( .C1(n13223), .C2(n13489), .A(n13356), .B(n13355), .ZN(
        n13357) );
  AOI21_X1 U15515 ( .B1(n13570), .B2(n13534), .A(n13357), .ZN(n13358) );
  OAI21_X1 U15516 ( .B1(n13574), .B2(n13512), .A(n13358), .ZN(P2_U3240) );
  OAI21_X1 U15517 ( .B1(n13360), .B2(n13363), .A(n13359), .ZN(n13362) );
  AOI21_X1 U15518 ( .B1(n13362), .B2(n13526), .A(n13361), .ZN(n13580) );
  NAND2_X1 U15519 ( .A1(n13364), .A2(n13363), .ZN(n13576) );
  NAND3_X1 U15520 ( .A1(n6898), .A2(n13534), .A3(n13576), .ZN(n13371) );
  INV_X1 U15521 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13365) );
  OAI22_X1 U15522 ( .A1(n13366), .A2(n13466), .B1(n13365), .B2(n13527), .ZN(
        n13367) );
  AOI21_X1 U15523 ( .B1(n13578), .B2(n13530), .A(n13367), .ZN(n13370) );
  AOI21_X1 U15524 ( .B1(n13578), .B2(n13382), .A(n10602), .ZN(n13368) );
  AND2_X1 U15525 ( .A1(n13368), .A2(n6545), .ZN(n13577) );
  NAND2_X1 U15526 ( .A1(n13577), .A2(n13538), .ZN(n13369) );
  AND3_X1 U15527 ( .A1(n13371), .A2(n13370), .A3(n13369), .ZN(n13372) );
  OAI21_X1 U15528 ( .B1(n13580), .B2(n13512), .A(n13372), .ZN(P2_U3241) );
  INV_X1 U15529 ( .A(n13583), .ZN(n13378) );
  OAI21_X1 U15530 ( .B1(n13375), .B2(n13374), .A(n13373), .ZN(n13376) );
  NAND2_X1 U15531 ( .A1(n13376), .A2(n13526), .ZN(n13589) );
  INV_X1 U15532 ( .A(n13589), .ZN(n13377) );
  AOI211_X1 U15533 ( .C1(n13529), .C2(n13379), .A(n13378), .B(n13377), .ZN(
        n13387) );
  OAI21_X1 U15534 ( .B1(n6606), .B2(n13381), .A(n13380), .ZN(n13587) );
  OAI211_X1 U15535 ( .C1(n13396), .C2(n13585), .A(n13510), .B(n13382), .ZN(
        n13584) );
  AOI22_X1 U15536 ( .A1(n13383), .A2(n13530), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13512), .ZN(n13384) );
  OAI21_X1 U15537 ( .B1(n13584), .B2(n13515), .A(n13384), .ZN(n13385) );
  AOI21_X1 U15538 ( .B1(n13587), .B2(n13534), .A(n13385), .ZN(n13386) );
  OAI21_X1 U15539 ( .B1(n13387), .B2(n13512), .A(n13386), .ZN(P2_U3242) );
  XNOR2_X1 U15540 ( .A(n13389), .B(n13388), .ZN(n13392) );
  INV_X1 U15541 ( .A(n13390), .ZN(n13391) );
  AOI21_X1 U15542 ( .B1(n13392), .B2(n13526), .A(n13391), .ZN(n13595) );
  INV_X1 U15543 ( .A(n13393), .ZN(n13394) );
  AOI21_X1 U15544 ( .B1(n7241), .B2(n13395), .A(n13394), .ZN(n13590) );
  INV_X1 U15545 ( .A(n13396), .ZN(n13398) );
  AOI21_X1 U15546 ( .B1(n13411), .B2(n13591), .A(n13470), .ZN(n13397) );
  NAND2_X1 U15547 ( .A1(n13398), .A2(n13397), .ZN(n13594) );
  INV_X1 U15548 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13399) );
  OAI22_X1 U15549 ( .A1(n13400), .A2(n13466), .B1(n13399), .B2(n13527), .ZN(
        n13401) );
  AOI21_X1 U15550 ( .B1(n13591), .B2(n13530), .A(n13401), .ZN(n13402) );
  OAI21_X1 U15551 ( .B1(n13594), .B2(n13515), .A(n13402), .ZN(n13403) );
  AOI21_X1 U15552 ( .B1(n13590), .B2(n13534), .A(n13403), .ZN(n13404) );
  OAI21_X1 U15553 ( .B1(n13595), .B2(n13512), .A(n13404), .ZN(P2_U3243) );
  XNOR2_X1 U15554 ( .A(n13405), .B(n13408), .ZN(n13407) );
  AOI21_X1 U15555 ( .B1(n13407), .B2(n13526), .A(n13406), .ZN(n13599) );
  XOR2_X1 U15556 ( .A(n13409), .B(n13408), .Z(n13600) );
  INV_X1 U15557 ( .A(n13600), .ZN(n13417) );
  AOI21_X1 U15558 ( .B1(n13597), .B2(n13422), .A(n10602), .ZN(n13412) );
  AND2_X1 U15559 ( .A1(n13412), .A2(n13411), .ZN(n13596) );
  NAND2_X1 U15560 ( .A1(n13596), .A2(n13538), .ZN(n13415) );
  AOI22_X1 U15561 ( .A1(n13413), .A2(n13529), .B1(n13512), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13414) );
  OAI211_X1 U15562 ( .C1(n13222), .C2(n13489), .A(n13415), .B(n13414), .ZN(
        n13416) );
  AOI21_X1 U15563 ( .B1(n13417), .B2(n13534), .A(n13416), .ZN(n13418) );
  OAI21_X1 U15564 ( .B1(n13599), .B2(n13512), .A(n13418), .ZN(P2_U3244) );
  XNOR2_X1 U15565 ( .A(n13419), .B(n13427), .ZN(n13421) );
  AOI21_X1 U15566 ( .B1(n13421), .B2(n13526), .A(n13420), .ZN(n13604) );
  AOI211_X1 U15567 ( .C1(n13602), .C2(n13437), .A(n10602), .B(n13410), .ZN(
        n13601) );
  INV_X1 U15568 ( .A(n13423), .ZN(n13424) );
  AOI22_X1 U15569 ( .A1(n13424), .A2(n13529), .B1(n13512), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n13425) );
  OAI21_X1 U15570 ( .B1(n13426), .B2(n13489), .A(n13425), .ZN(n13430) );
  XOR2_X1 U15571 ( .A(n13428), .B(n13427), .Z(n13605) );
  NOR2_X1 U15572 ( .A1(n13605), .A2(n13475), .ZN(n13429) );
  AOI211_X1 U15573 ( .C1(n13601), .C2(n13538), .A(n13430), .B(n13429), .ZN(
        n13431) );
  OAI21_X1 U15574 ( .B1(n13604), .B2(n13512), .A(n13431), .ZN(P2_U3245) );
  XNOR2_X1 U15575 ( .A(n13432), .B(n13433), .ZN(n13610) );
  XNOR2_X1 U15576 ( .A(n13434), .B(n13433), .ZN(n13436) );
  OAI21_X1 U15577 ( .B1(n13436), .B2(n13500), .A(n13435), .ZN(n13606) );
  INV_X1 U15578 ( .A(n13437), .ZN(n13438) );
  AOI211_X1 U15579 ( .C1(n13608), .C2(n13447), .A(n10602), .B(n13438), .ZN(
        n13607) );
  NAND2_X1 U15580 ( .A1(n13607), .A2(n13538), .ZN(n13442) );
  INV_X1 U15581 ( .A(n13439), .ZN(n13440) );
  AOI22_X1 U15582 ( .A1(n13512), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13440), 
        .B2(n13529), .ZN(n13441) );
  OAI211_X1 U15583 ( .C1(n6977), .C2(n13489), .A(n13442), .B(n13441), .ZN(
        n13443) );
  AOI21_X1 U15584 ( .B1(n13606), .B2(n13527), .A(n13443), .ZN(n13444) );
  OAI21_X1 U15585 ( .B1(n13475), .B2(n13610), .A(n13444), .ZN(P2_U3246) );
  XOR2_X1 U15586 ( .A(n13455), .B(n6548), .Z(n13446) );
  AOI21_X1 U15587 ( .B1(n13446), .B2(n13526), .A(n13445), .ZN(n13614) );
  AOI211_X1 U15588 ( .C1(n13612), .C2(n13471), .A(n10602), .B(n6978), .ZN(
        n13611) );
  INV_X1 U15589 ( .A(n13448), .ZN(n13449) );
  AOI22_X1 U15590 ( .A1(n13512), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13449), 
        .B2(n13529), .ZN(n13450) );
  OAI21_X1 U15591 ( .B1(n13451), .B2(n13489), .A(n13450), .ZN(n13457) );
  INV_X1 U15592 ( .A(n13452), .ZN(n13453) );
  AOI21_X1 U15593 ( .B1(n13455), .B2(n13454), .A(n13453), .ZN(n13615) );
  NOR2_X1 U15594 ( .A1(n13615), .A2(n13475), .ZN(n13456) );
  AOI211_X1 U15595 ( .C1(n13611), .C2(n13538), .A(n13457), .B(n13456), .ZN(
        n13458) );
  OAI21_X1 U15596 ( .B1(n13512), .B2(n13614), .A(n13458), .ZN(P2_U3247) );
  AOI21_X1 U15597 ( .B1(n13464), .B2(n13460), .A(n13459), .ZN(n13461) );
  OAI222_X1 U15598 ( .A1(n13505), .A2(n13502), .B1(n13503), .B2(n13462), .C1(
        n13500), .C2(n13461), .ZN(n13616) );
  OAI21_X1 U15599 ( .B1(n13465), .B2(n13464), .A(n13463), .ZN(n13620) );
  OAI22_X1 U15600 ( .A1(n13527), .A2(n13170), .B1(n13467), .B2(n13466), .ZN(
        n13468) );
  AOI21_X1 U15601 ( .B1(n13618), .B2(n13530), .A(n13468), .ZN(n13474) );
  INV_X1 U15602 ( .A(n13469), .ZN(n13486) );
  AOI21_X1 U15603 ( .B1(n13486), .B2(n13618), .A(n13470), .ZN(n13472) );
  AND2_X1 U15604 ( .A1(n13472), .A2(n13471), .ZN(n13617) );
  NAND2_X1 U15605 ( .A1(n13617), .A2(n13538), .ZN(n13473) );
  OAI211_X1 U15606 ( .C1(n13620), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13476) );
  AOI21_X1 U15607 ( .B1(n13616), .B2(n13527), .A(n13476), .ZN(n13477) );
  INV_X1 U15608 ( .A(n13477), .ZN(P2_U3248) );
  OAI211_X1 U15609 ( .C1(n13479), .C2(n13494), .A(n13478), .B(n13526), .ZN(
        n13483) );
  AOI22_X1 U15610 ( .A1(n13481), .A2(n13521), .B1(n13480), .B2(n13523), .ZN(
        n13482) );
  NAND2_X1 U15611 ( .A1(n13483), .A2(n13482), .ZN(n13626) );
  AOI21_X1 U15612 ( .B1(n13484), .B2(n13529), .A(n13626), .ZN(n13497) );
  INV_X1 U15613 ( .A(n13509), .ZN(n13487) );
  INV_X1 U15614 ( .A(n13485), .ZN(n13624) );
  OAI211_X1 U15615 ( .C1(n13487), .C2(n13624), .A(n13510), .B(n13486), .ZN(
        n13622) );
  INV_X1 U15616 ( .A(n13622), .ZN(n13491) );
  OAI22_X1 U15617 ( .A1(n13624), .A2(n13489), .B1(n13527), .B2(n13488), .ZN(
        n13490) );
  AOI21_X1 U15618 ( .B1(n13491), .B2(n13538), .A(n13490), .ZN(n13496) );
  NAND2_X1 U15619 ( .A1(n13493), .A2(n13494), .ZN(n13621) );
  NAND3_X1 U15620 ( .A1(n13492), .A2(n13534), .A3(n13621), .ZN(n13495) );
  OAI211_X1 U15621 ( .C1(n13497), .C2(n13512), .A(n13496), .B(n13495), .ZN(
        P2_U3249) );
  INV_X1 U15622 ( .A(n13498), .ZN(n13506) );
  XNOR2_X1 U15623 ( .A(n13499), .B(n13508), .ZN(n13501) );
  OAI222_X1 U15624 ( .A1(n13505), .A2(n13504), .B1(n13503), .B2(n13502), .C1(
        n13501), .C2(n13500), .ZN(n13630) );
  AOI21_X1 U15625 ( .B1(n13506), .B2(n13529), .A(n13630), .ZN(n13518) );
  OAI21_X1 U15626 ( .B1(n7452), .B2(n13508), .A(n13507), .ZN(n13632) );
  OAI211_X1 U15627 ( .C1(n13511), .C2(n13629), .A(n13510), .B(n13509), .ZN(
        n13628) );
  AOI22_X1 U15628 ( .A1(n13513), .A2(n13530), .B1(P2_REG2_REG_15__SCAN_IN), 
        .B2(n13512), .ZN(n13514) );
  OAI21_X1 U15629 ( .B1(n13628), .B2(n13515), .A(n13514), .ZN(n13516) );
  AOI21_X1 U15630 ( .B1(n13632), .B2(n13534), .A(n13516), .ZN(n13517) );
  OAI21_X1 U15631 ( .B1(n13518), .B2(n13512), .A(n13517), .ZN(P2_U3250) );
  OAI21_X1 U15632 ( .B1(n13520), .B2(n13533), .A(n13519), .ZN(n13525) );
  AOI222_X1 U15633 ( .A1(n13526), .A2(n13525), .B1(n13524), .B2(n13523), .C1(
        n13522), .C2(n13521), .ZN(n14916) );
  MUX2_X1 U15634 ( .A(n10017), .B(n14916), .S(n13527), .Z(n13542) );
  AOI22_X1 U15635 ( .A1(n14912), .A2(n13530), .B1(n13529), .B2(n13528), .ZN(
        n13541) );
  NAND2_X1 U15636 ( .A1(n13532), .A2(n13533), .ZN(n14913) );
  NAND3_X1 U15637 ( .A1(n13531), .A2(n14913), .A3(n13534), .ZN(n13540) );
  XNOR2_X1 U15638 ( .A(n13536), .B(n13535), .ZN(n13537) );
  NOR2_X1 U15639 ( .A1(n13537), .A2(n10602), .ZN(n14911) );
  NAND2_X1 U15640 ( .A1(n14911), .A2(n13538), .ZN(n13539) );
  NAND4_X1 U15641 ( .A1(n13542), .A2(n13541), .A3(n13540), .A4(n13539), .ZN(
        P2_U3259) );
  INV_X1 U15642 ( .A(n13543), .ZN(n13545) );
  OAI211_X1 U15643 ( .C1(n13545), .C2(n14927), .A(n13544), .B(n13546), .ZN(
        n13649) );
  MUX2_X1 U15644 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13649), .S(n14960), .Z(
        P2_U3530) );
  OAI211_X1 U15645 ( .C1(n13548), .C2(n14927), .A(n13547), .B(n13546), .ZN(
        n13650) );
  MUX2_X1 U15646 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13650), .S(n14960), .Z(
        P2_U3529) );
  OAI21_X1 U15647 ( .B1(n13550), .B2(n14927), .A(n13549), .ZN(n13551) );
  MUX2_X1 U15648 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13651), .S(n14960), .Z(
        P2_U3528) );
  AOI21_X1 U15649 ( .B1(n14936), .B2(n13555), .A(n7460), .ZN(n13556) );
  OAI211_X1 U15650 ( .C1(n14922), .C2(n13558), .A(n13557), .B(n13556), .ZN(
        n13652) );
  MUX2_X1 U15651 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13652), .S(n14960), .Z(
        P2_U3527) );
  INV_X1 U15652 ( .A(n13559), .ZN(n13560) );
  AOI21_X1 U15653 ( .B1(n14936), .B2(n13561), .A(n13560), .ZN(n13562) );
  OAI211_X1 U15654 ( .C1(n14922), .C2(n13564), .A(n13563), .B(n13562), .ZN(
        n13653) );
  MUX2_X1 U15655 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13653), .S(n14960), .Z(
        P2_U3526) );
  AOI21_X1 U15656 ( .B1(n14936), .B2(n13566), .A(n13565), .ZN(n13567) );
  OAI211_X1 U15657 ( .C1(n14922), .C2(n13569), .A(n13568), .B(n13567), .ZN(
        n13654) );
  MUX2_X1 U15658 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13654), .S(n14960), .Z(
        P2_U3525) );
  INV_X1 U15659 ( .A(n13570), .ZN(n13575) );
  AOI21_X1 U15660 ( .B1(n14936), .B2(n13572), .A(n13571), .ZN(n13573) );
  OAI211_X1 U15661 ( .C1(n14922), .C2(n13575), .A(n13574), .B(n13573), .ZN(
        n13655) );
  MUX2_X1 U15662 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13655), .S(n14960), .Z(
        P2_U3524) );
  NAND2_X1 U15663 ( .A1(n13576), .A2(n14934), .ZN(n13581) );
  AOI21_X1 U15664 ( .B1(n14936), .B2(n13578), .A(n13577), .ZN(n13579) );
  OAI211_X1 U15665 ( .C1(n13582), .C2(n13581), .A(n13580), .B(n13579), .ZN(
        n13656) );
  MUX2_X1 U15666 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13656), .S(n14960), .Z(
        P2_U3523) );
  OAI211_X1 U15667 ( .C1(n13585), .C2(n14927), .A(n13584), .B(n13583), .ZN(
        n13586) );
  AOI21_X1 U15668 ( .B1(n13587), .B2(n14934), .A(n13586), .ZN(n13588) );
  NAND2_X1 U15669 ( .A1(n13589), .A2(n13588), .ZN(n13657) );
  MUX2_X1 U15670 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13657), .S(n14960), .Z(
        P2_U3522) );
  NAND2_X1 U15671 ( .A1(n13590), .A2(n14934), .ZN(n13593) );
  NAND2_X1 U15672 ( .A1(n13591), .A2(n14936), .ZN(n13592) );
  NAND4_X1 U15673 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13658) );
  MUX2_X1 U15674 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13658), .S(n14960), .Z(
        P2_U3521) );
  AOI21_X1 U15675 ( .B1(n14936), .B2(n13597), .A(n13596), .ZN(n13598) );
  OAI211_X1 U15676 ( .C1(n14922), .C2(n13600), .A(n13599), .B(n13598), .ZN(
        n13659) );
  MUX2_X1 U15677 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13659), .S(n14960), .Z(
        P2_U3520) );
  AOI21_X1 U15678 ( .B1(n14936), .B2(n13602), .A(n13601), .ZN(n13603) );
  OAI211_X1 U15679 ( .C1(n14922), .C2(n13605), .A(n13604), .B(n13603), .ZN(
        n13660) );
  MUX2_X1 U15680 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13660), .S(n14960), .Z(
        P2_U3519) );
  AOI211_X1 U15681 ( .C1(n14936), .C2(n13608), .A(n13607), .B(n13606), .ZN(
        n13609) );
  OAI21_X1 U15682 ( .B1(n14922), .B2(n13610), .A(n13609), .ZN(n13661) );
  MUX2_X1 U15683 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13661), .S(n14960), .Z(
        P2_U3518) );
  AOI21_X1 U15684 ( .B1(n14936), .B2(n13612), .A(n13611), .ZN(n13613) );
  OAI211_X1 U15685 ( .C1(n14922), .C2(n13615), .A(n13614), .B(n13613), .ZN(
        n13662) );
  MUX2_X1 U15686 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13662), .S(n14960), .Z(
        P2_U3517) );
  AOI211_X1 U15687 ( .C1(n14936), .C2(n13618), .A(n13617), .B(n13616), .ZN(
        n13619) );
  OAI21_X1 U15688 ( .B1(n14922), .B2(n13620), .A(n13619), .ZN(n13663) );
  MUX2_X1 U15689 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13663), .S(n14960), .Z(
        P2_U3516) );
  NAND3_X1 U15690 ( .A1(n13492), .A2(n14934), .A3(n13621), .ZN(n13623) );
  OAI211_X1 U15691 ( .C1(n13624), .C2(n14927), .A(n13623), .B(n13622), .ZN(
        n13625) );
  NOR2_X1 U15692 ( .A1(n13626), .A2(n13625), .ZN(n13665) );
  NAND2_X1 U15693 ( .A1(n14957), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n13627) );
  OAI21_X1 U15694 ( .B1(n13665), .B2(n14957), .A(n13627), .ZN(P2_U3515) );
  OAI21_X1 U15695 ( .B1(n13629), .B2(n14927), .A(n13628), .ZN(n13631) );
  AOI211_X1 U15696 ( .C1(n14934), .C2(n13632), .A(n13631), .B(n13630), .ZN(
        n13667) );
  NAND2_X1 U15697 ( .A1(n14957), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n13633) );
  OAI21_X1 U15698 ( .B1(n13667), .B2(n14957), .A(n13633), .ZN(P2_U3514) );
  INV_X1 U15699 ( .A(n13634), .ZN(n13635) );
  AOI21_X1 U15700 ( .B1(n14936), .B2(n13636), .A(n13635), .ZN(n13637) );
  OAI211_X1 U15701 ( .C1(n14922), .C2(n13639), .A(n13638), .B(n13637), .ZN(
        n13668) );
  MUX2_X1 U15702 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13668), .S(n14960), .Z(
        P2_U3513) );
  AOI21_X1 U15703 ( .B1(n14936), .B2(n13641), .A(n13640), .ZN(n13643) );
  OAI211_X1 U15704 ( .C1(n14922), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        n13669) );
  MUX2_X1 U15705 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13669), .S(n14960), .Z(
        P2_U3512) );
  OAI211_X1 U15706 ( .C1(n13648), .C2(n13647), .A(n13646), .B(n13645), .ZN(
        n14891) );
  MUX2_X1 U15707 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14891), .S(n14960), .Z(
        P2_U3499) );
  MUX2_X1 U15708 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13649), .S(n14944), .Z(
        P2_U3498) );
  MUX2_X1 U15709 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13650), .S(n14944), .Z(
        P2_U3497) );
  MUX2_X1 U15710 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13652), .S(n14944), .Z(
        P2_U3495) );
  MUX2_X1 U15711 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13653), .S(n14944), .Z(
        P2_U3494) );
  MUX2_X1 U15712 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13654), .S(n14944), .Z(
        P2_U3493) );
  MUX2_X1 U15713 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13655), .S(n14944), .Z(
        P2_U3492) );
  MUX2_X1 U15714 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13656), .S(n14944), .Z(
        P2_U3491) );
  MUX2_X1 U15715 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13657), .S(n14944), .Z(
        P2_U3490) );
  MUX2_X1 U15716 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13658), .S(n14944), .Z(
        P2_U3489) );
  MUX2_X1 U15717 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13659), .S(n14944), .Z(
        P2_U3488) );
  MUX2_X1 U15718 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13660), .S(n14944), .Z(
        P2_U3487) );
  MUX2_X1 U15719 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13661), .S(n14944), .Z(
        P2_U3486) );
  MUX2_X1 U15720 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13662), .S(n14944), .Z(
        P2_U3484) );
  MUX2_X1 U15721 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13663), .S(n14944), .Z(
        P2_U3481) );
  NAND2_X1 U15722 ( .A1(n14942), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n13664) );
  OAI21_X1 U15723 ( .B1(n13665), .B2(n14942), .A(n13664), .ZN(P2_U3478) );
  NAND2_X1 U15724 ( .A1(n14942), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n13666) );
  OAI21_X1 U15725 ( .B1(n13667), .B2(n14942), .A(n13666), .ZN(P2_U3475) );
  MUX2_X1 U15726 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13668), .S(n14944), .Z(
        P2_U3472) );
  MUX2_X1 U15727 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13669), .S(n14944), .Z(
        P2_U3469) );
  INV_X1 U15728 ( .A(n13670), .ZN(n14356) );
  NOR4_X1 U15729 ( .A1(n13672), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3088), 
        .A4(n13671), .ZN(n13673) );
  AOI21_X1 U15730 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13683), .A(n13673), 
        .ZN(n13674) );
  OAI21_X1 U15731 ( .B1(n14356), .B2(n13685), .A(n13674), .ZN(P2_U3296) );
  OAI222_X1 U15732 ( .A1(n13685), .A2(n13677), .B1(n13676), .B2(P2_U3088), 
        .C1(n13675), .C2(n13688), .ZN(P2_U3297) );
  INV_X1 U15733 ( .A(n13678), .ZN(n14358) );
  OAI222_X1 U15734 ( .A1(n13685), .A2(n14358), .B1(P2_U3088), .B2(n13680), 
        .C1(n13679), .C2(n13688), .ZN(P2_U3298) );
  AOI21_X1 U15735 ( .B1(n13683), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13682), 
        .ZN(n13684) );
  OAI21_X1 U15736 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(P2_U3299) );
  INV_X1 U15737 ( .A(n13687), .ZN(n14365) );
  OAI222_X1 U15738 ( .A1(n13685), .A2(n14365), .B1(n13690), .B2(P2_U3088), 
        .C1(n13689), .C2(n13688), .ZN(P2_U3301) );
  MUX2_X1 U15739 ( .A(n13691), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15740 ( .A1(n13694), .A2(n13844), .ZN(n13699) );
  AOI22_X1 U15741 ( .A1(n13855), .A2(n13871), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13695) );
  OAI21_X1 U15742 ( .B1(n13696), .B2(n13857), .A(n13695), .ZN(n13697) );
  AOI21_X1 U15743 ( .B1(n13862), .B2(n14032), .A(n13697), .ZN(n13698) );
  OAI211_X1 U15744 ( .C1(n13700), .C2(n13858), .A(n13699), .B(n13698), .ZN(
        P1_U3214) );
  INV_X1 U15745 ( .A(n13701), .ZN(n13702) );
  AOI21_X1 U15746 ( .B1(n13704), .B2(n13703), .A(n13702), .ZN(n13711) );
  NAND2_X1 U15747 ( .A1(n13855), .A2(n13874), .ZN(n13705) );
  OAI211_X1 U15748 ( .C1(n13857), .C2(n14511), .A(n13706), .B(n13705), .ZN(
        n13707) );
  AOI21_X1 U15749 ( .B1(n13708), .B2(n13862), .A(n13707), .ZN(n13710) );
  NAND2_X1 U15750 ( .A1(n14513), .A2(n13817), .ZN(n13709) );
  OAI211_X1 U15751 ( .C1(n13711), .C2(n13864), .A(n13710), .B(n13709), .ZN(
        P1_U3215) );
  INV_X1 U15752 ( .A(n13712), .ZN(n13714) );
  NOR3_X1 U15753 ( .A1(n13715), .A2(n13714), .A3(n13713), .ZN(n13717) );
  INV_X1 U15754 ( .A(n13716), .ZN(n13794) );
  OAI21_X1 U15755 ( .B1(n13717), .B2(n13794), .A(n13844), .ZN(n13722) );
  NAND2_X1 U15756 ( .A1(n14134), .A2(n14498), .ZN(n14105) );
  NAND2_X1 U15757 ( .A1(n14112), .A2(n14642), .ZN(n13718) );
  AND2_X1 U15758 ( .A1(n14105), .A2(n13718), .ZN(n14287) );
  OAI22_X1 U15759 ( .A1(n14287), .A2(n13847), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13719), .ZN(n13720) );
  AOI21_X1 U15760 ( .B1(n14108), .B2(n13862), .A(n13720), .ZN(n13721) );
  OAI211_X1 U15761 ( .C1(n14115), .C2(n13858), .A(n13722), .B(n13721), .ZN(
        P1_U3216) );
  NAND2_X1 U15762 ( .A1(n13723), .A2(n13780), .ZN(n13783) );
  NAND2_X1 U15763 ( .A1(n13783), .A2(n13724), .ZN(n13834) );
  NAND2_X1 U15764 ( .A1(n13834), .A2(n13835), .ZN(n13833) );
  INV_X1 U15765 ( .A(n13833), .ZN(n13727) );
  OAI21_X1 U15766 ( .B1(n13727), .B2(n13726), .A(n13725), .ZN(n13729) );
  NAND3_X1 U15767 ( .A1(n13729), .A2(n13844), .A3(n13728), .ZN(n13733) );
  NOR2_X1 U15768 ( .A1(n13786), .A2(n14171), .ZN(n13731) );
  NAND2_X1 U15769 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14016)
         );
  OAI21_X1 U15770 ( .B1(n13828), .B2(n14175), .A(n14016), .ZN(n13730) );
  AOI211_X1 U15771 ( .C1(n13825), .C2(n14317), .A(n13731), .B(n13730), .ZN(
        n13732) );
  OAI211_X1 U15772 ( .C1(n14320), .C2(n13858), .A(n13733), .B(n13732), .ZN(
        P1_U3219) );
  OAI21_X1 U15773 ( .B1(n13736), .B2(n13735), .A(n13734), .ZN(n13737) );
  NAND2_X1 U15774 ( .A1(n13737), .A2(n13844), .ZN(n13741) );
  AOI22_X1 U15775 ( .A1(n13855), .A2(n10303), .B1(n13825), .B2(n8319), .ZN(
        n13740) );
  AOI22_X1 U15776 ( .A1(n14641), .A2(n13817), .B1(n13738), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n13739) );
  NAND3_X1 U15777 ( .A1(n13741), .A2(n13740), .A3(n13739), .ZN(P1_U3222) );
  AOI21_X1 U15778 ( .B1(n13743), .B2(n13742), .A(n6532), .ZN(n13748) );
  NAND2_X1 U15779 ( .A1(n14134), .A2(n13825), .ZN(n13745) );
  AOI22_X1 U15780 ( .A1(n13855), .A2(n14317), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13744) );
  OAI211_X1 U15781 ( .C1(n13786), .C2(n14139), .A(n13745), .B(n13744), .ZN(
        n13746) );
  AOI21_X1 U15782 ( .B1(n14301), .B2(n13817), .A(n13746), .ZN(n13747) );
  OAI21_X1 U15783 ( .B1(n13748), .B2(n13864), .A(n13747), .ZN(P1_U3223) );
  AND2_X1 U15784 ( .A1(n13749), .A2(n13750), .ZN(n13753) );
  OAI211_X1 U15785 ( .C1(n13753), .C2(n13752), .A(n13844), .B(n13751), .ZN(
        n13759) );
  NAND2_X1 U15786 ( .A1(n13855), .A2(n13876), .ZN(n13754) );
  OAI211_X1 U15787 ( .C1(n13857), .C2(n14510), .A(n13755), .B(n13754), .ZN(
        n13756) );
  AOI21_X1 U15788 ( .B1(n13757), .B2(n13862), .A(n13756), .ZN(n13758) );
  OAI211_X1 U15789 ( .C1(n13760), .C2(n13858), .A(n13759), .B(n13758), .ZN(
        P1_U3224) );
  NOR3_X1 U15790 ( .A1(n6533), .A2(n7315), .A3(n13762), .ZN(n13765) );
  INV_X1 U15791 ( .A(n13763), .ZN(n13764) );
  OAI21_X1 U15792 ( .B1(n13765), .B2(n13764), .A(n13844), .ZN(n13771) );
  NAND2_X1 U15793 ( .A1(n13871), .A2(n14642), .ZN(n13767) );
  NAND2_X1 U15794 ( .A1(n14112), .A2(n14498), .ZN(n13766) );
  AND2_X1 U15795 ( .A1(n13767), .A2(n13766), .ZN(n14275) );
  OAI22_X1 U15796 ( .A1(n13847), .A2(n14275), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13768), .ZN(n13769) );
  AOI21_X1 U15797 ( .B1(n13862), .B2(n14069), .A(n13769), .ZN(n13770) );
  OAI211_X1 U15798 ( .C1(n8653), .C2(n13858), .A(n13771), .B(n13770), .ZN(
        P1_U3225) );
  OAI21_X1 U15799 ( .B1(n13774), .B2(n13773), .A(n13772), .ZN(n13775) );
  NAND2_X1 U15800 ( .A1(n13775), .A2(n13844), .ZN(n13779) );
  AND2_X1 U15801 ( .A1(n13873), .A2(n14498), .ZN(n14231) );
  AOI21_X1 U15802 ( .B1(n14642), .B2(n13872), .A(n14231), .ZN(n14492) );
  OAI21_X1 U15803 ( .B1(n14492), .B2(n13847), .A(n13776), .ZN(n13777) );
  AOI21_X1 U15804 ( .B1(n13862), .B2(n7443), .A(n13777), .ZN(n13778) );
  OAI211_X1 U15805 ( .C1(n14494), .C2(n13858), .A(n13779), .B(n13778), .ZN(
        P1_U3226) );
  INV_X1 U15806 ( .A(n13772), .ZN(n13782) );
  NOR3_X1 U15807 ( .A1(n13782), .A2(n13781), .A3(n13780), .ZN(n13785) );
  INV_X1 U15808 ( .A(n13783), .ZN(n13784) );
  OAI21_X1 U15809 ( .B1(n13785), .B2(n13784), .A(n13844), .ZN(n13791) );
  NOR2_X1 U15810 ( .A1(n13786), .A2(n14207), .ZN(n13789) );
  OAI21_X1 U15811 ( .B1(n13828), .B2(n14209), .A(n13787), .ZN(n13788) );
  AOI211_X1 U15812 ( .C1(n13825), .C2(n14485), .A(n13789), .B(n13788), .ZN(
        n13790) );
  OAI211_X1 U15813 ( .C1(n14488), .C2(n13858), .A(n13791), .B(n13790), .ZN(
        P1_U3228) );
  NOR3_X1 U15814 ( .A1(n13794), .A2(n7316), .A3(n13793), .ZN(n13795) );
  OAI21_X1 U15815 ( .B1(n13795), .B2(n6533), .A(n13844), .ZN(n13800) );
  AOI22_X1 U15816 ( .A1(n13855), .A2(n14079), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13796) );
  OAI21_X1 U15817 ( .B1(n13797), .B2(n13857), .A(n13796), .ZN(n13798) );
  AOI21_X1 U15818 ( .B1(n14088), .B2(n13862), .A(n13798), .ZN(n13799) );
  OAI211_X1 U15819 ( .C1(n14341), .C2(n13858), .A(n13800), .B(n13799), .ZN(
        P1_U3229) );
  XNOR2_X1 U15820 ( .A(n13802), .B(n13801), .ZN(n13811) );
  NAND2_X1 U15821 ( .A1(n14152), .A2(n14642), .ZN(n13804) );
  NAND2_X1 U15822 ( .A1(n14199), .A2(n14498), .ZN(n13803) );
  NAND2_X1 U15823 ( .A1(n13804), .A2(n13803), .ZN(n14307) );
  NAND2_X1 U15824 ( .A1(n14307), .A2(n13805), .ZN(n13807) );
  NAND2_X1 U15825 ( .A1(n13862), .A2(n14151), .ZN(n13806) );
  OAI211_X1 U15826 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n13808), .A(n13807), .B(
        n13806), .ZN(n13809) );
  AOI21_X1 U15827 ( .B1(n14160), .B2(n13817), .A(n13809), .ZN(n13810) );
  OAI21_X1 U15828 ( .B1(n13811), .B2(n13864), .A(n13810), .ZN(P1_U3233) );
  XNOR2_X1 U15829 ( .A(n13812), .B(n13813), .ZN(n13820) );
  NAND2_X1 U15830 ( .A1(n13855), .A2(n13875), .ZN(n13814) );
  NAND2_X1 U15831 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14594)
         );
  OAI211_X1 U15832 ( .C1(n13857), .C2(n14523), .A(n13814), .B(n14594), .ZN(
        n13815) );
  AOI21_X1 U15833 ( .B1(n13816), .B2(n13862), .A(n13815), .ZN(n13819) );
  NAND2_X1 U15834 ( .A1(n14525), .A2(n13817), .ZN(n13818) );
  OAI211_X1 U15835 ( .C1(n13820), .C2(n13864), .A(n13819), .B(n13818), .ZN(
        P1_U3234) );
  INV_X1 U15836 ( .A(n13749), .ZN(n13824) );
  AOI21_X1 U15837 ( .B1(n11551), .B2(n13822), .A(n13821), .ZN(n13823) );
  OAI21_X1 U15838 ( .B1(n13824), .B2(n13823), .A(n13844), .ZN(n13832) );
  NAND2_X1 U15839 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n13985)
         );
  NAND2_X1 U15840 ( .A1(n13825), .A2(n13875), .ZN(n13826) );
  OAI211_X1 U15841 ( .C1(n13828), .C2(n13827), .A(n13985), .B(n13826), .ZN(
        n13829) );
  AOI21_X1 U15842 ( .B1(n13830), .B2(n13862), .A(n13829), .ZN(n13831) );
  OAI211_X1 U15843 ( .C1(n14531), .C2(n13858), .A(n13832), .B(n13831), .ZN(
        P1_U3236) );
  INV_X1 U15844 ( .A(n14182), .ZN(n14481) );
  OAI21_X1 U15845 ( .B1(n13835), .B2(n13834), .A(n13833), .ZN(n13836) );
  NAND2_X1 U15846 ( .A1(n13836), .A2(n13844), .ZN(n13840) );
  INV_X1 U15847 ( .A(n14194), .ZN(n13838) );
  NOR2_X1 U15848 ( .A1(n14233), .A2(n14520), .ZN(n14193) );
  AOI21_X1 U15849 ( .B1(n14642), .B2(n14199), .A(n14193), .ZN(n14479) );
  NAND2_X1 U15850 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14635)
         );
  OAI21_X1 U15851 ( .B1(n14479), .B2(n13847), .A(n14635), .ZN(n13837) );
  AOI21_X1 U15852 ( .B1(n13838), .B2(n13862), .A(n13837), .ZN(n13839) );
  OAI211_X1 U15853 ( .C1(n14481), .C2(n13858), .A(n13840), .B(n13839), .ZN(
        P1_U3238) );
  INV_X1 U15854 ( .A(n14046), .ZN(n14269) );
  OAI21_X1 U15855 ( .B1(n13843), .B2(n13842), .A(n13841), .ZN(n13845) );
  NAND2_X1 U15856 ( .A1(n13845), .A2(n13844), .ZN(n13850) );
  AOI22_X1 U15857 ( .A1(n14498), .A2(n14078), .B1(n13870), .B2(n14642), .ZN(
        n14268) );
  OAI22_X1 U15858 ( .A1(n13847), .A2(n14268), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13846), .ZN(n13848) );
  AOI21_X1 U15859 ( .B1(n13862), .B2(n14050), .A(n13848), .ZN(n13849) );
  OAI211_X1 U15860 ( .C1(n14269), .C2(n13858), .A(n13850), .B(n13849), .ZN(
        P1_U3240) );
  INV_X1 U15861 ( .A(n13851), .ZN(n13852) );
  AOI21_X1 U15862 ( .B1(n13854), .B2(n13853), .A(n13852), .ZN(n13865) );
  NAND2_X1 U15863 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14620)
         );
  NAND2_X1 U15864 ( .A1(n13855), .A2(n14499), .ZN(n13856) );
  OAI211_X1 U15865 ( .C1(n13857), .C2(n14209), .A(n14620), .B(n13856), .ZN(
        n13860) );
  NOR2_X1 U15866 ( .A1(n14503), .A2(n13858), .ZN(n13859) );
  AOI211_X1 U15867 ( .C1(n13862), .C2(n13861), .A(n13860), .B(n13859), .ZN(
        n13863) );
  OAI21_X1 U15868 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(P1_U3241) );
  MUX2_X1 U15869 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13866), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15870 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13867), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15871 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13868), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15872 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13869), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15873 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13870), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15874 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13871), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15875 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14078), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15876 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14112), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15877 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14079), .S(n13881), .Z(
        P1_U3583) );
  MUX2_X1 U15878 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14134), .S(n13881), .Z(
        P1_U3582) );
  MUX2_X1 U15879 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14152), .S(n13881), .Z(
        P1_U3581) );
  MUX2_X1 U15880 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14317), .S(n13881), .Z(
        P1_U3580) );
  MUX2_X1 U15881 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14199), .S(n13881), .Z(
        P1_U3579) );
  MUX2_X1 U15882 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14485), .S(n13881), .Z(
        P1_U3578) );
  MUX2_X1 U15883 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13872), .S(n13881), .Z(
        P1_U3577) );
  MUX2_X1 U15884 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14500), .S(n13881), .Z(
        P1_U3576) );
  MUX2_X1 U15885 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13873), .S(n13881), .Z(
        P1_U3575) );
  MUX2_X1 U15886 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14499), .S(n13881), .Z(
        P1_U3574) );
  MUX2_X1 U15887 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13874), .S(n13881), .Z(
        P1_U3573) );
  MUX2_X1 U15888 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13875), .S(n13881), .Z(
        P1_U3572) );
  MUX2_X1 U15889 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13876), .S(n13881), .Z(
        P1_U3571) );
  MUX2_X1 U15890 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13877), .S(n13881), .Z(
        P1_U3570) );
  MUX2_X1 U15891 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13878), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15892 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13879), .S(n13881), .Z(
        P1_U3568) );
  MUX2_X1 U15893 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13880), .S(n13881), .Z(
        P1_U3567) );
  MUX2_X1 U15894 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13882), .S(n13881), .Z(
        P1_U3566) );
  MUX2_X1 U15895 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13883), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15896 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13884), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15897 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13885), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15898 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8319), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15899 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14248), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15900 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10303), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15901 ( .C1(n13887), .C2(n13886), .A(n14600), .B(n13902), .ZN(
        n13893) );
  NAND2_X1 U15902 ( .A1(n14634), .A2(n13888), .ZN(n13892) );
  OAI211_X1 U15903 ( .C1(n13895), .C2(n13889), .A(n14628), .B(n13910), .ZN(
        n13891) );
  AOI22_X1 U15904 ( .A1(n14596), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13890) );
  NAND4_X1 U15905 ( .A1(n13893), .A2(n13892), .A3(n13891), .A4(n13890), .ZN(
        P1_U3244) );
  MUX2_X1 U15906 ( .A(n13895), .B(n13894), .S(n14362), .Z(n13897) );
  NAND2_X1 U15907 ( .A1(n13897), .A2(n13896), .ZN(n13899) );
  OAI211_X1 U15908 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n13900), .A(n13899), .B(
        P1_U4016), .ZN(n14592) );
  AOI22_X1 U15909 ( .A1(n14596), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13915) );
  MUX2_X1 U15910 ( .A(n10099), .B(P1_REG1_REG_2__SCAN_IN), .S(n13907), .Z(
        n13903) );
  NAND3_X1 U15911 ( .A1(n13903), .A2(n13902), .A3(n13901), .ZN(n13904) );
  NAND2_X1 U15912 ( .A1(n13904), .A2(n13922), .ZN(n13905) );
  OAI22_X1 U15913 ( .A1(n8316), .A2(n14618), .B1(n14626), .B2(n13905), .ZN(
        n13906) );
  INV_X1 U15914 ( .A(n13906), .ZN(n13914) );
  MUX2_X1 U15915 ( .A(n13908), .B(P1_REG2_REG_2__SCAN_IN), .S(n13907), .Z(
        n13911) );
  NAND3_X1 U15916 ( .A1(n13911), .A2(n13910), .A3(n13909), .ZN(n13912) );
  NAND3_X1 U15917 ( .A1(n14628), .A2(n13928), .A3(n13912), .ZN(n13913) );
  NAND4_X1 U15918 ( .A1(n14592), .A2(n13915), .A3(n13914), .A4(n13913), .ZN(
        P1_U3245) );
  OAI22_X1 U15919 ( .A1(n14637), .A2(n13916), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8322), .ZN(n13917) );
  AOI21_X1 U15920 ( .B1(n13924), .B2(n14634), .A(n13917), .ZN(n13932) );
  INV_X1 U15921 ( .A(n13918), .ZN(n13921) );
  MUX2_X1 U15922 ( .A(n13919), .B(P1_REG1_REG_3__SCAN_IN), .S(n13924), .Z(
        n13920) );
  NAND3_X1 U15923 ( .A1(n13922), .A2(n13921), .A3(n13920), .ZN(n13923) );
  NAND3_X1 U15924 ( .A1(n14600), .A2(n14577), .A3(n13923), .ZN(n13931) );
  MUX2_X1 U15925 ( .A(n13925), .B(P1_REG2_REG_3__SCAN_IN), .S(n13924), .Z(
        n13927) );
  NAND3_X1 U15926 ( .A1(n13928), .A2(n13927), .A3(n13926), .ZN(n13929) );
  NAND3_X1 U15927 ( .A1(n14628), .A2(n14585), .A3(n13929), .ZN(n13930) );
  NAND3_X1 U15928 ( .A1(n13932), .A2(n13931), .A3(n13930), .ZN(P1_U3246) );
  INV_X1 U15929 ( .A(n13933), .ZN(n13938) );
  NAND3_X1 U15930 ( .A1(n13936), .A2(n13935), .A3(n13934), .ZN(n13937) );
  NAND3_X1 U15931 ( .A1(n14600), .A2(n13938), .A3(n13937), .ZN(n13948) );
  NAND2_X1 U15932 ( .A1(n14634), .A2(n13939), .ZN(n13947) );
  MUX2_X1 U15933 ( .A(n10906), .B(P1_REG2_REG_7__SCAN_IN), .S(n13939), .Z(
        n13942) );
  NAND3_X1 U15934 ( .A1(n13942), .A2(n13941), .A3(n13940), .ZN(n13943) );
  NAND3_X1 U15935 ( .A1(n14628), .A2(n13958), .A3(n13943), .ZN(n13946) );
  AOI21_X1 U15936 ( .B1(n14596), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n13944), .ZN(
        n13945) );
  NAND4_X1 U15937 ( .A1(n13948), .A2(n13947), .A3(n13946), .A4(n13945), .ZN(
        P1_U3250) );
  OAI21_X1 U15938 ( .B1(n14637), .B2(n13950), .A(n13949), .ZN(n13951) );
  AOI21_X1 U15939 ( .B1(n13955), .B2(n14634), .A(n13951), .ZN(n13962) );
  NOR2_X1 U15940 ( .A1(n13953), .A2(n13952), .ZN(n13954) );
  OAI21_X1 U15941 ( .B1(n13954), .B2(n13969), .A(n14600), .ZN(n13961) );
  MUX2_X1 U15942 ( .A(n11144), .B(P1_REG2_REG_8__SCAN_IN), .S(n13955), .Z(
        n13956) );
  NAND3_X1 U15943 ( .A1(n13958), .A2(n13957), .A3(n13956), .ZN(n13959) );
  NAND3_X1 U15944 ( .A1(n14628), .A2(n13975), .A3(n13959), .ZN(n13960) );
  NAND3_X1 U15945 ( .A1(n13962), .A2(n13961), .A3(n13960), .ZN(P1_U3251) );
  NOR2_X1 U15946 ( .A1(n14618), .A2(n13963), .ZN(n13964) );
  AOI211_X1 U15947 ( .C1(n14596), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n13965), .B(
        n13964), .ZN(n13980) );
  INV_X1 U15948 ( .A(n13966), .ZN(n13971) );
  NOR3_X1 U15949 ( .A1(n13969), .A2(n13968), .A3(n13967), .ZN(n13970) );
  OAI21_X1 U15950 ( .B1(n13971), .B2(n13970), .A(n14600), .ZN(n13979) );
  MUX2_X1 U15951 ( .A(n10211), .B(P1_REG2_REG_9__SCAN_IN), .S(n13972), .Z(
        n13973) );
  NAND3_X1 U15952 ( .A1(n13975), .A2(n13974), .A3(n13973), .ZN(n13976) );
  NAND3_X1 U15953 ( .A1(n14628), .A2(n13977), .A3(n13976), .ZN(n13978) );
  NAND3_X1 U15954 ( .A1(n13980), .A2(n13979), .A3(n13978), .ZN(P1_U3252) );
  OAI21_X1 U15955 ( .B1(n13983), .B2(n13982), .A(n13981), .ZN(n13984) );
  NAND2_X1 U15956 ( .A1(n13984), .A2(n14600), .ZN(n13996) );
  OAI21_X1 U15957 ( .B1(n14637), .B2(n13986), .A(n13985), .ZN(n13987) );
  AOI21_X1 U15958 ( .B1(n14634), .B2(n13988), .A(n13987), .ZN(n13995) );
  MUX2_X1 U15959 ( .A(n10308), .B(P1_REG2_REG_11__SCAN_IN), .S(n13988), .Z(
        n13989) );
  NAND3_X1 U15960 ( .A1(n13991), .A2(n13990), .A3(n13989), .ZN(n13992) );
  NAND3_X1 U15961 ( .A1(n14628), .A2(n13993), .A3(n13992), .ZN(n13994) );
  NAND3_X1 U15962 ( .A1(n13996), .A2(n13995), .A3(n13994), .ZN(P1_U3254) );
  OAI21_X1 U15963 ( .B1(n11224), .B2(n13998), .A(n13997), .ZN(n14000) );
  INV_X1 U15964 ( .A(n14000), .ZN(n13999) );
  XNOR2_X1 U15965 ( .A(n14633), .B(n13999), .ZN(n14624) );
  NAND2_X1 U15966 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14624), .ZN(n14623) );
  NAND2_X1 U15967 ( .A1(n14633), .A2(n14000), .ZN(n14001) );
  NAND2_X1 U15968 ( .A1(n14623), .A2(n14001), .ZN(n14002) );
  XOR2_X1 U15969 ( .A(n14002), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14013) );
  NAND2_X1 U15970 ( .A1(n14003), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14005) );
  NAND2_X1 U15971 ( .A1(n14005), .A2(n14004), .ZN(n14006) );
  XOR2_X1 U15972 ( .A(n14633), .B(n14006), .Z(n14629) );
  NAND2_X1 U15973 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14629), .ZN(n14627) );
  NAND2_X1 U15974 ( .A1(n14633), .A2(n14006), .ZN(n14007) );
  NAND2_X1 U15975 ( .A1(n14627), .A2(n14007), .ZN(n14008) );
  INV_X1 U15976 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14172) );
  XOR2_X1 U15977 ( .A(n14008), .B(n14172), .Z(n14011) );
  NAND2_X1 U15978 ( .A1(n14011), .A2(n14628), .ZN(n14009) );
  OAI211_X1 U15979 ( .C1(n14013), .C2(n14626), .A(n14009), .B(n14618), .ZN(
        n14010) );
  INV_X1 U15980 ( .A(n14010), .ZN(n14015) );
  INV_X1 U15981 ( .A(n14011), .ZN(n14012) );
  AOI22_X1 U15982 ( .A1(n14013), .A2(n14600), .B1(n14628), .B2(n14012), .ZN(
        n14014) );
  MUX2_X1 U15983 ( .A(n14015), .B(n14014), .S(n6857), .Z(n14017) );
  OAI211_X1 U15984 ( .C1(n14018), .C2(n14637), .A(n14017), .B(n14016), .ZN(
        P1_U3262) );
  NAND2_X1 U15985 ( .A1(n14333), .A2(n14027), .ZN(n14020) );
  XOR2_X1 U15986 ( .A(n14020), .B(n14019), .Z(n14261) );
  NAND2_X1 U15987 ( .A1(n14261), .A2(n14244), .ZN(n14026) );
  INV_X1 U15988 ( .A(n14021), .ZN(n14022) );
  NOR2_X1 U15989 ( .A1(n14023), .A2(n14022), .ZN(n14264) );
  INV_X1 U15990 ( .A(n14264), .ZN(n14024) );
  NOR2_X1 U15991 ( .A1(n14147), .A2(n14024), .ZN(n14029) );
  AOI21_X1 U15992 ( .B1(n14147), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14029), 
        .ZN(n14025) );
  OAI211_X1 U15993 ( .C1(n14329), .C2(n14196), .A(n14026), .B(n14025), .ZN(
        P1_U3263) );
  XNOR2_X1 U15994 ( .A(n14333), .B(n14027), .ZN(n14028) );
  NAND2_X1 U15995 ( .A1(n14265), .A2(n14124), .ZN(n14031) );
  AOI21_X1 U15996 ( .B1(n14147), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14029), 
        .ZN(n14030) );
  OAI211_X1 U15997 ( .C1(n14333), .C2(n14196), .A(n14031), .B(n14030), .ZN(
        P1_U3264) );
  AOI22_X1 U15998 ( .A1(n14147), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14243), 
        .B2(n14032), .ZN(n14035) );
  NAND2_X1 U15999 ( .A1(n14033), .A2(n14246), .ZN(n14034) );
  OAI211_X1 U16000 ( .C1(n14036), .C2(n14239), .A(n14035), .B(n14034), .ZN(
        n14037) );
  INV_X1 U16001 ( .A(n14037), .ZN(n14038) );
  OAI21_X1 U16002 ( .B1(n14039), .B2(n14147), .A(n14038), .ZN(P1_U3266) );
  XNOR2_X1 U16003 ( .A(n14041), .B(n14040), .ZN(n14274) );
  NAND2_X1 U16004 ( .A1(n14063), .A2(n14042), .ZN(n14044) );
  XNOR2_X1 U16005 ( .A(n14044), .B(n14043), .ZN(n14272) );
  NAND2_X1 U16006 ( .A1(n14046), .A2(n14045), .ZN(n14047) );
  NAND2_X1 U16007 ( .A1(n14047), .A2(n14302), .ZN(n14048) );
  NOR2_X1 U16008 ( .A1(n14049), .A2(n14048), .ZN(n14271) );
  NAND2_X1 U16009 ( .A1(n14271), .A2(n14124), .ZN(n14054) );
  INV_X1 U16010 ( .A(n14050), .ZN(n14051) );
  OAI22_X1 U16011 ( .A1(n14147), .A2(n14268), .B1(n14051), .B2(n14206), .ZN(
        n14052) );
  AOI21_X1 U16012 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n14147), .A(n14052), 
        .ZN(n14053) );
  OAI211_X1 U16013 ( .C1(n14269), .C2(n14196), .A(n14054), .B(n14053), .ZN(
        n14055) );
  AOI21_X1 U16014 ( .B1(n14272), .B2(n14180), .A(n14055), .ZN(n14056) );
  OAI21_X1 U16015 ( .B1(n14274), .B2(n14219), .A(n14056), .ZN(P1_U3267) );
  XNOR2_X1 U16016 ( .A(n14058), .B(n14086), .ZN(n14059) );
  NAND2_X1 U16017 ( .A1(n14061), .A2(n14060), .ZN(n14062) );
  NAND2_X1 U16018 ( .A1(n14063), .A2(n14062), .ZN(n14064) );
  NAND2_X1 U16019 ( .A1(n14064), .A2(n14676), .ZN(n14280) );
  OAI211_X1 U16020 ( .C1(n14106), .C2(n14276), .A(n14280), .B(n14275), .ZN(
        n14073) );
  NAND2_X1 U16021 ( .A1(n14066), .A2(n14065), .ZN(n14067) );
  AND2_X1 U16022 ( .A1(n14068), .A2(n14067), .ZN(n14278) );
  NAND2_X1 U16023 ( .A1(n14278), .A2(n14256), .ZN(n14071) );
  AOI22_X1 U16024 ( .A1(n14147), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n14069), 
        .B2(n14243), .ZN(n14070) );
  OAI211_X1 U16025 ( .C1(n8653), .C2(n14196), .A(n14071), .B(n14070), .ZN(
        n14072) );
  AOI21_X1 U16026 ( .B1(n14073), .B2(n14253), .A(n14072), .ZN(n14074) );
  INV_X1 U16027 ( .A(n14074), .ZN(P1_U3268) );
  INV_X1 U16028 ( .A(n14075), .ZN(n14076) );
  AOI21_X1 U16029 ( .B1(n14081), .B2(n14077), .A(n14076), .ZN(n14085) );
  AOI22_X1 U16030 ( .A1(n14498), .A2(n14079), .B1(n14078), .B2(n14642), .ZN(
        n14084) );
  OAI211_X1 U16031 ( .C1(n14082), .C2(n14081), .A(n14080), .B(n14676), .ZN(
        n14083) );
  OAI211_X1 U16032 ( .C1(n14085), .C2(n14672), .A(n14084), .B(n14083), .ZN(
        n14284) );
  INV_X1 U16033 ( .A(n14284), .ZN(n14092) );
  AOI211_X1 U16034 ( .C1(n14087), .C2(n14095), .A(n14644), .B(n14057), .ZN(
        n14283) );
  AOI22_X1 U16035 ( .A1(n14147), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14088), 
        .B2(n14243), .ZN(n14089) );
  OAI21_X1 U16036 ( .B1(n14341), .B2(n14196), .A(n14089), .ZN(n14090) );
  AOI21_X1 U16037 ( .B1(n14283), .B2(n14124), .A(n14090), .ZN(n14091) );
  OAI21_X1 U16038 ( .B1(n14092), .B2(n14147), .A(n14091), .ZN(P1_U3269) );
  INV_X1 U16039 ( .A(n14122), .ZN(n14093) );
  AOI21_X1 U16040 ( .B1(n14093), .B2(n14289), .A(n14644), .ZN(n14094) );
  NAND2_X1 U16041 ( .A1(n14095), .A2(n14094), .ZN(n14291) );
  XNOR2_X1 U16042 ( .A(n14096), .B(n14099), .ZN(n14104) );
  INV_X1 U16043 ( .A(n14097), .ZN(n14098) );
  NAND2_X1 U16044 ( .A1(n14119), .A2(n14098), .ZN(n14100) );
  NAND2_X1 U16045 ( .A1(n14100), .A2(n14099), .ZN(n14101) );
  AND3_X1 U16046 ( .A1(n14102), .A2(n14684), .A3(n14101), .ZN(n14103) );
  AOI21_X1 U16047 ( .B1(n14104), .B2(n14676), .A(n14103), .ZN(n14293) );
  OAI211_X1 U16048 ( .C1(n14106), .C2(n14291), .A(n14293), .B(n14105), .ZN(
        n14107) );
  NAND2_X1 U16049 ( .A1(n14107), .A2(n14253), .ZN(n14114) );
  INV_X1 U16050 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14110) );
  INV_X1 U16051 ( .A(n14108), .ZN(n14109) );
  OAI22_X1 U16052 ( .A1(n14253), .A2(n14110), .B1(n14109), .B2(n14206), .ZN(
        n14111) );
  AOI21_X1 U16053 ( .B1(n14245), .B2(n14112), .A(n14111), .ZN(n14113) );
  OAI211_X1 U16054 ( .C1(n14115), .C2(n14196), .A(n14114), .B(n14113), .ZN(
        P1_U3270) );
  INV_X1 U16055 ( .A(n14116), .ZN(n14117) );
  AOI21_X1 U16056 ( .B1(n14120), .B2(n14118), .A(n14117), .ZN(n14300) );
  OAI21_X1 U16057 ( .B1(n14121), .B2(n14120), .A(n14119), .ZN(n14298) );
  AOI211_X1 U16058 ( .C1(n14123), .C2(n14137), .A(n14644), .B(n14122), .ZN(
        n14297) );
  NAND2_X1 U16059 ( .A1(n14297), .A2(n14124), .ZN(n14128) );
  OAI22_X1 U16060 ( .A1(n14294), .A2(n14147), .B1(n14125), .B2(n14206), .ZN(
        n14126) );
  AOI21_X1 U16061 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n14147), .A(n14126), 
        .ZN(n14127) );
  OAI211_X1 U16062 ( .C1(n14196), .C2(n14295), .A(n14128), .B(n14127), .ZN(
        n14129) );
  AOI21_X1 U16063 ( .B1(n14298), .B2(n14256), .A(n14129), .ZN(n14130) );
  OAI21_X1 U16064 ( .B1(n14300), .B2(n14131), .A(n14130), .ZN(P1_U3271) );
  OAI211_X1 U16065 ( .C1(n14133), .C2(n14144), .A(n14132), .B(n14676), .ZN(
        n14136) );
  AOI22_X1 U16066 ( .A1(n14134), .A2(n14642), .B1(n14498), .B2(n14317), .ZN(
        n14135) );
  AND2_X1 U16067 ( .A1(n14136), .A2(n14135), .ZN(n14305) );
  INV_X1 U16068 ( .A(n14137), .ZN(n14138) );
  AOI21_X1 U16069 ( .B1(n14301), .B2(n14156), .A(n14138), .ZN(n14303) );
  NOR2_X1 U16070 ( .A1(n6960), .A2(n14196), .ZN(n14142) );
  INV_X1 U16071 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14140) );
  OAI22_X1 U16072 ( .A1(n14253), .A2(n14140), .B1(n14139), .B2(n14206), .ZN(
        n14141) );
  AOI211_X1 U16073 ( .C1(n14303), .C2(n14244), .A(n14142), .B(n14141), .ZN(
        n14146) );
  XOR2_X1 U16074 ( .A(n14143), .B(n14144), .Z(n14306) );
  OR2_X1 U16075 ( .A1(n14306), .A2(n14219), .ZN(n14145) );
  OAI211_X1 U16076 ( .C1(n14305), .C2(n14147), .A(n14146), .B(n14145), .ZN(
        P1_U3272) );
  OAI211_X1 U16077 ( .C1(n14150), .C2(n14149), .A(n14676), .B(n14148), .ZN(
        n14313) );
  AOI22_X1 U16078 ( .A1(n14147), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14151), 
        .B2(n14243), .ZN(n14154) );
  NAND2_X1 U16079 ( .A1(n14152), .A2(n14245), .ZN(n14153) );
  OAI211_X1 U16080 ( .C1(n14155), .C2(n14210), .A(n14154), .B(n14153), .ZN(
        n14159) );
  AOI21_X1 U16081 ( .B1(n14160), .B2(n14170), .A(n14644), .ZN(n14157) );
  NAND2_X1 U16082 ( .A1(n14157), .A2(n14156), .ZN(n14309) );
  NOR2_X1 U16083 ( .A1(n14309), .A2(n14239), .ZN(n14158) );
  AOI211_X1 U16084 ( .C1(n14246), .C2(n14160), .A(n14159), .B(n14158), .ZN(
        n14166) );
  OR2_X1 U16085 ( .A1(n14162), .A2(n14161), .ZN(n14163) );
  NAND2_X1 U16086 ( .A1(n14164), .A2(n14163), .ZN(n14310) );
  OR2_X1 U16087 ( .A1(n14310), .A2(n14219), .ZN(n14165) );
  OAI211_X1 U16088 ( .C1(n14313), .C2(n14147), .A(n14166), .B(n14165), .ZN(
        P1_U3273) );
  XOR2_X1 U16089 ( .A(n14167), .B(n14168), .Z(n14324) );
  OAI21_X1 U16090 ( .B1(n6627), .B2(n7071), .A(n7070), .ZN(n14322) );
  OAI211_X1 U16091 ( .C1(n14185), .C2(n14320), .A(n14302), .B(n14170), .ZN(
        n14319) );
  OAI22_X1 U16092 ( .A1(n14253), .A2(n14172), .B1(n14171), .B2(n14206), .ZN(
        n14173) );
  AOI21_X1 U16093 ( .B1(n14245), .B2(n14317), .A(n14173), .ZN(n14174) );
  OAI21_X1 U16094 ( .B1(n14175), .B2(n14210), .A(n14174), .ZN(n14176) );
  AOI21_X1 U16095 ( .B1(n8544), .B2(n14246), .A(n14176), .ZN(n14177) );
  OAI21_X1 U16096 ( .B1(n14319), .B2(n14178), .A(n14177), .ZN(n14179) );
  AOI21_X1 U16097 ( .B1(n14322), .B2(n14180), .A(n14179), .ZN(n14181) );
  OAI21_X1 U16098 ( .B1(n14324), .B2(n14219), .A(n14181), .ZN(P1_U3274) );
  NAND2_X1 U16099 ( .A1(n14205), .A2(n14182), .ZN(n14183) );
  NAND2_X1 U16100 ( .A1(n14183), .A2(n14302), .ZN(n14184) );
  OR2_X1 U16101 ( .A1(n14185), .A2(n14184), .ZN(n14480) );
  XNOR2_X1 U16102 ( .A(n14187), .B(n14186), .ZN(n14192) );
  OAI211_X1 U16103 ( .C1(n14190), .C2(n14189), .A(n14188), .B(n14676), .ZN(
        n14191) );
  OAI21_X1 U16104 ( .B1(n14192), .B2(n14672), .A(n14191), .ZN(n14483) );
  OAI21_X1 U16105 ( .B1(n14483), .B2(n14193), .A(n14253), .ZN(n14201) );
  OAI22_X1 U16106 ( .A1(n14253), .A2(n14195), .B1(n14194), .B2(n14206), .ZN(
        n14198) );
  NOR2_X1 U16107 ( .A1(n14481), .A2(n14196), .ZN(n14197) );
  AOI211_X1 U16108 ( .C1(n14245), .C2(n14199), .A(n14198), .B(n14197), .ZN(
        n14200) );
  OAI211_X1 U16109 ( .C1(n14239), .C2(n14480), .A(n14201), .B(n14200), .ZN(
        P1_U3275) );
  XNOR2_X1 U16110 ( .A(n14202), .B(n14204), .ZN(n14491) );
  INV_X1 U16111 ( .A(n14491), .ZN(n14218) );
  AOI211_X1 U16112 ( .C1(n14204), .C2(n14203), .A(n14661), .B(n6630), .ZN(
        n14489) );
  OAI211_X1 U16113 ( .C1(n14221), .C2(n14488), .A(n14205), .B(n14302), .ZN(
        n14487) );
  OAI22_X1 U16114 ( .A1(n14253), .A2(n14208), .B1(n14207), .B2(n14206), .ZN(
        n14212) );
  NOR2_X1 U16115 ( .A1(n14210), .A2(n14209), .ZN(n14211) );
  AOI211_X1 U16116 ( .C1(n14245), .C2(n14485), .A(n14212), .B(n14211), .ZN(
        n14215) );
  NAND2_X1 U16117 ( .A1(n14213), .A2(n14246), .ZN(n14214) );
  OAI211_X1 U16118 ( .C1(n14487), .C2(n14239), .A(n14215), .B(n14214), .ZN(
        n14216) );
  AOI21_X1 U16119 ( .B1(n14489), .B2(n14253), .A(n14216), .ZN(n14217) );
  OAI21_X1 U16120 ( .B1(n14219), .B2(n14218), .A(n14217), .ZN(P1_U3276) );
  INV_X1 U16121 ( .A(n14220), .ZN(n14223) );
  INV_X1 U16122 ( .A(n14221), .ZN(n14222) );
  OAI211_X1 U16123 ( .C1(n14494), .C2(n14223), .A(n14222), .B(n14302), .ZN(
        n14493) );
  XNOR2_X1 U16124 ( .A(n14224), .B(n14227), .ZN(n14229) );
  OAI21_X1 U16125 ( .B1(n14227), .B2(n14226), .A(n14225), .ZN(n14228) );
  AOI22_X1 U16126 ( .A1(n14229), .A2(n14676), .B1(n14228), .B2(n14684), .ZN(
        n14230) );
  INV_X1 U16127 ( .A(n14230), .ZN(n14496) );
  OAI21_X1 U16128 ( .B1(n14496), .B2(n14231), .A(n14253), .ZN(n14238) );
  INV_X1 U16129 ( .A(n14245), .ZN(n14234) );
  AOI22_X1 U16130 ( .A1(n14147), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7443), 
        .B2(n14243), .ZN(n14232) );
  OAI21_X1 U16131 ( .B1(n14234), .B2(n14233), .A(n14232), .ZN(n14235) );
  AOI21_X1 U16132 ( .B1(n14236), .B2(n14246), .A(n14235), .ZN(n14237) );
  OAI211_X1 U16133 ( .C1(n14239), .C2(n14493), .A(n14238), .B(n14237), .ZN(
        P1_U3277) );
  AND2_X1 U16134 ( .A1(n14240), .A2(n14641), .ZN(n14241) );
  NOR2_X1 U16135 ( .A1(n14242), .A2(n14241), .ZN(n14640) );
  AOI22_X1 U16136 ( .A1(n14244), .A2(n14640), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14243), .ZN(n14260) );
  AOI22_X1 U16137 ( .A1(n14246), .A2(n14641), .B1(n14245), .B2(n8319), .ZN(
        n14259) );
  INV_X1 U16138 ( .A(n11987), .ZN(n14247) );
  AOI21_X1 U16139 ( .B1(n14247), .B2(n10303), .A(n14661), .ZN(n14252) );
  XNOR2_X1 U16140 ( .A(n14640), .B(n14248), .ZN(n14250) );
  OAI21_X1 U16141 ( .B1(n14250), .B2(n14661), .A(n14249), .ZN(n14251) );
  OAI21_X1 U16142 ( .B1(n14252), .B2(n14498), .A(n14251), .ZN(n14646) );
  MUX2_X1 U16143 ( .A(n14254), .B(n14646), .S(n14253), .Z(n14258) );
  XNOR2_X1 U16144 ( .A(n11987), .B(n14255), .ZN(n14649) );
  NAND2_X1 U16145 ( .A1(n14256), .A2(n14649), .ZN(n14257) );
  NAND4_X1 U16146 ( .A1(n14260), .A2(n14259), .A3(n14258), .A4(n14257), .ZN(
        P1_U3292) );
  INV_X1 U16147 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14262) );
  AOI21_X1 U16148 ( .B1(n14261), .B2(n14302), .A(n14264), .ZN(n14326) );
  MUX2_X1 U16149 ( .A(n14262), .B(n14326), .S(n14698), .Z(n14263) );
  OAI21_X1 U16150 ( .B1(n14329), .B2(n14316), .A(n14263), .ZN(P1_U3559) );
  INV_X1 U16151 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14266) );
  NOR2_X1 U16152 ( .A1(n14265), .A2(n14264), .ZN(n14330) );
  MUX2_X1 U16153 ( .A(n14266), .B(n14330), .S(n14698), .Z(n14267) );
  OAI21_X1 U16154 ( .B1(n14333), .B2(n14316), .A(n14267), .ZN(P1_U3558) );
  OAI21_X1 U16155 ( .B1(n14269), .B2(n14680), .A(n14268), .ZN(n14270) );
  AOI211_X1 U16156 ( .C1(n14272), .C2(n14676), .A(n14271), .B(n14270), .ZN(
        n14273) );
  OAI21_X1 U16157 ( .B1(n14274), .B2(n14672), .A(n14273), .ZN(n14334) );
  MUX2_X1 U16158 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14334), .S(n14698), .Z(
        P1_U3554) );
  NAND2_X1 U16159 ( .A1(n14276), .A2(n14275), .ZN(n14277) );
  AOI21_X1 U16160 ( .B1(n14278), .B2(n14684), .A(n14277), .ZN(n14279) );
  NAND2_X1 U16161 ( .A1(n14280), .A2(n14279), .ZN(n14335) );
  MUX2_X1 U16162 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14335), .S(n14698), .Z(
        n14281) );
  INV_X1 U16163 ( .A(n14281), .ZN(n14282) );
  OAI21_X1 U16164 ( .B1(n8653), .B2(n14316), .A(n14282), .ZN(P1_U3553) );
  INV_X1 U16165 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14285) );
  NOR2_X1 U16166 ( .A1(n14284), .A2(n14283), .ZN(n14338) );
  MUX2_X1 U16167 ( .A(n14285), .B(n14338), .S(n14698), .Z(n14286) );
  OAI21_X1 U16168 ( .B1(n14341), .B2(n14316), .A(n14286), .ZN(P1_U3552) );
  INV_X1 U16169 ( .A(n14287), .ZN(n14288) );
  AOI21_X1 U16170 ( .B1(n14289), .B2(n14669), .A(n14288), .ZN(n14290) );
  AND2_X1 U16171 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  NAND2_X1 U16172 ( .A1(n14293), .A2(n14292), .ZN(n14342) );
  MUX2_X1 U16173 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14342), .S(n14698), .Z(
        P1_U3551) );
  OAI21_X1 U16174 ( .B1(n14295), .B2(n14680), .A(n14294), .ZN(n14296) );
  AOI211_X1 U16175 ( .C1(n14298), .C2(n14684), .A(n14297), .B(n14296), .ZN(
        n14299) );
  OAI21_X1 U16176 ( .B1(n14300), .B2(n14661), .A(n14299), .ZN(n14343) );
  MUX2_X1 U16177 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14343), .S(n14698), .Z(
        P1_U3550) );
  AOI22_X1 U16178 ( .A1(n14303), .A2(n14302), .B1(n14669), .B2(n14301), .ZN(
        n14304) );
  OAI211_X1 U16179 ( .C1(n14306), .C2(n14672), .A(n14305), .B(n14304), .ZN(
        n14344) );
  MUX2_X1 U16180 ( .A(n14344), .B(P1_REG1_REG_21__SCAN_IN), .S(n14695), .Z(
        P1_U3549) );
  INV_X1 U16181 ( .A(n14307), .ZN(n14308) );
  AND2_X1 U16182 ( .A1(n14309), .A2(n14308), .ZN(n14312) );
  OR2_X1 U16183 ( .A1(n14310), .A2(n14672), .ZN(n14311) );
  MUX2_X1 U16184 ( .A(n14314), .B(n14345), .S(n14698), .Z(n14315) );
  OAI21_X1 U16185 ( .B1(n14349), .B2(n14316), .A(n14315), .ZN(P1_U3548) );
  AOI22_X1 U16186 ( .A1(n14317), .A2(n14642), .B1(n14498), .B2(n14485), .ZN(
        n14318) );
  OAI211_X1 U16187 ( .C1(n14320), .C2(n14680), .A(n14319), .B(n14318), .ZN(
        n14321) );
  AOI21_X1 U16188 ( .B1(n14322), .B2(n14676), .A(n14321), .ZN(n14323) );
  OAI21_X1 U16189 ( .B1(n14324), .B2(n14672), .A(n14323), .ZN(n14350) );
  MUX2_X1 U16190 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14350), .S(n14698), .Z(
        P1_U3547) );
  MUX2_X1 U16191 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14325), .S(n14698), .Z(
        P1_U3528) );
  INV_X1 U16192 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14327) );
  MUX2_X1 U16193 ( .A(n14327), .B(n14326), .S(n14687), .Z(n14328) );
  OAI21_X1 U16194 ( .B1(n14329), .B2(n14348), .A(n14328), .ZN(P1_U3527) );
  INV_X1 U16195 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14331) );
  MUX2_X1 U16196 ( .A(n14331), .B(n14330), .S(n14687), .Z(n14332) );
  OAI21_X1 U16197 ( .B1(n14333), .B2(n14348), .A(n14332), .ZN(P1_U3526) );
  MUX2_X1 U16198 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14334), .S(n14687), .Z(
        P1_U3522) );
  MUX2_X1 U16199 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14335), .S(n14687), .Z(
        n14336) );
  INV_X1 U16200 ( .A(n14336), .ZN(n14337) );
  OAI21_X1 U16201 ( .B1(n8653), .B2(n14348), .A(n14337), .ZN(P1_U3521) );
  INV_X1 U16202 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14339) );
  MUX2_X1 U16203 ( .A(n14339), .B(n14338), .S(n14687), .Z(n14340) );
  OAI21_X1 U16204 ( .B1(n14341), .B2(n14348), .A(n14340), .ZN(P1_U3520) );
  MUX2_X1 U16205 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14342), .S(n14687), .Z(
        P1_U3519) );
  MUX2_X1 U16206 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14343), .S(n14687), .Z(
        P1_U3518) );
  MUX2_X1 U16207 ( .A(n14344), .B(P1_REG0_REG_21__SCAN_IN), .S(n14685), .Z(
        P1_U3517) );
  INV_X1 U16208 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14346) );
  MUX2_X1 U16209 ( .A(n14346), .B(n14345), .S(n14687), .Z(n14347) );
  OAI21_X1 U16210 ( .B1(n14349), .B2(n14348), .A(n14347), .ZN(P1_U3516) );
  MUX2_X1 U16211 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14350), .S(n14687), .Z(
        P1_U3515) );
  NOR4_X1 U16212 ( .A1(n14352), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14351), .ZN(n14353) );
  AOI21_X1 U16213 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14354), .A(n14353), 
        .ZN(n14355) );
  OAI21_X1 U16214 ( .B1(n14356), .B2(n14366), .A(n14355), .ZN(P1_U3324) );
  INV_X1 U16215 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14357) );
  OAI222_X1 U16216 ( .A1(P1_U3086), .A2(n14359), .B1(n14366), .B2(n14358), 
        .C1(n14357), .C2(n14363), .ZN(P1_U3326) );
  OAI222_X1 U16217 ( .A1(P1_U3086), .A2(n14362), .B1(n14366), .B2(n14361), 
        .C1(n14360), .C2(n14363), .ZN(P1_U3328) );
  OAI222_X1 U16218 ( .A1(n14367), .A2(P1_U3086), .B1(n14366), .B2(n14365), 
        .C1(n14364), .C2(n14363), .ZN(P1_U3329) );
  MUX2_X1 U16219 ( .A(n6858), .B(n14368), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16220 ( .A(n14369), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U16221 ( .B1(n14372), .B2(n14371), .A(n14370), .ZN(n14373) );
  XNOR2_X1 U16222 ( .A(n14373), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16223 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14374) );
  OAI21_X1 U16224 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14374), 
        .ZN(U28) );
  OAI221_X1 U16225 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n7507), .C2(n7506), .A(n14375), .ZN(U29) );
  OAI21_X1 U16226 ( .B1(n14378), .B2(n14377), .A(n14376), .ZN(n14379) );
  XNOR2_X1 U16227 ( .A(n14379), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI22_X1 U16228 ( .A1(n14382), .A2(n14381), .B1(SI_11_), .B2(n14380), .ZN(
        n14383) );
  OAI21_X1 U16229 ( .B1(P3_U3151), .B2(n15036), .A(n14383), .ZN(P3_U3284) );
  AOI21_X1 U16230 ( .B1(n14386), .B2(n14385), .A(n14384), .ZN(SUB_1596_U57) );
  OAI21_X1 U16231 ( .B1(n14389), .B2(n14388), .A(n14387), .ZN(SUB_1596_U55) );
  AOI21_X1 U16232 ( .B1(n14392), .B2(n14391), .A(n14390), .ZN(SUB_1596_U54) );
  AOI21_X1 U16233 ( .B1(n14395), .B2(n14394), .A(n14393), .ZN(SUB_1596_U70) );
  AOI21_X1 U16234 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n14399) );
  XOR2_X1 U16235 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14399), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16236 ( .B1(n14402), .B2(n14401), .A(n14400), .ZN(n14417) );
  OAI21_X1 U16237 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14404), .A(n14403), 
        .ZN(n14410) );
  NOR2_X1 U16238 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14405), .ZN(n14406) );
  AOI21_X1 U16239 ( .B1(n15089), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14406), 
        .ZN(n14407) );
  OAI21_X1 U16240 ( .B1(n15092), .B2(n14408), .A(n14407), .ZN(n14409) );
  AOI21_X1 U16241 ( .B1(n14410), .B2(n15094), .A(n14409), .ZN(n14416) );
  NOR2_X1 U16242 ( .A1(n14412), .A2(n14411), .ZN(n14413) );
  OAI21_X1 U16243 ( .B1(n14414), .B2(n14413), .A(n15096), .ZN(n14415) );
  OAI211_X1 U16244 ( .C1(n14417), .C2(n15102), .A(n14416), .B(n14415), .ZN(
        P3_U3197) );
  AOI22_X1 U16245 ( .A1(n15002), .A2(n14418), .B1(n15089), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14432) );
  NAND2_X1 U16246 ( .A1(n14419), .A2(n6647), .ZN(n14420) );
  XNOR2_X1 U16247 ( .A(n14421), .B(n14420), .ZN(n14426) );
  OAI21_X1 U16248 ( .B1(n14424), .B2(n14423), .A(n14422), .ZN(n14425) );
  AOI22_X1 U16249 ( .A1(n14426), .A2(n15096), .B1(n15094), .B2(n14425), .ZN(
        n14431) );
  NAND2_X1 U16250 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14430)
         );
  OAI221_X1 U16251 ( .B1(n14428), .B2(n6570), .C1(n14428), .C2(n14427), .A(
        n14441), .ZN(n14429) );
  NAND4_X1 U16252 ( .A1(n14432), .A2(n14431), .A3(n14430), .A4(n14429), .ZN(
        P3_U3198) );
  AOI22_X1 U16253 ( .A1(n15002), .A2(n14433), .B1(n15089), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14448) );
  OAI21_X1 U16254 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14435), .A(n14434), 
        .ZN(n14440) );
  AOI211_X1 U16255 ( .C1(n14438), .C2(n14437), .A(n14436), .B(n15076), .ZN(
        n14439) );
  AOI21_X1 U16256 ( .B1(n15094), .B2(n14440), .A(n14439), .ZN(n14447) );
  NAND2_X1 U16257 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14446)
         );
  OAI221_X1 U16258 ( .B1(n14444), .B2(n14443), .C1(n14444), .C2(n14442), .A(
        n14441), .ZN(n14445) );
  NAND4_X1 U16259 ( .A1(n14448), .A2(n14447), .A3(n14446), .A4(n14445), .ZN(
        P3_U3199) );
  NAND2_X1 U16260 ( .A1(n14449), .A2(n15190), .ZN(n14452) );
  OR2_X1 U16261 ( .A1(n14450), .A2(n15185), .ZN(n14451) );
  AOI22_X1 U16262 ( .A1(n15205), .A2(n14455), .B1(n9077), .B2(n15203), .ZN(
        P3_U3472) );
  INV_X1 U16263 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U16264 ( .A1(n15193), .A2(n14455), .B1(n14454), .B2(n15191), .ZN(
        P3_U3429) );
  OAI22_X1 U16265 ( .A1(n14459), .A2(n14458), .B1(n14457), .B2(n14456), .ZN(
        n14466) );
  NAND2_X1 U16266 ( .A1(n14461), .A2(n14460), .ZN(n14463) );
  AOI21_X1 U16267 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(n14465) );
  AOI211_X1 U16268 ( .C1(n14937), .C2(n14467), .A(n14466), .B(n14465), .ZN(
        n14468) );
  NAND2_X1 U16269 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14794)
         );
  OAI211_X1 U16270 ( .C1(n14470), .C2(n14469), .A(n14468), .B(n14794), .ZN(
        P2_U3208) );
  AND2_X1 U16271 ( .A1(n14471), .A2(n14934), .ZN(n14476) );
  OAI21_X1 U16272 ( .B1(n14473), .B2(n14927), .A(n14472), .ZN(n14474) );
  NOR3_X1 U16273 ( .A1(n14476), .A2(n14475), .A3(n14474), .ZN(n14478) );
  AOI22_X1 U16274 ( .A1(n14960), .A2(n14478), .B1(n13198), .B2(n14957), .ZN(
        P2_U3511) );
  INV_X1 U16275 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U16276 ( .A1(n14944), .A2(n14478), .B1(n14477), .B2(n14942), .ZN(
        P2_U3466) );
  OAI211_X1 U16277 ( .C1(n14481), .C2(n14680), .A(n14480), .B(n14479), .ZN(
        n14482) );
  NOR2_X1 U16278 ( .A1(n14483), .A2(n14482), .ZN(n14537) );
  INV_X1 U16279 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14484) );
  AOI22_X1 U16280 ( .A1(n14698), .A2(n14537), .B1(n14484), .B2(n14695), .ZN(
        P1_U3546) );
  AOI22_X1 U16281 ( .A1(n14485), .A2(n14642), .B1(n14498), .B2(n14500), .ZN(
        n14486) );
  OAI211_X1 U16282 ( .C1(n14488), .C2(n14680), .A(n14487), .B(n14486), .ZN(
        n14490) );
  AOI211_X1 U16283 ( .C1(n14491), .C2(n14684), .A(n14490), .B(n14489), .ZN(
        n14539) );
  AOI22_X1 U16284 ( .A1(n14698), .A2(n14539), .B1(n11224), .B2(n14695), .ZN(
        P1_U3545) );
  OAI211_X1 U16285 ( .C1(n14494), .C2(n14680), .A(n14493), .B(n14492), .ZN(
        n14495) );
  NOR2_X1 U16286 ( .A1(n14496), .A2(n14495), .ZN(n14541) );
  AOI22_X1 U16287 ( .A1(n14698), .A2(n14541), .B1(n14497), .B2(n14695), .ZN(
        P1_U3544) );
  AOI22_X1 U16288 ( .A1(n14642), .A2(n14500), .B1(n14499), .B2(n14498), .ZN(
        n14501) );
  OAI211_X1 U16289 ( .C1(n14503), .C2(n14680), .A(n14502), .B(n14501), .ZN(
        n14507) );
  AND3_X1 U16290 ( .A1(n14505), .A2(n14676), .A3(n14504), .ZN(n14506) );
  AOI211_X1 U16291 ( .C1(n14684), .C2(n14508), .A(n14507), .B(n14506), .ZN(
        n14543) );
  INV_X1 U16292 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14509) );
  AOI22_X1 U16293 ( .A1(n14698), .A2(n14543), .B1(n14509), .B2(n14695), .ZN(
        P1_U3543) );
  OAI22_X1 U16294 ( .A1(n14511), .A2(n14522), .B1(n14510), .B2(n14520), .ZN(
        n14512) );
  AOI21_X1 U16295 ( .B1(n14513), .B2(n14669), .A(n14512), .ZN(n14515) );
  OAI211_X1 U16296 ( .C1(n14516), .C2(n14672), .A(n14515), .B(n14514), .ZN(
        n14517) );
  AOI21_X1 U16297 ( .B1(n14676), .B2(n14518), .A(n14517), .ZN(n14545) );
  AOI22_X1 U16298 ( .A1(n14698), .A2(n14545), .B1(n14519), .B2(n14695), .ZN(
        P1_U3542) );
  OAI22_X1 U16299 ( .A1(n14523), .A2(n14522), .B1(n14521), .B2(n14520), .ZN(
        n14524) );
  AOI21_X1 U16300 ( .B1(n14525), .B2(n14669), .A(n14524), .ZN(n14527) );
  AOI22_X1 U16301 ( .A1(n14698), .A2(n14547), .B1(n14529), .B2(n14695), .ZN(
        P1_U3541) );
  OAI21_X1 U16302 ( .B1(n14531), .B2(n14680), .A(n14530), .ZN(n14533) );
  AOI211_X1 U16303 ( .C1(n14684), .C2(n14534), .A(n14533), .B(n14532), .ZN(
        n14549) );
  AOI22_X1 U16304 ( .A1(n14698), .A2(n14549), .B1(n14535), .B2(n14695), .ZN(
        P1_U3539) );
  INV_X1 U16305 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14536) );
  AOI22_X1 U16306 ( .A1(n14687), .A2(n14537), .B1(n14536), .B2(n14685), .ZN(
        P1_U3513) );
  INV_X1 U16307 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14538) );
  AOI22_X1 U16308 ( .A1(n14687), .A2(n14539), .B1(n14538), .B2(n14685), .ZN(
        P1_U3510) );
  INV_X1 U16309 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14540) );
  AOI22_X1 U16310 ( .A1(n14687), .A2(n14541), .B1(n14540), .B2(n14685), .ZN(
        P1_U3507) );
  INV_X1 U16311 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14542) );
  AOI22_X1 U16312 ( .A1(n14687), .A2(n14543), .B1(n14542), .B2(n14685), .ZN(
        P1_U3504) );
  INV_X1 U16313 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U16314 ( .A1(n14687), .A2(n14545), .B1(n14544), .B2(n14685), .ZN(
        P1_U3501) );
  INV_X1 U16315 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U16316 ( .A1(n14687), .A2(n14547), .B1(n14546), .B2(n14685), .ZN(
        P1_U3498) );
  INV_X1 U16317 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14548) );
  AOI22_X1 U16318 ( .A1(n14687), .A2(n14549), .B1(n14548), .B2(n14685), .ZN(
        P1_U3492) );
  OAI21_X1 U16319 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n14553) );
  XNOR2_X1 U16320 ( .A(n14553), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16321 ( .B1(n14556), .B2(n14555), .A(n14554), .ZN(SUB_1596_U68) );
  OAI222_X1 U16322 ( .A1(n14561), .A2(n14560), .B1(n14561), .B2(n14559), .C1(
        n14558), .C2(n14557), .ZN(SUB_1596_U67) );
  OAI222_X1 U16323 ( .A1(n14566), .A2(n14565), .B1(n14566), .B2(n14564), .C1(
        n14563), .C2(n14562), .ZN(SUB_1596_U66) );
  AOI21_X1 U16324 ( .B1(n14568), .B2(n14567), .A(n6567), .ZN(n14569) );
  XOR2_X1 U16325 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14569), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16326 ( .B1(n14572), .B2(n14571), .A(n14570), .ZN(n14573) );
  XOR2_X1 U16327 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14573), .Z(SUB_1596_U64)
         );
  INV_X1 U16328 ( .A(n14574), .ZN(n14579) );
  NAND3_X1 U16329 ( .A1(n14577), .A2(n14576), .A3(n14575), .ZN(n14578) );
  NAND3_X1 U16330 ( .A1(n14600), .A2(n14579), .A3(n14578), .ZN(n14591) );
  NAND2_X1 U16331 ( .A1(n14634), .A2(n14582), .ZN(n14590) );
  AND2_X1 U16332 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14581) );
  AOI21_X1 U16333 ( .B1(n14596), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14581), .ZN(
        n14589) );
  MUX2_X1 U16334 ( .A(n10753), .B(P1_REG2_REG_4__SCAN_IN), .S(n14582), .Z(
        n14583) );
  NAND3_X1 U16335 ( .A1(n14585), .A2(n14584), .A3(n14583), .ZN(n14586) );
  NAND3_X1 U16336 ( .A1(n14628), .A2(n14587), .A3(n14586), .ZN(n14588) );
  AND4_X1 U16337 ( .A1(n14591), .A2(n14590), .A3(n14589), .A4(n14588), .ZN(
        n14593) );
  NAND2_X1 U16338 ( .A1(n14593), .A2(n14592), .ZN(P1_U3247) );
  INV_X1 U16339 ( .A(n14594), .ZN(n14595) );
  AOI21_X1 U16340 ( .B1(n14596), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n14595), 
        .ZN(n14597) );
  OAI21_X1 U16341 ( .B1(n14618), .B2(n14598), .A(n14597), .ZN(n14599) );
  INV_X1 U16342 ( .A(n14599), .ZN(n14609) );
  OAI211_X1 U16343 ( .C1(n14603), .C2(n14602), .A(n14601), .B(n14600), .ZN(
        n14608) );
  OAI211_X1 U16344 ( .C1(n14606), .C2(n14605), .A(n14628), .B(n14604), .ZN(
        n14607) );
  NAND3_X1 U16345 ( .A1(n14609), .A2(n14608), .A3(n14607), .ZN(P1_U3256) );
  AOI21_X1 U16346 ( .B1(n14611), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14610), 
        .ZN(n14615) );
  AOI21_X1 U16347 ( .B1(n14613), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14612), 
        .ZN(n14614) );
  OAI222_X1 U16348 ( .A1(n14618), .A2(n14617), .B1(n14616), .B2(n14615), .C1(
        n14626), .C2(n14614), .ZN(n14619) );
  INV_X1 U16349 ( .A(n14619), .ZN(n14621) );
  OAI211_X1 U16350 ( .C1(n14622), .C2(n14637), .A(n14621), .B(n14620), .ZN(
        P1_U3258) );
  OAI21_X1 U16351 ( .B1(n14624), .B2(P1_REG1_REG_18__SCAN_IN), .A(n14623), 
        .ZN(n14625) );
  NOR2_X1 U16352 ( .A1(n14626), .A2(n14625), .ZN(n14632) );
  OAI211_X1 U16353 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14629), .A(n14628), 
        .B(n14627), .ZN(n14630) );
  INV_X1 U16354 ( .A(n14630), .ZN(n14631) );
  AOI211_X1 U16355 ( .C1(n14634), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        n14636) );
  OAI211_X1 U16356 ( .C1(n14638), .C2(n14637), .A(n14636), .B(n14635), .ZN(
        P1_U3261) );
  AND2_X1 U16357 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14639), .ZN(P1_U3294) );
  AND2_X1 U16358 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14639), .ZN(P1_U3295) );
  AND2_X1 U16359 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14639), .ZN(P1_U3296) );
  AND2_X1 U16360 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14639), .ZN(P1_U3297) );
  AND2_X1 U16361 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14639), .ZN(P1_U3298) );
  AND2_X1 U16362 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14639), .ZN(P1_U3299) );
  AND2_X1 U16363 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14639), .ZN(P1_U3300) );
  AND2_X1 U16364 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14639), .ZN(P1_U3301) );
  AND2_X1 U16365 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14639), .ZN(P1_U3302) );
  AND2_X1 U16366 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14639), .ZN(P1_U3303) );
  AND2_X1 U16367 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14639), .ZN(P1_U3304) );
  AND2_X1 U16368 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14639), .ZN(P1_U3305) );
  AND2_X1 U16369 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14639), .ZN(P1_U3306) );
  AND2_X1 U16370 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14639), .ZN(P1_U3307) );
  AND2_X1 U16371 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14639), .ZN(P1_U3308) );
  AND2_X1 U16372 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14639), .ZN(P1_U3309) );
  AND2_X1 U16373 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14639), .ZN(P1_U3310) );
  AND2_X1 U16374 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14639), .ZN(P1_U3311) );
  AND2_X1 U16375 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14639), .ZN(P1_U3312) );
  AND2_X1 U16376 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14639), .ZN(P1_U3313) );
  AND2_X1 U16377 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14639), .ZN(P1_U3314) );
  AND2_X1 U16378 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14639), .ZN(P1_U3315) );
  AND2_X1 U16379 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14639), .ZN(P1_U3316) );
  AND2_X1 U16380 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14639), .ZN(P1_U3317) );
  AND2_X1 U16381 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14639), .ZN(P1_U3318) );
  AND2_X1 U16382 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14639), .ZN(P1_U3319) );
  AND2_X1 U16383 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14639), .ZN(P1_U3320) );
  AND2_X1 U16384 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14639), .ZN(P1_U3321) );
  AND2_X1 U16385 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14639), .ZN(P1_U3322) );
  AND2_X1 U16386 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14639), .ZN(P1_U3323) );
  INV_X1 U16387 ( .A(n14640), .ZN(n14645) );
  AOI22_X1 U16388 ( .A1(n8319), .A2(n14642), .B1(n14669), .B2(n14641), .ZN(
        n14643) );
  OAI21_X1 U16389 ( .B1(n14645), .B2(n14644), .A(n14643), .ZN(n14648) );
  INV_X1 U16390 ( .A(n14646), .ZN(n14647) );
  AOI211_X1 U16391 ( .C1(n14684), .C2(n14649), .A(n14648), .B(n14647), .ZN(
        n14688) );
  INV_X1 U16392 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14650) );
  AOI22_X1 U16393 ( .A1(n14687), .A2(n14688), .B1(n14650), .B2(n14685), .ZN(
        P1_U3462) );
  AOI21_X1 U16394 ( .B1(n14669), .B2(n14652), .A(n14651), .ZN(n14653) );
  OAI21_X1 U16395 ( .B1(n14672), .B2(n14654), .A(n14653), .ZN(n14656) );
  NOR2_X1 U16396 ( .A1(n14656), .A2(n14655), .ZN(n14690) );
  INV_X1 U16397 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14657) );
  AOI22_X1 U16398 ( .A1(n14687), .A2(n14690), .B1(n14657), .B2(n14685), .ZN(
        P1_U3471) );
  OAI211_X1 U16399 ( .C1(n14660), .C2(n14680), .A(n14659), .B(n14658), .ZN(
        n14664) );
  NOR2_X1 U16400 ( .A1(n14662), .A2(n14661), .ZN(n14663) );
  AOI211_X1 U16401 ( .C1(n14684), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14692) );
  INV_X1 U16402 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14666) );
  AOI22_X1 U16403 ( .A1(n14687), .A2(n14692), .B1(n14666), .B2(n14685), .ZN(
        P1_U3477) );
  AOI21_X1 U16404 ( .B1(n14669), .B2(n14668), .A(n14667), .ZN(n14670) );
  OAI211_X1 U16405 ( .C1(n14673), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n14674) );
  INV_X1 U16406 ( .A(n14674), .ZN(n14694) );
  INV_X1 U16407 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14675) );
  AOI22_X1 U16408 ( .A1(n14687), .A2(n14694), .B1(n14675), .B2(n14685), .ZN(
        P1_U3483) );
  NAND2_X1 U16409 ( .A1(n14677), .A2(n14676), .ZN(n14679) );
  OAI211_X1 U16410 ( .C1(n14681), .C2(n14680), .A(n14679), .B(n14678), .ZN(
        n14682) );
  AOI21_X1 U16411 ( .B1(n14684), .B2(n14683), .A(n14682), .ZN(n14697) );
  INV_X1 U16412 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14686) );
  AOI22_X1 U16413 ( .A1(n14687), .A2(n14697), .B1(n14686), .B2(n14685), .ZN(
        P1_U3489) );
  AOI22_X1 U16414 ( .A1(n14698), .A2(n14688), .B1(n10100), .B2(n14695), .ZN(
        P1_U3529) );
  AOI22_X1 U16415 ( .A1(n14698), .A2(n14690), .B1(n14689), .B2(n14695), .ZN(
        P1_U3532) );
  AOI22_X1 U16416 ( .A1(n14698), .A2(n14692), .B1(n14691), .B2(n14695), .ZN(
        P1_U3534) );
  AOI22_X1 U16417 ( .A1(n14698), .A2(n14694), .B1(n14693), .B2(n14695), .ZN(
        P1_U3536) );
  AOI22_X1 U16418 ( .A1(n14698), .A2(n14697), .B1(n14696), .B2(n14695), .ZN(
        P1_U3538) );
  NOR2_X1 U16419 ( .A1(n14849), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16420 ( .A1(n14849), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n14823), 
        .B2(n14699), .ZN(n14710) );
  NAND2_X1 U16421 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14709) );
  OAI211_X1 U16422 ( .C1(n14702), .C2(n14701), .A(n14851), .B(n14700), .ZN(
        n14708) );
  AOI211_X1 U16423 ( .C1(n14705), .C2(n14704), .A(n14703), .B(n14805), .ZN(
        n14706) );
  INV_X1 U16424 ( .A(n14706), .ZN(n14707) );
  NAND4_X1 U16425 ( .A1(n14710), .A2(n14709), .A3(n14708), .A4(n14707), .ZN(
        P2_U3217) );
  AOI22_X1 U16426 ( .A1(n14849), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n14823), 
        .B2(n14711), .ZN(n14722) );
  OAI211_X1 U16427 ( .C1(n14714), .C2(n14713), .A(n14851), .B(n14712), .ZN(
        n14720) );
  AOI211_X1 U16428 ( .C1(n14717), .C2(n14716), .A(n14805), .B(n14715), .ZN(
        n14718) );
  INV_X1 U16429 ( .A(n14718), .ZN(n14719) );
  NAND4_X1 U16430 ( .A1(n14722), .A2(n14721), .A3(n14720), .A4(n14719), .ZN(
        P2_U3218) );
  AOI22_X1 U16431 ( .A1(n14849), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n14823), 
        .B2(n14723), .ZN(n14734) );
  NAND2_X1 U16432 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14733) );
  OAI211_X1 U16433 ( .C1(n14726), .C2(n14725), .A(n14851), .B(n14724), .ZN(
        n14732) );
  AOI211_X1 U16434 ( .C1(n14729), .C2(n14728), .A(n14805), .B(n14727), .ZN(
        n14730) );
  INV_X1 U16435 ( .A(n14730), .ZN(n14731) );
  NAND4_X1 U16436 ( .A1(n14734), .A2(n14733), .A3(n14732), .A4(n14731), .ZN(
        P2_U3219) );
  AOI22_X1 U16437 ( .A1(n14849), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(n14823), 
        .B2(n14735), .ZN(n14746) );
  OAI211_X1 U16438 ( .C1(n14738), .C2(n14737), .A(n14851), .B(n14736), .ZN(
        n14744) );
  AOI211_X1 U16439 ( .C1(n14741), .C2(n14740), .A(n14805), .B(n14739), .ZN(
        n14742) );
  INV_X1 U16440 ( .A(n14742), .ZN(n14743) );
  NAND4_X1 U16441 ( .A1(n14746), .A2(n14745), .A3(n14744), .A4(n14743), .ZN(
        P2_U3220) );
  AOI22_X1 U16442 ( .A1(n14849), .A2(P2_ADDR_REG_8__SCAN_IN), .B1(n14823), 
        .B2(n14747), .ZN(n14758) );
  NAND2_X1 U16443 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14757) );
  AOI211_X1 U16444 ( .C1(n14750), .C2(n14749), .A(n14881), .B(n14748), .ZN(
        n14751) );
  INV_X1 U16445 ( .A(n14751), .ZN(n14756) );
  OAI211_X1 U16446 ( .C1(n14754), .C2(n14753), .A(n14752), .B(n14877), .ZN(
        n14755) );
  NAND4_X1 U16447 ( .A1(n14758), .A2(n14757), .A3(n14756), .A4(n14755), .ZN(
        P2_U3222) );
  AOI22_X1 U16448 ( .A1(n14849), .A2(P2_ADDR_REG_9__SCAN_IN), .B1(n14823), 
        .B2(n14759), .ZN(n14771) );
  OAI21_X1 U16449 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14763) );
  NAND2_X1 U16450 ( .A1(n14763), .A2(n14851), .ZN(n14769) );
  AOI21_X1 U16451 ( .B1(n14766), .B2(n14765), .A(n14764), .ZN(n14767) );
  OR2_X1 U16452 ( .A1(n14767), .A2(n14805), .ZN(n14768) );
  NAND4_X1 U16453 ( .A1(n14771), .A2(n14770), .A3(n14769), .A4(n14768), .ZN(
        P2_U3223) );
  AOI22_X1 U16454 ( .A1(n14849), .A2(P2_ADDR_REG_10__SCAN_IN), .B1(n14823), 
        .B2(n14772), .ZN(n14783) );
  OAI211_X1 U16455 ( .C1(n14775), .C2(n14774), .A(n14773), .B(n14877), .ZN(
        n14781) );
  AOI21_X1 U16456 ( .B1(n14777), .B2(n14776), .A(n14881), .ZN(n14779) );
  NAND2_X1 U16457 ( .A1(n14779), .A2(n14778), .ZN(n14780) );
  NAND4_X1 U16458 ( .A1(n14783), .A2(n14782), .A3(n14781), .A4(n14780), .ZN(
        P2_U3224) );
  AOI22_X1 U16459 ( .A1(n14849), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n14823), 
        .B2(n14784), .ZN(n14795) );
  AOI21_X1 U16460 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(n14788) );
  OR2_X1 U16461 ( .A1(n14788), .A2(n14881), .ZN(n14793) );
  OAI211_X1 U16462 ( .C1(n14791), .C2(n14790), .A(n14789), .B(n14877), .ZN(
        n14792) );
  NAND4_X1 U16463 ( .A1(n14795), .A2(n14794), .A3(n14793), .A4(n14792), .ZN(
        P2_U3225) );
  INV_X1 U16464 ( .A(n14796), .ZN(n14797) );
  AOI22_X1 U16465 ( .A1(n14849), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n14823), 
        .B2(n14797), .ZN(n14810) );
  NAND2_X1 U16466 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14809)
         );
  AOI21_X1 U16467 ( .B1(n14800), .B2(n14799), .A(n14798), .ZN(n14801) );
  OR2_X1 U16468 ( .A1(n14801), .A2(n14881), .ZN(n14808) );
  AOI21_X1 U16469 ( .B1(n14804), .B2(n14803), .A(n14802), .ZN(n14806) );
  OR2_X1 U16470 ( .A1(n14806), .A2(n14805), .ZN(n14807) );
  NAND4_X1 U16471 ( .A1(n14810), .A2(n14809), .A3(n14808), .A4(n14807), .ZN(
        P2_U3226) );
  AOI22_X1 U16472 ( .A1(n14849), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14821) );
  OAI211_X1 U16473 ( .C1(n14813), .C2(n14812), .A(n14851), .B(n14811), .ZN(
        n14820) );
  OAI211_X1 U16474 ( .C1(n14816), .C2(n14815), .A(n14877), .B(n14814), .ZN(
        n14819) );
  NAND2_X1 U16475 ( .A1(n14823), .A2(n14817), .ZN(n14818) );
  NAND4_X1 U16476 ( .A1(n14821), .A2(n14820), .A3(n14819), .A4(n14818), .ZN(
        P2_U3227) );
  AOI22_X1 U16477 ( .A1(n14849), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n14823), 
        .B2(n14822), .ZN(n14832) );
  NAND2_X1 U16478 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14831)
         );
  OAI211_X1 U16479 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n14825), .A(n14851), 
        .B(n14824), .ZN(n14830) );
  OAI211_X1 U16480 ( .C1(n14828), .C2(n14827), .A(n14877), .B(n14826), .ZN(
        n14829) );
  NAND4_X1 U16481 ( .A1(n14832), .A2(n14831), .A3(n14830), .A4(n14829), .ZN(
        P2_U3228) );
  OAI21_X1 U16482 ( .B1(n14834), .B2(n14873), .A(n14833), .ZN(n14835) );
  AOI21_X1 U16483 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n14849), .A(n14835), 
        .ZN(n14842) );
  OAI211_X1 U16484 ( .C1(n14837), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14877), 
        .B(n14836), .ZN(n14841) );
  OAI211_X1 U16485 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14839), .A(n14851), 
        .B(n14838), .ZN(n14840) );
  NAND3_X1 U16486 ( .A1(n14842), .A2(n14841), .A3(n14840), .ZN(P2_U3229) );
  OAI211_X1 U16487 ( .C1(n14845), .C2(n14844), .A(n14877), .B(n14843), .ZN(
        n14846) );
  NAND2_X1 U16488 ( .A1(n14847), .A2(n14846), .ZN(n14848) );
  AOI21_X1 U16489 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n14849), .A(n14848), 
        .ZN(n14855) );
  OAI211_X1 U16490 ( .C1(n14853), .C2(n14852), .A(n14851), .B(n14850), .ZN(
        n14854) );
  OAI211_X1 U16491 ( .C1(n14873), .C2(n14856), .A(n14855), .B(n14854), .ZN(
        P2_U3230) );
  OAI21_X1 U16492 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14868) );
  OAI211_X1 U16493 ( .C1(n14862), .C2(n14861), .A(n14877), .B(n14860), .ZN(
        n14864) );
  OAI211_X1 U16494 ( .C1(n14865), .C2(n14873), .A(n14864), .B(n14863), .ZN(
        n14866) );
  AOI21_X1 U16495 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n14849), .A(n14866), 
        .ZN(n14867) );
  OAI21_X1 U16496 ( .B1(n14881), .B2(n14868), .A(n14867), .ZN(P2_U3231) );
  AOI21_X1 U16497 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14870), .A(n14869), 
        .ZN(n14882) );
  NOR2_X1 U16498 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14871), .ZN(n14875) );
  NOR2_X1 U16499 ( .A1(n14873), .A2(n14872), .ZN(n14874) );
  AOI211_X1 U16500 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n14849), .A(n14875), 
        .B(n14874), .ZN(n14880) );
  OAI211_X1 U16501 ( .C1(n14878), .C2(P2_REG1_REG_18__SCAN_IN), .A(n14877), 
        .B(n14876), .ZN(n14879) );
  OAI211_X1 U16502 ( .C1(n14882), .C2(n14881), .A(n14880), .B(n14879), .ZN(
        P2_U3232) );
  AND2_X1 U16503 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14884), .ZN(P2_U3266) );
  AND2_X1 U16504 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14884), .ZN(P2_U3267) );
  AND2_X1 U16505 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14884), .ZN(P2_U3268) );
  AND2_X1 U16506 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14884), .ZN(P2_U3269) );
  AND2_X1 U16507 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14884), .ZN(P2_U3270) );
  AND2_X1 U16508 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14884), .ZN(P2_U3271) );
  AND2_X1 U16509 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14884), .ZN(P2_U3272) );
  AND2_X1 U16510 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14884), .ZN(P2_U3273) );
  AND2_X1 U16511 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14884), .ZN(P2_U3274) );
  AND2_X1 U16512 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14884), .ZN(P2_U3275) );
  AND2_X1 U16513 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14884), .ZN(P2_U3276) );
  AND2_X1 U16514 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14884), .ZN(P2_U3277) );
  AND2_X1 U16515 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14884), .ZN(P2_U3278) );
  AND2_X1 U16516 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14884), .ZN(P2_U3279) );
  AND2_X1 U16517 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14884), .ZN(P2_U3280) );
  AND2_X1 U16518 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14884), .ZN(P2_U3281) );
  AND2_X1 U16519 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14884), .ZN(P2_U3282) );
  AND2_X1 U16520 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14884), .ZN(P2_U3283) );
  AND2_X1 U16521 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14884), .ZN(P2_U3284) );
  AND2_X1 U16522 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14884), .ZN(P2_U3285) );
  AND2_X1 U16523 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14884), .ZN(P2_U3286) );
  AND2_X1 U16524 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14884), .ZN(P2_U3287) );
  AND2_X1 U16525 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14884), .ZN(P2_U3288) );
  AND2_X1 U16526 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14884), .ZN(P2_U3289) );
  AND2_X1 U16527 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14884), .ZN(P2_U3290) );
  AND2_X1 U16528 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14884), .ZN(P2_U3291) );
  AND2_X1 U16529 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14884), .ZN(P2_U3292) );
  AND2_X1 U16530 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14884), .ZN(P2_U3293) );
  AND2_X1 U16531 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14884), .ZN(P2_U3294) );
  AND2_X1 U16532 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14884), .ZN(P2_U3295) );
  AOI22_X1 U16533 ( .A1(n14887), .A2(n14886), .B1(n14885), .B2(n14889), .ZN(
        P2_U3416) );
  AOI21_X1 U16534 ( .B1(n14890), .B2(n14889), .A(n14888), .ZN(P2_U3417) );
  INV_X1 U16535 ( .A(n14891), .ZN(n14893) );
  INV_X1 U16536 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14892) );
  AOI22_X1 U16537 ( .A1(n14944), .A2(n14893), .B1(n14892), .B2(n14942), .ZN(
        P2_U3430) );
  OAI21_X1 U16538 ( .B1(n8191), .B2(n14927), .A(n14894), .ZN(n14896) );
  AOI211_X1 U16539 ( .C1(n14932), .C2(n14897), .A(n14896), .B(n14895), .ZN(
        n14946) );
  INV_X1 U16540 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14898) );
  AOI22_X1 U16541 ( .A1(n14944), .A2(n14946), .B1(n14898), .B2(n14942), .ZN(
        P2_U3436) );
  OAI21_X1 U16542 ( .B1(n6979), .B2(n14927), .A(n14899), .ZN(n14901) );
  AOI211_X1 U16543 ( .C1(n14934), .C2(n14902), .A(n14901), .B(n14900), .ZN(
        n14948) );
  INV_X1 U16544 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14903) );
  AOI22_X1 U16545 ( .A1(n14944), .A2(n14948), .B1(n14903), .B2(n14942), .ZN(
        P2_U3442) );
  INV_X1 U16546 ( .A(n14904), .ZN(n14906) );
  OAI21_X1 U16547 ( .B1(n14906), .B2(n14927), .A(n14905), .ZN(n14908) );
  AOI211_X1 U16548 ( .C1(n14932), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        n14950) );
  INV_X1 U16549 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14910) );
  AOI22_X1 U16550 ( .A1(n14944), .A2(n14950), .B1(n14910), .B2(n14942), .ZN(
        P2_U3445) );
  AOI21_X1 U16551 ( .B1(n14936), .B2(n14912), .A(n14911), .ZN(n14915) );
  NAND3_X1 U16552 ( .A1(n13531), .A2(n14913), .A3(n14934), .ZN(n14914) );
  AND3_X1 U16553 ( .A1(n14916), .A2(n14915), .A3(n14914), .ZN(n14952) );
  INV_X1 U16554 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14917) );
  AOI22_X1 U16555 ( .A1(n14944), .A2(n14952), .B1(n14917), .B2(n14942), .ZN(
        P2_U3448) );
  AOI21_X1 U16556 ( .B1(n14936), .B2(n14919), .A(n14918), .ZN(n14920) );
  OAI211_X1 U16557 ( .C1(n14923), .C2(n14922), .A(n14921), .B(n14920), .ZN(
        n14924) );
  INV_X1 U16558 ( .A(n14924), .ZN(n14954) );
  INV_X1 U16559 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U16560 ( .A1(n14944), .A2(n14954), .B1(n14925), .B2(n14942), .ZN(
        P2_U3451) );
  OAI21_X1 U16561 ( .B1(n14928), .B2(n14927), .A(n14926), .ZN(n14930) );
  AOI211_X1 U16562 ( .C1(n14932), .C2(n14931), .A(n14930), .B(n14929), .ZN(
        n14956) );
  INV_X1 U16563 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14933) );
  AOI22_X1 U16564 ( .A1(n14944), .A2(n14956), .B1(n14933), .B2(n14942), .ZN(
        P2_U3460) );
  AND2_X1 U16565 ( .A1(n14935), .A2(n14934), .ZN(n14940) );
  AND2_X1 U16566 ( .A1(n14937), .A2(n14936), .ZN(n14938) );
  NOR4_X1 U16567 ( .A1(n14941), .A2(n14940), .A3(n14939), .A4(n14938), .ZN(
        n14959) );
  INV_X1 U16568 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U16569 ( .A1(n14944), .A2(n14959), .B1(n14943), .B2(n14942), .ZN(
        P2_U3463) );
  AOI22_X1 U16570 ( .A1(n14960), .A2(n14946), .B1(n14945), .B2(n14957), .ZN(
        P2_U3501) );
  AOI22_X1 U16571 ( .A1(n14960), .A2(n14948), .B1(n14947), .B2(n14957), .ZN(
        P2_U3503) );
  AOI22_X1 U16572 ( .A1(n14960), .A2(n14950), .B1(n14949), .B2(n14957), .ZN(
        P2_U3504) );
  AOI22_X1 U16573 ( .A1(n14960), .A2(n14952), .B1(n14951), .B2(n14957), .ZN(
        P2_U3505) );
  AOI22_X1 U16574 ( .A1(n14960), .A2(n14954), .B1(n14953), .B2(n14957), .ZN(
        P2_U3506) );
  AOI22_X1 U16575 ( .A1(n14960), .A2(n14956), .B1(n14955), .B2(n14957), .ZN(
        P2_U3509) );
  AOI22_X1 U16576 ( .A1(n14960), .A2(n14959), .B1(n14958), .B2(n14957), .ZN(
        P2_U3510) );
  NOR2_X1 U16577 ( .A1(P3_U3897), .A2(n15089), .ZN(P3_U3150) );
  OAI22_X1 U16578 ( .A1(n14973), .A2(n14962), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14961), .ZN(n14968) );
  OAI211_X1 U16579 ( .C1(n14965), .C2(n14964), .A(n14963), .B(n14974), .ZN(
        n14966) );
  INV_X1 U16580 ( .A(n14966), .ZN(n14967) );
  AOI211_X1 U16581 ( .C1(n14982), .C2(n14969), .A(n14968), .B(n14967), .ZN(
        n14970) );
  OAI21_X1 U16582 ( .B1(n14985), .B2(n14971), .A(n14970), .ZN(P3_U3153) );
  OAI21_X1 U16583 ( .B1(n14973), .B2(n15170), .A(n14972), .ZN(n14980) );
  OAI211_X1 U16584 ( .C1(n14977), .C2(n14976), .A(n14975), .B(n14974), .ZN(
        n14978) );
  INV_X1 U16585 ( .A(n14978), .ZN(n14979) );
  AOI211_X1 U16586 ( .C1(n14982), .C2(n14981), .A(n14980), .B(n14979), .ZN(
        n14983) );
  OAI21_X1 U16587 ( .B1(n14985), .B2(n14984), .A(n14983), .ZN(P3_U3161) );
  AOI22_X1 U16588 ( .A1(n15002), .A2(P3_IR_REG_0__SCAN_IN), .B1(n15089), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n14992) );
  INV_X1 U16589 ( .A(n15094), .ZN(n14986) );
  NAND3_X1 U16590 ( .A1(n14986), .A2(n15102), .A3(n15076), .ZN(n14990) );
  OAI21_X1 U16591 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n14988), .A(n14987), .ZN(
        n14989) );
  NAND2_X1 U16592 ( .A1(n14990), .A2(n14989), .ZN(n14991) );
  OAI211_X1 U16593 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n14993), .A(n14992), .B(
        n14991), .ZN(P3_U3182) );
  INV_X1 U16594 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15012) );
  NAND2_X1 U16595 ( .A1(n6649), .A2(n14994), .ZN(n14995) );
  XNOR2_X1 U16596 ( .A(n14996), .B(n14995), .ZN(n14997) );
  NOR2_X1 U16597 ( .A1(n14997), .A2(n15076), .ZN(n15008) );
  AOI21_X1 U16598 ( .B1(n14999), .B2(n9016), .A(n14998), .ZN(n15006) );
  OAI21_X1 U16599 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15001), .A(n15000), .ZN(
        n15004) );
  AOI22_X1 U16600 ( .A1(n15004), .A2(n15094), .B1(n15003), .B2(n15002), .ZN(
        n15005) );
  OAI21_X1 U16601 ( .B1(n15006), .B2(n15102), .A(n15005), .ZN(n15007) );
  NOR2_X1 U16602 ( .A1(n15008), .A2(n15007), .ZN(n15010) );
  OAI211_X1 U16603 ( .C1(n15012), .C2(n15011), .A(n15010), .B(n15009), .ZN(
        P3_U3191) );
  AOI21_X1 U16604 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15029) );
  OAI21_X1 U16605 ( .B1(n15018), .B2(n15017), .A(n15016), .ZN(n15027) );
  NAND2_X1 U16606 ( .A1(n15089), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n15019) );
  OAI211_X1 U16607 ( .C1(n15092), .C2(n15021), .A(n15020), .B(n15019), .ZN(
        n15026) );
  AOI21_X1 U16608 ( .B1(n15023), .B2(n15022), .A(n6641), .ZN(n15024) );
  NOR2_X1 U16609 ( .A1(n15024), .A2(n15076), .ZN(n15025) );
  AOI211_X1 U16610 ( .C1(n15094), .C2(n15027), .A(n15026), .B(n15025), .ZN(
        n15028) );
  OAI21_X1 U16611 ( .B1(n15029), .B2(n15102), .A(n15028), .ZN(P3_U3192) );
  AOI21_X1 U16612 ( .B1(n12839), .B2(n15031), .A(n15030), .ZN(n15045) );
  OAI21_X1 U16613 ( .B1(n15033), .B2(P3_REG1_REG_11__SCAN_IN), .A(n15032), 
        .ZN(n15034) );
  AND2_X1 U16614 ( .A1(n15034), .A2(n15094), .ZN(n15038) );
  OAI21_X1 U16615 ( .B1(n15092), .B2(n15036), .A(n15035), .ZN(n15037) );
  AOI211_X1 U16616 ( .C1(P3_ADDR_REG_11__SCAN_IN), .C2(n15089), .A(n15038), 
        .B(n15037), .ZN(n15044) );
  AOI21_X1 U16617 ( .B1(n15041), .B2(n15040), .A(n15039), .ZN(n15042) );
  OR2_X1 U16618 ( .A1(n15042), .A2(n15076), .ZN(n15043) );
  OAI211_X1 U16619 ( .C1(n15045), .C2(n15102), .A(n15044), .B(n15043), .ZN(
        P3_U3193) );
  AOI21_X1 U16620 ( .B1(n15048), .B2(n15047), .A(n15046), .ZN(n15062) );
  OAI21_X1 U16621 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(n15052) );
  AND2_X1 U16622 ( .A1(n15052), .A2(n15094), .ZN(n15056) );
  OAI21_X1 U16623 ( .B1(n15092), .B2(n15054), .A(n15053), .ZN(n15055) );
  AOI211_X1 U16624 ( .C1(P3_ADDR_REG_12__SCAN_IN), .C2(n15089), .A(n15056), 
        .B(n15055), .ZN(n15061) );
  OAI211_X1 U16625 ( .C1(n15059), .C2(n15058), .A(n15057), .B(n15096), .ZN(
        n15060) );
  OAI211_X1 U16626 ( .C1(n15062), .C2(n15102), .A(n15061), .B(n15060), .ZN(
        P3_U3194) );
  AOI21_X1 U16627 ( .B1(n9076), .B2(n15064), .A(n15063), .ZN(n15080) );
  OAI21_X1 U16628 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15066), .A(n15065), 
        .ZN(n15072) );
  NOR2_X1 U16629 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15067), .ZN(n15068) );
  AOI21_X1 U16630 ( .B1(n15089), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15068), 
        .ZN(n15069) );
  OAI21_X1 U16631 ( .B1(n15092), .B2(n15070), .A(n15069), .ZN(n15071) );
  AOI21_X1 U16632 ( .B1(n15072), .B2(n15094), .A(n15071), .ZN(n15079) );
  AOI21_X1 U16633 ( .B1(n15075), .B2(n15074), .A(n15073), .ZN(n15077) );
  OR2_X1 U16634 ( .A1(n15077), .A2(n15076), .ZN(n15078) );
  OAI211_X1 U16635 ( .C1(n15080), .C2(n15102), .A(n15079), .B(n15078), .ZN(
        P3_U3195) );
  AOI21_X1 U16636 ( .B1(n15083), .B2(n15082), .A(n15081), .ZN(n15103) );
  OAI21_X1 U16637 ( .B1(n15086), .B2(n15085), .A(n15084), .ZN(n15095) );
  NOR2_X1 U16638 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15087), .ZN(n15088) );
  AOI21_X1 U16639 ( .B1(n15089), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n15088), 
        .ZN(n15090) );
  OAI21_X1 U16640 ( .B1(n15092), .B2(n15091), .A(n15090), .ZN(n15093) );
  AOI21_X1 U16641 ( .B1(n15095), .B2(n15094), .A(n15093), .ZN(n15101) );
  OAI211_X1 U16642 ( .C1(n15099), .C2(n15098), .A(n15097), .B(n15096), .ZN(
        n15100) );
  OAI211_X1 U16643 ( .C1(n15103), .C2(n15102), .A(n15101), .B(n15100), .ZN(
        P3_U3196) );
  INV_X1 U16644 ( .A(n15119), .ZN(n15114) );
  XNOR2_X1 U16645 ( .A(n15105), .B(n15104), .ZN(n15138) );
  NOR2_X1 U16646 ( .A1(n15106), .A2(n15185), .ZN(n15137) );
  INV_X1 U16647 ( .A(n15137), .ZN(n15108) );
  OAI22_X1 U16648 ( .A1(n15108), .A2(n15122), .B1(n15121), .B2(n15107), .ZN(
        n15113) );
  XNOR2_X1 U16649 ( .A(n15109), .B(n15104), .ZN(n15112) );
  NAND2_X1 U16650 ( .A1(n15138), .A2(n15175), .ZN(n15111) );
  OAI211_X1 U16651 ( .C1(n15117), .C2(n15112), .A(n15111), .B(n15110), .ZN(
        n15136) );
  AOI211_X1 U16652 ( .C1(n15114), .C2(n15138), .A(n15113), .B(n15136), .ZN(
        n15115) );
  AOI22_X1 U16653 ( .A1(n15128), .A2(n6655), .B1(n15115), .B2(n15126), .ZN(
        P3_U3231) );
  XOR2_X1 U16654 ( .A(n15116), .B(n10775), .Z(n15118) );
  NOR2_X1 U16655 ( .A1(n15118), .A2(n15117), .ZN(n15134) );
  XNOR2_X1 U16656 ( .A(n12138), .B(n10775), .ZN(n15130) );
  AOI21_X1 U16657 ( .B1(n15164), .B2(n15119), .A(n15130), .ZN(n15125) );
  NOR2_X1 U16658 ( .A1(n6535), .A2(n15185), .ZN(n15132) );
  INV_X1 U16659 ( .A(n15132), .ZN(n15123) );
  OAI22_X1 U16660 ( .A1(n15123), .A2(n15122), .B1(n15121), .B2(n15120), .ZN(
        n15124) );
  NOR4_X1 U16661 ( .A1(n15134), .A2(n15125), .A3(n15131), .A4(n15124), .ZN(
        n15127) );
  AOI22_X1 U16662 ( .A1(n15128), .A2(n8852), .B1(n15127), .B2(n15126), .ZN(
        P3_U3232) );
  INV_X1 U16663 ( .A(n15190), .ZN(n15129) );
  NOR2_X1 U16664 ( .A1(n15130), .A2(n15129), .ZN(n15133) );
  NOR4_X1 U16665 ( .A1(n15134), .A2(n15133), .A3(n15132), .A4(n15131), .ZN(
        n15194) );
  INV_X1 U16666 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15135) );
  AOI22_X1 U16667 ( .A1(n15193), .A2(n15194), .B1(n15135), .B2(n15191), .ZN(
        P3_U3393) );
  AOI211_X1 U16668 ( .C1(n15138), .C2(n15182), .A(n15137), .B(n15136), .ZN(
        n15195) );
  INV_X1 U16669 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15139) );
  AOI22_X1 U16670 ( .A1(n15193), .A2(n15195), .B1(n15139), .B2(n15191), .ZN(
        P3_U3396) );
  INV_X1 U16671 ( .A(n15182), .ZN(n15171) );
  OAI22_X1 U16672 ( .A1(n15141), .A2(n15171), .B1(n15140), .B2(n15185), .ZN(
        n15144) );
  INV_X1 U16673 ( .A(n15142), .ZN(n15143) );
  AOI211_X1 U16674 ( .C1(n15175), .C2(n15145), .A(n15144), .B(n15143), .ZN(
        n15196) );
  INV_X1 U16675 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15146) );
  AOI22_X1 U16676 ( .A1(n15193), .A2(n15196), .B1(n15146), .B2(n15191), .ZN(
        P3_U3399) );
  OAI22_X1 U16677 ( .A1(n15148), .A2(n15171), .B1(n15147), .B2(n15185), .ZN(
        n15149) );
  NOR2_X1 U16678 ( .A1(n15150), .A2(n15149), .ZN(n15197) );
  INV_X1 U16679 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15151) );
  AOI22_X1 U16680 ( .A1(n15193), .A2(n15197), .B1(n15151), .B2(n15191), .ZN(
        P3_U3402) );
  INV_X1 U16681 ( .A(n15152), .ZN(n15156) );
  OAI21_X1 U16682 ( .B1(n15154), .B2(n15185), .A(n15153), .ZN(n15155) );
  AOI21_X1 U16683 ( .B1(n15156), .B2(n15190), .A(n15155), .ZN(n15198) );
  INV_X1 U16684 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15157) );
  AOI22_X1 U16685 ( .A1(n15193), .A2(n15198), .B1(n15157), .B2(n15191), .ZN(
        P3_U3405) );
  NOR2_X1 U16686 ( .A1(n15158), .A2(n15185), .ZN(n15160) );
  AOI211_X1 U16687 ( .C1(n15182), .C2(n15161), .A(n15160), .B(n15159), .ZN(
        n15199) );
  INV_X1 U16688 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15162) );
  AOI22_X1 U16689 ( .A1(n15193), .A2(n15199), .B1(n15162), .B2(n15191), .ZN(
        P3_U3408) );
  AOI21_X1 U16690 ( .B1(n15164), .B2(n15171), .A(n15163), .ZN(n15165) );
  AOI211_X1 U16691 ( .C1(n15168), .C2(n15167), .A(n15166), .B(n15165), .ZN(
        n15200) );
  INV_X1 U16692 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U16693 ( .A1(n15193), .A2(n15200), .B1(n15169), .B2(n15191), .ZN(
        P3_U3411) );
  INV_X1 U16694 ( .A(n15172), .ZN(n15176) );
  OAI22_X1 U16695 ( .A1(n15172), .A2(n15171), .B1(n15170), .B2(n15185), .ZN(
        n15174) );
  AOI211_X1 U16696 ( .C1(n15176), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15201) );
  INV_X1 U16697 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15177) );
  AOI22_X1 U16698 ( .A1(n15193), .A2(n15201), .B1(n15177), .B2(n15191), .ZN(
        P3_U3414) );
  INV_X1 U16699 ( .A(n15178), .ZN(n15183) );
  NOR2_X1 U16700 ( .A1(n15179), .A2(n15185), .ZN(n15181) );
  AOI211_X1 U16701 ( .C1(n15183), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15202) );
  INV_X1 U16702 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15184) );
  AOI22_X1 U16703 ( .A1(n15193), .A2(n15202), .B1(n15184), .B2(n15191), .ZN(
        P3_U3417) );
  NOR2_X1 U16704 ( .A1(n15186), .A2(n15185), .ZN(n15188) );
  AOI211_X1 U16705 ( .C1(n15190), .C2(n15189), .A(n15188), .B(n15187), .ZN(
        n15204) );
  INV_X1 U16706 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15192) );
  AOI22_X1 U16707 ( .A1(n15193), .A2(n15204), .B1(n15192), .B2(n15191), .ZN(
        P3_U3420) );
  AOI22_X1 U16708 ( .A1(n15205), .A2(n15194), .B1(n11107), .B2(n15203), .ZN(
        P3_U3460) );
  AOI22_X1 U16709 ( .A1(n15205), .A2(n15195), .B1(n9863), .B2(n15203), .ZN(
        P3_U3461) );
  AOI22_X1 U16710 ( .A1(n15205), .A2(n15196), .B1(n9889), .B2(n15203), .ZN(
        P3_U3462) );
  AOI22_X1 U16711 ( .A1(n15205), .A2(n15197), .B1(n8915), .B2(n15203), .ZN(
        P3_U3463) );
  AOI22_X1 U16712 ( .A1(n15205), .A2(n15198), .B1(n8943), .B2(n15203), .ZN(
        P3_U3464) );
  AOI22_X1 U16713 ( .A1(n15205), .A2(n15199), .B1(n8962), .B2(n15203), .ZN(
        P3_U3465) );
  AOI22_X1 U16714 ( .A1(n15205), .A2(n15200), .B1(n8972), .B2(n15203), .ZN(
        P3_U3466) );
  AOI22_X1 U16715 ( .A1(n15205), .A2(n15201), .B1(n8996), .B2(n15203), .ZN(
        P3_U3467) );
  AOI22_X1 U16716 ( .A1(n15205), .A2(n15202), .B1(n9019), .B2(n15203), .ZN(
        P3_U3468) );
  AOI22_X1 U16717 ( .A1(n15205), .A2(n15204), .B1(n9030), .B2(n15203), .ZN(
        P3_U3469) );
  AOI21_X1 U16718 ( .B1(n15208), .B2(n15207), .A(n15206), .ZN(SUB_1596_U59) );
  OAI21_X1 U16719 ( .B1(n15211), .B2(n15210), .A(n15209), .ZN(SUB_1596_U58) );
  XOR2_X1 U16720 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15212), .Z(SUB_1596_U53) );
  AOI21_X1 U16721 ( .B1(n15215), .B2(n15214), .A(n15213), .ZN(SUB_1596_U56) );
  AOI21_X1 U16722 ( .B1(n15218), .B2(n15217), .A(n15216), .ZN(n15219) );
  XOR2_X1 U16723 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15219), .Z(SUB_1596_U60) );
  AOI21_X1 U16724 ( .B1(n15222), .B2(n15221), .A(n15220), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7267 ( .A(n11835), .Z(n11961) );
  OAI21_X1 U7282 ( .B1(n12873), .B2(n9700), .A(n12698), .ZN(n9702) );
  CLKBUF_X2 U7309 ( .A(n8984), .Z(n9714) );
  XNOR2_X1 U9784 ( .A(n7498), .B(n7497), .ZN(n7500) );
  CLKBUF_X1 U14394 ( .A(n10148), .Z(n6469) );
endmodule

