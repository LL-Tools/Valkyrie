

module b17_C_AntiSAT_k_128_4 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9622, n9623, n9625, n9626, n9627, n9628, n9629, n9631, n9632, n9633,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152;

  NOR2_X1 U11066 ( .A1(n13418), .A2(n13417), .ZN(n13441) );
  NOR2_X1 U11067 ( .A1(n12622), .A2(n12621), .ZN(n15118) );
  AND2_X1 U11068 ( .A1(n10028), .A2(n10027), .ZN(n12622) );
  OAI21_X1 U11069 ( .B1(n15131), .B2(n10697), .A(n10029), .ZN(n10028) );
  AOI21_X1 U11070 ( .B1(n15131), .B2(n12626), .A(n15130), .ZN(n10027) );
  NOR2_X1 U11071 ( .A1(n17594), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17593) );
  INV_X1 U11072 ( .A(n15943), .ZN(n14761) );
  INV_X1 U11074 ( .A(n18892), .ZN(n18268) );
  OR2_X1 U11075 ( .A1(n10318), .A2(n10309), .ZN(n19404) );
  OR2_X1 U11076 ( .A1(n10318), .A2(n10313), .ZN(n15552) );
  OR2_X2 U11077 ( .A1(n10314), .A2(n10320), .ZN(n19469) );
  NAND2_X1 U11078 ( .A1(n11538), .A2(n11537), .ZN(n11609) );
  OR2_X1 U11079 ( .A1(n20378), .A2(n11443), .ZN(n20315) );
  XNOR2_X1 U11080 ( .A(n10273), .B(n10274), .ZN(n10287) );
  INV_X2 U11081 ( .A(n17233), .ZN(n17244) );
  AND2_X1 U11082 ( .A1(n12890), .A2(n10330), .ZN(n12929) );
  AND2_X1 U11083 ( .A1(n10222), .A2(n10221), .ZN(n10254) );
  AND2_X1 U11084 ( .A1(n10327), .A2(n12890), .ZN(n12930) );
  CLKBUF_X2 U11085 ( .A(n13433), .Z(n13419) );
  CLKBUF_X2 U11086 ( .A(n11286), .Z(n12239) );
  CLKBUF_X1 U11087 ( .A(n11349), .Z(n12211) );
  AND2_X1 U11088 ( .A1(n13621), .A2(n11404), .ZN(n15770) );
  AND2_X1 U11089 ( .A1(n10210), .A2(n9987), .ZN(n10247) );
  NAND2_X1 U11090 ( .A1(n10217), .A2(n16384), .ZN(n10767) );
  BUF_X2 U11091 ( .A(n11403), .Z(n20261) );
  BUF_X1 U11092 ( .A(n10203), .Z(n15558) );
  CLKBUF_X2 U11093 ( .A(n11402), .Z(n20295) );
  AND4_X1 U11094 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n10096) );
  NAND4_X2 U11095 ( .A1(n11281), .A2(n11280), .A3(n11279), .A4(n11278), .ZN(
        n11541) );
  INV_X1 U11096 ( .A(n11379), .ZN(n12238) );
  BUF_X2 U11097 ( .A(n11340), .Z(n12212) );
  AND2_X1 U11098 ( .A1(n13957), .A2(n9845), .ZN(n11286) );
  INV_X1 U11099 ( .A(n12184), .ZN(n11779) );
  CLKBUF_X1 U11100 ( .A(n20305), .Z(n9622) );
  NOR2_X1 U11101 ( .A1(n20256), .A2(n20258), .ZN(n20305) );
  CLKBUF_X1 U11102 ( .A(n20304), .Z(n9623) );
  NOR2_X1 U11103 ( .A1(n20258), .A2(n20257), .ZN(n20304) );
  INV_X1 U11105 ( .A(n21152), .ZN(n9625) );
  INV_X1 U11106 ( .A(n10497), .ZN(n10751) );
  AND2_X1 U11107 ( .A1(n12890), .A2(n10328), .ZN(n12924) );
  NOR2_X1 U11108 ( .A1(n10582), .A2(n10581), .ZN(n10036) );
  INV_X1 U11109 ( .A(n10204), .ZN(n11200) );
  NOR2_X1 U11110 ( .A1(n11356), .A2(n11355), .ZN(n11413) );
  AND2_X1 U11111 ( .A1(n12890), .A2(n10329), .ZN(n12923) );
  AND2_X1 U11112 ( .A1(n10735), .A2(n14169), .ZN(n12913) );
  INV_X1 U11113 ( .A(n11130), .ZN(n12909) );
  NAND2_X1 U11114 ( .A1(n10391), .A2(n9655), .ZN(n10582) );
  NAND2_X1 U11115 ( .A1(n19364), .A2(n10203), .ZN(n10213) );
  INV_X1 U11117 ( .A(n12555), .ZN(n12584) );
  NAND2_X1 U11118 ( .A1(n11443), .A2(n20378), .ZN(n11478) );
  INV_X1 U11119 ( .A(n12238), .ZN(n12175) );
  XNOR2_X1 U11120 ( .A(n13012), .B(n13013), .ZN(n14983) );
  OAI21_X1 U11121 ( .B1(n15191), .B2(n15192), .A(n15453), .ZN(n16248) );
  OAI21_X1 U11123 ( .B1(n14166), .B2(n13088), .A(n12764), .ZN(n13597) );
  NOR2_X1 U11124 ( .A1(n17581), .A2(n16462), .ZN(n15721) );
  NAND2_X1 U11125 ( .A1(n17721), .A2(n17834), .ZN(n17676) );
  AOI211_X2 U11126 ( .C1(n9639), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n13275), .B(n13274), .ZN(n18281) );
  CLKBUF_X3 U11127 ( .A(n11426), .Z(n12555) );
  INV_X1 U11128 ( .A(n13549), .ZN(n19284) );
  BUF_X1 U11129 ( .A(n12769), .Z(n14127) );
  INV_X1 U11130 ( .A(n17226), .ZN(n17252) );
  INV_X2 U11131 ( .A(n13156), .ZN(n17246) );
  NAND2_X1 U11132 ( .A1(n17715), .A2(n17784), .ZN(n17919) );
  NAND2_X1 U11133 ( .A1(n16466), .A2(n16464), .ZN(n17834) );
  INV_X1 U11134 ( .A(n15877), .ZN(n20101) );
  OR2_X2 U11135 ( .A1(n18740), .A2(n18750), .ZN(n16579) );
  AOI211_X1 U11136 ( .C1(n9632), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n13125), .B(n13124), .ZN(n17428) );
  INV_X2 U11137 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18879) );
  INV_X1 U11138 ( .A(n13141), .ZN(n17219) );
  BUF_X1 U11139 ( .A(n15595), .Z(n9626) );
  AOI211_X1 U11140 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n13265), .B(n13264), .ZN(n15595) );
  NAND2_X2 U11141 ( .A1(n20195), .A2(n12357), .ZN(n12358) );
  INV_X2 U11142 ( .A(n16984), .ZN(n17264) );
  NAND2_X2 U11143 ( .A1(n15515), .A2(n14169), .ZN(n13428) );
  AND2_X2 U11144 ( .A1(n15504), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15515) );
  NAND2_X2 U11145 ( .A1(n9988), .A2(n10495), .ZN(n10969) );
  INV_X2 U11146 ( .A(n11270), .ZN(n9627) );
  INV_X1 U11147 ( .A(n9627), .ZN(n9628) );
  NAND2_X1 U11149 ( .A1(n13957), .A2(n14918), .ZN(n11270) );
  AOI21_X2 U11150 ( .B1(n9880), .B2(n9662), .A(n18160), .ZN(n13354) );
  NAND2_X1 U11151 ( .A1(n14282), .A2(n18879), .ZN(n17233) );
  NAND2_X2 U11154 ( .A1(n10200), .A2(n10199), .ZN(n10205) );
  NOR2_X2 U11155 ( .A1(n15711), .A2(n18075), .ZN(n17940) );
  NAND2_X2 U11156 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18076), .ZN(
        n18075) );
  NAND2_X2 U11158 ( .A1(n10277), .A2(n10276), .ZN(n10840) );
  AND2_X4 U11159 ( .A1(n10330), .A2(n16364), .ZN(n10342) );
  AND2_X4 U11160 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10330) );
  XNOR2_X2 U11161 ( .A(n12366), .B(n20220), .ZN(n13911) );
  NAND2_X2 U11162 ( .A1(n13785), .A2(n12359), .ZN(n12366) );
  NAND2_X1 U11163 ( .A1(n14136), .A2(n14137), .ZN(n10812) );
  NAND2_X1 U11164 ( .A1(n9767), .A2(n9881), .ZN(n16458) );
  AND2_X1 U11165 ( .A1(n15381), .A2(n9721), .ZN(n14312) );
  INV_X1 U11166 ( .A(n17789), .ZN(n17784) );
  OR2_X1 U11168 ( .A1(n11538), .A2(n11537), .ZN(n11539) );
  INV_X4 U11169 ( .A(n17927), .ZN(n17884) );
  NAND2_X1 U11170 ( .A1(n11598), .A2(n11597), .ZN(n14910) );
  NOR2_X2 U11171 ( .A1(n18691), .A2(n18712), .ZN(n18129) );
  NOR3_X1 U11172 ( .A1(n15805), .A2(n18262), .A3(n18268), .ZN(n15808) );
  OAI21_X1 U11173 ( .B1(n11442), .B2(n11441), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11446) );
  CLKBUF_X2 U11174 ( .A(n10261), .Z(n10956) );
  INV_X1 U11175 ( .A(n11425), .ZN(n9631) );
  CLKBUF_X2 U11176 ( .A(n10995), .Z(n11187) );
  AOI211_X1 U11177 ( .C1(n17246), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n13114), .B(n13113), .ZN(n17419) );
  CLKBUF_X2 U11178 ( .A(n10978), .Z(n11184) );
  INV_X4 U11179 ( .A(n14029), .ZN(n9930) );
  NOR2_X1 U11180 ( .A1(n15543), .A2(n10495), .ZN(n10220) );
  NAND2_X1 U11181 ( .A1(n20261), .A2(n20275), .ZN(n14036) );
  NAND2_X1 U11182 ( .A1(n11473), .A2(n11402), .ZN(n12586) );
  BUF_X2 U11183 ( .A(n11473), .Z(n20290) );
  AND2_X1 U11184 ( .A1(n11413), .A2(n12342), .ZN(n11405) );
  INV_X1 U11185 ( .A(n12342), .ZN(n13404) );
  NAND2_X2 U11186 ( .A1(n11336), .A2(n10096), .ZN(n12342) );
  AOI211_X1 U11187 ( .C1(n17255), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n13301), .B(n13300), .ZN(n13302) );
  INV_X1 U11188 ( .A(n11422), .ZN(n9948) );
  BUF_X1 U11189 ( .A(n11413), .Z(n20280) );
  NAND4_X2 U11190 ( .A1(n11323), .A2(n11322), .A3(n11321), .A4(n11320), .ZN(
        n11402) );
  NAND4_X2 U11191 ( .A1(n11303), .A2(n11301), .A3(n11302), .A4(n11300), .ZN(
        n11422) );
  AND4_X1 U11192 ( .A1(n11269), .A2(n11268), .A3(n11267), .A4(n11266), .ZN(
        n11280) );
  AND4_X1 U11193 ( .A1(n11311), .A2(n11310), .A3(n11309), .A4(n11308), .ZN(
        n11322) );
  AND4_X1 U11194 ( .A1(n11295), .A2(n11294), .A3(n11293), .A4(n11292), .ZN(
        n11301) );
  AND4_X1 U11195 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(
        n11323) );
  INV_X4 U11196 ( .A(n17199), .ZN(n17230) );
  INV_X1 U11197 ( .A(n10126), .ZN(n9636) );
  INV_X4 U11198 ( .A(n12182), .ZN(n11794) );
  INV_X4 U11199 ( .A(n13126), .ZN(n9632) );
  INV_X1 U11200 ( .A(n17251), .ZN(n17199) );
  CLKBUF_X2 U11201 ( .A(n10341), .Z(n13431) );
  INV_X4 U11202 ( .A(n17058), .ZN(n13196) );
  AND2_X2 U11203 ( .A1(n14918), .A2(n11249), .ZN(n11367) );
  INV_X2 U11204 ( .A(n18229), .ZN(n9633) );
  NOR2_X1 U11205 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16942) );
  INV_X1 U11206 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11241) );
  NOR2_X2 U11207 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11249) );
  AND2_X1 U11208 ( .A1(n11239), .A2(n9942), .ZN(n9941) );
  OR2_X1 U11209 ( .A1(n14795), .A2(n20016), .ZN(n9755) );
  AND2_X1 U11210 ( .A1(n10079), .A2(n13474), .ZN(n9754) );
  OAI21_X1 U11211 ( .B1(n13094), .B2(n19297), .A(n13093), .ZN(n13095) );
  OR2_X1 U11212 ( .A1(n15148), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15300) );
  OR2_X1 U11213 ( .A1(n14328), .A2(n20258), .ZN(n10079) );
  AOI21_X1 U11214 ( .B1(n13401), .B2(n13402), .A(n9945), .ZN(n14658) );
  OR2_X1 U11215 ( .A1(n14651), .A2(n14650), .ZN(n14652) );
  OAI21_X1 U11216 ( .B1(n14378), .B2(n14379), .A(n14365), .ZN(n14675) );
  CLKBUF_X1 U11217 ( .A(n13471), .Z(n14366) );
  NAND2_X1 U11218 ( .A1(n9772), .A2(n9773), .ZN(n15407) );
  NAND2_X1 U11219 ( .A1(n10055), .A2(n14966), .ZN(n14976) );
  NOR2_X1 U11220 ( .A1(n14671), .A2(n12606), .ZN(n12438) );
  AND2_X1 U11221 ( .A1(n9887), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12436) );
  CLKBUF_X1 U11222 ( .A(n14497), .Z(n14503) );
  AOI21_X2 U11223 ( .B1(n15439), .B2(n15437), .A(n15194), .ZN(n15231) );
  NAND2_X1 U11224 ( .A1(n12433), .A2(n14761), .ZN(n9887) );
  NAND2_X1 U11225 ( .A1(n12433), .A2(n15896), .ZN(n14709) );
  AOI21_X1 U11226 ( .B1(n16248), .B2(n16245), .A(n15193), .ZN(n15439) );
  OR2_X1 U11227 ( .A1(n13014), .A2(n13013), .ZN(n10065) );
  NAND2_X1 U11228 ( .A1(n9901), .A2(n14862), .ZN(n15895) );
  OR2_X1 U11229 ( .A1(n12988), .A2(n12989), .ZN(n12990) );
  NAND2_X1 U11230 ( .A1(n12414), .A2(n12413), .ZN(n14772) );
  AND2_X1 U11231 ( .A1(n12724), .A2(n12723), .ZN(n15278) );
  XNOR2_X1 U11232 ( .A(n12724), .B(n11188), .ZN(n16115) );
  OAI211_X1 U11233 ( .C1(n10812), .C2(n10813), .A(n10811), .B(n10042), .ZN(
        n14246) );
  OR2_X1 U11234 ( .A1(n12629), .A2(n12631), .ZN(n16124) );
  AOI21_X1 U11235 ( .B1(n17745), .B2(n17581), .A(n16463), .ZN(n17570) );
  NAND2_X1 U11236 ( .A1(n16458), .A2(n17944), .ZN(n17580) );
  OR2_X1 U11237 ( .A1(n16458), .A2(n17944), .ZN(n17581) );
  XNOR2_X1 U11238 ( .A(n10792), .B(n11003), .ZN(n19292) );
  NAND2_X1 U11239 ( .A1(n20184), .A2(n12374), .ZN(n15964) );
  XNOR2_X1 U11240 ( .A(n12580), .B(n12579), .ZN(n12659) );
  AND2_X1 U11241 ( .A1(n11671), .A2(n11670), .ZN(n13905) );
  OAI211_X1 U11242 ( .C1(n13911), .C2(n9891), .A(n20185), .B(n9890), .ZN(
        n20184) );
  NAND2_X1 U11243 ( .A1(n12406), .A2(n12405), .ZN(n12419) );
  AND2_X1 U11244 ( .A1(n10580), .A2(n10579), .ZN(n10808) );
  NOR2_X1 U11245 ( .A1(n19599), .A2(n19600), .ZN(n19651) );
  XNOR2_X1 U11246 ( .A(n12406), .B(n11700), .ZN(n12395) );
  NAND2_X1 U11247 ( .A1(n9847), .A2(n11696), .ZN(n12406) );
  NAND2_X1 U11248 ( .A1(n12366), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12367) );
  AND2_X1 U11249 ( .A1(n9765), .A2(n9764), .ZN(n17607) );
  NOR2_X1 U11250 ( .A1(n17759), .A2(n18072), .ZN(n18065) );
  NAND2_X1 U11251 ( .A1(n11659), .A2(n11660), .ZN(n11694) );
  AOI22_X1 U11252 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19538), .B1(
        n10443), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U11253 ( .A1(n17676), .A2(n17662), .ZN(n17710) );
  NAND2_X1 U11254 ( .A1(n12778), .A2(n12777), .ZN(n13692) );
  NAND2_X1 U11255 ( .A1(n11610), .A2(n9846), .ZN(n11662) );
  NAND2_X1 U11256 ( .A1(n10298), .A2(n10302), .ZN(n10553) );
  INV_X1 U11257 ( .A(n10319), .ZN(n10298) );
  INV_X1 U11258 ( .A(n11609), .ZN(n11610) );
  OR2_X2 U11259 ( .A1(n10318), .A2(n10317), .ZN(n19435) );
  NAND2_X1 U11260 ( .A1(n9643), .A2(n10302), .ZN(n19692) );
  OR2_X2 U11261 ( .A1(n10318), .A2(n10320), .ZN(n10544) );
  OR2_X1 U11262 ( .A1(n10319), .A2(n10313), .ZN(n10540) );
  XNOR2_X1 U11263 ( .A(n11609), .B(n14910), .ZN(n20260) );
  NAND2_X1 U11264 ( .A1(n12756), .A2(n12755), .ZN(n12779) );
  NOR2_X1 U11265 ( .A1(n18220), .A2(n18235), .ZN(n18246) );
  AND2_X1 U11266 ( .A1(n12349), .A2(n11564), .ZN(n11537) );
  XNOR2_X1 U11267 ( .A(n13970), .B(n20415), .ZN(n20536) );
  XNOR2_X1 U11268 ( .A(n13597), .B(n12765), .ZN(n13860) );
  OR2_X1 U11269 ( .A1(n13527), .A2(n19320), .ZN(n10320) );
  NOR2_X1 U11270 ( .A1(n17300), .A2(n17437), .ZN(n17357) );
  OAI21_X1 U11271 ( .B1(n14906), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11495), 
        .ZN(n12349) );
  OAI21_X1 U11272 ( .B1(n11556), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11552), 
        .ZN(n11550) );
  XNOR2_X1 U11273 ( .A(n10841), .B(n10842), .ZN(n10839) );
  NOR2_X1 U11274 ( .A1(n13593), .A2(n19166), .ZN(n19160) );
  INV_X1 U11275 ( .A(n11220), .ZN(n11211) );
  AND2_X1 U11276 ( .A1(n9865), .A2(n9864), .ZN(n17858) );
  NAND2_X1 U11277 ( .A1(n10284), .A2(n10283), .ZN(n10841) );
  AOI21_X1 U11278 ( .B1(n10286), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10285), .ZN(n10842) );
  NOR2_X1 U11279 ( .A1(n9914), .A2(n9913), .ZN(n9912) );
  OAI221_X1 U11280 ( .B1(n15808), .B2(n15807), .C1(n15808), .C2(n15806), .A(
        n18902), .ZN(n17441) );
  CLKBUF_X1 U11281 ( .A(n10290), .Z(n10293) );
  NOR2_X1 U11282 ( .A1(n9916), .A2(n16320), .ZN(n9915) );
  OR2_X1 U11283 ( .A1(n10994), .A2(n10998), .ZN(n13667) );
  OR2_X1 U11284 ( .A1(n9803), .A2(n9802), .ZN(n9800) );
  NAND2_X1 U11285 ( .A1(n10615), .A2(n10690), .ZN(n10614) );
  OR2_X1 U11286 ( .A1(n11446), .A2(n11445), .ZN(n11447) );
  OR2_X1 U11287 ( .A1(n16114), .A2(n12738), .ZN(n19146) );
  NAND2_X1 U11288 ( .A1(n18725), .A2(n13488), .ZN(n18712) );
  AOI21_X1 U11289 ( .B1(n13609), .B2(n10993), .A(n10992), .ZN(n10998) );
  OAI21_X1 U11290 ( .B1(n10251), .B2(n10250), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10252) );
  NOR2_X1 U11291 ( .A1(n17896), .A2(n13210), .ZN(n13211) );
  AOI21_X1 U11292 ( .B1(n14249), .B2(n9921), .A(n9920), .ZN(n9919) );
  INV_X2 U11293 ( .A(n17524), .ZN(n17542) );
  AND3_X1 U11294 ( .A1(n10246), .A2(n10245), .A3(n10244), .ZN(n10253) );
  NAND2_X1 U11295 ( .A1(n13605), .A2(n10987), .ZN(n13609) );
  NAND2_X1 U11296 ( .A1(n17512), .A2(n14286), .ZN(n13489) );
  OR2_X1 U11297 ( .A1(n13352), .A2(n16578), .ZN(n14286) );
  OR2_X1 U11298 ( .A1(n11191), .A2(n19994), .ZN(n10245) );
  NOR2_X1 U11299 ( .A1(n17904), .A2(n13207), .ZN(n17898) );
  AND2_X1 U11300 ( .A1(n13601), .A2(n13600), .ZN(n13598) );
  AND3_X1 U11301 ( .A1(n11006), .A2(n11005), .A3(n11004), .ZN(n14053) );
  AND2_X1 U11302 ( .A1(n13333), .A2(n13351), .ZN(n9752) );
  NAND2_X1 U11303 ( .A1(n13338), .A2(n13349), .ZN(n16578) );
  NOR2_X1 U11304 ( .A1(n17906), .A2(n17905), .ZN(n17904) );
  NOR2_X1 U11305 ( .A1(n13336), .A2(n13339), .ZN(n13353) );
  OAI21_X1 U11306 ( .B1(n10261), .B2(n10242), .A(n10073), .ZN(n10243) );
  NOR2_X1 U11307 ( .A1(n13330), .A2(n15709), .ZN(n13336) );
  NAND2_X1 U11308 ( .A1(n15591), .A2(n9753), .ZN(n13351) );
  AND2_X1 U11309 ( .A1(n13329), .A2(n9668), .ZN(n13338) );
  AND4_X1 U11310 ( .A1(n11430), .A2(n13702), .A3(n11429), .A4(n11428), .ZN(
        n11434) );
  AND2_X4 U11311 ( .A1(n13448), .A2(n10963), .ZN(n11160) );
  INV_X1 U11312 ( .A(n12277), .ZN(n12287) );
  XNOR2_X1 U11313 ( .A(n13193), .B(n18227), .ZN(n17905) );
  NAND2_X1 U11314 ( .A1(n11411), .A2(n11410), .ZN(n14922) );
  OR2_X1 U11315 ( .A1(n11424), .A2(n11414), .ZN(n11415) );
  OR2_X1 U11316 ( .A1(n13331), .A2(n18296), .ZN(n9753) );
  AND3_X1 U11317 ( .A1(n10207), .A2(n10037), .A3(n10206), .ZN(n10217) );
  NOR2_X1 U11318 ( .A1(n17448), .A2(n10083), .ZN(n13208) );
  NOR2_X1 U11319 ( .A1(n12696), .A2(n18985), .ZN(n12698) );
  AND2_X1 U11320 ( .A1(n9930), .A2(n15558), .ZN(n13448) );
  NAND2_X1 U11321 ( .A1(n9749), .A2(n11579), .ZN(n12277) );
  NAND2_X1 U11322 ( .A1(n10157), .A2(n10220), .ZN(n10228) );
  XNOR2_X1 U11323 ( .A(n10083), .B(n17448), .ZN(n13193) );
  OR2_X2 U11324 ( .A1(n10493), .A2(n10492), .ZN(n15135) );
  INV_X1 U11325 ( .A(n17300), .ZN(n18285) );
  AND2_X1 U11326 ( .A1(n10751), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10760) );
  INV_X1 U11327 ( .A(n13350), .ZN(n18289) );
  NAND4_X1 U11328 ( .A1(n13305), .A2(n13304), .A3(n13303), .A4(n13302), .ZN(
        n13349) );
  OAI211_X1 U11329 ( .C1(n13194), .C2(n13168), .A(n13167), .B(n13166), .ZN(
        n17432) );
  INV_X1 U11330 ( .A(n10184), .ZN(n15543) );
  INV_X2 U11331 ( .A(n10205), .ZN(n10218) );
  OR2_X1 U11332 ( .A1(n10495), .A2(n10184), .ZN(n10771) );
  NAND3_X1 U11333 ( .A1(n9873), .A2(n9868), .A3(n13205), .ZN(n17926) );
  BUF_X2 U11334 ( .A(n10495), .Z(n14029) );
  AND3_X1 U11335 ( .A1(n13154), .A2(n13153), .A3(n13152), .ZN(n10083) );
  INV_X1 U11336 ( .A(n19364), .ZN(n10774) );
  OR2_X2 U11337 ( .A1(n10962), .A2(n16384), .ZN(n10497) );
  BUF_X4 U11338 ( .A(n10962), .Z(n19348) );
  NAND2_X1 U11339 ( .A1(n10170), .A2(n10169), .ZN(n10962) );
  AND4_X1 U11340 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11279) );
  NAND4_X1 U11341 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11376) );
  AND4_X1 U11342 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11335) );
  AND4_X1 U11343 ( .A1(n11327), .A2(n11326), .A3(n11325), .A4(n11324), .ZN(
        n11336) );
  AND2_X1 U11344 ( .A1(n10194), .A2(n10193), .ZN(n10195) );
  AND4_X1 U11345 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11281) );
  AND4_X1 U11346 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11374) );
  AND4_X1 U11347 ( .A1(n11383), .A2(n11382), .A3(n11381), .A4(n11380), .ZN(
        n11399) );
  AND4_X1 U11348 ( .A1(n11316), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(
        n11321) );
  CLKBUF_X1 U11349 ( .A(n12065), .Z(n12186) );
  NAND2_X1 U11350 ( .A1(n10343), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12882) );
  CLKBUF_X3 U11351 ( .A(n12887), .Z(n12991) );
  NAND2_X2 U11352 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19916), .ZN(n19924) );
  NAND2_X2 U11353 ( .A1(n18843), .A2(n18776), .ZN(n18826) );
  INV_X2 U11354 ( .A(n16563), .ZN(U215) );
  INV_X4 U11355 ( .A(n20244), .ZN(n20209) );
  INV_X4 U11356 ( .A(n17208), .ZN(n17253) );
  INV_X2 U11357 ( .A(n13098), .ZN(n17245) );
  NAND2_X2 U11358 ( .A1(n14282), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17250) );
  INV_X4 U11359 ( .A(n13131), .ZN(n17255) );
  INV_X2 U11360 ( .A(n17226), .ZN(n9639) );
  CLKBUF_X1 U11361 ( .A(n12170), .Z(n12242) );
  NAND2_X2 U11362 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13099), .ZN(
        n17229) );
  INV_X2 U11363 ( .A(n15640), .ZN(n9635) );
  INV_X2 U11364 ( .A(n20005), .ZN(n19916) );
  INV_X2 U11365 ( .A(n16567), .ZN(n16569) );
  NAND2_X1 U11366 ( .A1(n18879), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13105) );
  AND2_X1 U11367 ( .A1(n13752), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11248) );
  AND2_X1 U11368 ( .A1(n9996), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10327) );
  AND2_X2 U11369 ( .A1(n10098), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10121) );
  NAND3_X2 U11370 ( .A1(n18911), .A2(n18898), .A3(n18910), .ZN(n18229) );
  AND2_X1 U11371 ( .A1(n13752), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11246) );
  INV_X2 U11372 ( .A(n19217), .ZN(n9637) );
  NAND3_X1 U11373 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n16942), .ZN(n17058) );
  NOR2_X2 U11374 ( .A1(n11241), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13960) );
  OR3_X2 U11375 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18701), .ZN(n13156) );
  AND2_X1 U11376 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11254) );
  NOR2_X1 U11377 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10098) );
  INV_X1 U11378 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13752) );
  INV_X2 U11379 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16364) );
  INV_X1 U11380 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18873) );
  AND2_X1 U11381 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18722) );
  NAND2_X1 U11382 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18701) );
  AOI22_X1 U11383 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12212), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11364) );
  AND2_X4 U11384 ( .A1(n11247), .A2(n13954), .ZN(n9638) );
  OR2_X1 U11385 ( .A1(n13105), .A2(n9884), .ZN(n17208) );
  INV_X1 U11386 ( .A(n10121), .ZN(n10126) );
  NOR2_X2 U11387 ( .A1(n11377), .A2(n11376), .ZN(n11403) );
  OR2_X1 U11388 ( .A1(n13106), .A2(n13105), .ZN(n17226) );
  AND2_X2 U11390 ( .A1(n10062), .A2(n10061), .ZN(n9717) );
  XNOR2_X2 U11391 ( .A(n10254), .B(n10255), .ZN(n10294) );
  NOR4_X2 U11392 ( .A1(n17625), .A2(n17949), .A3(n17624), .A4(n17738), .ZN(
        n17592) );
  INV_X2 U11393 ( .A(n15640), .ZN(n9640) );
  OR2_X1 U11394 ( .A1(n13106), .A2(n13103), .ZN(n15640) );
  NOR2_X2 U11395 ( .A1(n15015), .A2(n15018), .ZN(n12939) );
  NOR2_X2 U11396 ( .A1(n14457), .A2(n14547), .ZN(n14444) );
  NOR2_X4 U11397 ( .A1(n13104), .A2(n18701), .ZN(n13141) );
  XNOR2_X1 U11398 ( .A(n10292), .B(n10295), .ZN(n13527) );
  OAI21_X2 U11399 ( .B1(n10293), .B2(n10291), .A(n10292), .ZN(n14166) );
  NOR2_X2 U11400 ( .A1(n15000), .A2(n15002), .ZN(n15001) );
  NOR2_X2 U11401 ( .A1(n15007), .A2(n12940), .ZN(n15000) );
  NOR2_X2 U11402 ( .A1(n13906), .A2(n13905), .ZN(n13907) );
  NOR2_X2 U11403 ( .A1(n13073), .A2(n13072), .ZN(n13418) );
  NOR2_X2 U11404 ( .A1(n14001), .A2(n14076), .ZN(n14075) );
  AND2_X4 U11406 ( .A1(n13945), .A2(n12782), .ZN(n14025) );
  NOR2_X4 U11407 ( .A1(n13892), .A2(n12781), .ZN(n13945) );
  AND2_X2 U11408 ( .A1(n14406), .A2(n9702), .ZN(n13471) );
  NOR2_X4 U11409 ( .A1(n14497), .A2(n14498), .ZN(n14406) );
  INV_X1 U11410 ( .A(n14367), .ZN(n9957) );
  BUF_X1 U11411 ( .A(n11367), .Z(n12148) );
  INV_X1 U11412 ( .A(n11662), .ZN(n11659) );
  NAND2_X1 U11413 ( .A1(n10497), .A2(n10729), .ZN(n10744) );
  INV_X1 U11414 ( .A(n10260), .ZN(n10830) );
  NOR2_X1 U11415 ( .A1(n19348), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10978) );
  OAI211_X1 U11416 ( .C1(n11448), .C2(n11241), .A(n11450), .B(n11449), .ZN(
        n11451) );
  NAND2_X1 U11417 ( .A1(n14445), .A2(n9691), .ZN(n14497) );
  NOR2_X1 U11419 ( .A1(n9907), .A2(n9904), .ZN(n9903) );
  INV_X1 U11420 ( .A(n12427), .ZN(n9906) );
  NOR2_X1 U11421 ( .A1(n9812), .A2(n10676), .ZN(n9811) );
  INV_X1 U11422 ( .A(n10684), .ZN(n9812) );
  NAND2_X1 U11423 ( .A1(n10827), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10260) );
  AND2_X1 U11424 ( .A1(n10059), .A2(n15037), .ZN(n10058) );
  OR2_X1 U11425 ( .A1(n9934), .A2(n15413), .ZN(n9933) );
  INV_X1 U11426 ( .A(n10228), .ZN(n11203) );
  NAND2_X1 U11427 ( .A1(n10695), .A2(n10694), .ZN(n10696) );
  INV_X1 U11428 ( .A(n15158), .ZN(n10695) );
  AND2_X1 U11429 ( .A1(n10587), .A2(n9689), .ZN(n10034) );
  INV_X1 U11430 ( .A(n9919), .ZN(n9916) );
  INV_X1 U11431 ( .A(n10830), .ZN(n10896) );
  NAND3_X1 U11432 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19938), .A3(n19788), 
        .ZN(n14017) );
  NAND3_X1 U11433 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18873), .ZN(n13100) );
  NOR3_X1 U11434 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n18879), .ZN(n13099) );
  NOR2_X1 U11435 ( .A1(n13215), .A2(n17858), .ZN(n13217) );
  AND2_X1 U11436 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13214), .ZN(
        n13215) );
  XOR2_X1 U11437 ( .A(n13191), .B(n17419), .Z(n13214) );
  AOI21_X1 U11438 ( .B1(n9876), .B2(n9878), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U11439 ( .A1(n13341), .A2(n13338), .ZN(n13488) );
  NAND2_X1 U11440 ( .A1(n20536), .A2(n9758), .ZN(n11598) );
  NAND2_X1 U11441 ( .A1(n10765), .A2(n10764), .ZN(n16389) );
  NAND2_X1 U11442 ( .A1(n10763), .A2(n13552), .ZN(n10764) );
  OR2_X1 U11443 ( .A1(n19977), .A2(n10740), .ZN(n10741) );
  NAND2_X1 U11444 ( .A1(n15135), .A2(n10967), .ZN(n9921) );
  AND2_X1 U11445 ( .A1(n15159), .A2(n10043), .ZN(n10826) );
  AND2_X1 U11446 ( .A1(n10044), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10043) );
  NAND2_X1 U11447 ( .A1(n14145), .A2(n16359), .ZN(n15473) );
  NAND2_X1 U11448 ( .A1(n15427), .A2(n11219), .ZN(n11235) );
  AOI22_X1 U11449 ( .A1(n18692), .A2(n15702), .B1(n18696), .B2(n18171), .ZN(
        n18740) );
  XNOR2_X1 U11450 ( .A(n13217), .B(n13216), .ZN(n17850) );
  NAND2_X1 U11451 ( .A1(n12577), .A2(n12576), .ZN(n12580) );
  AOI21_X1 U11452 ( .B1(n18988), .B2(n19338), .A(n15430), .ZN(n9779) );
  AND2_X2 U11453 ( .A1(n9946), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9845) );
  INV_X1 U11454 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9946) );
  AND2_X1 U11455 ( .A1(n12277), .A2(n12276), .ZN(n12296) );
  AND2_X1 U11456 ( .A1(n11401), .A2(n11541), .ZN(n10097) );
  OAI21_X1 U11457 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(n10265) );
  AND2_X1 U11458 ( .A1(n12284), .A2(n12261), .ZN(n12273) );
  AND2_X1 U11459 ( .A1(n14910), .A2(n11627), .ZN(n9846) );
  INV_X1 U11460 ( .A(n11628), .ZN(n11627) );
  NAND2_X1 U11461 ( .A1(n9888), .A2(n11417), .ZN(n11440) );
  INV_X1 U11462 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U11463 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11363) );
  NOR2_X1 U11464 ( .A1(n12270), .A2(n12271), .ZN(n12269) );
  NAND2_X1 U11465 ( .A1(n10097), .A2(n20290), .ZN(n11425) );
  NOR2_X1 U11466 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12890) );
  NOR2_X1 U11467 ( .A1(n10774), .A2(n10203), .ZN(n10157) );
  BUF_X1 U11468 ( .A(n10271), .Z(n10286) );
  NAND2_X1 U11469 ( .A1(n10183), .A2(n10182), .ZN(n10223) );
  NAND2_X1 U11470 ( .A1(n12444), .A2(n11404), .ZN(n12581) );
  NOR2_X1 U11471 ( .A1(n9693), .A2(n9953), .ZN(n9952) );
  INV_X1 U11472 ( .A(n9954), .ZN(n9953) );
  OR2_X1 U11473 ( .A1(n14922), .A2(n9758), .ZN(n12255) );
  INV_X1 U11474 ( .A(n12220), .ZN(n12259) );
  INV_X1 U11475 ( .A(n11602), .ZN(n12220) );
  NOR2_X1 U11476 ( .A1(n11541), .A2(n20780), .ZN(n11602) );
  NAND2_X1 U11477 ( .A1(n9760), .A2(n9727), .ZN(n14844) );
  INV_X1 U11478 ( .A(n15916), .ZN(n9760) );
  AND2_X1 U11479 ( .A1(n9854), .A2(n9853), .ZN(n9852) );
  INV_X1 U11480 ( .A(n14535), .ZN(n9853) );
  AND2_X1 U11481 ( .A1(n14543), .A2(n14447), .ZN(n9854) );
  OR2_X1 U11482 ( .A1(n14855), .A2(n12421), .ZN(n14739) );
  OR2_X1 U11483 ( .A1(n12424), .A2(n14724), .ZN(n14737) );
  NAND2_X1 U11484 ( .A1(n14235), .A2(n12412), .ZN(n12414) );
  INV_X1 U11485 ( .A(n12393), .ZN(n9896) );
  INV_X1 U11486 ( .A(n15952), .ZN(n9895) );
  INV_X1 U11487 ( .A(n15951), .ZN(n9898) );
  AND2_X1 U11488 ( .A1(n14071), .A2(n14005), .ZN(n9862) );
  INV_X1 U11489 ( .A(n11694), .ZN(n9847) );
  NAND2_X1 U11490 ( .A1(n12573), .A2(n12555), .ZN(n12534) );
  INV_X1 U11491 ( .A(n12534), .ZN(n12568) );
  NAND2_X1 U11492 ( .A1(n12462), .A2(n12573), .ZN(n12533) );
  NAND2_X1 U11493 ( .A1(n12584), .A2(n13573), .ZN(n12567) );
  AND2_X1 U11494 ( .A1(n11515), .A2(n11514), .ZN(n12351) );
  OR2_X1 U11495 ( .A1(n11472), .A2(n11471), .ZN(n11475) );
  OR2_X1 U11496 ( .A1(n11452), .A2(n11451), .ZN(n11453) );
  NAND2_X1 U11497 ( .A1(n20261), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11579) );
  NAND2_X1 U11498 ( .A1(n20290), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9749) );
  AOI21_X1 U11499 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20590), .A(
        n12269), .ZN(n12266) );
  AND3_X1 U11500 ( .A1(n11474), .A2(n11412), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12302) );
  NAND2_X1 U11501 ( .A1(n10762), .A2(n10761), .ZN(n10765) );
  AND2_X1 U11502 ( .A1(n10626), .A2(n15035), .ZN(n9809) );
  INV_X1 U11503 ( .A(n10643), .ZN(n9819) );
  NAND2_X1 U11504 ( .A1(n10609), .A2(n13948), .ZN(n10615) );
  INV_X1 U11505 ( .A(n10516), .ZN(n9816) );
  INV_X1 U11506 ( .A(n11143), .ZN(n12910) );
  INV_X1 U11507 ( .A(n11138), .ZN(n12912) );
  NAND2_X1 U11508 ( .A1(n12991), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U11509 ( .A1(n10735), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U11510 ( .A1(n12999), .A2(n10138), .ZN(n11137) );
  NAND2_X1 U11511 ( .A1(n12991), .A2(n10138), .ZN(n11143) );
  OR2_X1 U11512 ( .A1(n12888), .A2(n10138), .ZN(n11141) );
  NAND2_X1 U11513 ( .A1(n13419), .A2(n10138), .ZN(n11131) );
  NAND2_X1 U11514 ( .A1(n13431), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11133) );
  AND2_X1 U11515 ( .A1(n9929), .A2(n15095), .ZN(n9928) );
  INV_X1 U11516 ( .A(n15360), .ZN(n9929) );
  INV_X1 U11517 ( .A(n13779), .ZN(n12922) );
  NOR2_X1 U11518 ( .A1(n12826), .A2(n10060), .ZN(n10059) );
  INV_X1 U11519 ( .A(n12783), .ZN(n10060) );
  NAND2_X1 U11520 ( .A1(n12757), .A2(n15543), .ZN(n13031) );
  AND2_X1 U11521 ( .A1(n10003), .A2(n10002), .ZN(n10001) );
  INV_X1 U11522 ( .A(n10078), .ZN(n10002) );
  NOR2_X1 U11523 ( .A1(n14062), .A2(n10010), .ZN(n10009) );
  INV_X1 U11524 ( .A(n14026), .ZN(n10010) );
  NOR2_X1 U11525 ( .A1(n16284), .A2(n9985), .ZN(n9984) );
  INV_X1 U11526 ( .A(n15065), .ZN(n9911) );
  AND2_X1 U11527 ( .A1(n16165), .A2(n15135), .ZN(n10700) );
  NAND2_X1 U11528 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  INV_X1 U11529 ( .A(n14089), .ZN(n10008) );
  INV_X1 U11530 ( .A(n13898), .ZN(n9994) );
  AND2_X1 U11531 ( .A1(n13746), .A2(n13889), .ZN(n9995) );
  OR2_X1 U11532 ( .A1(n10816), .A2(n11013), .ZN(n10820) );
  INV_X1 U11533 ( .A(n13931), .ZN(n9926) );
  NAND2_X1 U11534 ( .A1(n10830), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10284) );
  INV_X1 U11535 ( .A(n10956), .ZN(n10909) );
  NAND2_X1 U11536 ( .A1(n16383), .A2(n9669), .ZN(n10024) );
  NAND2_X1 U11537 ( .A1(n10254), .A2(n10257), .ZN(n10258) );
  NAND2_X1 U11538 ( .A1(n10977), .A2(n10976), .ZN(n13601) );
  NAND2_X1 U11539 ( .A1(n10973), .A2(n10972), .ZN(n13600) );
  NAND2_X1 U11540 ( .A1(n12751), .A2(n19986), .ZN(n12770) );
  AND2_X1 U11541 ( .A1(n13085), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12768) );
  INV_X1 U11542 ( .A(n10320), .ZN(n10302) );
  AND2_X1 U11543 ( .A1(n9626), .A2(n17340), .ZN(n13329) );
  NOR2_X1 U11544 ( .A1(n16877), .A2(n9826), .ZN(n9824) );
  NOR2_X1 U11545 ( .A1(n17428), .A2(n13212), .ZN(n13192) );
  AND2_X1 U11546 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13209), .ZN(
        n13210) );
  NOR2_X1 U11547 ( .A1(n9671), .A2(n9877), .ZN(n9876) );
  NAND2_X1 U11548 ( .A1(n13137), .A2(n13136), .ZN(n9877) );
  AOI21_X1 U11549 ( .B1(n13171), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n13130), .ZN(n13136) );
  NAND4_X1 U11550 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13337) );
  NAND2_X1 U11551 ( .A1(n9789), .A2(n9788), .ZN(n9787) );
  NAND2_X1 U11552 ( .A1(n18735), .A2(n18736), .ZN(n9788) );
  NAND2_X1 U11553 ( .A1(n9786), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n9785) );
  INV_X1 U11554 ( .A(n18736), .ZN(n9786) );
  CLKBUF_X1 U11555 ( .A(n12581), .Z(n13575) );
  AND2_X1 U11556 ( .A1(n12502), .A2(n12501), .ZN(n15883) );
  OR2_X1 U11557 ( .A1(n15774), .A2(n13403), .ZN(n13727) );
  INV_X1 U11558 ( .A(n13944), .ZN(n11638) );
  INV_X1 U11559 ( .A(n20256), .ZN(n20257) );
  NAND2_X1 U11560 ( .A1(n12164), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12226) );
  NOR2_X1 U11561 ( .A1(n12012), .A2(n12011), .ZN(n12013) );
  NAND2_X1 U11562 ( .A1(n12013), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12076) );
  AND2_X1 U11563 ( .A1(n15774), .A2(n13407), .ZN(n13630) );
  AND2_X1 U11564 ( .A1(n14397), .A2(n9722), .ZN(n14330) );
  INV_X1 U11565 ( .A(n14329), .ZN(n9849) );
  NOR2_X1 U11566 ( .A1(n15969), .A2(n9740), .ZN(n12610) );
  NAND2_X1 U11567 ( .A1(n15916), .A2(n9902), .ZN(n9901) );
  AND2_X1 U11568 ( .A1(n15915), .A2(n9729), .ZN(n9902) );
  AND2_X1 U11569 ( .A1(n14522), .A2(n14521), .ZN(n14524) );
  NOR2_X1 U11570 ( .A1(n14556), .A2(n12519), .ZN(n14544) );
  OR2_X1 U11571 ( .A1(n14162), .A2(n14163), .ZN(n14216) );
  AND2_X1 U11572 ( .A1(n12599), .A2(n20253), .ZN(n16044) );
  XNOR2_X1 U11573 ( .A(n12355), .B(n12354), .ZN(n20196) );
  AOI21_X1 U11574 ( .B1(n12456), .B2(n12455), .A(n20010), .ZN(n12598) );
  INV_X1 U11575 ( .A(n9747), .ZN(n12455) );
  OAI21_X1 U11576 ( .B1(n15774), .B2(n12450), .A(n12454), .ZN(n9747) );
  CLKBUF_X1 U11577 ( .A(n13697), .Z(n13698) );
  OR2_X1 U11578 ( .A1(n20260), .A2(n20259), .ZN(n20373) );
  AND2_X1 U11579 ( .A1(n20421), .A2(n20595), .ZN(n20737) );
  AOI22_X2 U11580 ( .A1(n16106), .A2(n20931), .B1(n9758), .B2(n14930), .ZN(
        n20317) );
  OAI21_X1 U11581 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16100), .A(n12303), 
        .ZN(n12306) );
  NAND2_X1 U11582 ( .A1(n9733), .A2(n9732), .ZN(n12303) );
  OR2_X1 U11583 ( .A1(n12302), .A2(n12314), .ZN(n9732) );
  OR2_X1 U11584 ( .A1(n9735), .A2(n9734), .ZN(n9733) );
  AND2_X1 U11585 ( .A1(n10732), .A2(n10731), .ZN(n13514) );
  OR2_X1 U11586 ( .A1(n15134), .A2(n10703), .ZN(n10706) );
  NAND2_X1 U11587 ( .A1(n10690), .A2(n15132), .ZN(n10710) );
  NAND2_X1 U11588 ( .A1(n10674), .A2(n9713), .ZN(n10689) );
  NOR2_X1 U11589 ( .A1(n10689), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10693) );
  OR2_X1 U11590 ( .A1(n10599), .A2(n9930), .ZN(n10690) );
  AND2_X1 U11591 ( .A1(n15030), .A2(n15024), .ZN(n10003) );
  AND2_X1 U11592 ( .A1(n14272), .A2(n15038), .ZN(n15040) );
  INV_X1 U11593 ( .A(n11141), .ZN(n12915) );
  INV_X1 U11594 ( .A(n11131), .ZN(n12914) );
  INV_X1 U11595 ( .A(n11133), .ZN(n12916) );
  INV_X1 U11596 ( .A(n11137), .ZN(n12911) );
  INV_X1 U11597 ( .A(n11132), .ZN(n12931) );
  OR2_X1 U11598 ( .A1(n9659), .A2(n10050), .ZN(n10049) );
  INV_X1 U11599 ( .A(n10053), .ZN(n10050) );
  NAND2_X1 U11600 ( .A1(n15381), .A2(n9708), .ZN(n15088) );
  NAND2_X1 U11601 ( .A1(n9932), .A2(n15106), .ZN(n9931) );
  INV_X1 U11602 ( .A(n9933), .ZN(n9932) );
  AND3_X1 U11603 ( .A1(n11067), .A2(n11066), .A3(n11065), .ZN(n16311) );
  NOR2_X1 U11604 ( .A1(n13510), .A2(n19348), .ZN(n13521) );
  NAND2_X1 U11605 ( .A1(n12693), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12696) );
  NOR2_X1 U11606 ( .A1(n12692), .A2(n16256), .ZN(n12681) );
  NAND2_X1 U11607 ( .A1(n12682), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12692) );
  NOR2_X2 U11608 ( .A1(n12687), .A2(n15268), .ZN(n12689) );
  AND2_X1 U11609 ( .A1(n15331), .A2(n11232), .ZN(n15302) );
  INV_X1 U11610 ( .A(n15137), .ZN(n15136) );
  XNOR2_X1 U11611 ( .A(n9805), .B(n15323), .ZN(n15158) );
  NAND2_X1 U11612 ( .A1(n16155), .A2(n15135), .ZN(n9805) );
  OR2_X1 U11613 ( .A1(n10018), .A2(n15178), .ZN(n10015) );
  AOI21_X1 U11614 ( .B1(n10094), .B2(n10673), .A(n9688), .ZN(n10018) );
  NOR2_X1 U11615 ( .A1(n10017), .A2(n15178), .ZN(n10016) );
  INV_X1 U11616 ( .A(n10673), .ZN(n10017) );
  OAI21_X1 U11617 ( .B1(n15231), .B2(n9770), .A(n9768), .ZN(n15211) );
  AOI21_X1 U11618 ( .B1(n9771), .B2(n9769), .A(n9695), .ZN(n9768) );
  INV_X1 U11619 ( .A(n9771), .ZN(n9770) );
  OR2_X1 U11620 ( .A1(n15211), .A2(n15212), .ZN(n15215) );
  NAND2_X1 U11621 ( .A1(n15231), .A2(n9775), .ZN(n9772) );
  AOI211_X1 U11622 ( .C1(n15429), .C2(n10874), .A(n15443), .B(n15428), .ZN(
        n15730) );
  NAND2_X1 U11623 ( .A1(n15239), .A2(n10041), .ZN(n16249) );
  AND2_X1 U11624 ( .A1(n11128), .A2(n11127), .ZN(n16285) );
  NAND2_X1 U11625 ( .A1(n15474), .A2(n9937), .ZN(n15456) );
  NOR2_X1 U11626 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  INV_X1 U11627 ( .A(n15457), .ZN(n9938) );
  NOR2_X1 U11628 ( .A1(n15468), .A2(n10612), .ZN(n10023) );
  NAND2_X1 U11629 ( .A1(n15468), .A2(n10612), .ZN(n10022) );
  NAND2_X1 U11630 ( .A1(n10607), .A2(n10606), .ZN(n15467) );
  NAND2_X1 U11631 ( .A1(n10033), .A2(n10030), .ZN(n10607) );
  AND2_X1 U11632 ( .A1(n16276), .A2(n10031), .ZN(n10030) );
  NOR2_X1 U11633 ( .A1(n10032), .A2(n15250), .ZN(n10031) );
  INV_X1 U11634 ( .A(n10595), .ZN(n10032) );
  AND2_X1 U11635 ( .A1(n10605), .A2(n15493), .ZN(n15250) );
  INV_X1 U11636 ( .A(n16340), .ZN(n9920) );
  NOR2_X1 U11637 ( .A1(n14254), .A2(n14248), .ZN(n16334) );
  NAND2_X1 U11638 ( .A1(n14245), .A2(n10815), .ZN(n14264) );
  AND2_X1 U11639 ( .A1(n13930), .A2(n13928), .ZN(n14145) );
  NOR2_X1 U11640 ( .A1(n19947), .A2(n19970), .ZN(n19400) );
  NOR2_X1 U11641 ( .A1(n14104), .A2(n19970), .ZN(n19682) );
  NAND2_X1 U11642 ( .A1(n19947), .A2(n19970), .ZN(n19599) );
  NOR2_X2 U11643 ( .A1(n19166), .A2(n14017), .ZN(n19362) );
  OR2_X1 U11644 ( .A1(n16404), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14013) );
  INV_X1 U11645 ( .A(n19788), .ZN(n19601) );
  NOR2_X1 U11646 ( .A1(n16617), .A2(n9829), .ZN(n16608) );
  OAI21_X1 U11647 ( .B1(n16630), .B2(n9834), .A(n9832), .ZN(n16617) );
  NAND2_X1 U11648 ( .A1(n9829), .A2(n9833), .ZN(n9832) );
  OR2_X1 U11649 ( .A1(n17563), .A2(n16619), .ZN(n9834) );
  INV_X1 U11650 ( .A(n16619), .ZN(n9833) );
  NOR2_X1 U11651 ( .A1(n16630), .A2(n17563), .ZN(n16629) );
  NOR2_X1 U11652 ( .A1(n16596), .A2(n9829), .ZN(n16639) );
  INV_X1 U11653 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17218) );
  OR2_X1 U11654 ( .A1(n9629), .A2(n13159), .ZN(n13160) );
  NOR2_X1 U11655 ( .A1(n15640), .A2(n13147), .ZN(n13148) );
  NOR2_X1 U11656 ( .A1(n15594), .A2(n15593), .ZN(n15805) );
  OR2_X1 U11657 ( .A1(n13204), .A2(n9875), .ZN(n9874) );
  NOR2_X1 U11658 ( .A1(n9629), .A2(n21110), .ZN(n9875) );
  NOR2_X1 U11659 ( .A1(n13360), .A2(n17923), .ZN(n16426) );
  NOR2_X1 U11660 ( .A1(n17419), .A2(n13191), .ZN(n16466) );
  NOR2_X1 U11661 ( .A1(n17629), .A2(n17986), .ZN(n9764) );
  INV_X1 U11662 ( .A(n17615), .ZN(n9765) );
  AND2_X1 U11663 ( .A1(n13219), .A2(n21117), .ZN(n9879) );
  AOI211_X1 U11664 ( .C1(n13244), .C2(n13243), .A(n13348), .B(n13345), .ZN(
        n18692) );
  INV_X1 U11665 ( .A(n17859), .ZN(n9864) );
  XNOR2_X1 U11666 ( .A(n13211), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9762) );
  NAND2_X1 U11667 ( .A1(n9762), .A2(n17883), .ZN(n17882) );
  NOR2_X1 U11668 ( .A1(n17925), .A2(n17918), .ZN(n17917) );
  NOR2_X1 U11669 ( .A1(n15708), .A2(n14285), .ZN(n18171) );
  NAND2_X1 U11670 ( .A1(n17926), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17925) );
  INV_X1 U11671 ( .A(n18732), .ZN(n18742) );
  NAND2_X1 U11672 ( .A1(n12656), .A2(n12655), .ZN(n20092) );
  AOI211_X1 U11673 ( .C1(P1_STATE2_REG_0__SCAN_IN), .C2(n15775), .A(n20209), 
        .B(n20935), .ZN(n12656) );
  AND2_X1 U11674 ( .A1(n12661), .A2(n12660), .ZN(n20099) );
  OR2_X1 U11675 ( .A1(n14366), .A2(n13472), .ZN(n13473) );
  NOR2_X2 U11676 ( .A1(n12336), .A2(n20256), .ZN(n14633) );
  NAND2_X1 U11677 ( .A1(n9667), .A2(n9746), .ZN(n9745) );
  INV_X1 U11678 ( .A(n12647), .ZN(n9746) );
  XNOR2_X1 U11679 ( .A(n13469), .B(n9686), .ZN(n14795) );
  INV_X1 U11680 ( .A(n16013), .ZN(n20242) );
  AND2_X1 U11681 ( .A1(n15774), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14930) );
  AOI21_X1 U11682 ( .B1(n9704), .B2(n16216), .A(n9962), .ZN(n9961) );
  INV_X1 U11683 ( .A(n16183), .ZN(n9962) );
  NAND2_X1 U11684 ( .A1(n16190), .A2(n16191), .ZN(n16189) );
  AND2_X1 U11685 ( .A1(n18920), .A2(n16397), .ZN(n19098) );
  NAND2_X1 U11686 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n9971), .ZN(n9970) );
  NOR2_X1 U11687 ( .A1(n14990), .A2(n9997), .ZN(n10961) );
  OR2_X1 U11688 ( .A1(n16125), .A2(n15042), .ZN(n13078) );
  INV_X1 U11689 ( .A(n19970), .ZN(n14110) );
  NAND2_X2 U11690 ( .A1(n13075), .A2(n19843), .ZN(n15042) );
  OAI21_X1 U11691 ( .B1(n13481), .B2(n19323), .A(n9993), .ZN(n9992) );
  NAND2_X1 U11692 ( .A1(n13480), .A2(n19290), .ZN(n9993) );
  AOI21_X1 U11693 ( .B1(n13092), .B2(n19290), .A(n13091), .ZN(n13093) );
  AND2_X1 U11694 ( .A1(n13084), .A2(n19997), .ZN(n19318) );
  AND2_X1 U11695 ( .A1(n12634), .A2(n10076), .ZN(n12635) );
  OR2_X1 U11696 ( .A1(n16125), .A2(n16341), .ZN(n12634) );
  OR2_X1 U11697 ( .A1(n15368), .A2(n11231), .ZN(n14311) );
  OR2_X1 U11698 ( .A1(n15431), .A2(n19330), .ZN(n9780) );
  NAND2_X1 U11699 ( .A1(n15730), .A2(n9782), .ZN(n9781) );
  OR2_X1 U11700 ( .A1(n16359), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9782) );
  AOI21_X1 U11701 ( .B1(n15231), .B2(n15232), .A(n15196), .ZN(n15224) );
  INV_X1 U11702 ( .A(n19330), .ZN(n16350) );
  CLKBUF_X1 U11703 ( .A(n10827), .Z(n10828) );
  INV_X1 U11704 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19973) );
  INV_X1 U11705 ( .A(n19532), .ZN(n19520) );
  AND2_X1 U11706 ( .A1(n12730), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19843) );
  NOR2_X1 U11707 ( .A1(n16672), .A2(n9829), .ZN(n16665) );
  INV_X1 U11708 ( .A(n16955), .ZN(n16954) );
  OAI211_X1 U11709 ( .C1(n17264), .C2(n13180), .A(n13179), .B(n13178), .ZN(
        n17422) );
  INV_X1 U11710 ( .A(n17437), .ZN(n17425) );
  NAND2_X1 U11711 ( .A1(n15811), .A2(n17340), .ZN(n17437) );
  INV_X1 U11712 ( .A(n17441), .ZN(n15811) );
  NAND2_X1 U11713 ( .A1(n13395), .A2(n17916), .ZN(n13396) );
  NOR2_X2 U11714 ( .A1(n17416), .A2(n17931), .ZN(n17829) );
  NAND2_X1 U11715 ( .A1(n9647), .A2(n9766), .ZN(n13232) );
  OR2_X1 U11716 ( .A1(n13238), .A2(n13239), .ZN(n13234) );
  NAND2_X1 U11717 ( .A1(n12264), .A2(n12263), .ZN(n12274) );
  AND2_X1 U11718 ( .A1(n20701), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12286) );
  CLKBUF_X1 U11719 ( .A(n11779), .Z(n12200) );
  NAND2_X1 U11720 ( .A1(n9908), .A2(n12427), .ZN(n9907) );
  INV_X1 U11721 ( .A(n12413), .ZN(n9904) );
  OR2_X1 U11722 ( .A1(n11656), .A2(n11655), .ZN(n12388) );
  NOR2_X1 U11723 ( .A1(n11435), .A2(n9758), .ZN(n9757) );
  OAI211_X1 U11724 ( .C1(n12238), .C2(n11257), .A(n11256), .B(n11255), .ZN(
        n11258) );
  INV_X1 U11725 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11485) );
  OR2_X1 U11726 ( .A1(n12182), .A2(n11312), .ZN(n11316) );
  OAI22_X1 U11727 ( .A1(n12300), .A2(n12299), .B1(n12310), .B2(n12375), .ZN(
        n9738) );
  NOR2_X1 U11728 ( .A1(n9818), .A2(n10583), .ZN(n9817) );
  INV_X1 U11729 ( .A(n10519), .ZN(n9818) );
  OR2_X1 U11730 ( .A1(n18984), .A2(n11013), .ZN(n10662) );
  OR2_X1 U11731 ( .A1(n10956), .A2(n13921), .ZN(n10280) );
  AOI22_X1 U11732 ( .A1(n13762), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19987), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U11733 ( .A1(n10830), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10270) );
  OR2_X1 U11734 ( .A1(n10350), .A2(n10349), .ZN(n10968) );
  AOI22_X1 U11735 ( .A1(n10173), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13433), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10102) );
  OR2_X1 U11736 ( .A1(n13329), .A2(n13337), .ZN(n13333) );
  INV_X1 U11737 ( .A(n13328), .ZN(n13334) );
  NOR3_X1 U11738 ( .A1(n18700), .A2(n13326), .A3(n13349), .ZN(n13330) );
  NAND2_X1 U11739 ( .A1(n9793), .A2(n9792), .ZN(n9791) );
  OR2_X1 U11740 ( .A1(n18733), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n9793) );
  AOI21_X1 U11741 ( .B1(n18718), .B2(n18732), .A(n18717), .ZN(n9792) );
  NAND2_X1 U11742 ( .A1(n18733), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n9790) );
  AND2_X1 U11743 ( .A1(n14393), .A2(n12105), .ZN(n9958) );
  NOR2_X1 U11744 ( .A1(n11971), .A2(n9955), .ZN(n9954) );
  NAND2_X1 U11745 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  AND2_X1 U11746 ( .A1(n14859), .A2(n12417), .ZN(n12422) );
  AND2_X1 U11747 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11688), .ZN(
        n11701) );
  NOR2_X1 U11748 ( .A1(n11665), .A2(n11668), .ZN(n11688) );
  INV_X1 U11749 ( .A(n14370), .ZN(n9850) );
  AND2_X1 U11750 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  INV_X1 U11751 ( .A(n14505), .ZN(n9858) );
  NOR2_X1 U11752 ( .A1(n14514), .A2(n9860), .ZN(n9859) );
  INV_X1 U11753 ( .A(n14424), .ZN(n9860) );
  OR2_X1 U11754 ( .A1(n11687), .A2(n11686), .ZN(n12397) );
  AND2_X1 U11755 ( .A1(n13573), .A2(n12555), .ZN(n12553) );
  OAI21_X1 U11756 ( .B1(n12349), .B2(n13621), .A(n12348), .ZN(n12355) );
  INV_X1 U11757 ( .A(n9749), .ZN(n11531) );
  OR2_X1 U11758 ( .A1(n11530), .A2(n11529), .ZN(n12407) );
  AOI21_X1 U11759 ( .B1(n11431), .B2(n14922), .A(n11415), .ZN(n11418) );
  NAND2_X1 U11760 ( .A1(n11536), .A2(n11535), .ZN(n11564) );
  INV_X1 U11761 ( .A(n11550), .ZN(n11536) );
  OR2_X1 U11762 ( .A1(n11596), .A2(n11595), .ZN(n12378) );
  AOI22_X1 U11763 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11366) );
  AOI21_X1 U11764 ( .B1(n9739), .B2(n9737), .A(n9736), .ZN(n9735) );
  NOR2_X1 U11765 ( .A1(n12302), .A2(n12310), .ZN(n9736) );
  INV_X1 U11766 ( .A(n9738), .ZN(n9737) );
  OR2_X1 U11767 ( .A1(n12298), .A2(n12297), .ZN(n9739) );
  NOR2_X1 U11768 ( .A1(n12301), .A2(n12314), .ZN(n9734) );
  NAND2_X1 U11769 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12267), .ZN(
        n12314) );
  AND2_X1 U11770 ( .A1(n16100), .A2(n12266), .ZN(n12267) );
  AND2_X1 U11771 ( .A1(n19973), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10728) );
  AND2_X1 U11772 ( .A1(n10501), .A2(n10744), .ZN(n10717) );
  AND2_X1 U11773 ( .A1(n10724), .A2(n10723), .ZN(n10763) );
  AND2_X1 U11774 ( .A1(n9809), .A2(n10633), .ZN(n9806) );
  AND2_X1 U11775 ( .A1(n10632), .A2(n10633), .ZN(n10635) );
  OR2_X1 U11776 ( .A1(n10599), .A2(n10596), .ZN(n10598) );
  NOR2_X1 U11777 ( .A1(n9814), .A2(n9813), .ZN(n10593) );
  INV_X1 U11778 ( .A(n9817), .ZN(n9813) );
  OR2_X1 U11779 ( .A1(n10516), .A2(n9815), .ZN(n9814) );
  INV_X1 U11780 ( .A(n10520), .ZN(n9815) );
  MUX2_X1 U11781 ( .A(n10717), .B(P2_EBX_REG_2__SCAN_IN), .S(n9930), .Z(n10521) );
  OR2_X1 U11782 ( .A1(n14975), .A2(n10054), .ZN(n10053) );
  NOR2_X1 U11783 ( .A1(n10052), .A2(n10053), .ZN(n10051) );
  INV_X1 U11784 ( .A(n13033), .ZN(n10052) );
  INV_X1 U11785 ( .A(n13031), .ZN(n12983) );
  OR2_X1 U11786 ( .A1(n15728), .A2(n9935), .ZN(n9934) );
  INV_X1 U11787 ( .A(n14196), .ZN(n9935) );
  AND3_X1 U11788 ( .A1(n10578), .A2(n10577), .A3(n10576), .ZN(n10966) );
  NOR2_X1 U11789 ( .A1(n12705), .A2(n9979), .ZN(n9978) );
  NAND2_X1 U11790 ( .A1(n9999), .A2(n12632), .ZN(n9998) );
  INV_X1 U11791 ( .A(n14978), .ZN(n9999) );
  AND2_X1 U11792 ( .A1(n10045), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10044) );
  INV_X1 U11793 ( .A(n15139), .ZN(n10029) );
  NOR2_X1 U11794 ( .A1(n15288), .A2(n15323), .ZN(n10045) );
  INV_X1 U11795 ( .A(n14313), .ZN(n9927) );
  NOR2_X1 U11796 ( .A1(n9774), .A2(n15199), .ZN(n9771) );
  INV_X1 U11797 ( .A(n9775), .ZN(n9769) );
  NOR2_X1 U11798 ( .A1(n15223), .A2(n9776), .ZN(n9775) );
  INV_X1 U11799 ( .A(n15232), .ZN(n9776) );
  NAND2_X1 U11800 ( .A1(n10041), .A2(n11226), .ZN(n10039) );
  NOR2_X1 U11801 ( .A1(n10039), .A2(n15417), .ZN(n10038) );
  AND2_X1 U11802 ( .A1(n11213), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10041) );
  NAND2_X1 U11803 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  NAND2_X1 U11804 ( .A1(n9940), .A2(n15476), .ZN(n9939) );
  INV_X1 U11805 ( .A(n16297), .ZN(n9940) );
  NAND2_X1 U11806 ( .A1(n10518), .A2(n19114), .ZN(n10536) );
  NAND2_X1 U11807 ( .A1(n10391), .A2(n10390), .ZN(n10793) );
  INV_X1 U11808 ( .A(n10968), .ZN(n10794) );
  NOR2_X1 U11809 ( .A1(n10372), .A2(n10371), .ZN(n10982) );
  INV_X1 U11810 ( .A(n10184), .ZN(n9988) );
  INV_X1 U11811 ( .A(n10223), .ZN(n10226) );
  NOR2_X2 U11812 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10329) );
  NOR2_X1 U11813 ( .A1(n10217), .A2(n19996), .ZN(n10208) );
  AND2_X1 U11814 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12891) );
  NAND2_X1 U11815 ( .A1(n10298), .A2(n10310), .ZN(n19630) );
  AND2_X1 U11816 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10120) );
  NAND2_X1 U11817 ( .A1(n13419), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11138) );
  NOR2_X1 U11818 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18879), .ZN(
        n13343) );
  AOI22_X1 U11819 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14282), .B2(n9672), .ZN(n13257) );
  INV_X1 U11820 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21120) );
  INV_X1 U11821 ( .A(n16942), .ZN(n13103) );
  NAND2_X1 U11822 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18856), .ZN(
        n13106) );
  NOR2_X1 U11823 ( .A1(n14289), .A2(n14288), .ZN(n15593) );
  INV_X1 U11824 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17119) );
  AND2_X1 U11825 ( .A1(n17638), .A2(n9701), .ZN(n13359) );
  INV_X1 U11826 ( .A(n17575), .ZN(n9841) );
  INV_X1 U11827 ( .A(n17695), .ZN(n9838) );
  NOR2_X1 U11828 ( .A1(n17731), .A2(n9840), .ZN(n9839) );
  NOR2_X1 U11829 ( .A1(n17885), .A2(n9822), .ZN(n9821) );
  NOR2_X1 U11830 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NAND2_X1 U11831 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13249) );
  NAND2_X1 U11832 ( .A1(n13192), .A2(n17422), .ZN(n13191) );
  INV_X1 U11833 ( .A(n17937), .ZN(n9883) );
  AOI21_X1 U11834 ( .B1(n13239), .B2(n13238), .A(n13237), .ZN(n13348) );
  NOR2_X1 U11835 ( .A1(n18115), .A2(n18067), .ZN(n17760) );
  NOR2_X1 U11836 ( .A1(n13380), .A2(n17872), .ZN(n13382) );
  AND2_X1 U11837 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13379), .ZN(
        n13380) );
  NOR2_X1 U11838 ( .A1(n18281), .A2(n13350), .ZN(n18700) );
  NOR2_X1 U11839 ( .A1(n13106), .A2(n18701), .ZN(n13195) );
  NAND2_X1 U11840 ( .A1(n20261), .A2(n13621), .ZN(n14033) );
  OR2_X1 U11841 ( .A1(n14330), .A2(n12555), .ZN(n12577) );
  NAND2_X1 U11842 ( .A1(n14330), .A2(n13410), .ZN(n12576) );
  OR2_X1 U11843 ( .A1(n13869), .A2(n12446), .ZN(n12336) );
  OR2_X1 U11844 ( .A1(n12226), .A2(n14332), .ZN(n12645) );
  AND2_X1 U11845 ( .A1(n12163), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12164) );
  AND2_X1 U11846 ( .A1(n14678), .A2(n12654), .ZN(n12159) );
  NAND2_X1 U11847 ( .A1(n12131), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12162) );
  OR2_X1 U11848 ( .A1(n12083), .A2(n12082), .ZN(n14498) );
  AND2_X1 U11849 ( .A1(n12654), .A2(n15822), .ZN(n12049) );
  AND2_X1 U11850 ( .A1(n12015), .A2(n12014), .ZN(n14511) );
  AND2_X1 U11851 ( .A1(n11992), .A2(n11991), .ZN(n14512) );
  NOR2_X1 U11852 ( .A1(n11923), .A2(n14731), .ZN(n11924) );
  NAND2_X1 U11853 ( .A1(n11924), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11966) );
  CLKBUF_X1 U11854 ( .A(n14455), .Z(n14456) );
  NAND2_X1 U11855 ( .A1(n11829), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11830) );
  INV_X1 U11856 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21078) );
  NOR2_X1 U11857 ( .A1(n11813), .A2(n11793), .ZN(n11829) );
  INV_X1 U11858 ( .A(n9951), .ZN(n9950) );
  OAI21_X1 U11859 ( .B1(n9641), .B2(n9658), .A(n9714), .ZN(n9951) );
  AND2_X1 U11860 ( .A1(n11773), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11774) );
  NOR2_X1 U11861 ( .A1(n11768), .A2(n14179), .ZN(n11773) );
  NAND2_X1 U11862 ( .A1(n11730), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11768) );
  AND2_X1 U11863 ( .A1(n11701), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11730) );
  AOI21_X1 U11864 ( .B1(n12395), .B2(n11857), .A(n11708), .ZN(n14002) );
  OAI211_X1 U11865 ( .C1(n12220), .C2(n14069), .A(n11693), .B(n11692), .ZN(
        n14068) );
  INV_X1 U11866 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11668) );
  AOI21_X1 U11867 ( .B1(n12368), .B2(n11857), .A(n11637), .ZN(n13944) );
  NAND2_X1 U11868 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11599) );
  NOR2_X1 U11869 ( .A1(n11599), .A2(n14045), .ZN(n11633) );
  NAND2_X1 U11870 ( .A1(n13788), .A2(n11571), .ZN(n13876) );
  NAND2_X1 U11871 ( .A1(n13786), .A2(n13787), .ZN(n13785) );
  AND2_X1 U11872 ( .A1(n14397), .A2(n14400), .ZN(n14398) );
  NAND2_X1 U11873 ( .A1(n14397), .A2(n9707), .ZN(n14386) );
  AND2_X1 U11874 ( .A1(n12607), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9886) );
  AND2_X1 U11875 ( .A1(n14524), .A2(n9855), .ZN(n14499) );
  AND2_X1 U11876 ( .A1(n9857), .A2(n9856), .ZN(n9855) );
  INV_X1 U11877 ( .A(n14500), .ZN(n9856) );
  CLKBUF_X1 U11878 ( .A(n9887), .Z(n9885) );
  OR2_X1 U11879 ( .A1(n14709), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14691) );
  NAND2_X1 U11880 ( .A1(n14524), .A2(n9857), .ZN(n14507) );
  NAND2_X1 U11881 ( .A1(n14524), .A2(n9859), .ZN(n14517) );
  NAND2_X1 U11882 ( .A1(n14524), .A2(n14424), .ZN(n14515) );
  NAND2_X1 U11883 ( .A1(n14544), .A2(n9852), .ZN(n14538) );
  AND2_X1 U11884 ( .A1(n14544), .A2(n9720), .ZN(n14522) );
  INV_X1 U11885 ( .A(n14434), .ZN(n9851) );
  NOR2_X1 U11886 ( .A1(n14737), .A2(n15922), .ZN(n12425) );
  NAND2_X1 U11887 ( .A1(n14544), .A2(n9854), .ZN(n14536) );
  AND2_X1 U11888 ( .A1(n14544), .A2(n14543), .ZN(n14546) );
  OR2_X1 U11889 ( .A1(n12419), .A2(n12613), .ZN(n14859) );
  OR2_X1 U11890 ( .A1(n14476), .A2(n12511), .ZN(n14556) );
  AND3_X1 U11891 ( .A1(n12498), .A2(n12533), .A3(n12497), .ZN(n14217) );
  NOR2_X1 U11892 ( .A1(n14216), .A2(n14217), .ZN(n15884) );
  AOI21_X1 U11893 ( .B1(n15952), .B2(n9899), .A(n9898), .ZN(n9897) );
  INV_X1 U11894 ( .A(n12394), .ZN(n9899) );
  AND2_X1 U11895 ( .A1(n9862), .A2(n10084), .ZN(n9861) );
  NAND2_X1 U11896 ( .A1(n14070), .A2(n9862), .ZN(n14078) );
  NAND2_X1 U11897 ( .A1(n12481), .A2(n12480), .ZN(n16087) );
  INV_X1 U11898 ( .A(n13941), .ZN(n12480) );
  INV_X1 U11899 ( .A(n13942), .ZN(n12481) );
  INV_X1 U11900 ( .A(n12367), .ZN(n9891) );
  INV_X1 U11901 ( .A(n13910), .ZN(n9892) );
  NAND2_X1 U11902 ( .A1(n13855), .A2(n13886), .ZN(n13942) );
  NAND2_X1 U11903 ( .A1(n12598), .A2(n13706), .ZN(n20229) );
  OR2_X1 U11904 ( .A1(n20226), .A2(n20206), .ZN(n16013) );
  OR2_X1 U11905 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15798), .ZN(
        n20240) );
  NAND2_X1 U11906 ( .A1(n20196), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20195) );
  OAI21_X1 U11907 ( .B1(n12353), .B2(n12375), .A(n12352), .ZN(n13662) );
  CLKBUF_X1 U11908 ( .A(n12523), .Z(n12524) );
  INV_X1 U11909 ( .A(n20229), .ZN(n20206) );
  AND2_X1 U11910 ( .A1(n12598), .A2(n12593), .ZN(n14902) );
  XNOR2_X1 U11911 ( .A(n9761), .B(n11477), .ZN(n11538) );
  AND2_X1 U11912 ( .A1(n11378), .A2(n11408), .ZN(n13580) );
  INV_X1 U11913 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U11914 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20421), .ZN(n20289) );
  AND2_X1 U11915 ( .A1(n20338), .A2(n20339), .ZN(n20700) );
  INV_X1 U11916 ( .A(n20289), .ZN(n20306) );
  NOR2_X1 U11917 ( .A1(n13980), .A2(n14909), .ZN(n20732) );
  INV_X1 U11918 ( .A(n20372), .ZN(n20630) );
  AOI21_X1 U11919 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20701), .A(n20317), 
        .ZN(n20789) );
  AND2_X1 U11920 ( .A1(n12639), .A2(n12638), .ZN(n15759) );
  NOR2_X1 U11921 ( .A1(n11195), .A2(n11194), .ZN(n16385) );
  AND2_X1 U11922 ( .A1(n12712), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12713) );
  OR2_X1 U11923 ( .A1(n10706), .A2(n10705), .ZN(n10709) );
  NAND2_X1 U11924 ( .A1(n10710), .A2(n10698), .ZN(n15134) );
  NAND2_X1 U11925 ( .A1(n10674), .A2(n9811), .ZN(n10685) );
  NAND2_X1 U11926 ( .A1(n10632), .A2(n9807), .ZN(n10677) );
  AND2_X1 U11927 ( .A1(n9809), .A2(n9808), .ZN(n9807) );
  AND2_X1 U11928 ( .A1(n10633), .A2(n18942), .ZN(n9808) );
  NAND2_X1 U11929 ( .A1(n10635), .A2(n10626), .ZN(n10656) );
  AND2_X1 U11930 ( .A1(n10614), .A2(n9700), .ZN(n10651) );
  NAND2_X1 U11931 ( .A1(n10614), .A2(n9653), .ZN(n10646) );
  NAND2_X1 U11932 ( .A1(n10614), .A2(n10613), .ZN(n10644) );
  NOR2_X1 U11933 ( .A1(n10598), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10601) );
  AND2_X1 U11934 ( .A1(n10601), .A2(n13994), .ZN(n10609) );
  NAND2_X1 U11935 ( .A1(n10520), .A2(n10519), .ZN(n10533) );
  OR2_X1 U11936 ( .A1(n10516), .A2(n10533), .ZN(n10584) );
  INV_X1 U11937 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14953) );
  OR3_X1 U11938 ( .A1(n14969), .A2(n9998), .A3(n12742), .ZN(n9997) );
  OR2_X1 U11939 ( .A1(n11049), .A2(n11048), .ZN(n13896) );
  OAI211_X1 U11940 ( .C1(n10260), .C2(n16351), .A(n10253), .B(n10252), .ZN(
        n10290) );
  AND2_X1 U11941 ( .A1(n10248), .A2(n10249), .ZN(n10250) );
  NOR2_X1 U11942 ( .A1(n10777), .A2(n10497), .ZN(n10229) );
  NAND2_X1 U11943 ( .A1(n9910), .A2(n9909), .ZN(n15054) );
  INV_X1 U11944 ( .A(n15052), .ZN(n9909) );
  XNOR2_X1 U11945 ( .A(n12939), .B(n12963), .ZN(n15009) );
  NOR2_X1 U11946 ( .A1(n15009), .A2(n15008), .ZN(n15007) );
  NAND2_X1 U11947 ( .A1(n15381), .A2(n15095), .ZN(n15359) );
  CLKBUF_X1 U11948 ( .A(n15015), .Z(n15016) );
  AND2_X1 U11949 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  INV_X1 U11950 ( .A(n15028), .ZN(n10057) );
  AND2_X1 U11951 ( .A1(n11164), .A2(n11163), .ZN(n15413) );
  OR2_X1 U11952 ( .A1(n15729), .A2(n9934), .ZN(n15412) );
  INV_X1 U11953 ( .A(n19994), .ZN(n13552) );
  INV_X1 U11954 ( .A(n13458), .ZN(n19167) );
  OR2_X1 U11955 ( .A1(n12712), .A2(n9967), .ZN(n9965) );
  NAND2_X1 U11956 ( .A1(n9969), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9966) );
  NOR2_X1 U11957 ( .A1(n12710), .A2(n15143), .ZN(n12712) );
  NAND2_X1 U11958 ( .A1(n12703), .A2(n9977), .ZN(n12710) );
  AND2_X1 U11959 ( .A1(n9656), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9977) );
  OR2_X1 U11960 ( .A1(n14987), .A2(n14988), .ZN(n14990) );
  NAND2_X1 U11961 ( .A1(n12703), .A2(n9656), .ZN(n12708) );
  AND2_X1 U11962 ( .A1(n10917), .A2(n10916), .ZN(n14310) );
  NAND2_X1 U11963 ( .A1(n15040), .A2(n10000), .ZN(n15011) );
  AND2_X1 U11964 ( .A1(n10001), .A2(n15012), .ZN(n10000) );
  AND2_X1 U11965 ( .A1(n15040), .A2(n15030), .ZN(n15032) );
  NAND2_X1 U11966 ( .A1(n12698), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12699) );
  AND2_X1 U11967 ( .A1(n14229), .A2(n14228), .ZN(n14273) );
  AND3_X1 U11968 ( .A1(n10873), .A2(n10872), .A3(n10871), .ZN(n14089) );
  NOR2_X1 U11969 ( .A1(n14061), .A2(n10007), .ZN(n14185) );
  NAND2_X1 U11970 ( .A1(n10004), .A2(n10009), .ZN(n14088) );
  AND2_X1 U11971 ( .A1(n9652), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9983) );
  AND2_X1 U11972 ( .A1(n13745), .A2(n9676), .ZN(n13991) );
  NAND2_X1 U11973 ( .A1(n12689), .A2(n9652), .ZN(n12690) );
  AND2_X1 U11974 ( .A1(n12689), .A2(n9984), .ZN(n12691) );
  NAND2_X1 U11975 ( .A1(n12689), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U11976 ( .A1(n9973), .A2(n9646), .ZN(n12687) );
  NAND2_X1 U11977 ( .A1(n9973), .A2(n9974), .ZN(n12685) );
  NOR2_X1 U11978 ( .A1(n12684), .A2(n19301), .ZN(n12686) );
  OR2_X1 U11979 ( .A1(n14990), .A2(n14978), .ZN(n14980) );
  OR2_X1 U11980 ( .A1(n10701), .A2(n15322), .ZN(n15168) );
  CLKBUF_X1 U11981 ( .A(n14305), .Z(n15171) );
  CLKBUF_X1 U11982 ( .A(n15180), .Z(n15181) );
  CLKBUF_X1 U11983 ( .A(n15205), .Z(n15206) );
  NAND2_X1 U11984 ( .A1(n15444), .A2(n15445), .ZN(n15729) );
  NOR2_X1 U11985 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  INV_X1 U11986 ( .A(n14186), .ZN(n10006) );
  NOR2_X1 U11987 ( .A1(n14208), .A2(n14209), .ZN(n14229) );
  OR2_X1 U11988 ( .A1(n19007), .A2(n10665), .ZN(n15437) );
  NOR2_X1 U11989 ( .A1(n14061), .A2(n14062), .ZN(n14060) );
  NOR2_X1 U11990 ( .A1(n9939), .A2(n9936), .ZN(n15455) );
  INV_X1 U11991 ( .A(n15474), .ZN(n9936) );
  AND2_X1 U11992 ( .A1(n10860), .A2(n10859), .ZN(n13898) );
  INV_X1 U11993 ( .A(n15490), .ZN(n9913) );
  INV_X1 U11994 ( .A(n9915), .ZN(n9914) );
  CLKBUF_X1 U11995 ( .A(n15239), .Z(n15240) );
  OAI22_X1 U11996 ( .A1(n14264), .A2(n10047), .B1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n10046), .ZN(n15265) );
  NOR2_X1 U11997 ( .A1(n14265), .A2(n16337), .ZN(n10047) );
  INV_X1 U11998 ( .A(n14265), .ZN(n10046) );
  NAND2_X1 U11999 ( .A1(n13745), .A2(n9995), .ZN(n13897) );
  AND2_X1 U12000 ( .A1(n13688), .A2(n13739), .ZN(n13850) );
  NAND2_X1 U12001 ( .A1(n10812), .A2(n10074), .ZN(n10042) );
  NAND2_X1 U12002 ( .A1(n9925), .A2(n9924), .ZN(n9923) );
  INV_X1 U12003 ( .A(n14053), .ZN(n9924) );
  NAND2_X1 U12004 ( .A1(n10807), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14139) );
  NAND2_X1 U12005 ( .A1(n9777), .A2(n10831), .ZN(n14137) );
  INV_X1 U12006 ( .A(n10807), .ZN(n9777) );
  NAND2_X1 U12007 ( .A1(n9922), .A2(n9925), .ZN(n14054) );
  NAND2_X1 U12008 ( .A1(n10845), .A2(n10844), .ZN(n13741) );
  NAND2_X1 U12009 ( .A1(n10843), .A2(n10842), .ZN(n10844) );
  NOR2_X1 U12010 ( .A1(n13741), .A2(n13740), .ZN(n13739) );
  AND2_X1 U12011 ( .A1(n13676), .A2(n11223), .ZN(n13930) );
  NAND2_X1 U12012 ( .A1(n10790), .A2(n19843), .ZN(n11220) );
  OR3_X1 U12013 ( .A1(n13082), .A2(n10789), .A3(n10788), .ZN(n10790) );
  XNOR2_X1 U12014 ( .A(n13598), .B(n10981), .ZN(n13605) );
  AOI21_X1 U12015 ( .B1(n13527), .B2(n12768), .A(n12763), .ZN(n13861) );
  NAND2_X1 U12016 ( .A1(n10339), .A2(n10138), .ZN(n13779) );
  OR2_X1 U12017 ( .A1(n12779), .A2(n12759), .ZN(n12760) );
  AND2_X1 U12018 ( .A1(n12891), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10735) );
  NOR2_X1 U12019 ( .A1(n19947), .A2(n14110), .ZN(n19548) );
  AND2_X1 U12020 ( .A1(n19955), .A2(n19960), .ZN(n19723) );
  INV_X1 U12021 ( .A(n19723), .ZN(n15577) );
  INV_X1 U12022 ( .A(n19682), .ZN(n19569) );
  INV_X1 U12023 ( .A(n19363), .ZN(n19352) );
  NAND2_X1 U12024 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19788), .ZN(n19363) );
  AND2_X1 U12025 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19537) );
  INV_X1 U12026 ( .A(n19361), .ZN(n19366) );
  INV_X1 U12027 ( .A(n19362), .ZN(n19368) );
  NAND2_X1 U12028 ( .A1(n16389), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16404) );
  AND3_X1 U12029 ( .A1(n13774), .A2(n13773), .A3(n13772), .ZN(n16392) );
  NOR2_X1 U12030 ( .A1(n16639), .A2(n16640), .ZN(n16638) );
  NOR2_X1 U12031 ( .A1(n16685), .A2(n17653), .ZN(n16684) );
  NOR2_X1 U12032 ( .A1(n16703), .A2(n17681), .ZN(n16702) );
  NOR2_X1 U12033 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16843), .ZN(n16820) );
  INV_X2 U12034 ( .A(n17250), .ZN(n17236) );
  NAND2_X1 U12035 ( .A1(n18856), .A2(n18865), .ZN(n9884) );
  NAND2_X1 U12036 ( .A1(n18721), .A2(n9670), .ZN(n15806) );
  AOI21_X1 U12037 ( .B1(n14286), .B2(n18746), .A(n18891), .ZN(n17449) );
  NOR2_X1 U12038 ( .A1(n18750), .A2(n16576), .ZN(n17450) );
  NAND2_X1 U12039 ( .A1(n17638), .A2(n9654), .ZN(n17574) );
  NOR2_X1 U12040 ( .A1(n17995), .A2(n15711), .ZN(n17565) );
  NOR2_X1 U12041 ( .A1(n17611), .A2(n9843), .ZN(n9842) );
  NAND2_X1 U12042 ( .A1(n17638), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17610) );
  NAND2_X1 U12043 ( .A1(n9837), .A2(n9835), .ZN(n17648) );
  NOR2_X1 U12044 ( .A1(n9683), .A2(n9836), .ZN(n9835) );
  NOR2_X1 U12045 ( .A1(n17730), .A2(n9683), .ZN(n17678) );
  NAND2_X1 U12046 ( .A1(n9837), .A2(n9839), .ZN(n17694) );
  NOR2_X1 U12047 ( .A1(n17730), .A2(n17731), .ZN(n17716) );
  INV_X1 U12048 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17772) );
  INV_X1 U12049 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17773) );
  AOI21_X1 U12050 ( .B1(n17680), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18636), .ZN(n17769) );
  NOR2_X1 U12051 ( .A1(n16772), .A2(n16773), .ZN(n17800) );
  INV_X1 U12052 ( .A(n18115), .ZN(n17777) );
  NAND2_X1 U12053 ( .A1(n9825), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17857) );
  NOR2_X1 U12054 ( .A1(n17885), .A2(n9826), .ZN(n9825) );
  NAND2_X1 U12055 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17885) );
  INV_X1 U12056 ( .A(n13228), .ZN(n13229) );
  NAND2_X1 U12057 ( .A1(n15784), .A2(n17834), .ZN(n9766) );
  NAND2_X1 U12058 ( .A1(n15721), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15783) );
  NOR2_X1 U12059 ( .A1(n13226), .A2(n9882), .ZN(n9881) );
  INV_X1 U12060 ( .A(n17593), .ZN(n9767) );
  NOR2_X1 U12061 ( .A1(n9883), .A2(n17834), .ZN(n9882) );
  OAI211_X1 U12062 ( .C1(n17607), .C2(n17949), .A(n17606), .B(n9763), .ZN(
        n17594) );
  OR2_X1 U12063 ( .A1(n17834), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9763) );
  NAND2_X1 U12064 ( .A1(n13224), .A2(n10072), .ZN(n13225) );
  NAND2_X1 U12065 ( .A1(n17710), .A2(n17958), .ZN(n17629) );
  NOR2_X1 U12066 ( .A1(n17745), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17709) );
  NOR2_X1 U12067 ( .A1(n18285), .A2(n13349), .ZN(n15709) );
  INV_X1 U12068 ( .A(n18695), .ZN(n16576) );
  AND2_X1 U12069 ( .A1(n17746), .A2(n17811), .ZN(n17785) );
  INV_X1 U12070 ( .A(n18698), .ZN(n9801) );
  INV_X1 U12071 ( .A(n18699), .ZN(n9802) );
  NAND2_X1 U12072 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17833), .ZN(
        n18115) );
  NOR2_X1 U12073 ( .A1(n17841), .A2(n18160), .ZN(n17840) );
  NOR2_X1 U12074 ( .A1(n18155), .A2(n17862), .ZN(n17861) );
  NOR2_X1 U12075 ( .A1(n17874), .A2(n17873), .ZN(n17872) );
  NOR2_X2 U12076 ( .A1(n18912), .A2(n14288), .ZN(n18691) );
  NAND2_X1 U12077 ( .A1(n9876), .A2(n9870), .ZN(n9869) );
  INV_X1 U12078 ( .A(n9872), .ZN(n9871) );
  AND2_X1 U12079 ( .A1(n9878), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9870) );
  OR2_X1 U12080 ( .A1(n9803), .A2(n13488), .ZN(n18721) );
  INV_X1 U12081 ( .A(n18721), .ZN(n14287) );
  NOR2_X1 U12082 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18261), .ZN(n18547) );
  INV_X1 U12083 ( .A(n9626), .ZN(n18262) );
  NAND2_X1 U12084 ( .A1(n9784), .A2(n9783), .ZN(n18741) );
  AND2_X1 U12085 ( .A1(n18740), .A2(n9698), .ZN(n9783) );
  NAND2_X1 U12086 ( .A1(n9787), .A2(n9785), .ZN(n9784) );
  INV_X1 U12087 ( .A(n20935), .ZN(n14035) );
  OR2_X1 U12088 ( .A1(n12670), .A2(n12669), .ZN(n20071) );
  INV_X1 U12089 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14045) );
  AND2_X2 U12090 ( .A1(n13408), .A2(n13407), .ZN(n20116) );
  INV_X1 U12091 ( .A(n20112), .ZN(n14568) );
  OR2_X1 U12092 ( .A1(n12336), .A2(n20257), .ZN(n14628) );
  NAND2_X1 U12093 ( .A1(n14637), .A2(n13872), .ZN(n14645) );
  AND2_X1 U12094 ( .A1(n13630), .A2(n13629), .ZN(n20121) );
  BUF_X1 U12095 ( .A(n20120), .Z(n20141) );
  INV_X1 U12096 ( .A(n15846), .ZN(n15908) );
  AND2_X1 U12097 ( .A1(n16104), .A2(n20791), .ZN(n20189) );
  INV_X1 U12098 ( .A(n15913), .ZN(n20194) );
  INV_X1 U12099 ( .A(n20189), .ZN(n20258) );
  XNOR2_X1 U12100 ( .A(n14654), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14787) );
  NAND2_X1 U12101 ( .A1(n14653), .A2(n14652), .ZN(n14654) );
  OR2_X1 U12102 ( .A1(n14331), .A2(n14330), .ZN(n14791) );
  NAND2_X1 U12103 ( .A1(n9742), .A2(n9741), .ZN(n15969) );
  NAND2_X1 U12104 ( .A1(n16066), .A2(n12604), .ZN(n9741) );
  INV_X1 U12105 ( .A(n15983), .ZN(n9742) );
  AND2_X1 U12106 ( .A1(n16066), .A2(n9743), .ZN(n15983) );
  OR2_X1 U12107 ( .A1(n15988), .A2(n15797), .ZN(n9743) );
  AND2_X1 U12108 ( .A1(n12598), .A2(n15750), .ZN(n15798) );
  NAND2_X1 U12109 ( .A1(n9900), .A2(n12394), .ZN(n15954) );
  NAND2_X1 U12110 ( .A1(n15959), .A2(n12393), .ZN(n9900) );
  OR2_X1 U12111 ( .A1(n15798), .A2(n14902), .ZN(n20226) );
  AND2_X1 U12112 ( .A1(n20226), .A2(n20240), .ZN(n20222) );
  OR2_X1 U12113 ( .A1(n12641), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20244) );
  AND2_X1 U12114 ( .A1(n12598), .A2(n12583), .ZN(n20235) );
  INV_X1 U12115 ( .A(n20791), .ZN(n20782) );
  OAI21_X1 U12116 ( .B1(n14911), .B2(n20782), .A(n20666), .ZN(n20787) );
  OR3_X1 U12117 ( .A1(n13995), .A2(n15766), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n13979) );
  INV_X1 U12118 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16100) );
  OR2_X1 U12119 ( .A1(n20373), .A2(n20469), .ZN(n20413) );
  OAI21_X1 U12120 ( .B1(n10070), .B2(n20422), .A(n20737), .ZN(n20440) );
  INV_X1 U12121 ( .A(n20529), .ZN(n20558) );
  INV_X1 U12122 ( .A(n20796), .ZN(n20600) );
  INV_X1 U12123 ( .A(n20816), .ZN(n20614) );
  INV_X1 U12124 ( .A(n20822), .ZN(n20618) );
  INV_X1 U12125 ( .A(n20828), .ZN(n20622) );
  NAND2_X1 U12126 ( .A1(n20631), .A2(n20731), .ZN(n20648) );
  AND2_X1 U12127 ( .A1(n20732), .A2(n20661), .ZN(n20724) );
  INV_X1 U12128 ( .A(n20679), .ZN(n20802) );
  INV_X1 U12129 ( .A(n20686), .ZN(n21140) );
  AND2_X1 U12130 ( .A1(n20295), .A2(n20306), .ZN(n20816) );
  AND2_X1 U12131 ( .A1(n20732), .A2(n20731), .ZN(n20833) );
  AND2_X1 U12132 ( .A1(n11541), .A2(n20306), .ZN(n20828) );
  OAI21_X1 U12133 ( .B1(n12306), .B2(n12305), .A(n12304), .ZN(n9748) );
  OR2_X1 U12134 ( .A1(n12315), .A2(n12307), .ZN(n12308) );
  CLKBUF_X1 U12135 ( .A(n20893), .Z(n20928) );
  OR2_X1 U12136 ( .A1(n12727), .A2(n12728), .ZN(n13510) );
  NOR2_X1 U12137 ( .A1(n16383), .A2(n10497), .ZN(n19978) );
  NAND2_X1 U12138 ( .A1(n16128), .A2(n16129), .ZN(n16127) );
  NOR2_X1 U12139 ( .A1(n10710), .A2(n10688), .ZN(n16155) );
  NAND2_X1 U12140 ( .A1(n9960), .A2(n9959), .ZN(n16170) );
  AOI21_X1 U12141 ( .B1(n9961), .B2(n9963), .A(n9963), .ZN(n9959) );
  NAND2_X1 U12142 ( .A1(n18955), .A2(n9704), .ZN(n18947) );
  NAND2_X1 U12143 ( .A1(n18967), .A2(n9704), .ZN(n18956) );
  NAND2_X1 U12144 ( .A1(n18956), .A2(n18957), .ZN(n18955) );
  AND2_X1 U12145 ( .A1(n13521), .A2(n12729), .ZN(n19089) );
  NAND2_X1 U12146 ( .A1(n18968), .A2(n18969), .ZN(n18967) );
  NAND2_X1 U12147 ( .A1(n9704), .A2(n10071), .ZN(n18991) );
  OR2_X1 U12148 ( .A1(n14250), .A2(n14249), .ZN(n9918) );
  INV_X1 U12149 ( .A(n19098), .ZN(n19144) );
  INV_X1 U12150 ( .A(n19142), .ZN(n19130) );
  INV_X1 U12151 ( .A(n19139), .ZN(n19127) );
  NAND2_X1 U12152 ( .A1(n15040), .A2(n10003), .ZN(n15019) );
  OR2_X1 U12153 ( .A1(n11126), .A2(n11125), .ZN(n14086) );
  OR2_X1 U12154 ( .A1(n11096), .A2(n11095), .ZN(n14063) );
  OR2_X1 U12155 ( .A1(n11080), .A2(n11079), .ZN(n14064) );
  OR2_X1 U12156 ( .A1(n11064), .A2(n11063), .ZN(n13987) );
  AND2_X1 U12157 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10061) );
  CLKBUF_X1 U12158 ( .A(n13892), .Z(n13893) );
  NAND2_X1 U12159 ( .A1(n10062), .A2(n13734), .ZN(n13846) );
  INV_X1 U12160 ( .A(n19947), .ZN(n14104) );
  CLKBUF_X1 U12161 ( .A(n14983), .Z(n14986) );
  OR2_X1 U12162 ( .A1(n13766), .A2(n13444), .ZN(n13445) );
  NOR2_X1 U12163 ( .A1(n19191), .A2(n19206), .ZN(n19197) );
  INV_X1 U12164 ( .A(n19187), .ZN(n19205) );
  INV_X1 U12165 ( .A(n19210), .ZN(n19191) );
  INV_X1 U12166 ( .A(n19189), .ZN(n19214) );
  NOR2_X1 U12167 ( .A1(n16249), .A2(n15226), .ZN(n15426) );
  INV_X1 U12168 ( .A(n12681), .ZN(n12694) );
  INV_X1 U12169 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15268) );
  INV_X1 U12170 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19301) );
  CLKBUF_X1 U12171 ( .A(n12750), .Z(n14948) );
  AND2_X1 U12172 ( .A1(n19312), .A2(n19958), .ZN(n19319) );
  INV_X1 U12173 ( .A(n19323), .ZN(n16265) );
  INV_X1 U12174 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19311) );
  AND2_X1 U12175 ( .A1(n10064), .A2(n9680), .ZN(n9942) );
  XNOR2_X1 U12176 ( .A(n9804), .B(n15140), .ZN(n15299) );
  NAND2_X1 U12177 ( .A1(n15301), .A2(n9661), .ZN(n9804) );
  CLKBUF_X1 U12178 ( .A(n15159), .Z(n15160) );
  INV_X1 U12179 ( .A(n15316), .ZN(n15321) );
  AND2_X1 U12180 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  INV_X1 U12181 ( .A(n15350), .ZN(n10014) );
  NAND2_X1 U12182 ( .A1(n10012), .A2(n10015), .ZN(n15351) );
  AND2_X1 U12183 ( .A1(n11228), .A2(n15473), .ZN(n15368) );
  XOR2_X1 U12184 ( .A(n15201), .B(n15200), .Z(n15377) );
  NAND2_X1 U12185 ( .A1(n15215), .A2(n15210), .ZN(n15200) );
  NOR2_X1 U12186 ( .A1(n16287), .A2(n11214), .ZN(n15442) );
  XNOR2_X1 U12187 ( .A(n15191), .B(n9711), .ZN(n16259) );
  OR2_X1 U12188 ( .A1(n15467), .A2(n10023), .ZN(n10020) );
  AND2_X1 U12189 ( .A1(n10033), .A2(n10031), .ZN(n16274) );
  NAND2_X1 U12190 ( .A1(n10033), .A2(n10595), .ZN(n15252) );
  NAND2_X1 U12191 ( .A1(n9917), .A2(n9919), .ZN(n16319) );
  NOR3_X1 U12192 ( .A1(n16359), .A2(n20944), .A3(n13929), .ZN(n19336) );
  INV_X1 U12193 ( .A(n19343), .ZN(n16329) );
  INV_X1 U12194 ( .A(n19331), .ZN(n16344) );
  INV_X1 U12195 ( .A(n11235), .ZN(n16359) );
  NOR2_X1 U12196 ( .A1(n13597), .A2(n13596), .ZN(n19970) );
  INV_X1 U12197 ( .A(n19963), .ZN(n19960) );
  INV_X1 U12198 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19957) );
  CLKBUF_X1 U12200 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n15516) );
  XNOR2_X1 U12201 ( .A(n13861), .B(n13860), .ZN(n19963) );
  XNOR2_X1 U12202 ( .A(n13757), .B(n13756), .ZN(n19955) );
  INV_X1 U12203 ( .A(n13755), .ZN(n13756) );
  AND2_X1 U12204 ( .A1(n13694), .A2(n13693), .ZN(n19947) );
  OR2_X1 U12205 ( .A1(n13692), .A2(n13691), .ZN(n13694) );
  INV_X1 U12206 ( .A(n19480), .ZN(n19490) );
  OR3_X1 U12207 ( .A1(n15568), .A2(n19601), .A3(n15567), .ZN(n19533) );
  INV_X1 U12208 ( .A(n19598), .ZN(n19588) );
  OAI21_X1 U12209 ( .B1(n19593), .B2(n19572), .A(n19788), .ZN(n19595) );
  OAI21_X1 U12210 ( .B1(n19577), .B2(n19576), .A(n19575), .ZN(n19594) );
  NOR2_X1 U12211 ( .A1(n19569), .A2(n19600), .ZN(n19617) );
  INV_X1 U12212 ( .A(n19671), .ZN(n19677) );
  INV_X1 U12213 ( .A(n19749), .ZN(n19730) );
  INV_X1 U12214 ( .A(n19793), .ZN(n19695) );
  NOR2_X2 U12215 ( .A1(n19599), .A2(n15577), .ZN(n19771) );
  OAI21_X1 U12216 ( .B1(n15587), .B2(n15586), .A(n15585), .ZN(n19772) );
  NOR2_X1 U12217 ( .A1(n19569), .A2(n19543), .ZN(n19797) );
  INV_X1 U12218 ( .A(n19347), .ZN(n19796) );
  AND2_X1 U12219 ( .A1(n14029), .A2(n19352), .ZN(n19820) );
  INV_X1 U12220 ( .A(n19529), .ZN(n19828) );
  AND2_X1 U12221 ( .A1(n19537), .A2(n19719), .ZN(n19833) );
  NOR2_X2 U12222 ( .A1(n19599), .A2(n19543), .ZN(n19837) );
  INV_X1 U12223 ( .A(n19372), .ZN(n19832) );
  NOR2_X1 U12224 ( .A1(n18694), .A2(n17511), .ZN(n18913) );
  INV_X1 U12225 ( .A(n17450), .ZN(n17511) );
  NOR2_X1 U12226 ( .A1(n16629), .A2(n9829), .ZN(n16618) );
  OAI21_X1 U12227 ( .B1(n16652), .B2(n9710), .A(n9830), .ZN(n16596) );
  NAND2_X1 U12228 ( .A1(n9829), .A2(n9831), .ZN(n9830) );
  INV_X1 U12229 ( .A(n17591), .ZN(n9831) );
  NOR2_X1 U12230 ( .A1(n16651), .A2(n9829), .ZN(n13502) );
  NOR2_X1 U12231 ( .A1(n16652), .A2(n17603), .ZN(n16651) );
  OAI21_X1 U12232 ( .B1(n16685), .B2(n9712), .A(n9827), .ZN(n16672) );
  NAND2_X1 U12233 ( .A1(n9829), .A2(n9828), .ZN(n9827) );
  INV_X1 U12234 ( .A(n17632), .ZN(n9828) );
  NOR2_X1 U12235 ( .A1(n16684), .A2(n9829), .ZN(n16673) );
  NOR2_X1 U12236 ( .A1(n16692), .A2(n17671), .ZN(n16691) );
  NOR2_X1 U12237 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16763), .ZN(n16749) );
  INV_X1 U12238 ( .A(n16925), .ZN(n16948) );
  NOR2_X1 U12239 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16862), .ZN(n16847) );
  NAND4_X1 U12240 ( .A1(n18229), .A2(n18900), .A3(n18757), .A4(n18749), .ZN(
        n16958) );
  NOR2_X1 U12241 ( .A1(n21056), .A2(n17012), .ZN(n17017) );
  NOR2_X1 U12242 ( .A1(n16679), .A2(n17022), .ZN(n17028) );
  AND2_X1 U12243 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17285), .ZN(n17282) );
  AND2_X1 U12244 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17287), .ZN(n17285) );
  AOI22_X1 U12245 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n13171), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17245), .ZN(n13315) );
  AOI211_X1 U12246 ( .C1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .C2(n17244), .A(
        n13313), .B(n13312), .ZN(n13314) );
  INV_X1 U12247 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17291) );
  NOR4_X2 U12248 ( .A1(n18892), .A2(n9626), .A3(n15805), .A4(n18750), .ZN(
        n17298) );
  NOR2_X1 U12249 ( .A1(n17458), .A2(n17321), .ZN(n17315) );
  NAND2_X1 U12250 ( .A1(n17326), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17321) );
  NOR2_X1 U12251 ( .A1(n17330), .A2(n17462), .ZN(n17326) );
  NOR2_X1 U12252 ( .A1(n17336), .A2(n17340), .ZN(n17331) );
  NAND2_X1 U12253 ( .A1(n17331), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17330) );
  NOR4_X1 U12254 ( .A1(n17468), .A2(n17477), .A3(n17375), .A4(n17346), .ZN(
        n17337) );
  NOR2_X1 U12255 ( .A1(n17473), .A2(n17364), .ZN(n17358) );
  NAND2_X1 U12256 ( .A1(n17379), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17375) );
  NAND2_X1 U12257 ( .A1(n17385), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n17380) );
  NOR2_X1 U12258 ( .A1(n17380), .A2(n17560), .ZN(n17379) );
  NOR2_X1 U12259 ( .A1(n17441), .A2(n17384), .ZN(n17385) );
  AOI211_X1 U12260 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n13165), .B(n13164), .ZN(n13166) );
  AOI211_X1 U12261 ( .C1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .C2(n17254), .A(
        n13149), .B(n13148), .ZN(n13153) );
  NAND2_X1 U12262 ( .A1(n17425), .A2(n18708), .ZN(n17440) );
  NAND2_X1 U12263 ( .A1(n15809), .A2(n15811), .ZN(n17447) );
  NAND2_X1 U12264 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n9868) );
  NOR2_X1 U12265 ( .A1(n13203), .A2(n9874), .ZN(n9873) );
  INV_X1 U12266 ( .A(n17440), .ZN(n17442) );
  INV_X1 U12267 ( .A(n17447), .ZN(n17423) );
  AND2_X1 U12269 ( .A1(n17524), .A2(n18268), .ZN(n17557) );
  NOR2_X1 U12270 ( .A1(n17942), .A2(n16445), .ZN(n16437) );
  NOR2_X1 U12271 ( .A1(n17648), .A2(n17649), .ZN(n17638) );
  NOR2_X1 U12272 ( .A1(n17773), .A2(n17772), .ZN(n17771) );
  INV_X1 U12273 ( .A(n17829), .ZN(n17845) );
  INV_X1 U12274 ( .A(n17919), .ZN(n17910) );
  INV_X1 U12275 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18859) );
  INV_X1 U12276 ( .A(n17580), .ZN(n16463) );
  AND3_X1 U12277 ( .A1(n13220), .A2(n13222), .A3(n13219), .ZN(n17722) );
  NOR2_X1 U12278 ( .A1(n13354), .A2(n13355), .ZN(n18164) );
  INV_X1 U12279 ( .A(n18145), .ZN(n18168) );
  INV_X1 U12280 ( .A(n9880), .ZN(n17849) );
  INV_X1 U12281 ( .A(n9865), .ZN(n17860) );
  NAND2_X1 U12282 ( .A1(n17882), .A2(n13213), .ZN(n17870) );
  INV_X1 U12283 ( .A(n18250), .ZN(n18233) );
  INV_X1 U12284 ( .A(n18877), .ZN(n18880) );
  OR2_X1 U12285 ( .A1(n18748), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9796) );
  OR2_X1 U12286 ( .A1(n18751), .A2(n18750), .ZN(n9797) );
  INV_X1 U12287 ( .A(n16935), .ZN(n18757) );
  NAND2_X1 U12288 ( .A1(n18849), .A2(n9799), .ZN(n18753) );
  NAND2_X1 U12289 ( .A1(n18895), .A2(n18910), .ZN(n9799) );
  CLKBUF_X1 U12290 ( .A(n18836), .Z(n18830) );
  AND2_X1 U12291 ( .A1(n12334), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20256)
         );
  OAI21_X1 U12293 ( .B1(n12659), .B2(n20088), .A(n12677), .ZN(n12678) );
  NAND2_X1 U12294 ( .A1(n9755), .A2(n9754), .ZN(P1_U2970) );
  NAND2_X1 U12295 ( .A1(n9889), .A2(n9744), .ZN(P1_U3000) );
  NOR3_X1 U12296 ( .A1(n12620), .A2(n12619), .A3(n9745), .ZN(n9744) );
  NAND2_X1 U12297 ( .A1(n12717), .A2(n12716), .ZN(n12718) );
  OAI21_X1 U12298 ( .B1(n16190), .B2(n9963), .A(n9961), .ZN(n16181) );
  NAND2_X1 U12299 ( .A1(n13076), .A2(n10066), .ZN(n13080) );
  INV_X1 U12300 ( .A(n9992), .ZN(n9991) );
  INV_X1 U12301 ( .A(n13095), .ZN(n13096) );
  NOR2_X1 U12302 ( .A1(n12628), .A2(n12627), .ZN(n12637) );
  AND2_X1 U12303 ( .A1(n15295), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12627) );
  AOI21_X1 U12304 ( .B1(n9781), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n9778), .ZN(n15435) );
  NAND2_X1 U12305 ( .A1(n9780), .A2(n9779), .ZN(n9778) );
  OR2_X1 U12306 ( .A1(n16626), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9820) );
  AOI211_X1 U12307 ( .C1(n16613), .C2(n16935), .A(n16612), .B(n16611), .ZN(
        n16616) );
  OAI21_X1 U12308 ( .B1(n17301), .B2(P3_EAX_REG_31__SCAN_IN), .A(n9750), .ZN(
        P3_U2704) );
  OAI22_X1 U12309 ( .A1(n17306), .A2(n17425), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n17414), .ZN(n9751) );
  AOI21_X1 U12310 ( .B1(n16453), .B2(n17842), .A(n13398), .ZN(n13399) );
  NAND2_X1 U12311 ( .A1(n13397), .A2(n13396), .ZN(n13398) );
  OAI21_X1 U12312 ( .B1(n9798), .B2(n18898), .A(n9794), .ZN(P3_U2996) );
  AND2_X1 U12313 ( .A1(n9797), .A2(n9795), .ZN(n9794) );
  NOR2_X1 U12314 ( .A1(n18747), .A2(n18753), .ZN(n9798) );
  AND2_X1 U12315 ( .A1(n9796), .A2(n18749), .ZN(n9795) );
  AND2_X2 U12316 ( .A1(n9972), .A2(n9970), .ZN(n9704) );
  INV_X2 U12317 ( .A(n10186), .ZN(n12973) );
  INV_X2 U12318 ( .A(n10186), .ZN(n12999) );
  NOR2_X1 U12319 ( .A1(n12702), .A2(n16224), .ZN(n12703) );
  AND2_X1 U12320 ( .A1(n14212), .A2(n11778), .ZN(n9641) );
  INV_X1 U12321 ( .A(n11403), .ZN(n11412) );
  INV_X1 U12322 ( .A(n20261), .ZN(n11404) );
  NAND2_X2 U12323 ( .A1(n10181), .A2(n10180), .ZN(n16384) );
  INV_X1 U12324 ( .A(n16384), .ZN(n19996) );
  AND2_X1 U12325 ( .A1(n14159), .A2(n14212), .ZN(n9642) );
  AND2_X1 U12326 ( .A1(n14127), .A2(n12750), .ZN(n9643) );
  NAND2_X1 U12327 ( .A1(n18722), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14294) );
  INV_X1 U12328 ( .A(n14294), .ZN(n14282) );
  OR2_X1 U12329 ( .A1(n10040), .A2(n16286), .ZN(n9644) );
  NAND3_X1 U12330 ( .A1(n9996), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10186) );
  INV_X1 U12331 ( .A(n17869), .ZN(n9866) );
  AND2_X1 U12332 ( .A1(n13734), .A2(n9715), .ZN(n9645) );
  AND2_X1 U12333 ( .A1(n9696), .A2(n9974), .ZN(n9646) );
  AND2_X1 U12334 ( .A1(n15783), .A2(n9730), .ZN(n9647) );
  INV_X1 U12335 ( .A(n15239), .ZN(n10040) );
  AND2_X1 U12336 ( .A1(n13213), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9648) );
  INV_X1 U12337 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19104) );
  NAND2_X1 U12338 ( .A1(n9866), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9649) );
  NOR2_X1 U12339 ( .A1(n20536), .A2(n20265), .ZN(n9650) );
  INV_X1 U12340 ( .A(n12684), .ZN(n9973) );
  NAND2_X1 U12341 ( .A1(n14025), .A2(n10058), .ZN(n15027) );
  AND2_X1 U12342 ( .A1(n9917), .A2(n9915), .ZN(n15488) );
  AND2_X1 U12343 ( .A1(n12681), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12693) );
  AND2_X1 U12344 ( .A1(n9973), .A2(n9692), .ZN(n9651) );
  AND2_X1 U12345 ( .A1(n9984), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9652) );
  AND2_X1 U12346 ( .A1(n10613), .A2(n9819), .ZN(n9653) );
  AND2_X1 U12347 ( .A1(n9842), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9654) );
  AND2_X1 U12348 ( .A1(n10390), .A2(n9694), .ZN(n9655) );
  INV_X1 U12349 ( .A(n16884), .ZN(n13498) );
  INV_X2 U12350 ( .A(n12889), .ZN(n10343) );
  AND2_X1 U12351 ( .A1(n13850), .A2(n13849), .ZN(n13745) );
  NOR2_X1 U12352 ( .A1(n12699), .A2(n9981), .ZN(n12701) );
  AND2_X1 U12353 ( .A1(n9978), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9656) );
  OR2_X1 U12354 ( .A1(n13668), .A2(n10998), .ZN(n9657) );
  AND2_X1 U12355 ( .A1(n14212), .A2(n11792), .ZN(n9658) );
  AND2_X1 U12356 ( .A1(n13033), .A2(n14967), .ZN(n9659) );
  NAND2_X1 U12357 ( .A1(n12703), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12704) );
  INV_X1 U12358 ( .A(n13155), .ZN(n13194) );
  NOR2_X4 U12359 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13100), .ZN(
        n13155) );
  NAND2_X1 U12360 ( .A1(n14445), .A2(n14532), .ZN(n14430) );
  NAND2_X1 U12361 ( .A1(n15916), .A2(n15915), .ZN(n14714) );
  AND2_X1 U12362 ( .A1(n15045), .A2(n12630), .ZN(n12629) );
  AND2_X1 U12363 ( .A1(n14406), .A2(n12105), .ZN(n14391) );
  NAND2_X1 U12364 ( .A1(n14445), .A2(n9954), .ZN(n9956) );
  NAND2_X1 U12365 ( .A1(n12779), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9660) );
  OR2_X1 U12366 ( .A1(n15138), .A2(n15137), .ZN(n9661) );
  OR2_X1 U12367 ( .A1(n13217), .A2(n13216), .ZN(n9662) );
  AND2_X1 U12368 ( .A1(n9995), .A2(n9994), .ZN(n9663) );
  NOR2_X1 U12370 ( .A1(n10039), .A2(n10040), .ZN(n15227) );
  OAI21_X1 U12371 ( .B1(n15191), .B2(n10094), .A(n10673), .ZN(n15177) );
  NOR2_X1 U12372 ( .A1(n13103), .A2(n13104), .ZN(n13140) );
  INV_X1 U12373 ( .A(n13140), .ZN(n13126) );
  NAND2_X1 U12374 ( .A1(n14918), .A2(n11254), .ZN(n9664) );
  NAND2_X1 U12375 ( .A1(n9876), .A2(n9878), .ZN(n13363) );
  INV_X1 U12376 ( .A(n13363), .ZN(n17448) );
  NAND2_X1 U12377 ( .A1(n10020), .A2(n10022), .ZN(n15241) );
  AND2_X1 U12378 ( .A1(n13213), .A2(n9866), .ZN(n9665) );
  INV_X1 U12379 ( .A(n17340), .ZN(n18296) );
  OR3_X1 U12380 ( .A1(n13401), .A2(n13402), .A3(n9944), .ZN(n9666) );
  NAND2_X1 U12381 ( .A1(n10495), .A2(n10184), .ZN(n10770) );
  AND2_X1 U12382 ( .A1(n14406), .A2(n9958), .ZN(n14378) );
  OR2_X1 U12383 ( .A1(n12659), .A2(n20246), .ZN(n9667) );
  AND2_X1 U12384 ( .A1(n12760), .A2(n13736), .ZN(n13691) );
  AND3_X1 U12385 ( .A1(n13331), .A2(n18277), .A3(n18281), .ZN(n9668) );
  NAND2_X1 U12386 ( .A1(n10013), .A2(n10012), .ZN(n15349) );
  NOR2_X1 U12387 ( .A1(n14976), .A2(n14975), .ZN(n14974) );
  AND2_X1 U12388 ( .A1(n10218), .A2(n19997), .ZN(n9669) );
  OR2_X1 U12389 ( .A1(n17512), .A2(n18892), .ZN(n9670) );
  NAND4_X1 U12390 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        n9671) );
  NAND2_X1 U12391 ( .A1(n9949), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11448) );
  AND2_X1 U12392 ( .A1(n14445), .A2(n9952), .ZN(n14502) );
  AND2_X1 U12393 ( .A1(n18879), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n9672) );
  INV_X2 U12394 ( .A(n12419), .ZN(n15943) );
  AND2_X1 U12395 ( .A1(n10651), .A2(n10621), .ZN(n10632) );
  INV_X1 U12396 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15504) );
  NAND2_X1 U12397 ( .A1(n10632), .A2(n9806), .ZN(n9673) );
  AOI21_X1 U12398 ( .B1(n13327), .B2(n13329), .A(n13489), .ZN(n18725) );
  INV_X1 U12399 ( .A(n18725), .ZN(n9803) );
  NAND2_X1 U12400 ( .A1(n14159), .A2(n9641), .ZN(n14472) );
  AND2_X1 U12401 ( .A1(n13699), .A2(n12320), .ZN(n11438) );
  INV_X1 U12402 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18856) );
  AND2_X1 U12403 ( .A1(n14029), .A2(n19986), .ZN(n9674) );
  OR2_X1 U12404 ( .A1(n13334), .A2(n13331), .ZN(n9675) );
  AND2_X1 U12405 ( .A1(n9663), .A2(n13989), .ZN(n9676) );
  AND2_X1 U12406 ( .A1(n10220), .A2(n15558), .ZN(n9677) );
  AND2_X1 U12407 ( .A1(n9662), .A2(n18160), .ZN(n9678) );
  NAND2_X1 U12408 ( .A1(n11496), .A2(n11497), .ZN(n11500) );
  AND2_X1 U12409 ( .A1(n11405), .A2(n14340), .ZN(n9679) );
  OAI21_X1 U12410 ( .B1(n12416), .B2(n9906), .A(n15943), .ZN(n9905) );
  OR2_X1 U12411 ( .A1(n11238), .A2(n16341), .ZN(n9680) );
  AND2_X1 U12412 ( .A1(n13479), .A2(n13478), .ZN(n9681) );
  INV_X1 U12413 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9996) );
  INV_X1 U12414 ( .A(n11287), .ZN(n12018) );
  INV_X1 U12415 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U12416 ( .A1(n14025), .A2(n12783), .ZN(n14085) );
  NOR2_X1 U12417 ( .A1(n19301), .A2(n9975), .ZN(n9974) );
  NOR2_X1 U12418 ( .A1(n15456), .A2(n16285), .ZN(n15444) );
  AND2_X1 U12419 ( .A1(n14159), .A2(n9950), .ZN(n14474) );
  AND2_X1 U12420 ( .A1(n14025), .A2(n10056), .ZN(n15022) );
  AND2_X1 U12421 ( .A1(n14025), .A2(n10059), .ZN(n14276) );
  AND2_X1 U12422 ( .A1(n12689), .A2(n9983), .ZN(n12682) );
  AND2_X1 U12423 ( .A1(n15040), .A2(n10001), .ZN(n9682) );
  NAND2_X1 U12424 ( .A1(n9839), .A2(n9838), .ZN(n9683) );
  NOR2_X1 U12425 ( .A1(n15011), .A2(n14310), .ZN(n14309) );
  NOR2_X1 U12426 ( .A1(n15729), .A2(n15728), .ZN(n14195) );
  AND2_X1 U12427 ( .A1(n15381), .A2(n9928), .ZN(n9684) );
  NAND2_X1 U12428 ( .A1(n9893), .A2(n9897), .ZN(n14235) );
  AND2_X1 U12429 ( .A1(n9958), .A2(n14379), .ZN(n9685) );
  AND2_X1 U12430 ( .A1(n14650), .A2(n13468), .ZN(n9686) );
  NOR2_X1 U12431 ( .A1(n15729), .A2(n9931), .ZN(n15105) );
  AND2_X1 U12432 ( .A1(n14273), .A2(n14274), .ZN(n14272) );
  NAND2_X1 U12433 ( .A1(n13991), .A2(n13946), .ZN(n14061) );
  NOR2_X1 U12434 ( .A1(n15729), .A2(n9933), .ZN(n9687) );
  AND2_X1 U12435 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12683) );
  AND2_X1 U12436 ( .A1(n10679), .A2(n15357), .ZN(n9688) );
  AND2_X1 U12437 ( .A1(n15260), .A2(n15257), .ZN(n9689) );
  OR2_X1 U12438 ( .A1(n14029), .A2(n10620), .ZN(n9690) );
  AND2_X1 U12439 ( .A1(n9952), .A2(n14504), .ZN(n9691) );
  INV_X1 U12440 ( .A(n12581), .ZN(n9888) );
  AND2_X1 U12441 ( .A1(n9974), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9692) );
  NAND2_X1 U12442 ( .A1(n9911), .A2(n11177), .ZN(n15066) );
  INV_X1 U12443 ( .A(n15066), .ZN(n9910) );
  INV_X1 U12444 ( .A(n9774), .ZN(n9773) );
  OAI21_X1 U12445 ( .B1(n15223), .B2(n15195), .A(n15198), .ZN(n9774) );
  NAND2_X1 U12446 ( .A1(n14512), .A2(n14511), .ZN(n9693) );
  INV_X1 U12447 ( .A(n20275), .ZN(n13621) );
  AND2_X1 U12448 ( .A1(n11003), .A2(n10999), .ZN(n9694) );
  AND2_X1 U12449 ( .A1(n14499), .A2(n14415), .ZN(n14397) );
  NAND2_X1 U12450 ( .A1(n15405), .A2(n15392), .ZN(n9695) );
  AND2_X1 U12451 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9696) );
  AND2_X1 U12452 ( .A1(n15242), .A2(n10021), .ZN(n9697) );
  AND2_X1 U12453 ( .A1(n18739), .A2(n18738), .ZN(n9698) );
  AND2_X1 U12454 ( .A1(n10219), .A2(n11204), .ZN(n9699) );
  AND2_X1 U12455 ( .A1(n9653), .A2(n9690), .ZN(n9700) );
  AND2_X1 U12456 ( .A1(n9654), .A2(n9841), .ZN(n9701) );
  AND2_X1 U12457 ( .A1(n9685), .A2(n9957), .ZN(n9702) );
  AND2_X1 U12458 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9703) );
  INV_X1 U12459 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15244) );
  INV_X1 U12460 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11435) );
  INV_X1 U12461 ( .A(n13824), .ZN(n20151) );
  INV_X1 U12462 ( .A(n9704), .ZN(n9963) );
  NAND2_X1 U12463 ( .A1(n12727), .A2(n10767), .ZN(n11189) );
  INV_X1 U12464 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9836) );
  INV_X1 U12465 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U12466 ( .A1(n13693), .A2(n9660), .ZN(n10062) );
  AND2_X1 U12467 ( .A1(n10062), .A2(n9645), .ZN(n13744) );
  NOR2_X1 U12468 ( .A1(n16087), .A2(n16086), .ZN(n14070) );
  AND2_X1 U12469 ( .A1(n13745), .A2(n9663), .ZN(n9705) );
  NAND2_X1 U12470 ( .A1(n9917), .A2(n9912), .ZN(n15489) );
  NAND2_X1 U12471 ( .A1(n13745), .A2(n13746), .ZN(n9706) );
  AND2_X1 U12472 ( .A1(n14400), .A2(n14387), .ZN(n9707) );
  AND2_X1 U12473 ( .A1(n9928), .A2(n15086), .ZN(n9708) );
  AND2_X1 U12474 ( .A1(n13858), .A2(n13857), .ZN(n13855) );
  NAND2_X1 U12475 ( .A1(n9918), .A2(n9921), .ZN(n16339) );
  AND2_X1 U12476 ( .A1(n9707), .A2(n9850), .ZN(n9709) );
  INV_X1 U12477 ( .A(n11771), .ZN(n11857) );
  OR2_X1 U12478 ( .A1(n17591), .A2(n17603), .ZN(n9710) );
  AND2_X1 U12479 ( .A1(n15453), .A2(n15452), .ZN(n9711) );
  OR2_X1 U12480 ( .A1(n17632), .A2(n17653), .ZN(n9712) );
  NAND2_X1 U12481 ( .A1(n12701), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12702) );
  AND2_X1 U12482 ( .A1(n9811), .A2(n9810), .ZN(n9713) );
  AND2_X1 U12483 ( .A1(n14473), .A2(n14563), .ZN(n9714) );
  AND2_X1 U12484 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9715) );
  AND2_X1 U12485 ( .A1(n12703), .A2(n9978), .ZN(n9716) );
  NOR2_X1 U12486 ( .A1(n15489), .A2(n16311), .ZN(n15474) );
  OR3_X1 U12487 ( .A1(n12699), .A2(n9982), .A3(n18963), .ZN(n9718) );
  AND2_X1 U12488 ( .A1(n14070), .A2(n14071), .ZN(n9719) );
  NOR2_X1 U12489 ( .A1(n13667), .A2(n13666), .ZN(n13668) );
  INV_X1 U12490 ( .A(n13668), .ZN(n9922) );
  OR2_X1 U12491 ( .A1(n17850), .A2(n18154), .ZN(n9880) );
  AND2_X1 U12492 ( .A1(n9852), .A2(n9851), .ZN(n9720) );
  AND2_X1 U12493 ( .A1(n9708), .A2(n9927), .ZN(n9721) );
  AND2_X1 U12494 ( .A1(n9709), .A2(n9849), .ZN(n9722) );
  AND2_X1 U12495 ( .A1(n9665), .A2(n17882), .ZN(n9723) );
  AND2_X1 U12496 ( .A1(n9968), .A2(n9967), .ZN(n9724) );
  INV_X1 U12497 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9844) );
  INV_X1 U12498 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9843) );
  INV_X1 U12499 ( .A(n13573), .ZN(n12573) );
  AND2_X1 U12500 ( .A1(n11926), .A2(n11925), .ZN(n14532) );
  INV_X1 U12501 ( .A(n14532), .ZN(n9955) );
  INV_X1 U12502 ( .A(n14967), .ZN(n10054) );
  INV_X1 U12503 ( .A(n9969), .ZN(n9968) );
  NAND2_X1 U12504 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9969) );
  INV_X1 U12505 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9979) );
  INV_X1 U12506 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9967) );
  INV_X1 U12507 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9976) );
  INV_X1 U12508 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n9810) );
  INV_X1 U12509 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9971) );
  AND2_X1 U12510 ( .A1(n9823), .A2(n9824), .ZN(n9725) );
  NAND2_X1 U12511 ( .A1(n17800), .A2(n10067), .ZN(n17730) );
  INV_X1 U12512 ( .A(n17730), .ZN(n9837) );
  AND2_X1 U12513 ( .A1(n17638), .A2(n9842), .ZN(n9726) );
  AND2_X1 U12514 ( .A1(n14716), .A2(n15994), .ZN(n9727) );
  OR2_X1 U12515 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n12432), .ZN(
        n9728) );
  AND2_X1 U12516 ( .A1(n12616), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9729) );
  INV_X1 U12517 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21095) );
  INV_X1 U12518 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9867) );
  INV_X1 U12519 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U12520 ( .A1(n17887), .A2(n17885), .ZN(n9823) );
  OR2_X1 U12521 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16444), .ZN(
        n9730) );
  INV_X1 U12522 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9822) );
  INV_X1 U12523 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n9985) );
  INV_X1 U12524 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18910) );
  INV_X1 U12525 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9980) );
  INV_X1 U12526 ( .A(n15265), .ZN(n10819) );
  NOR2_X2 U12527 ( .A1(n18289), .A2(n17437), .ZN(n17374) );
  AOI22_X2 U12528 ( .A1(DATAI_17_), .A2(n9622), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n9623), .ZN(n20801) );
  AOI22_X2 U12529 ( .A1(DATAI_31_), .A2(n9622), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9623), .ZN(n20774) );
  AOI22_X2 U12530 ( .A1(DATAI_16_), .A2(n9622), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n9623), .ZN(n20795) );
  AOI22_X2 U12531 ( .A1(DATAI_18_), .A2(n9622), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n9623), .ZN(n20807) );
  AOI22_X2 U12532 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n9623), .B1(DATAI_21_), 
        .B2(n9622), .ZN(n20821) );
  AOI22_X2 U12533 ( .A1(DATAI_22_), .A2(n9622), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n9623), .ZN(n20827) );
  AOI22_X2 U12534 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9623), .B1(DATAI_27_), 
        .B2(n9622), .ZN(n20754) );
  NAND2_X1 U12535 ( .A1(n18547), .A2(n18604), .ZN(n18363) );
  AOI22_X2 U12536 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19361), .ZN(n19831) );
  NOR2_X2 U12537 ( .A1(n19167), .A2(n14017), .ZN(n19361) );
  AOI22_X1 U12538 ( .A1(n9751), .A2(P3_EAX_REG_31__SCAN_IN), .B1(n17374), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n9750) );
  AOI22_X2 U12539 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9623), .B1(DATAI_20_), 
        .B2(n9622), .ZN(n21149) );
  NOR2_X1 U12540 ( .A1(n19364), .A2(n19363), .ZN(n9731) );
  NAND2_X2 U12541 ( .A1(n10133), .A2(n10132), .ZN(n19364) );
  NOR2_X4 U12542 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14918) );
  AND2_X1 U12543 ( .A1(n14902), .A2(n12605), .ZN(n9740) );
  AND2_X2 U12544 ( .A1(n12308), .A2(n9748), .ZN(n15774) );
  OAI211_X1 U12545 ( .C1(n11579), .C2(n12341), .A(n11533), .B(n9749), .ZN(
        n11534) );
  NOR2_X1 U12546 ( .A1(n12404), .A2(n9749), .ZN(n12405) );
  OAI22_X1 U12547 ( .A1(n13697), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12360), 
        .B2(n9749), .ZN(n9761) );
  NOR2_X2 U12548 ( .A1(n17311), .A2(n17454), .ZN(n17306) );
  NAND3_X1 U12549 ( .A1(n9675), .A2(n13332), .A3(n9752), .ZN(n14284) );
  AND2_X1 U12550 ( .A1(n11422), .A2(n11402), .ZN(n11357) );
  NAND2_X1 U12551 ( .A1(n11400), .A2(n11422), .ZN(n11401) );
  AOI21_X2 U12552 ( .B1(n14651), .B2(n15943), .A(n12438), .ZN(n13469) );
  NAND2_X1 U12553 ( .A1(n9756), .A2(n11437), .ZN(n9759) );
  NAND2_X1 U12554 ( .A1(n9949), .A2(n9757), .ZN(n9756) );
  NAND2_X2 U12556 ( .A1(n14764), .A2(n12416), .ZN(n14723) );
  OR2_X2 U12557 ( .A1(n14772), .A2(n12415), .ZN(n14764) );
  NOR2_X2 U12558 ( .A1(n14709), .A2(n9728), .ZN(n14684) );
  OAI21_X2 U12559 ( .B1(n14844), .B2(n12430), .A(n15943), .ZN(n15896) );
  OAI21_X1 U12560 ( .B1(n17883), .B2(n9762), .A(n17882), .ZN(n18197) );
  AND2_X4 U12561 ( .A1(n15515), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13433) );
  XNOR2_X2 U12562 ( .A(n10475), .B(n10582), .ZN(n10807) );
  NAND2_X2 U12563 ( .A1(n15267), .A2(n10822), .ZN(n15239) );
  INV_X2 U12564 ( .A(n10962), .ZN(n19997) );
  NAND3_X1 U12565 ( .A1(n9791), .A2(n21095), .A3(n9790), .ZN(n9789) );
  INV_X2 U12566 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18865) );
  INV_X2 U12567 ( .A(n18723), .ZN(n17934) );
  NAND2_X2 U12568 ( .A1(n9801), .A2(n9800), .ZN(n18723) );
  NAND2_X1 U12569 ( .A1(n13342), .A2(n13341), .ZN(n18698) );
  NAND2_X1 U12570 ( .A1(n18723), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n18724) );
  NAND2_X1 U12571 ( .A1(n15148), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15301) );
  XNOR2_X1 U12572 ( .A(n15138), .B(n15136), .ZN(n15148) );
  NAND2_X1 U12573 ( .A1(n10674), .A2(n10675), .ZN(n10683) );
  NAND4_X1 U12574 ( .A1(n9816), .A2(n9817), .A3(n10520), .A4(n10591), .ZN(
        n10599) );
  MUX2_X1 U12575 ( .A(n10999), .B(n10719), .S(n10497), .Z(n10507) );
  MUX2_X1 U12576 ( .A(n11003), .B(n10720), .S(n10497), .Z(n10512) );
  MUX2_X1 U12577 ( .A(n10794), .B(n10752), .S(n10497), .Z(n10718) );
  NAND3_X1 U12578 ( .A1(n16616), .A2(n16615), .A3(n9820), .ZN(P3_U2641) );
  NAND3_X1 U12579 ( .A1(n9824), .A2(n9821), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16772) );
  CLKBUF_X1 U12580 ( .A(n16884), .Z(n9829) );
  AND2_X2 U12581 ( .A1(n9845), .A2(n11254), .ZN(n11340) );
  AND2_X2 U12582 ( .A1(n9845), .A2(n11249), .ZN(n11287) );
  AND2_X4 U12583 ( .A1(n13960), .A2(n9845), .ZN(n12170) );
  NAND3_X1 U12584 ( .A1(n11378), .A2(n11408), .A3(n13621), .ZN(n13699) );
  NAND2_X1 U12585 ( .A1(n12435), .A2(n14684), .ZN(n14651) );
  OAI211_X2 U12586 ( .C1(n12426), .C2(n14723), .A(n12425), .B(n12429), .ZN(
        n15916) );
  AND2_X4 U12587 ( .A1(n9848), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13957) );
  INV_X2 U12588 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U12589 ( .A1(n14397), .A2(n9709), .ZN(n14368) );
  NAND2_X1 U12590 ( .A1(n14070), .A2(n9861), .ZN(n14162) );
  OAI21_X1 U12591 ( .B1(n9648), .B2(n9665), .A(n17882), .ZN(n9863) );
  NAND2_X1 U12592 ( .A1(n9863), .A2(n9649), .ZN(n9865) );
  NAND2_X1 U12593 ( .A1(n9871), .A2(n9869), .ZN(n17918) );
  INV_X1 U12594 ( .A(n13129), .ZN(n9878) );
  NAND3_X1 U12595 ( .A1(n13220), .A2(n9879), .A3(n13222), .ZN(n17721) );
  NAND2_X1 U12596 ( .A1(n13225), .A2(n17676), .ZN(n17616) );
  NAND2_X1 U12597 ( .A1(n9880), .A2(n9678), .ZN(n17744) );
  NAND2_X1 U12598 ( .A1(n9887), .A2(n9886), .ZN(n14671) );
  AND2_X2 U12599 ( .A1(n9679), .A2(n9631), .ZN(n12444) );
  NAND2_X1 U12600 ( .A1(n12640), .A2(n20249), .ZN(n9889) );
  XNOR2_X1 U12601 ( .A(n12441), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12640) );
  NAND2_X1 U12602 ( .A1(n12367), .A2(n9892), .ZN(n9890) );
  NAND2_X1 U12603 ( .A1(n13909), .A2(n12367), .ZN(n20186) );
  NAND2_X1 U12604 ( .A1(n13911), .A2(n13910), .ZN(n13909) );
  NAND2_X1 U12605 ( .A1(n15959), .A2(n9894), .ZN(n9893) );
  NOR2_X1 U12606 ( .A1(n9895), .A2(n9896), .ZN(n9894) );
  NAND4_X4 U12607 ( .A1(n9848), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12184) );
  AND2_X2 U12608 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13707) );
  NAND2_X1 U12609 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11309) );
  AOI21_X1 U12610 ( .B1(n12414), .B2(n9903), .A(n9905), .ZN(n12428) );
  INV_X1 U12611 ( .A(n12415), .ZN(n9908) );
  NAND2_X2 U12612 ( .A1(n20315), .A2(n11478), .ZN(n14906) );
  NOR2_X2 U12613 ( .A1(n15054), .A2(n15046), .ZN(n15045) );
  NAND2_X1 U12614 ( .A1(n14250), .A2(n9921), .ZN(n9917) );
  NOR2_X2 U12615 ( .A1(n13668), .A2(n9923), .ZN(n14143) );
  NOR2_X1 U12616 ( .A1(n10998), .A2(n9926), .ZN(n9925) );
  MUX2_X1 U12617 ( .A(n10496), .B(n10982), .S(n14029), .Z(n10525) );
  NAND2_X1 U12618 ( .A1(n15474), .A2(n15476), .ZN(n15475) );
  NAND3_X1 U12619 ( .A1(n11240), .A2(n11237), .A3(n9941), .ZN(P2_U3015) );
  AND4_X2 U12620 ( .A1(n11337), .A2(n11358), .A3(n11427), .A4(n11359), .ZN(
        n11408) );
  NOR2_X1 U12621 ( .A1(n13401), .A2(n13402), .ZN(n9945) );
  NAND2_X1 U12622 ( .A1(n9666), .A2(n9943), .ZN(n12658) );
  OAI21_X1 U12623 ( .B1(n13401), .B2(n13402), .A(n9944), .ZN(n9943) );
  INV_X1 U12624 ( .A(n12260), .ZN(n9944) );
  CLKBUF_X1 U12625 ( .A(n9948), .Z(n9947) );
  NAND2_X2 U12626 ( .A1(n9948), .A2(n11402), .ZN(n13870) );
  NAND2_X1 U12627 ( .A1(n9947), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11771) );
  AOI21_X1 U12628 ( .B1(n12403), .B2(n9947), .A(n20261), .ZN(n11407) );
  AOI21_X1 U12629 ( .B1(n12353), .B2(n9947), .A(n20780), .ZN(n13659) );
  NAND2_X1 U12630 ( .A1(n11610), .A2(n14910), .ZN(n11629) );
  NAND4_X1 U12631 ( .A1(n11438), .A2(n11440), .A3(n12590), .A4(n11418), .ZN(
        n9949) );
  NAND2_X1 U12632 ( .A1(n9949), .A2(n9703), .ZN(n11421) );
  INV_X1 U12633 ( .A(n11448), .ZN(n11572) );
  INV_X1 U12634 ( .A(n9956), .ZN(n14420) );
  NAND2_X1 U12635 ( .A1(n14406), .A2(n9685), .ZN(n14365) );
  NAND2_X1 U12636 ( .A1(n16190), .A2(n9961), .ZN(n9960) );
  NAND2_X1 U12637 ( .A1(n16189), .A2(n9704), .ZN(n16182) );
  NAND2_X1 U12638 ( .A1(n12712), .A2(n9724), .ZN(n9964) );
  NAND3_X1 U12639 ( .A1(n9965), .A2(n9964), .A3(n9966), .ZN(n13480) );
  NAND4_X1 U12640 ( .A1(n9965), .A2(n9964), .A3(n9966), .A4(n13085), .ZN(n9972) );
  INV_X1 U12641 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9975) );
  NAND3_X1 U12642 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U12643 ( .A1(n12699), .A2(n18963), .ZN(n12700) );
  INV_X1 U12644 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9982) );
  NAND3_X1 U12645 ( .A1(n11208), .A2(n11206), .A3(n9986), .ZN(n14165) );
  AND2_X1 U12646 ( .A1(n11207), .A2(n9987), .ZN(n9986) );
  NAND2_X1 U12647 ( .A1(n10209), .A2(n10208), .ZN(n9987) );
  NAND2_X2 U12648 ( .A1(n9990), .A2(n9989), .ZN(n10184) );
  NAND2_X1 U12649 ( .A1(n10119), .A2(n10138), .ZN(n9989) );
  NAND2_X1 U12650 ( .A1(n10114), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9990) );
  NAND3_X1 U12651 ( .A1(n9681), .A2(n13482), .A3(n9991), .ZN(P2_U2983) );
  OR3_X1 U12652 ( .A1(n14990), .A2(n9998), .A3(n14969), .ZN(n12743) );
  NOR3_X1 U12653 ( .A1(n14990), .A2(n14978), .A3(n14969), .ZN(n14970) );
  INV_X1 U12654 ( .A(n14061), .ZN(n10004) );
  NAND2_X1 U12655 ( .A1(n10004), .A2(n10005), .ZN(n14208) );
  NAND2_X2 U12656 ( .A1(n10011), .A2(n10109), .ZN(n10495) );
  NAND2_X1 U12657 ( .A1(n10103), .A2(n10138), .ZN(n10011) );
  NAND2_X1 U12658 ( .A1(n15191), .A2(n10016), .ZN(n10012) );
  NAND2_X1 U12659 ( .A1(n15349), .A2(n10682), .ZN(n14303) );
  NAND2_X1 U12660 ( .A1(n15467), .A2(n10022), .ZN(n10019) );
  NAND2_X1 U12661 ( .A1(n10019), .A2(n9697), .ZN(n10619) );
  NAND2_X1 U12662 ( .A1(n10025), .A2(n10024), .ZN(n11191) );
  NAND2_X1 U12663 ( .A1(n10026), .A2(n10037), .ZN(n16383) );
  INV_X1 U12664 ( .A(n10782), .ZN(n10025) );
  AND2_X2 U12665 ( .A1(n10215), .A2(n10026), .ZN(n10782) );
  NOR2_X2 U12666 ( .A1(n10214), .A2(n10213), .ZN(n10026) );
  NAND2_X1 U12667 ( .A1(n10588), .A2(n10034), .ZN(n10033) );
  NAND2_X1 U12668 ( .A1(n10588), .A2(n10587), .ZN(n14267) );
  NAND2_X1 U12669 ( .A1(n10816), .A2(n10035), .ZN(n10806) );
  OR2_X1 U12670 ( .A1(n10036), .A2(n10808), .ZN(n10035) );
  NAND2_X1 U12671 ( .A1(n10036), .A2(n10808), .ZN(n10816) );
  INV_X1 U12672 ( .A(n10770), .ZN(n10037) );
  NAND2_X1 U12673 ( .A1(n15239), .A2(n10038), .ZN(n15205) );
  AND2_X1 U12674 ( .A1(n15159), .A2(n10045), .ZN(n12624) );
  NAND2_X1 U12675 ( .A1(n15159), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15141) );
  NAND2_X1 U12676 ( .A1(n15159), .A2(n10044), .ZN(n12625) );
  XNOR2_X1 U12677 ( .A(n10793), .B(n10999), .ZN(n13917) );
  OR2_X1 U12678 ( .A1(n13034), .A2(n10051), .ZN(n10048) );
  NAND2_X1 U12679 ( .A1(n13034), .A2(n13033), .ZN(n14966) );
  OR2_X1 U12680 ( .A1(n13034), .A2(n13033), .ZN(n10055) );
  NAND2_X1 U12681 ( .A1(n10048), .A2(n10049), .ZN(n13073) );
  NAND3_X1 U12682 ( .A1(n10219), .A2(n11204), .A3(n9677), .ZN(n10063) );
  NAND3_X1 U12683 ( .A1(n12727), .A2(n10767), .A3(n10063), .ZN(n13762) );
  NAND2_X1 U12684 ( .A1(n10782), .A2(n19996), .ZN(n12727) );
  NAND2_X1 U12685 ( .A1(n13870), .A2(n12342), .ZN(n11427) );
  AND2_X1 U12686 ( .A1(n12438), .A2(n12437), .ZN(n14649) );
  AOI22_X1 U12687 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11243) );
  CLKBUF_X1 U12688 ( .A(n15156), .Z(n15170) );
  INV_X1 U12689 ( .A(n13874), .ZN(n11639) );
  XNOR2_X1 U12690 ( .A(n12349), .B(n11564), .ZN(n20338) );
  NAND2_X1 U12691 ( .A1(n13471), .A2(n13472), .ZN(n13401) );
  NOR2_X1 U12692 ( .A1(n19364), .A2(n19363), .ZN(n19814) );
  AND2_X1 U12693 ( .A1(n10969), .A2(n19348), .ZN(n11202) );
  NAND2_X1 U12694 ( .A1(n10969), .A2(n11200), .ZN(n10183) );
  CLKBUF_X1 U12695 ( .A(n10782), .Z(n16398) );
  NAND2_X1 U12696 ( .A1(n10782), .A2(n10760), .ZN(n10261) );
  AND2_X1 U12697 ( .A1(n20275), .A2(n20306), .ZN(n20796) );
  NAND2_X1 U12698 ( .A1(n16116), .A2(n19319), .ZN(n13479) );
  NAND2_X1 U12699 ( .A1(n10840), .A2(n10839), .ZN(n10845) );
  BUF_X1 U12700 ( .A(n10255), .Z(n10256) );
  AND2_X1 U12701 ( .A1(n10770), .A2(n10218), .ZN(n10201) );
  NAND2_X1 U12702 ( .A1(n12658), .A2(n12324), .ZN(n12340) );
  NAND2_X1 U12703 ( .A1(n11501), .A2(n11500), .ZN(n11556) );
  AND3_X1 U12704 ( .A1(n10128), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10127), .ZN(n10129) );
  NAND2_X1 U12705 ( .A1(n10791), .A2(n10999), .ZN(n10792) );
  AND2_X1 U12706 ( .A1(n12671), .A2(n12670), .ZN(n20103) );
  OR2_X1 U12707 ( .A1(n11236), .A2(n9971), .ZN(n10064) );
  INV_X1 U12708 ( .A(n10264), .ZN(n10278) );
  NAND2_X1 U12709 ( .A1(n11209), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10264) );
  INV_X2 U12710 ( .A(n10959), .ZN(n10951) );
  AND2_X1 U12711 ( .A1(n14348), .A2(n15029), .ZN(n10066) );
  INV_X1 U12712 ( .A(n14557), .ZN(n20111) );
  NAND2_X1 U12713 ( .A1(n20116), .A2(n13412), .ZN(n14557) );
  AND2_X1 U12714 ( .A1(n13630), .A2(n15759), .ZN(n20200) );
  NOR2_X1 U12715 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12225) );
  INV_X1 U12716 ( .A(n14075), .ZN(n14157) );
  INV_X1 U12717 ( .A(n17916), .ZN(n17932) );
  NAND2_X2 U12718 ( .A1(n14637), .A2(n13871), .ZN(n14647) );
  AND2_X1 U12719 ( .A1(n17771), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10067) );
  NOR2_X1 U12720 ( .A1(n13227), .A2(n10091), .ZN(n10068) );
  AND2_X1 U12721 ( .A1(n12636), .A2(n12635), .ZN(n10069) );
  NOR2_X1 U12722 ( .A1(n20662), .A2(n20470), .ZN(n10070) );
  NAND2_X1 U12723 ( .A1(n17646), .A2(n17927), .ZN(n17715) );
  INV_X1 U12724 ( .A(n17715), .ZN(n17680) );
  OR2_X1 U12725 ( .A1(n18996), .A2(n12695), .ZN(n10071) );
  INV_X1 U12726 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10498) );
  OR3_X1 U12727 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17655), .ZN(n10072) );
  AND2_X1 U12728 ( .A1(n10241), .A2(n10240), .ZN(n10073) );
  AND2_X1 U12729 ( .A1(n10813), .A2(n14139), .ZN(n10074) );
  OR2_X1 U12730 ( .A1(n15124), .A2(n19305), .ZN(n10075) );
  NOR2_X1 U12731 ( .A1(n12633), .A2(n13089), .ZN(n10076) );
  NOR2_X1 U12732 ( .A1(n20662), .A2(n20632), .ZN(n10077) );
  AND2_X1 U12733 ( .A1(n10908), .A2(n10907), .ZN(n10078) );
  NAND2_X1 U12734 ( .A1(n13401), .A2(n13473), .ZN(n14328) );
  OR2_X1 U12735 ( .A1(n13126), .A2(n17225), .ZN(n10080) );
  AND3_X1 U12736 ( .A1(n10152), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10151), .ZN(n10081) );
  NOR2_X1 U12737 ( .A1(n15105), .A2(n15107), .ZN(n10082) );
  INV_X1 U12738 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14179) );
  INV_X1 U12739 ( .A(n13523), .ZN(n13542) );
  NAND3_X1 U12740 ( .A1(n12493), .A2(n12533), .A3(n12492), .ZN(n10084) );
  AND3_X1 U12741 ( .A1(n13248), .A2(n13247), .A3(n13246), .ZN(n10085) );
  INV_X1 U12742 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11793) );
  AND3_X1 U12743 ( .A1(n10123), .A2(n10122), .A3(n10138), .ZN(n10086) );
  BUF_X1 U12744 ( .A(n11794), .Z(n12210) );
  AND3_X1 U12745 ( .A1(n10177), .A2(n10176), .A3(n10138), .ZN(n10087) );
  AND3_X1 U12746 ( .A1(n10148), .A2(n10138), .A3(n10147), .ZN(n10088) );
  INV_X1 U12747 ( .A(n15044), .ZN(n15029) );
  AND3_X1 U12748 ( .A1(n10161), .A2(n10160), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10089) );
  INV_X1 U12749 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12440) );
  NOR2_X1 U12750 ( .A1(n18289), .A2(n18285), .ZN(n13331) );
  NAND3_X1 U12751 ( .A1(n11034), .A2(n11033), .A3(n11032), .ZN(n10090) );
  INV_X1 U12752 ( .A(n13195), .ZN(n16912) );
  INV_X1 U12753 ( .A(n14910), .ZN(n14909) );
  INV_X1 U12754 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12752) );
  AND2_X1 U12755 ( .A1(n17834), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10091) );
  INV_X2 U12756 ( .A(n15943), .ZN(n14862) );
  INV_X1 U12757 ( .A(n11204), .ZN(n10777) );
  AND3_X1 U12758 ( .A1(n10172), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10171), .ZN(n10092) );
  AND2_X1 U12759 ( .A1(n12963), .A2(n12962), .ZN(n10093) );
  OR2_X1 U12760 ( .A1(n10657), .A2(n15212), .ZN(n10094) );
  NOR2_X1 U12761 ( .A1(n10700), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15167) );
  OR2_X1 U12762 ( .A1(n13083), .A2(n19323), .ZN(n10095) );
  INV_X1 U12763 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19950) );
  NAND2_X1 U12764 ( .A1(n12750), .A2(n10289), .ZN(n10319) );
  INV_X1 U12765 ( .A(n11473), .ZN(n11474) );
  CLKBUF_X3 U12766 ( .A(n11367), .Z(n12240) );
  NAND2_X1 U12767 ( .A1(n14033), .A2(n12278), .ZN(n12295) );
  INV_X1 U12768 ( .A(n12442), .ZN(n11417) );
  NAND2_X1 U12769 ( .A1(n10228), .A2(n10204), .ZN(n10158) );
  OAI22_X1 U12770 ( .A1(n10540), .A2(n10353), .B1(n19692), .B2(n12803), .ZN(
        n10303) );
  AND2_X1 U12771 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10192) );
  INV_X1 U12772 ( .A(n12273), .ZN(n12264) );
  INV_X1 U12773 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11360) );
  AND2_X1 U12774 ( .A1(n12274), .A2(n12265), .ZN(n12270) );
  INV_X1 U12775 ( .A(n10265), .ZN(n10266) );
  AND2_X1 U12776 ( .A1(n10774), .A2(n10203), .ZN(n10182) );
  INV_X1 U12777 ( .A(n11454), .ZN(n12232) );
  OR2_X1 U12778 ( .A1(n11626), .A2(n11625), .ZN(n12377) );
  NAND2_X1 U12779 ( .A1(n11357), .A2(n11413), .ZN(n11358) );
  OAI21_X1 U12780 ( .B1(n10956), .B2(n10267), .A(n10266), .ZN(n10268) );
  INV_X1 U12781 ( .A(n10309), .ZN(n10310) );
  NAND2_X1 U12782 ( .A1(n13330), .A2(n9626), .ZN(n13332) );
  INV_X1 U12783 ( .A(n14526), .ZN(n11969) );
  BUF_X2 U12784 ( .A(n11466), .Z(n12234) );
  INV_X1 U12785 ( .A(n11270), .ZN(n12144) );
  INV_X1 U12786 ( .A(n14002), .ZN(n11709) );
  INV_X1 U12787 ( .A(n11695), .ZN(n11696) );
  NAND2_X1 U12788 ( .A1(n12566), .A2(n11426), .ZN(n12523) );
  AND4_X1 U12789 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n11261) );
  AND2_X1 U12790 ( .A1(n15017), .A2(n12963), .ZN(n12940) );
  OR2_X1 U12791 ( .A1(n13598), .A2(n10988), .ZN(n10993) );
  INV_X1 U12792 ( .A(n15167), .ZN(n10694) );
  AND2_X1 U12793 ( .A1(n10524), .A2(n10523), .ZN(n10747) );
  AOI22_X1 U12794 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10127) );
  INV_X1 U12795 ( .A(n10317), .ZN(n10305) );
  INV_X1 U12796 ( .A(n20295), .ZN(n14340) );
  INV_X1 U12797 ( .A(n14471), .ZN(n11778) );
  INV_X1 U12798 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12063) );
  INV_X1 U12799 ( .A(n14408), .ZN(n12105) );
  INV_X1 U12800 ( .A(n11475), .ZN(n12360) );
  INV_X1 U12801 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12431) );
  NAND2_X1 U12802 ( .A1(n11553), .A2(n11552), .ZN(n11554) );
  AND2_X1 U12803 ( .A1(n14064), .A2(n14063), .ZN(n12782) );
  AND2_X1 U12804 ( .A1(n19997), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12757) );
  OR2_X1 U12805 ( .A1(n13009), .A2(n13011), .ZN(n13032) );
  OR2_X1 U12806 ( .A1(n14278), .A2(n14193), .ZN(n12826) );
  AND2_X1 U12807 ( .A1(n19348), .A2(n19986), .ZN(n10963) );
  NAND2_X1 U12808 ( .A1(n10968), .A2(n10967), .ZN(n10973) );
  NAND2_X1 U12809 ( .A1(n9643), .A2(n10305), .ZN(n19776) );
  INV_X1 U12810 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17102) );
  INV_X1 U12811 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17101) );
  AND2_X1 U12812 ( .A1(n13344), .A2(n13343), .ZN(n13233) );
  NOR2_X1 U12813 ( .A1(n15592), .A2(n18268), .ZN(n13327) );
  AOI211_X1 U12814 ( .C1(n9640), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n13321), .B(n13320), .ZN(n13322) );
  INV_X1 U12815 ( .A(n12076), .ZN(n12077) );
  OR2_X1 U12816 ( .A1(n20033), .A2(n14100), .ZN(n14423) );
  OR2_X1 U12817 ( .A1(n20261), .A2(n14035), .ZN(n12669) );
  INV_X1 U12818 ( .A(n13790), .ZN(n11570) );
  AND2_X1 U12819 ( .A1(n20780), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12258) );
  NOR2_X1 U12820 ( .A1(n12130), .A2(n14696), .ZN(n12131) );
  NOR2_X1 U12821 ( .A1(n11966), .A2(n11927), .ZN(n11928) );
  AND2_X1 U12822 ( .A1(n11883), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11884) );
  AND3_X1 U12823 ( .A1(n11729), .A2(n11728), .A3(n11727), .ZN(n14076) );
  OAI21_X1 U12824 ( .B1(n13980), .B2(n11771), .A(n11545), .ZN(n11546) );
  OR2_X1 U12825 ( .A1(n14761), .A2(n12601), .ZN(n14741) );
  OR2_X1 U12826 ( .A1(n20229), .A2(n14869), .ZN(n14847) );
  NAND2_X1 U12827 ( .A1(n15884), .A2(n15883), .ZN(n14476) );
  INV_X1 U12828 ( .A(n12553), .ZN(n12564) );
  AND3_X1 U12829 ( .A1(n12479), .A2(n12533), .A3(n12478), .ZN(n13941) );
  NAND2_X1 U12830 ( .A1(n11578), .A2(n11577), .ZN(n20415) );
  INV_X1 U12831 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20537) );
  INV_X1 U12832 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20590) );
  INV_X1 U12833 ( .A(n12882), .ZN(n12921) );
  NOR2_X2 U12834 ( .A1(n15156), .A2(n10696), .ZN(n15131) );
  INV_X1 U12835 ( .A(n15135), .ZN(n11013) );
  INV_X1 U12836 ( .A(n15264), .ZN(n10818) );
  INV_X1 U12837 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14169) );
  NAND2_X1 U12838 ( .A1(n12775), .A2(n12774), .ZN(n12777) );
  NAND2_X1 U12839 ( .A1(n10298), .A2(n10305), .ZN(n14011) );
  INV_X1 U12840 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17122) );
  NOR2_X1 U12841 ( .A1(n17250), .A2(n17291), .ZN(n13130) );
  NAND2_X1 U12842 ( .A1(n17745), .A2(n18059), .ZN(n13219) );
  AOI21_X1 U12843 ( .B1(n18714), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13233), .ZN(n13239) );
  INV_X1 U12844 ( .A(n18064), .ZN(n18116) );
  INV_X1 U12845 ( .A(n13098), .ZN(n17215) );
  NOR2_X1 U12846 ( .A1(n13349), .A2(n13337), .ZN(n18699) );
  OAI211_X1 U12847 ( .C1(n17264), .C2(n21086), .A(n13285), .B(n13284), .ZN(
        n13350) );
  AND2_X1 U12848 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12077), .ZN(
        n12078) );
  INV_X1 U12849 ( .A(n20100), .ZN(n14486) );
  INV_X1 U12850 ( .A(n20071), .ZN(n20090) );
  INV_X1 U12851 ( .A(n20103), .ZN(n20034) );
  NAND2_X1 U12852 ( .A1(n11928), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12012) );
  NAND2_X1 U12853 ( .A1(n11884), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11923) );
  NOR2_X1 U12854 ( .A1(n21078), .A2(n11830), .ZN(n11883) );
  INV_X1 U12855 ( .A(n12403), .ZN(n12375) );
  INV_X1 U12856 ( .A(n15970), .ZN(n14836) );
  OR2_X1 U12857 ( .A1(n14847), .A2(n12613), .ZN(n12614) );
  INV_X1 U12858 ( .A(n20808), .ZN(n20607) );
  INV_X1 U12859 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20779) );
  INV_X1 U12860 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19986) );
  INV_X1 U12861 ( .A(n19089), .ZN(n19149) );
  OR2_X1 U12862 ( .A1(n12825), .A2(n14204), .ZN(n14193) );
  NAND2_X1 U12863 ( .A1(n19996), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19994) );
  INV_X1 U12864 ( .A(n15126), .ZN(n15127) );
  AND2_X1 U12865 ( .A1(n16123), .A2(n10708), .ZN(n15117) );
  NAND2_X1 U12866 ( .A1(n10681), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10682) );
  OR2_X1 U12867 ( .A1(n15418), .A2(n15417), .ZN(n15400) );
  AND2_X1 U12868 ( .A1(n11098), .A2(n11097), .ZN(n16297) );
  AND2_X1 U12869 ( .A1(n11036), .A2(n11035), .ZN(n16320) );
  OR2_X1 U12870 ( .A1(n19955), .A2(n19963), .ZN(n19600) );
  OR2_X1 U12871 ( .A1(n19955), .A2(n19960), .ZN(n19939) );
  INV_X1 U12872 ( .A(n19783), .ZN(n19543) );
  NOR2_X1 U12873 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16792), .ZN(n16770) );
  NOR2_X1 U12874 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16886), .ZN(n16871) );
  NAND2_X1 U12875 ( .A1(n18913), .A2(n18262), .ZN(n13503) );
  NAND2_X1 U12876 ( .A1(n10085), .A2(n13253), .ZN(n13254) );
  INV_X1 U12877 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17225) );
  INV_X1 U12878 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n21086) );
  INV_X1 U12879 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16877) );
  INV_X1 U12880 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17887) );
  INV_X1 U12881 ( .A(n17565), .ZN(n17942) );
  NAND2_X1 U12882 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17760), .ZN(
        n17759) );
  INV_X1 U12883 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n21110) );
  INV_X1 U12884 ( .A(n18691), .ZN(n18731) );
  INV_X1 U12885 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18714) );
  INV_X1 U12886 ( .A(n18272), .ZN(n18295) );
  NAND2_X1 U12887 ( .A1(n13620), .A2(n13525), .ZN(n20935) );
  NAND2_X1 U12888 ( .A1(n12078), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12130) );
  NOR2_X1 U12889 ( .A1(n14433), .A2(n14432), .ZN(n15888) );
  AND2_X1 U12890 ( .A1(n20092), .A2(n14044), .ZN(n15877) );
  AND2_X1 U12891 ( .A1(n20092), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20095) );
  AND2_X1 U12892 ( .A1(n20092), .A2(n12657), .ZN(n20052) );
  INV_X1 U12893 ( .A(n14542), .ZN(n20112) );
  INV_X1 U12894 ( .A(n14628), .ZN(n14625) );
  NAND2_X1 U12895 ( .A1(n12323), .A2(n13407), .ZN(n13869) );
  INV_X1 U12896 ( .A(n13795), .ZN(n20166) );
  INV_X2 U12897 ( .A(n13794), .ZN(n20181) );
  NAND2_X1 U12898 ( .A1(n11774), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11813) );
  NAND2_X1 U12899 ( .A1(n11633), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11665) );
  AND2_X1 U12900 ( .A1(n15913), .A2(n12643), .ZN(n20199) );
  AND2_X1 U12901 ( .A1(n16002), .A2(n12618), .ZN(n15970) );
  INV_X1 U12902 ( .A(n20230), .ZN(n20249) );
  INV_X1 U12903 ( .A(n20317), .ZN(n20421) );
  NOR2_X1 U12904 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16097) );
  OR2_X1 U12905 ( .A1(n20339), .A2(n20338), .ZN(n20469) );
  INV_X1 U12906 ( .A(n20423), .ZN(n20439) );
  NOR2_X1 U12907 ( .A1(n13980), .A2(n14910), .ZN(n20506) );
  INV_X1 U12908 ( .A(n20624), .ZN(n20582) );
  INV_X1 U12909 ( .A(n20414), .ZN(n20661) );
  INV_X1 U12910 ( .A(n20469), .ZN(n20731) );
  AND2_X1 U12911 ( .A1(n20260), .A2(n13980), .ZN(n20631) );
  OAI211_X1 U12912 ( .C1(n20767), .C2(n20738), .A(n20737), .B(n20736), .ZN(
        n20770) );
  INV_X1 U12913 ( .A(n20663), .ZN(n20783) );
  AND2_X1 U12914 ( .A1(n12342), .A2(n20306), .ZN(n20808) );
  AND2_X1 U12915 ( .A1(n11422), .A2(n20306), .ZN(n20822) );
  INV_X1 U12916 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20008) );
  NAND2_X1 U12917 ( .A1(n12745), .A2(n19151), .ZN(n12746) );
  NAND2_X1 U12918 ( .A1(n16149), .A2(n16150), .ZN(n16148) );
  NAND2_X1 U12919 ( .A1(n16170), .A2(n16171), .ZN(n16169) );
  NAND2_X1 U12920 ( .A1(n18947), .A2(n18948), .ZN(n18946) );
  OR2_X1 U12921 ( .A1(n18920), .A2(n12731), .ZN(n19142) );
  AND2_X1 U12922 ( .A1(n13521), .A2(n12744), .ZN(n19151) );
  AND3_X1 U12923 ( .A1(n11156), .A2(n11155), .A3(n11154), .ZN(n14204) );
  OR2_X1 U12924 ( .A1(n11111), .A2(n11110), .ZN(n14084) );
  NOR2_X1 U12925 ( .A1(n13593), .A2(n19167), .ZN(n19159) );
  AND2_X1 U12926 ( .A1(n19187), .A2(n13447), .ZN(n19206) );
  INV_X1 U12927 ( .A(n19287), .ZN(n13540) );
  INV_X1 U12928 ( .A(n13542), .ZN(n19285) );
  AND2_X1 U12929 ( .A1(n19312), .A2(n19314), .ZN(n19290) );
  AND2_X1 U12930 ( .A1(n16272), .A2(n16271), .ZN(n16316) );
  NAND2_X1 U12931 ( .A1(n10803), .A2(n10802), .ZN(n19294) );
  NAND2_X1 U12932 ( .A1(n14013), .A2(n14012), .ZN(n19788) );
  OAI21_X1 U12933 ( .B1(n15534), .B2(n15537), .A(n15533), .ZN(n19374) );
  NOR2_X2 U12934 ( .A1(n19600), .A2(n15530), .ZN(n19387) );
  INV_X1 U12935 ( .A(n19423), .ZN(n19426) );
  AND2_X1 U12936 ( .A1(n19400), .A2(n19430), .ZN(n19450) );
  OAI21_X1 U12937 ( .B1(n19473), .B2(n19472), .A(n19471), .ZN(n19491) );
  AND2_X1 U12938 ( .A1(n19400), .A2(n19723), .ZN(n19511) );
  NOR2_X2 U12939 ( .A1(n14111), .A2(n15577), .ZN(n19532) );
  NOR2_X1 U12940 ( .A1(n19541), .A2(n19540), .ZN(n19564) );
  AND2_X1 U12941 ( .A1(n19955), .A2(n19963), .ZN(n19783) );
  OAI21_X1 U12942 ( .B1(n19639), .B2(n19638), .A(n19788), .ZN(n19658) );
  INV_X1 U12943 ( .A(n19939), .ZN(n19430) );
  NOR2_X1 U12944 ( .A1(n19599), .A2(n19939), .ZN(n19707) );
  INV_X1 U12945 ( .A(n19842), .ZN(n19770) );
  INV_X1 U12946 ( .A(n15582), .ZN(n19781) );
  NAND2_X1 U12947 ( .A1(n18268), .A2(n9626), .ZN(n13352) );
  NOR2_X1 U12948 ( .A1(n14287), .A2(n13489), .ZN(n18694) );
  NOR2_X1 U12949 ( .A1(n18824), .A2(n16593), .ZN(n16637) );
  NOR2_X1 U12950 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16720), .ZN(n16704) );
  NOR2_X1 U12951 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16743), .ZN(n16728) );
  NOR2_X1 U12952 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16811), .ZN(n16797) );
  NOR2_X2 U12953 ( .A1(n18745), .A2(n13503), .ZN(n16925) );
  INV_X1 U12954 ( .A(n16944), .ZN(n16923) );
  NOR2_X1 U12955 ( .A1(n16696), .A2(n17056), .ZN(n17029) );
  NOR2_X1 U12956 ( .A1(n17113), .A2(n17086), .ZN(n17083) );
  INV_X1 U12957 ( .A(n17242), .ZN(n17202) );
  INV_X1 U12958 ( .A(n17298), .ZN(n17113) );
  OAI211_X2 U12959 ( .C1(n21077), .C2(n13194), .A(n13315), .B(n13314), .ZN(
        n17340) );
  NAND2_X1 U12960 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17315), .ZN(n17311) );
  NOR3_X1 U12961 ( .A1(n17340), .A2(n17477), .A3(n17375), .ZN(n17368) );
  INV_X1 U12962 ( .A(n17509), .ZN(n17451) );
  INV_X1 U12963 ( .A(n18065), .ZN(n17995) );
  NOR2_X1 U12964 ( .A1(n13392), .A2(n17840), .ZN(n18117) );
  INV_X1 U12965 ( .A(n17924), .ZN(n17868) );
  INV_X1 U12966 ( .A(n17834), .ZN(n17745) );
  INV_X1 U12967 ( .A(n18235), .ZN(n18242) );
  INV_X1 U12968 ( .A(n18547), .ZN(n18362) );
  NOR2_X1 U12969 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18850), .ZN(
        n18874) );
  INV_X1 U12970 ( .A(n18406), .ZN(n18399) );
  INV_X1 U12971 ( .A(n18429), .ZN(n18422) );
  INV_X1 U12972 ( .A(n18599), .ZN(n18589) );
  INV_X1 U12973 ( .A(n18629), .ZN(n18619) );
  NAND2_X1 U12974 ( .A1(n13630), .A2(n9888), .ZN(n13620) );
  INV_X1 U12975 ( .A(n20942), .ZN(n20893) );
  INV_X1 U12976 ( .A(n12678), .ZN(n12679) );
  INV_X1 U12977 ( .A(n20095), .ZN(n20102) );
  INV_X1 U12978 ( .A(n20052), .ZN(n15859) );
  INV_X1 U12979 ( .A(n20099), .ZN(n20088) );
  NAND2_X1 U12980 ( .A1(n20116), .A2(n11541), .ZN(n14542) );
  NOR2_X1 U12981 ( .A1(n12338), .A2(n12337), .ZN(n12339) );
  OR2_X1 U12982 ( .A1(n20121), .A2(n20141), .ZN(n20123) );
  INV_X1 U12983 ( .A(n20121), .ZN(n20143) );
  NOR2_X1 U12984 ( .A1(n13620), .A2(n13619), .ZN(n13824) );
  OR2_X1 U12985 ( .A1(n20200), .A2(n12642), .ZN(n15913) );
  INV_X1 U12986 ( .A(n20199), .ZN(n20193) );
  INV_X1 U12987 ( .A(n20200), .ZN(n20016) );
  OR2_X1 U12988 ( .A1(n12461), .A2(n12460), .ZN(n20230) );
  INV_X1 U12989 ( .A(n20235), .ZN(n20246) );
  INV_X1 U12990 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20701) );
  AOI21_X1 U12991 ( .B1(n13979), .B2(n13978), .A(n20421), .ZN(n20255) );
  OR2_X1 U12992 ( .A1(n20373), .A2(n20414), .ZN(n20337) );
  OR2_X1 U12993 ( .A1(n20373), .A2(n20314), .ZN(n21148) );
  OR2_X1 U12994 ( .A1(n20373), .A2(n20372), .ZN(n20423) );
  NAND2_X1 U12995 ( .A1(n20506), .A2(n20661), .ZN(n20468) );
  NAND2_X1 U12996 ( .A1(n20506), .A2(n20700), .ZN(n20500) );
  NAND2_X1 U12997 ( .A1(n20506), .A2(n20731), .ZN(n20535) );
  NAND2_X1 U12998 ( .A1(n20631), .A2(n20661), .ZN(n20586) );
  NAND2_X1 U12999 ( .A1(n20631), .A2(n20700), .ZN(n20624) );
  NAND2_X1 U13000 ( .A1(n20631), .A2(n20630), .ZN(n20699) );
  NAND2_X1 U13001 ( .A1(n20732), .A2(n20700), .ZN(n20773) );
  NAND2_X1 U13002 ( .A1(n20732), .A2(n20630), .ZN(n20837) );
  INV_X1 U13003 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16108) );
  NAND2_X1 U13004 ( .A1(n13082), .A2(n13081), .ZN(n13515) );
  AND2_X1 U13005 ( .A1(n12747), .A2(n12746), .ZN(n12748) );
  INV_X1 U13006 ( .A(n19151), .ZN(n19121) );
  AND2_X1 U13007 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  INV_X2 U13008 ( .A(n15042), .ZN(n15036) );
  AND2_X1 U13009 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  AND2_X1 U13010 ( .A1(n13445), .A2(n19843), .ZN(n19187) );
  NAND2_X1 U13011 ( .A1(n19187), .A2(n13446), .ZN(n19210) );
  NAND2_X1 U13012 ( .A1(n13551), .A2(n19995), .ZN(n19249) );
  NAND2_X1 U13013 ( .A1(n12733), .A2(n19348), .ZN(n13549) );
  INV_X1 U13014 ( .A(n19290), .ZN(n19304) );
  INV_X1 U13015 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16284) );
  INV_X1 U13016 ( .A(n19318), .ZN(n19297) );
  INV_X1 U13017 ( .A(n19319), .ZN(n19305) );
  OR2_X1 U13018 ( .A1(n18919), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19091) );
  NAND2_X1 U13019 ( .A1(n11211), .A2(n19978), .ZN(n19331) );
  INV_X1 U13020 ( .A(n19338), .ZN(n16341) );
  INV_X1 U13021 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16376) );
  INV_X1 U13022 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15700) );
  AOI21_X1 U13023 ( .B1(n15538), .B2(n15537), .A(n15536), .ZN(n19378) );
  INV_X1 U13024 ( .A(n19450), .ZN(n19460) );
  INV_X1 U13025 ( .A(n19511), .ZN(n19495) );
  AND2_X1 U13026 ( .A1(n14109), .A2(n14108), .ZN(n19515) );
  NAND2_X1 U13027 ( .A1(n19783), .A2(n19400), .ZN(n19563) );
  NAND2_X1 U13028 ( .A1(n19548), .A2(n19783), .ZN(n19598) );
  INV_X1 U13029 ( .A(n19617), .ZN(n19629) );
  INV_X1 U13030 ( .A(n19651), .ZN(n19661) );
  AND2_X1 U13031 ( .A1(n14016), .A2(n14015), .ZN(n19674) );
  INV_X1 U13032 ( .A(n19707), .ZN(n19718) );
  NAND2_X1 U13033 ( .A1(n19682), .A2(n19723), .ZN(n19749) );
  AOI211_X2 U13034 ( .C1(n15580), .C2(n15586), .A(n19601), .B(n15579), .ZN(
        n19775) );
  INV_X1 U13035 ( .A(n19797), .ZN(n19841) );
  INV_X1 U13036 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19777) );
  INV_X1 U13037 ( .A(n19937), .ZN(n19850) );
  INV_X1 U13038 ( .A(n16956), .ZN(n16947) );
  NAND2_X1 U13039 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16958), .ZN(n16944) );
  NOR2_X1 U13040 ( .A1(n16645), .A2(n17002), .ZN(n17007) );
  NOR2_X1 U13041 ( .A1(n17113), .A2(n15690), .ZN(n17272) );
  INV_X1 U13042 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17277) );
  AND2_X1 U13043 ( .A1(n17298), .A2(n17340), .ZN(n17296) );
  NOR2_X1 U13044 ( .A1(n17502), .A2(n17431), .ZN(n17435) );
  NAND2_X1 U13045 ( .A1(n17451), .A2(n18262), .ZN(n17479) );
  NAND2_X1 U13046 ( .A1(n17450), .A2(n17449), .ZN(n17509) );
  AOI211_X1 U13047 ( .C1(n18895), .C2(n18268), .A(n17512), .B(n17511), .ZN(
        n17524) );
  INV_X1 U13048 ( .A(n17557), .ZN(n17553) );
  OAI21_X2 U13049 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18901), .A(n16579), 
        .ZN(n17927) );
  NOR2_X1 U13050 ( .A1(n17884), .A2(n17886), .ZN(n17924) );
  OAI221_X2 U13051 ( .B1(n15710), .B2(n18692), .C1(n15710), .C2(n15709), .A(
        n18902), .ZN(n18235) );
  INV_X1 U13052 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18148) );
  INV_X1 U13053 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18713) );
  INV_X1 U13054 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18255) );
  INV_X1 U13055 ( .A(n18902), .ZN(n18750) );
  INV_X1 U13056 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18850) );
  INV_X1 U13057 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18768) );
  INV_X1 U13058 ( .A(n16523), .ZN(n16528) );
  OAI21_X1 U13059 ( .B1(n14574), .B2(n14542), .A(n13415), .ZN(P1_U2842) );
  NAND2_X1 U13060 ( .A1(n13080), .A2(n13079), .ZN(P2_U2858) );
  NAND2_X1 U13061 ( .A1(n10095), .A2(n13096), .ZN(P2_U2985) );
  INV_X1 U13062 ( .A(n13428), .ZN(n10173) );
  AOI22_X1 U13063 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10101) );
  AND2_X4 U13064 ( .A1(n10327), .A2(n16364), .ZN(n10341) );
  AND2_X4 U13065 ( .A1(n10329), .A2(n16364), .ZN(n10337) );
  AOI22_X1 U13066 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10100) );
  AND2_X4 U13067 ( .A1(n10330), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10339) );
  AOI22_X1 U13068 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10099) );
  NAND4_X1 U13069 ( .A1(n10102), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n10103) );
  AOI22_X1 U13070 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10173), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U13071 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U13072 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U13073 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10104) );
  NAND4_X1 U13074 ( .A1(n10107), .A2(n10106), .A3(n10105), .A4(n10104), .ZN(
        n10108) );
  NAND2_X1 U13075 ( .A1(n10108), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10109) );
  AOI22_X1 U13076 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10173), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10113) );
  AOI22_X1 U13077 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13433), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U13078 ( .A1(n10337), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U13079 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10110) );
  NAND4_X1 U13080 ( .A1(n10113), .A2(n10112), .A3(n10111), .A4(n10110), .ZN(
        n10114) );
  AOI22_X1 U13081 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U13082 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U13083 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13433), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U13084 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10115) );
  NAND4_X1 U13085 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10119) );
  AOI21_X1 U13086 ( .B1(n12887), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n10120), .ZN(n10125) );
  AOI22_X1 U13087 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U13088 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U13089 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10122) );
  NAND3_X1 U13090 ( .A1(n10125), .A2(n10124), .A3(n10086), .ZN(n10133) );
  INV_X2 U13091 ( .A(n13428), .ZN(n12887) );
  AOI22_X1 U13092 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12887), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13093 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U13094 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10128) );
  NAND3_X1 U13095 ( .A1(n10131), .A2(n10130), .A3(n10129), .ZN(n10132) );
  NAND3_X1 U13096 ( .A1(n10771), .A2(n19364), .A3(n10770), .ZN(n10778) );
  NAND2_X1 U13097 ( .A1(n10969), .A2(n10774), .ZN(n10768) );
  AOI22_X1 U13098 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10173), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13099 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n10121), .ZN(n10136) );
  AOI22_X1 U13100 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10341), .B1(
        n13433), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U13101 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10134) );
  NAND4_X1 U13102 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10139) );
  NAND2_X1 U13103 ( .A1(n10139), .A2(n10138), .ZN(n10146) );
  AOI22_X1 U13104 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U13105 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U13106 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13433), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13107 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10140) );
  NAND4_X1 U13108 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n10144) );
  NAND2_X1 U13109 ( .A1(n10144), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10145) );
  NAND2_X1 U13110 ( .A1(n10146), .A2(n10145), .ZN(n10203) );
  NAND3_X1 U13111 ( .A1(n10778), .A2(n10768), .A3(n15558), .ZN(n11198) );
  AOI22_X1 U13112 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12887), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13113 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13114 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U13115 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10147) );
  NAND3_X1 U13116 ( .A1(n10150), .A2(n10149), .A3(n10088), .ZN(n10156) );
  AOI22_X1 U13117 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10173), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13118 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U13119 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U13120 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10151) );
  NAND3_X1 U13121 ( .A1(n10154), .A2(n10153), .A3(n10081), .ZN(n10155) );
  NAND2_X2 U13122 ( .A1(n10156), .A2(n10155), .ZN(n10204) );
  NAND2_X1 U13123 ( .A1(n11198), .A2(n11200), .ZN(n10159) );
  NAND2_X1 U13124 ( .A1(n10159), .A2(n10158), .ZN(n10248) );
  AOI22_X1 U13125 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13126 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13127 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12887), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13128 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10162) );
  NAND3_X1 U13129 ( .A1(n10089), .A2(n10163), .A3(n10162), .ZN(n10170) );
  AOI22_X1 U13130 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13131 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10164) );
  AND3_X1 U13132 ( .A1(n10165), .A2(n10164), .A3(n10138), .ZN(n10168) );
  AOI22_X1 U13133 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12887), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13134 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10166) );
  NAND3_X1 U13135 ( .A1(n10168), .A2(n10167), .A3(n10166), .ZN(n10169) );
  AOI22_X1 U13136 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13137 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13138 ( .A1(n10173), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13139 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10341), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10174) );
  NAND3_X1 U13140 ( .A1(n10092), .A2(n10175), .A3(n10174), .ZN(n10181) );
  AOI22_X1 U13141 ( .A1(n12887), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13142 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13433), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13143 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U13144 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10176) );
  NAND3_X1 U13145 ( .A1(n10179), .A2(n10178), .A3(n10087), .ZN(n10180) );
  NAND2_X1 U13146 ( .A1(n10248), .A2(n10751), .ZN(n10211) );
  NAND3_X1 U13147 ( .A1(n10204), .A2(n19364), .A3(n10184), .ZN(n10185) );
  NAND2_X1 U13148 ( .A1(n10223), .A2(n10185), .ZN(n10202) );
  AOI22_X1 U13149 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12887), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13150 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13151 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13152 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10187) );
  NAND4_X1 U13153 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10191) );
  NAND2_X1 U13154 ( .A1(n10191), .A2(n10138), .ZN(n10200) );
  AOI21_X1 U13155 ( .B1(n12887), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n10192), .ZN(n10197) );
  AOI22_X1 U13156 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10121), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13157 ( .A1(n10341), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10337), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13158 ( .A1(n10342), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10339), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10193) );
  NAND3_X1 U13159 ( .A1(n10197), .A2(n10196), .A3(n10195), .ZN(n10198) );
  NAND2_X1 U13160 ( .A1(n10198), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10199) );
  NAND2_X1 U13161 ( .A1(n10202), .A2(n10201), .ZN(n10209) );
  INV_X1 U13162 ( .A(n10213), .ZN(n10207) );
  AND2_X1 U13163 ( .A1(n10204), .A2(n10205), .ZN(n10206) );
  NAND2_X1 U13164 ( .A1(n11202), .A2(n10228), .ZN(n10249) );
  NAND2_X1 U13165 ( .A1(n10249), .A2(n16384), .ZN(n10210) );
  NAND2_X1 U13166 ( .A1(n10211), .A2(n10247), .ZN(n10212) );
  NAND2_X1 U13167 ( .A1(n10212), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U13168 ( .A1(n10218), .A2(n11200), .ZN(n10214) );
  INV_X1 U13169 ( .A(n10771), .ZN(n10215) );
  NAND2_X1 U13170 ( .A1(n10216), .A2(n10245), .ZN(n10271) );
  NAND2_X1 U13171 ( .A1(n10271), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10222) );
  NAND2_X1 U13172 ( .A1(n19348), .A2(n16384), .ZN(n10224) );
  INV_X1 U13173 ( .A(n10224), .ZN(n10219) );
  AND2_X2 U13174 ( .A1(n10218), .A2(n10204), .ZN(n11204) );
  NOR2_X1 U13175 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19987) );
  NAND2_X1 U13176 ( .A1(n13762), .A2(n19348), .ZN(n10227) );
  NAND2_X2 U13177 ( .A1(n10497), .A2(n10224), .ZN(n11196) );
  OAI21_X1 U13178 ( .B1(n10771), .B2(n19996), .A(n10204), .ZN(n10225) );
  NAND3_X1 U13179 ( .A1(n10226), .A2(n11196), .A3(n10225), .ZN(n14167) );
  INV_X1 U13180 ( .A(n14167), .ZN(n11190) );
  NAND2_X1 U13181 ( .A1(n11190), .A2(n11204), .ZN(n13760) );
  NAND2_X1 U13182 ( .A1(n10227), .A2(n13760), .ZN(n10827) );
  INV_X1 U13183 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15508) );
  AND2_X2 U13184 ( .A1(n11203), .A2(n10229), .ZN(n11209) );
  INV_X1 U13185 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10494) );
  INV_X1 U13186 ( .A(n10261), .ZN(n10230) );
  NAND2_X1 U13187 ( .A1(n10230), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U13188 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10231) );
  OAI211_X1 U13189 ( .C1(n10264), .C2(n10494), .A(n10232), .B(n10231), .ZN(
        n10233) );
  INV_X1 U13190 ( .A(n10233), .ZN(n10234) );
  OAI21_X2 U13191 ( .B1(n10260), .B2(n15508), .A(n10234), .ZN(n10255) );
  INV_X1 U13192 ( .A(n10760), .ZN(n10235) );
  NOR2_X1 U13193 ( .A1(n10235), .A2(n10777), .ZN(n10236) );
  INV_X1 U13194 ( .A(n10264), .ZN(n10959) );
  OAI22_X1 U13195 ( .A1(n10271), .A2(n10236), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10959), .ZN(n10239) );
  INV_X1 U13196 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13085) );
  INV_X1 U13197 ( .A(n19987), .ZN(n10241) );
  OAI22_X1 U13198 ( .A1(n13760), .A2(n13085), .B1(n10241), .B2(n19973), .ZN(
        n10237) );
  INV_X1 U13199 ( .A(n10237), .ZN(n10238) );
  NAND2_X1 U13200 ( .A1(n10239), .A2(n10238), .ZN(n10291) );
  INV_X1 U13201 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16351) );
  INV_X1 U13202 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U13203 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10240) );
  INV_X1 U13204 ( .A(n10243), .ZN(n10246) );
  NAND2_X1 U13205 ( .A1(n10278), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10244) );
  INV_X1 U13206 ( .A(n10247), .ZN(n10251) );
  NAND2_X1 U13207 ( .A1(n10291), .A2(n10290), .ZN(n10292) );
  NAND2_X1 U13208 ( .A1(n10294), .A2(n10292), .ZN(n10259) );
  INV_X1 U13209 ( .A(n10256), .ZN(n10257) );
  NAND2_X2 U13210 ( .A1(n10259), .A2(n10258), .ZN(n10288) );
  INV_X1 U13211 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10267) );
  INV_X1 U13212 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U13213 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10262) );
  INV_X1 U13214 ( .A(n10268), .ZN(n10269) );
  NAND2_X1 U13215 ( .A1(n10270), .A2(n10269), .ZN(n10273) );
  OAI21_X1 U13216 ( .B1(n19957), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15803), 
        .ZN(n10272) );
  AOI21_X2 U13217 ( .B1(n10286), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10272), .ZN(n10274) );
  NAND2_X1 U13218 ( .A1(n10288), .A2(n10287), .ZN(n10277) );
  INV_X1 U13219 ( .A(n10273), .ZN(n10275) );
  NAND2_X1 U13220 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  INV_X1 U13221 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10281) );
  INV_X1 U13222 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13921) );
  NAND2_X1 U13223 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10279) );
  OAI211_X1 U13224 ( .C1(n10264), .C2(n10281), .A(n10280), .B(n10279), .ZN(
        n10282) );
  INV_X1 U13225 ( .A(n10282), .ZN(n10283) );
  AND2_X1 U13226 ( .A1(n19987), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10285) );
  XNOR2_X2 U13227 ( .A(n10840), .B(n10839), .ZN(n12750) );
  XNOR2_X2 U13228 ( .A(n10288), .B(n10287), .ZN(n12769) );
  INV_X1 U13229 ( .A(n12769), .ZN(n10289) );
  OR2_X2 U13230 ( .A1(n12750), .A2(n10289), .ZN(n10314) );
  OR2_X1 U13231 ( .A1(n14166), .A2(n10295), .ZN(n10313) );
  OR2_X2 U13232 ( .A1(n10314), .A2(n10313), .ZN(n14114) );
  INV_X1 U13233 ( .A(n10295), .ZN(n10296) );
  OR2_X1 U13234 ( .A1(n10296), .A2(n14166), .ZN(n10317) );
  NOR2_X1 U13235 ( .A1(n10314), .A2(n10317), .ZN(n10442) );
  NAND2_X1 U13236 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10297) );
  OAI211_X1 U13237 ( .C1(n19498), .C2(n14114), .A(n10297), .B(n19997), .ZN(
        n10300) );
  INV_X1 U13238 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12949) );
  NAND2_X1 U13239 ( .A1(n13527), .A2(n14166), .ZN(n10309) );
  INV_X1 U13241 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10351) );
  OAI22_X1 U13242 ( .A1(n14011), .A2(n12949), .B1(n15566), .B2(n10351), .ZN(
        n10299) );
  NOR2_X1 U13243 ( .A1(n10300), .A2(n10299), .ZN(n10326) );
  INV_X1 U13244 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10301) );
  OR2_X2 U13245 ( .A1(n12750), .A2(n14127), .ZN(n10318) );
  INV_X1 U13246 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10356) );
  OAI22_X1 U13247 ( .A1(n10301), .A2(n19404), .B1(n19630), .B2(n10356), .ZN(
        n10304) );
  INV_X1 U13248 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10353) );
  INV_X1 U13249 ( .A(n14166), .ZN(n19320) );
  INV_X1 U13250 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12803) );
  NOR2_X1 U13251 ( .A1(n10304), .A2(n10303), .ZN(n10325) );
  INV_X1 U13252 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10308) );
  INV_X1 U13253 ( .A(n10313), .ZN(n10306) );
  NAND2_X1 U13254 ( .A1(n9643), .A2(n10306), .ZN(n10550) );
  INV_X1 U13255 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10307) );
  OAI22_X1 U13256 ( .A1(n10308), .A2(n19776), .B1(n10550), .B2(n10307), .ZN(
        n10312) );
  INV_X1 U13257 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U13258 ( .A1(n9643), .A2(n10310), .ZN(n10431) );
  INV_X1 U13259 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10363) );
  OAI22_X1 U13260 ( .A1(n10362), .A2(n10544), .B1(n10431), .B2(n10363), .ZN(
        n10311) );
  NOR2_X1 U13261 ( .A1(n10312), .A2(n10311), .ZN(n10324) );
  INV_X1 U13262 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10316) );
  INV_X1 U13263 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10315) );
  OAI22_X1 U13264 ( .A1(n10316), .A2(n15552), .B1(n19469), .B2(n10315), .ZN(
        n10322) );
  INV_X1 U13265 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12942) );
  INV_X1 U13266 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10365) );
  OAI22_X1 U13267 ( .A1(n12942), .A2(n19435), .B1(n10553), .B2(n10365), .ZN(
        n10321) );
  NOR2_X1 U13268 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  NAND4_X1 U13269 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10391) );
  AND2_X1 U13270 ( .A1(n15504), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10328) );
  AOI22_X1 U13271 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12924), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13272 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10335) );
  INV_X1 U13273 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15590) );
  INV_X1 U13274 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19346) );
  OAI22_X1 U13275 ( .A1(n11138), .A2(n15590), .B1(n11132), .B2(n19346), .ZN(
        n10331) );
  INV_X1 U13276 ( .A(n10331), .ZN(n10334) );
  INV_X1 U13277 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15575) );
  INV_X1 U13278 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14121) );
  OAI22_X1 U13279 ( .A1(n11131), .A2(n15575), .B1(n11143), .B2(n14121), .ZN(
        n10332) );
  INV_X1 U13280 ( .A(n10332), .ZN(n10333) );
  NAND4_X1 U13281 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10350) );
  AOI22_X1 U13282 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12913), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10348) );
  INV_X1 U13283 ( .A(n10337), .ZN(n12888) );
  INV_X1 U13284 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13285 ( .A1(n10121), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11087) );
  INV_X1 U13286 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11021) );
  OAI22_X1 U13287 ( .A1(n11141), .A2(n11028), .B1(n11087), .B2(n11021), .ZN(
        n10338) );
  INV_X1 U13288 ( .A(n10338), .ZN(n10347) );
  INV_X1 U13289 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11029) );
  INV_X1 U13290 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11017) );
  OAI22_X1 U13291 ( .A1(n11130), .A2(n11029), .B1(n13779), .B2(n11017), .ZN(
        n10340) );
  INV_X1 U13292 ( .A(n10340), .ZN(n10346) );
  INV_X1 U13293 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14023) );
  INV_X1 U13294 ( .A(n10342), .ZN(n12889) );
  INV_X1 U13295 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12817) );
  OAI22_X1 U13296 ( .A1(n11133), .A2(n14023), .B1(n12882), .B2(n12817), .ZN(
        n10344) );
  INV_X1 U13297 ( .A(n10344), .ZN(n10345) );
  NAND4_X1 U13298 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10349) );
  OR2_X1 U13299 ( .A1(n10794), .A2(n19997), .ZN(n16355) );
  OAI22_X1 U13300 ( .A1(n11131), .A2(n10351), .B1(n12882), .B2(n12803), .ZN(
        n10352) );
  INV_X1 U13301 ( .A(n10352), .ZN(n10361) );
  AOI22_X1 U13302 ( .A1(n12909), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12913), .ZN(n10360) );
  INV_X1 U13303 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10354) );
  OAI22_X1 U13304 ( .A1(n11137), .A2(n10354), .B1(n11141), .B2(n10353), .ZN(
        n10355) );
  INV_X1 U13305 ( .A(n10355), .ZN(n10359) );
  OAI22_X1 U13306 ( .A1(n11133), .A2(n12949), .B1(n10356), .B2(n11087), .ZN(
        n10357) );
  INV_X1 U13307 ( .A(n10357), .ZN(n10358) );
  NAND4_X1 U13308 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10372) );
  AOI22_X1 U13309 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12924), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13310 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10369) );
  OAI22_X1 U13311 ( .A1(n11138), .A2(n10363), .B1(n11132), .B2(n10362), .ZN(
        n10364) );
  INV_X1 U13312 ( .A(n10364), .ZN(n10368) );
  OAI22_X1 U13313 ( .A1(n11143), .A2(n19498), .B1(n13779), .B2(n10365), .ZN(
        n10366) );
  INV_X1 U13314 ( .A(n10366), .ZN(n10367) );
  NAND4_X1 U13315 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10371) );
  NOR2_X1 U13316 ( .A1(n16355), .A2(n10982), .ZN(n10798) );
  INV_X1 U13317 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12784) );
  INV_X1 U13318 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10373) );
  OAI22_X1 U13319 ( .A1(n12784), .A2(n11131), .B1(n11130), .B2(n10373), .ZN(
        n10375) );
  INV_X1 U13320 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12975) );
  INV_X1 U13321 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12773) );
  OAI22_X1 U13322 ( .A1(n11133), .A2(n12975), .B1(n11132), .B2(n12773), .ZN(
        n10374) );
  NOR2_X1 U13323 ( .A1(n10375), .A2(n10374), .ZN(n10389) );
  INV_X1 U13324 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19756) );
  INV_X1 U13325 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10376) );
  OAI22_X1 U13326 ( .A1(n19756), .A2(n11138), .B1(n11137), .B2(n10376), .ZN(
        n10379) );
  INV_X1 U13327 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10377) );
  OAI22_X1 U13328 ( .A1(n11143), .A2(n19501), .B1(n11141), .B2(n10377), .ZN(
        n10378) );
  NOR2_X1 U13329 ( .A1(n10379), .A2(n10378), .ZN(n10388) );
  AOI22_X1 U13330 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12924), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13331 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10382) );
  INV_X1 U13332 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12793) );
  OR2_X1 U13333 ( .A1(n11087), .A2(n12793), .ZN(n10381) );
  NAND2_X1 U13334 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10380) );
  NAND4_X1 U13335 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10386) );
  INV_X1 U13336 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10384) );
  INV_X1 U13337 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12788) );
  OAI22_X1 U13338 ( .A1(n10384), .A2(n13779), .B1(n12882), .B2(n12788), .ZN(
        n10385) );
  NOR2_X1 U13339 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  NAND3_X1 U13340 ( .A1(n10389), .A2(n10388), .A3(n10387), .ZN(n10989) );
  OR2_X1 U13341 ( .A1(n10798), .A2(n10989), .ZN(n10390) );
  INV_X1 U13342 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12839) );
  INV_X1 U13343 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13023) );
  OAI22_X1 U13344 ( .A1(n12839), .A2(n11131), .B1(n11133), .B2(n13023), .ZN(
        n10394) );
  INV_X1 U13345 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10392) );
  INV_X1 U13346 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12780) );
  OAI22_X1 U13347 ( .A1(n11130), .A2(n10392), .B1(n11132), .B2(n12780), .ZN(
        n10393) );
  NOR2_X1 U13348 ( .A1(n10394), .A2(n10393), .ZN(n10408) );
  INV_X1 U13349 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10395) );
  INV_X1 U13350 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12849) );
  OAI22_X1 U13351 ( .A1(n10395), .A2(n11137), .B1(n11138), .B2(n12849), .ZN(
        n10398) );
  INV_X1 U13352 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12840) );
  INV_X1 U13353 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10396) );
  OAI22_X1 U13354 ( .A1(n11143), .A2(n12840), .B1(n11141), .B2(n10396), .ZN(
        n10397) );
  NOR2_X1 U13355 ( .A1(n10398), .A2(n10397), .ZN(n10407) );
  AOI22_X1 U13356 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12924), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13357 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12930), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10401) );
  INV_X1 U13358 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12850) );
  OR2_X1 U13359 ( .A1(n11087), .A2(n12850), .ZN(n10400) );
  NAND2_X1 U13360 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10399) );
  NAND4_X1 U13361 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10405) );
  INV_X1 U13362 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10403) );
  INV_X1 U13363 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12844) );
  OAI22_X1 U13364 ( .A1(n10403), .A2(n13779), .B1(n12882), .B2(n12844), .ZN(
        n10404) );
  NOR2_X1 U13365 ( .A1(n10405), .A2(n10404), .ZN(n10406) );
  NAND3_X1 U13366 ( .A1(n10408), .A2(n10407), .A3(n10406), .ZN(n11003) );
  INV_X1 U13367 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10409) );
  INV_X1 U13368 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13001) );
  OAI22_X1 U13369 ( .A1(n10409), .A2(n11138), .B1(n11133), .B2(n13001), .ZN(
        n10412) );
  INV_X1 U13370 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10410) );
  INV_X1 U13371 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12758) );
  OAI22_X1 U13372 ( .A1(n11137), .A2(n10410), .B1(n11132), .B2(n12758), .ZN(
        n10411) );
  NOR2_X1 U13373 ( .A1(n10412), .A2(n10411), .ZN(n10430) );
  INV_X1 U13374 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10414) );
  INV_X1 U13375 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10413) );
  OAI22_X1 U13376 ( .A1(n10414), .A2(n11131), .B1(n11130), .B2(n10413), .ZN(
        n10418) );
  INV_X1 U13377 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10416) );
  INV_X1 U13378 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10415) );
  OAI22_X1 U13379 ( .A1(n11143), .A2(n10416), .B1(n11141), .B2(n10415), .ZN(
        n10417) );
  NOR2_X1 U13380 ( .A1(n10418), .A2(n10417), .ZN(n10429) );
  AOI22_X1 U13381 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12924), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U13382 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10422) );
  INV_X1 U13383 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10419) );
  OR2_X1 U13384 ( .A1(n11087), .A2(n10419), .ZN(n10421) );
  NAND2_X1 U13385 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10420) );
  NAND4_X1 U13386 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n10427) );
  INV_X1 U13387 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10425) );
  INV_X1 U13388 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10424) );
  OAI22_X1 U13389 ( .A1(n10425), .A2(n13779), .B1(n12882), .B2(n10424), .ZN(
        n10426) );
  NOR2_X1 U13390 ( .A1(n10427), .A2(n10426), .ZN(n10428) );
  NAND3_X1 U13391 ( .A1(n10430), .A2(n10429), .A3(n10428), .ZN(n10999) );
  INV_X1 U13392 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10455) );
  INV_X1 U13393 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10449) );
  OAI22_X1 U13394 ( .A1(n10455), .A2(n10540), .B1(n10550), .B2(n10449), .ZN(
        n10434) );
  INV_X1 U13395 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10432) );
  INV_X1 U13396 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10453) );
  OAI22_X1 U13397 ( .A1(n10432), .A2(n19776), .B1(n10431), .B2(n10453), .ZN(
        n10433) );
  NOR2_X1 U13398 ( .A1(n10434), .A2(n10433), .ZN(n10441) );
  INV_X1 U13399 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12854) );
  INV_X1 U13400 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13038) );
  OAI22_X1 U13401 ( .A1(n12854), .A2(n19469), .B1(n19435), .B2(n13038), .ZN(
        n10436) );
  INV_X1 U13402 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13845) );
  INV_X1 U13403 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10464) );
  OAI22_X1 U13404 ( .A1(n13845), .A2(n10544), .B1(n10553), .B2(n10464), .ZN(
        n10435) );
  NOR2_X1 U13405 ( .A1(n10436), .A2(n10435), .ZN(n10440) );
  INV_X1 U13406 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10450) );
  INV_X1 U13407 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10448) );
  OAI22_X1 U13408 ( .A1(n10450), .A2(n15566), .B1(n14114), .B2(n10448), .ZN(
        n10438) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12858) );
  INV_X1 U13410 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14032) );
  OAI22_X1 U13411 ( .A1(n12858), .A2(n15552), .B1(n14011), .B2(n14032), .ZN(
        n10437) );
  NOR2_X1 U13412 ( .A1(n10438), .A2(n10437), .ZN(n10439) );
  NAND3_X1 U13413 ( .A1(n10441), .A2(n10440), .A3(n10439), .ZN(n10474) );
  INV_X1 U13414 ( .A(n19630), .ZN(n10443) );
  INV_X1 U13415 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10444) );
  INV_X1 U13416 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10465) );
  OAI22_X1 U13417 ( .A1(n10444), .A2(n19404), .B1(n19692), .B2(n10465), .ZN(
        n10445) );
  INV_X1 U13418 ( .A(n10445), .ZN(n10446) );
  NAND2_X1 U13419 ( .A1(n10447), .A2(n10446), .ZN(n10473) );
  OAI22_X1 U13420 ( .A1(n11130), .A2(n10449), .B1(n11143), .B2(n10448), .ZN(
        n10452) );
  OAI22_X1 U13421 ( .A1(n11131), .A2(n10450), .B1(n11132), .B2(n13845), .ZN(
        n10451) );
  NOR2_X1 U13422 ( .A1(n10452), .A2(n10451), .ZN(n10470) );
  INV_X1 U13423 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10454) );
  OAI22_X1 U13424 ( .A1(n11137), .A2(n10454), .B1(n11138), .B2(n10453), .ZN(
        n10457) );
  OAI22_X1 U13425 ( .A1(n11133), .A2(n14032), .B1(n11141), .B2(n10455), .ZN(
        n10456) );
  NOR2_X1 U13426 ( .A1(n10457), .A2(n10456), .ZN(n10469) );
  AOI22_X1 U13427 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12924), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13428 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10462) );
  INV_X1 U13429 ( .A(n11087), .ZN(n10458) );
  INV_X1 U13430 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10459) );
  OR2_X1 U13431 ( .A1(n11087), .A2(n10459), .ZN(n10461) );
  NAND2_X1 U13432 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10460) );
  NAND4_X1 U13433 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10467) );
  OAI22_X1 U13434 ( .A1(n12882), .A2(n10465), .B1(n13779), .B2(n10464), .ZN(
        n10466) );
  NOR2_X1 U13435 ( .A1(n10467), .A2(n10466), .ZN(n10468) );
  NAND3_X1 U13436 ( .A1(n10470), .A2(n10469), .A3(n10468), .ZN(n11007) );
  INV_X1 U13437 ( .A(n11007), .ZN(n10471) );
  NAND2_X1 U13438 ( .A1(n10471), .A2(n19348), .ZN(n10472) );
  OAI21_X2 U13439 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(n10581) );
  INV_X1 U13440 ( .A(n10581), .ZN(n10475) );
  INV_X1 U13441 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11142) );
  INV_X1 U13442 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11150) );
  OAI22_X1 U13443 ( .A1(n11142), .A2(n11131), .B1(n11130), .B2(n11150), .ZN(
        n10476) );
  INV_X1 U13444 ( .A(n10476), .ZN(n10483) );
  INV_X1 U13445 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13427) );
  INV_X1 U13446 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11129) );
  OAI22_X1 U13447 ( .A1(n13427), .A2(n11137), .B1(n11138), .B2(n11129), .ZN(
        n10477) );
  INV_X1 U13448 ( .A(n10477), .ZN(n10482) );
  INV_X1 U13449 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13424) );
  INV_X1 U13450 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19377) );
  OAI22_X1 U13451 ( .A1(n11133), .A2(n13424), .B1(n11132), .B2(n19377), .ZN(
        n10478) );
  INV_X1 U13452 ( .A(n10478), .ZN(n10481) );
  INV_X1 U13453 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13426) );
  INV_X1 U13454 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11151) );
  OAI22_X1 U13455 ( .A1(n11143), .A2(n13426), .B1(n11141), .B2(n11151), .ZN(
        n10479) );
  INV_X1 U13456 ( .A(n10479), .ZN(n10480) );
  NAND4_X1 U13457 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10493) );
  INV_X1 U13458 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12927) );
  INV_X1 U13459 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11136) );
  OAI22_X1 U13460 ( .A1(n12927), .A2(n12882), .B1(n13779), .B2(n11136), .ZN(
        n10484) );
  INV_X1 U13461 ( .A(n10484), .ZN(n10491) );
  INV_X1 U13462 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U13463 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10486) );
  NAND2_X1 U13464 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10485) );
  OAI211_X1 U13465 ( .C1(n11087), .C2(n11140), .A(n10486), .B(n10485), .ZN(
        n10487) );
  INV_X1 U13466 ( .A(n10487), .ZN(n10490) );
  AOI22_X1 U13467 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U13468 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10488) );
  NAND4_X1 U13469 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10492) );
  NAND2_X1 U13470 ( .A1(n10807), .A2(n11013), .ZN(n10518) );
  INV_X1 U13471 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13863) );
  NAND2_X1 U13472 ( .A1(n10494), .A2(n13863), .ZN(n10496) );
  NAND2_X1 U13473 ( .A1(n10751), .A2(n10989), .ZN(n10501) );
  MUX2_X1 U13474 ( .A(n10498), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10716) );
  NAND2_X1 U13475 ( .A1(n10716), .A2(n10728), .ZN(n10500) );
  NAND2_X1 U13476 ( .A1(n10498), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10499) );
  NAND2_X1 U13477 ( .A1(n10500), .A2(n10499), .ZN(n10503) );
  XNOR2_X1 U13478 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10502) );
  XNOR2_X1 U13479 ( .A(n10503), .B(n10502), .ZN(n10749) );
  INV_X1 U13480 ( .A(n10749), .ZN(n10729) );
  NOR2_X2 U13481 ( .A1(n10525), .A2(n10521), .ZN(n10520) );
  NAND2_X1 U13482 ( .A1(n10503), .A2(n10502), .ZN(n10505) );
  NAND2_X1 U13483 ( .A1(n19957), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13484 ( .A1(n10505), .A2(n10504), .ZN(n10510) );
  MUX2_X1 U13485 ( .A(n12752), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10509) );
  INV_X1 U13486 ( .A(n10509), .ZN(n10506) );
  XNOR2_X1 U13487 ( .A(n10510), .B(n10506), .ZN(n10719) );
  MUX2_X1 U13488 ( .A(n10507), .B(n10281), .S(n9930), .Z(n10519) );
  NOR2_X1 U13489 ( .A1(n10138), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10508) );
  AOI21_X1 U13490 ( .B1(n10510), .B2(n10509), .A(n10508), .ZN(n10722) );
  NOR2_X1 U13491 ( .A1(n16376), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10511) );
  NAND2_X1 U13492 ( .A1(n10722), .A2(n10511), .ZN(n10720) );
  INV_X1 U13493 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n20945) );
  MUX2_X1 U13494 ( .A(n10512), .B(n20945), .S(n9930), .Z(n10515) );
  INV_X1 U13495 ( .A(n10515), .ZN(n10532) );
  INV_X1 U13496 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10835) );
  MUX2_X1 U13497 ( .A(n10835), .B(n11007), .S(n14029), .Z(n10514) );
  INV_X1 U13498 ( .A(n10514), .ZN(n10513) );
  OAI21_X1 U13499 ( .B1(n10533), .B2(n10532), .A(n10513), .ZN(n10517) );
  NAND2_X1 U13500 ( .A1(n10515), .A2(n10514), .ZN(n10516) );
  NAND2_X1 U13501 ( .A1(n10517), .A2(n10584), .ZN(n19114) );
  INV_X1 U13502 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10831) );
  XNOR2_X1 U13503 ( .A(n10536), .B(n10831), .ZN(n14134) );
  XOR2_X1 U13504 ( .A(n10519), .B(n10520), .Z(n14943) );
  NOR2_X1 U13505 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14943), .ZN(
        n10531) );
  INV_X1 U13506 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11221) );
  AOI21_X1 U13507 ( .B1(n10521), .B2(n10525), .A(n10520), .ZN(n10522) );
  INV_X1 U13508 ( .A(n10522), .ZN(n14124) );
  NOR2_X1 U13509 ( .A1(n11221), .A2(n14124), .ZN(n10530) );
  INV_X1 U13510 ( .A(n10728), .ZN(n10524) );
  NAND2_X1 U13511 ( .A1(n14169), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10523) );
  INV_X1 U13512 ( .A(n10747), .ZN(n10752) );
  MUX2_X1 U13513 ( .A(n10718), .B(n13863), .S(n9930), .Z(n19148) );
  NOR2_X1 U13514 ( .A1(n19148), .A2(n16351), .ZN(n10528) );
  NAND2_X1 U13515 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10526) );
  OAI21_X1 U13516 ( .B1(n10526), .B2(n14029), .A(n10525), .ZN(n14956) );
  INV_X1 U13517 ( .A(n14956), .ZN(n10527) );
  NAND2_X1 U13518 ( .A1(n10528), .A2(n10527), .ZN(n13528) );
  INV_X1 U13519 ( .A(n13528), .ZN(n10529) );
  INV_X1 U13520 ( .A(n10528), .ZN(n16353) );
  NAND2_X1 U13521 ( .A1(n16353), .A2(n14956), .ZN(n13529) );
  OAI21_X1 U13522 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10529), .A(
        n13529), .ZN(n13672) );
  XNOR2_X1 U13523 ( .A(n11221), .B(n14124), .ZN(n13671) );
  NOR2_X1 U13524 ( .A1(n13672), .A2(n13671), .ZN(n13670) );
  NOR2_X1 U13525 ( .A1(n10530), .A2(n13670), .ZN(n13919) );
  NAND2_X1 U13526 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14943), .ZN(
        n13918) );
  OAI21_X1 U13527 ( .B1(n10531), .B2(n13919), .A(n13918), .ZN(n19296) );
  XNOR2_X1 U13528 ( .A(n10533), .B(n10532), .ZN(n19128) );
  XNOR2_X1 U13529 ( .A(n19128), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19295) );
  NAND2_X1 U13530 ( .A1(n19296), .A2(n19295), .ZN(n10535) );
  INV_X1 U13531 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19335) );
  OR2_X1 U13532 ( .A1(n19128), .A2(n19335), .ZN(n10534) );
  NAND2_X1 U13533 ( .A1(n10535), .A2(n10534), .ZN(n14135) );
  NAND2_X1 U13534 ( .A1(n14134), .A2(n14135), .ZN(n10538) );
  NAND2_X1 U13535 ( .A1(n10536), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10537) );
  NAND2_X1 U13536 ( .A1(n10538), .A2(n10537), .ZN(n14243) );
  INV_X1 U13537 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10539) );
  INV_X1 U13538 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12883) );
  OAI22_X1 U13539 ( .A1(n10539), .A2(n19404), .B1(n19630), .B2(n12883), .ZN(
        n10543) );
  INV_X1 U13540 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10541) );
  INV_X1 U13541 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10566) );
  OAI22_X1 U13542 ( .A1(n10541), .A2(n19776), .B1(n10540), .B2(n10566), .ZN(
        n10542) );
  NOR2_X1 U13543 ( .A1(n10543), .A2(n10542), .ZN(n10560) );
  INV_X1 U13544 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10562) );
  INV_X1 U13545 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10545) );
  OAI22_X1 U13546 ( .A1(n10562), .A2(n10544), .B1(n19435), .B2(n10545), .ZN(
        n10548) );
  INV_X1 U13547 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10546) );
  INV_X1 U13548 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12872) );
  OAI22_X1 U13549 ( .A1(n10546), .A2(n15552), .B1(n14114), .B2(n12872), .ZN(
        n10547) );
  NOR2_X1 U13550 ( .A1(n10548), .A2(n10547), .ZN(n10559) );
  INV_X1 U13551 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10565) );
  INV_X1 U13552 ( .A(n19538), .ZN(n10549) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12876) );
  OAI22_X1 U13554 ( .A1(n10565), .A2(n10549), .B1(n19692), .B2(n12876), .ZN(
        n10552) );
  INV_X1 U13555 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12881) );
  INV_X1 U13556 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10561) );
  OAI22_X1 U13557 ( .A1(n12881), .A2(n10431), .B1(n10550), .B2(n10561), .ZN(
        n10551) );
  NOR2_X1 U13558 ( .A1(n10552), .A2(n10551), .ZN(n10558) );
  INV_X1 U13559 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10554) );
  INV_X1 U13560 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10573) );
  OAI22_X1 U13561 ( .A1(n10554), .A2(n19469), .B1(n10553), .B2(n10573), .ZN(
        n10556) );
  INV_X1 U13562 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12869) );
  INV_X1 U13563 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13062) );
  OAI22_X1 U13564 ( .A1(n12869), .A2(n15566), .B1(n14011), .B2(n13062), .ZN(
        n10555) );
  NOR2_X1 U13565 ( .A1(n10556), .A2(n10555), .ZN(n10557) );
  NAND4_X1 U13566 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10580) );
  OAI22_X1 U13567 ( .A1(n12869), .A2(n11131), .B1(n11130), .B2(n10561), .ZN(
        n10564) );
  OAI22_X1 U13568 ( .A1(n11133), .A2(n13062), .B1(n11132), .B2(n10562), .ZN(
        n10563) );
  NOR2_X1 U13569 ( .A1(n10564), .A2(n10563), .ZN(n10578) );
  OAI22_X1 U13570 ( .A1(n10565), .A2(n11137), .B1(n11138), .B2(n12881), .ZN(
        n10568) );
  OAI22_X1 U13571 ( .A1(n11143), .A2(n12872), .B1(n11141), .B2(n10566), .ZN(
        n10567) );
  NOR2_X1 U13572 ( .A1(n10568), .A2(n10567), .ZN(n10577) );
  AOI22_X1 U13573 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12924), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13574 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10571) );
  OR2_X1 U13575 ( .A1(n11087), .A2(n12883), .ZN(n10570) );
  NAND2_X1 U13576 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10569) );
  NAND4_X1 U13577 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10575) );
  OAI22_X1 U13578 ( .A1(n10573), .A2(n13779), .B1(n12882), .B2(n12876), .ZN(
        n10574) );
  NOR2_X1 U13579 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  NAND2_X1 U13580 ( .A1(n10966), .A2(n19348), .ZN(n10579) );
  MUX2_X1 U13581 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n10966), .S(n14029), .Z(
        n10583) );
  AND2_X1 U13582 ( .A1(n10584), .A2(n10583), .ZN(n10585) );
  OR2_X1 U13583 ( .A1(n10585), .A2(n10593), .ZN(n19103) );
  OAI21_X1 U13584 ( .B1(n10806), .B2(n15135), .A(n19103), .ZN(n10586) );
  INV_X1 U13585 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14254) );
  XNOR2_X1 U13586 ( .A(n10586), .B(n14254), .ZN(n14244) );
  NAND2_X1 U13587 ( .A1(n14243), .A2(n14244), .ZN(n10588) );
  NAND2_X1 U13588 ( .A1(n10586), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10587) );
  INV_X1 U13589 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13747) );
  MUX2_X1 U13590 ( .A(n13747), .B(n15135), .S(n14029), .Z(n10591) );
  INV_X1 U13591 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10854) );
  NOR2_X1 U13592 ( .A1(n14029), .A2(n10854), .ZN(n10596) );
  INV_X1 U13593 ( .A(n10596), .ZN(n10589) );
  XNOR2_X1 U13594 ( .A(n10599), .B(n10589), .ZN(n19082) );
  AND2_X1 U13595 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10590) );
  NAND2_X1 U13596 ( .A1(n19082), .A2(n10590), .ZN(n15260) );
  INV_X1 U13597 ( .A(n10591), .ZN(n10592) );
  XNOR2_X1 U13598 ( .A(n10593), .B(n10592), .ZN(n19090) );
  NAND2_X1 U13599 ( .A1(n19090), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15257) );
  NAND2_X1 U13600 ( .A1(n19082), .A2(n15135), .ZN(n10594) );
  INV_X1 U13601 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16324) );
  NAND2_X1 U13602 ( .A1(n10594), .A2(n16324), .ZN(n15261) );
  OR2_X1 U13603 ( .A1(n19090), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15259) );
  AND2_X1 U13604 ( .A1(n15261), .A2(n15259), .ZN(n10595) );
  NAND2_X1 U13605 ( .A1(n9930), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10597) );
  XNOR2_X1 U13606 ( .A(n10598), .B(n10597), .ZN(n19072) );
  NAND2_X1 U13607 ( .A1(n19072), .A2(n15135), .ZN(n10605) );
  INV_X1 U13608 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15493) );
  INV_X1 U13609 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13994) );
  NAND2_X1 U13610 ( .A1(n9930), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10600) );
  OAI21_X1 U13611 ( .B1(n10601), .B2(n10600), .A(n10690), .ZN(n10602) );
  OR2_X1 U13612 ( .A1(n10609), .A2(n10602), .ZN(n19060) );
  INV_X1 U13613 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16269) );
  OAI21_X1 U13614 ( .B1(n19060), .B2(n11013), .A(n16269), .ZN(n16276) );
  INV_X1 U13615 ( .A(n19060), .ZN(n10604) );
  AND2_X1 U13616 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10603) );
  NAND2_X1 U13617 ( .A1(n10604), .A2(n10603), .ZN(n16275) );
  OR2_X1 U13618 ( .A1(n10605), .A2(n15493), .ZN(n15249) );
  AND2_X1 U13619 ( .A1(n16275), .A2(n15249), .ZN(n10606) );
  NAND2_X1 U13620 ( .A1(n9930), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10608) );
  OR2_X1 U13621 ( .A1(n10609), .A2(n10608), .ZN(n10611) );
  INV_X1 U13622 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13948) );
  INV_X1 U13623 ( .A(n10614), .ZN(n10610) );
  AND2_X1 U13624 ( .A1(n10611), .A2(n10610), .ZN(n19052) );
  NAND2_X1 U13625 ( .A1(n19052), .A2(n15135), .ZN(n15468) );
  INV_X1 U13626 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13627 ( .A1(n9930), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10613) );
  NAND3_X1 U13628 ( .A1(n9930), .A2(n10615), .A3(P2_EBX_REG_12__SCAN_IN), .ZN(
        n10616) );
  AND2_X1 U13629 ( .A1(n10644), .A2(n10616), .ZN(n19042) );
  NAND2_X1 U13630 ( .A1(n19042), .A2(n15135), .ZN(n10617) );
  XNOR2_X1 U13631 ( .A(n10617), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15242) );
  INV_X1 U13632 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16300) );
  NAND2_X1 U13633 ( .A1(n10617), .A2(n16300), .ZN(n10618) );
  NAND2_X1 U13634 ( .A1(n10619), .A2(n10618), .ZN(n15191) );
  INV_X1 U13635 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10870) );
  NOR2_X1 U13636 ( .A1(n14029), .A2(n10870), .ZN(n10643) );
  NOR2_X1 U13637 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n10620) );
  OAI21_X1 U13638 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(P2_EBX_REG_16__SCAN_IN), 
        .A(n9930), .ZN(n10621) );
  NAND2_X1 U13639 ( .A1(n9930), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U13640 ( .A1(n9930), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10626) );
  INV_X1 U13641 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n18942) );
  NAND2_X1 U13642 ( .A1(n9673), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10622) );
  OAI21_X1 U13643 ( .B1(n10622), .B2(n14029), .A(n10690), .ZN(n10623) );
  INV_X1 U13644 ( .A(n10623), .ZN(n10624) );
  NAND2_X1 U13645 ( .A1(n10677), .A2(n10624), .ZN(n18940) );
  OR2_X1 U13646 ( .A1(n18940), .A2(n11013), .ZN(n10625) );
  INV_X1 U13647 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21096) );
  NAND2_X1 U13648 ( .A1(n10625), .A2(n21096), .ZN(n15190) );
  OR2_X1 U13649 ( .A1(n10635), .A2(n10626), .ZN(n10627) );
  NAND2_X1 U13650 ( .A1(n10656), .A2(n10627), .ZN(n18962) );
  INV_X1 U13651 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20966) );
  OAI21_X1 U13652 ( .B1(n18962), .B2(n11013), .A(n20966), .ZN(n15392) );
  NAND2_X1 U13653 ( .A1(n10646), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10628) );
  MUX2_X1 U13654 ( .A(n10628), .B(n10646), .S(n14029), .Z(n10630) );
  INV_X1 U13655 ( .A(n10646), .ZN(n10629) );
  INV_X1 U13656 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14094) );
  NAND2_X1 U13657 ( .A1(n10629), .A2(n14094), .ZN(n10639) );
  NAND2_X1 U13658 ( .A1(n10630), .A2(n10639), .ZN(n19022) );
  INV_X1 U13659 ( .A(n19022), .ZN(n10631) );
  NAND2_X1 U13660 ( .A1(n10631), .A2(n15135), .ZN(n10670) );
  INV_X1 U13661 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16251) );
  NAND2_X1 U13662 ( .A1(n10670), .A2(n16251), .ZN(n16245) );
  AND2_X1 U13663 ( .A1(n15392), .A2(n16245), .ZN(n10654) );
  NOR2_X1 U13664 ( .A1(n10632), .A2(n10633), .ZN(n10634) );
  OR2_X1 U13665 ( .A1(n10635), .A2(n10634), .ZN(n18974) );
  INV_X1 U13666 ( .A(n18974), .ZN(n10636) );
  NAND2_X1 U13667 ( .A1(n10636), .A2(n15135), .ZN(n10658) );
  INV_X1 U13668 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15417) );
  NAND2_X1 U13669 ( .A1(n10658), .A2(n15417), .ZN(n15405) );
  INV_X1 U13670 ( .A(n10632), .ZN(n10638) );
  INV_X1 U13671 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10879) );
  NAND2_X1 U13672 ( .A1(n10651), .A2(n10879), .ZN(n10649) );
  NAND3_X1 U13673 ( .A1(n10649), .A2(n9930), .A3(P2_EBX_REG_17__SCAN_IN), .ZN(
        n10637) );
  NAND2_X1 U13674 ( .A1(n10638), .A2(n10637), .ZN(n18984) );
  INV_X1 U13675 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U13676 ( .A1(n10662), .A2(n10882), .ZN(n15197) );
  INV_X1 U13677 ( .A(n10651), .ZN(n10641) );
  NAND3_X1 U13678 ( .A1(n10639), .A2(n9930), .A3(P2_EBX_REG_15__SCAN_IN), .ZN(
        n10640) );
  NAND2_X1 U13679 ( .A1(n10641), .A2(n10640), .ZN(n19007) );
  OR2_X1 U13680 ( .A1(n19007), .A2(n11013), .ZN(n10642) );
  INV_X1 U13681 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U13682 ( .A1(n10642), .A2(n10874), .ZN(n15438) );
  NAND2_X1 U13683 ( .A1(n10644), .A2(n10643), .ZN(n10645) );
  NAND2_X1 U13684 ( .A1(n10646), .A2(n10645), .ZN(n19028) );
  INV_X1 U13685 ( .A(n19028), .ZN(n10647) );
  NAND2_X1 U13686 ( .A1(n10647), .A2(n15135), .ZN(n10666) );
  INV_X1 U13687 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10648) );
  NAND2_X1 U13688 ( .A1(n10666), .A2(n10648), .ZN(n15452) );
  AND4_X1 U13689 ( .A1(n15405), .A2(n15197), .A3(n15438), .A4(n15452), .ZN(
        n10653) );
  NAND2_X1 U13690 ( .A1(n9930), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10650) );
  OAI211_X1 U13691 ( .C1(n10651), .C2(n10650), .A(n10690), .B(n10649), .ZN(
        n19000) );
  OR2_X1 U13692 ( .A1(n19000), .A2(n11013), .ZN(n10652) );
  XNOR2_X1 U13693 ( .A(n10652), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15232) );
  NAND4_X1 U13694 ( .A1(n15190), .A2(n10654), .A3(n10653), .A4(n15232), .ZN(
        n10657) );
  NAND2_X1 U13695 ( .A1(n9930), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10655) );
  XNOR2_X1 U13696 ( .A(n10656), .B(n10655), .ZN(n18952) );
  AOI21_X1 U13697 ( .B1(n18952), .B2(n15135), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15212) );
  INV_X1 U13698 ( .A(n10658), .ZN(n10659) );
  NAND2_X1 U13699 ( .A1(n10659), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15406) );
  INV_X1 U13700 ( .A(n18962), .ZN(n10661) );
  AND2_X1 U13701 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10660) );
  NAND2_X1 U13702 ( .A1(n10661), .A2(n10660), .ZN(n15391) );
  NAND2_X1 U13703 ( .A1(n15406), .A2(n15391), .ZN(n15199) );
  INV_X1 U13704 ( .A(n10662), .ZN(n10663) );
  NAND2_X1 U13705 ( .A1(n10663), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15198) );
  NAND2_X1 U13706 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10664) );
  OR2_X1 U13707 ( .A1(n19000), .A2(n10664), .ZN(n15195) );
  NAND2_X1 U13708 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10665) );
  INV_X1 U13709 ( .A(n10666), .ZN(n10667) );
  NAND2_X1 U13710 ( .A1(n10667), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15453) );
  NAND4_X1 U13711 ( .A1(n15198), .A2(n15195), .A3(n15437), .A4(n15453), .ZN(
        n10668) );
  NOR2_X1 U13712 ( .A1(n15199), .A2(n10668), .ZN(n10672) );
  AND2_X1 U13713 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10669) );
  NAND2_X1 U13714 ( .A1(n18952), .A2(n10669), .ZN(n15210) );
  OR3_X1 U13715 ( .A1(n18940), .A2(n11013), .A3(n21096), .ZN(n15189) );
  INV_X1 U13716 ( .A(n10670), .ZN(n10671) );
  NAND2_X1 U13717 ( .A1(n10671), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16246) );
  AND4_X1 U13718 ( .A1(n10672), .A2(n15210), .A3(n15189), .A4(n16246), .ZN(
        n10673) );
  NAND2_X1 U13719 ( .A1(n10677), .A2(n10690), .ZN(n10674) );
  NAND2_X1 U13720 ( .A1(n9930), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10675) );
  INV_X1 U13721 ( .A(n10675), .ZN(n10676) );
  NAND2_X1 U13722 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  AND2_X1 U13723 ( .A1(n10683), .A2(n10678), .ZN(n15737) );
  NAND2_X1 U13724 ( .A1(n15737), .A2(n15135), .ZN(n10679) );
  INV_X1 U13725 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15357) );
  NOR2_X1 U13726 ( .A1(n10679), .A2(n15357), .ZN(n15178) );
  NAND2_X1 U13727 ( .A1(n9930), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10684) );
  XNOR2_X1 U13728 ( .A(n10683), .B(n10684), .ZN(n16186) );
  NAND2_X1 U13729 ( .A1(n16186), .A2(n15135), .ZN(n10680) );
  INV_X1 U13730 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15342) );
  XNOR2_X1 U13731 ( .A(n10680), .B(n15342), .ZN(n15350) );
  INV_X1 U13732 ( .A(n10680), .ZN(n10681) );
  NAND3_X1 U13733 ( .A1(n10685), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n9930), .ZN(
        n10686) );
  AND3_X1 U13734 ( .A1(n10689), .A2(n10690), .A3(n10686), .ZN(n16177) );
  NAND2_X1 U13735 ( .A1(n16177), .A2(n15135), .ZN(n10687) );
  INV_X1 U13736 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14308) );
  NOR2_X1 U13737 ( .A1(n10687), .A2(n14308), .ZN(n14301) );
  NAND2_X1 U13738 ( .A1(n10687), .A2(n14308), .ZN(n14299) );
  OAI21_X2 U13739 ( .B1(n14303), .B2(n14301), .A(n14299), .ZN(n15156) );
  INV_X1 U13740 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10925) );
  NOR3_X1 U13741 ( .A1(n10693), .A2(n10925), .A3(n14029), .ZN(n10688) );
  NAND2_X1 U13742 ( .A1(n10693), .A2(n10925), .ZN(n15132) );
  NAND3_X1 U13743 ( .A1(n10689), .A2(n9930), .A3(P2_EBX_REG_25__SCAN_IN), .ZN(
        n10691) );
  NAND2_X1 U13744 ( .A1(n10691), .A2(n10690), .ZN(n10692) );
  NOR2_X1 U13745 ( .A1(n10693), .A2(n10692), .ZN(n16165) );
  OR2_X1 U13746 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10697) );
  NAND2_X1 U13747 ( .A1(n9930), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10698) );
  INV_X1 U13748 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10937) );
  NOR2_X1 U13749 ( .A1(n14029), .A2(n10937), .ZN(n10703) );
  INV_X1 U13750 ( .A(n10703), .ZN(n10699) );
  XNOR2_X1 U13751 ( .A(n15134), .B(n10699), .ZN(n16134) );
  NAND2_X1 U13752 ( .A1(n16134), .A2(n15135), .ZN(n15139) );
  AND2_X1 U13753 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12626) );
  NAND3_X1 U13754 ( .A1(n16155), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15135), .ZN(n10702) );
  INV_X1 U13755 ( .A(n10700), .ZN(n10701) );
  INV_X1 U13756 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15322) );
  NAND2_X1 U13757 ( .A1(n10702), .A2(n15168), .ZN(n15130) );
  INV_X1 U13758 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10944) );
  NOR2_X1 U13759 ( .A1(n14029), .A2(n10944), .ZN(n10705) );
  INV_X1 U13760 ( .A(n10705), .ZN(n10704) );
  XNOR2_X1 U13761 ( .A(n10706), .B(n10704), .ZN(n16123) );
  AOI21_X1 U13762 ( .B1(n16123), .B2(n15135), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12621) );
  INV_X1 U13763 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10950) );
  NOR2_X1 U13764 ( .A1(n14029), .A2(n10950), .ZN(n10707) );
  XNOR2_X1 U13765 ( .A(n10709), .B(n10707), .ZN(n12732) );
  INV_X1 U13766 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15274) );
  OAI21_X1 U13767 ( .B1(n12732), .B2(n11013), .A(n15274), .ZN(n15120) );
  NOR3_X1 U13768 ( .A1(n12732), .A2(n11013), .A3(n15274), .ZN(n15119) );
  AND2_X1 U13769 ( .A1(n15135), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10708) );
  AOI211_X1 U13770 ( .C1(n15118), .C2(n15120), .A(n15119), .B(n15117), .ZN(
        n10715) );
  NOR2_X1 U13771 ( .A1(n10709), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10712) );
  INV_X1 U13772 ( .A(n10710), .ZN(n10711) );
  MUX2_X1 U13773 ( .A(n10712), .B(n10711), .S(n14029), .Z(n16113) );
  NAND2_X1 U13774 ( .A1(n16113), .A2(n15135), .ZN(n10713) );
  XNOR2_X1 U13775 ( .A(n10713), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10714) );
  XNOR2_X1 U13776 ( .A(n10715), .B(n10714), .ZN(n13475) );
  INV_X1 U13777 ( .A(n10716), .ZN(n10753) );
  OAI21_X1 U13778 ( .B1(n10718), .B2(n10753), .A(n10717), .ZN(n10726) );
  NAND2_X1 U13779 ( .A1(n10720), .A2(n10719), .ZN(n10759) );
  INV_X1 U13780 ( .A(n10759), .ZN(n10725) );
  NAND2_X1 U13781 ( .A1(n16376), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U13782 ( .A1(n10722), .A2(n10721), .ZN(n10724) );
  NAND2_X1 U13783 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15700), .ZN(
        n10723) );
  AOI21_X1 U13784 ( .B1(n10726), .B2(n10725), .A(n10763), .ZN(n19976) );
  AND2_X1 U13785 ( .A1(n19348), .A2(n19996), .ZN(n12726) );
  INV_X1 U13786 ( .A(n12726), .ZN(n10727) );
  NOR2_X1 U13787 ( .A1(n16383), .A2(n10727), .ZN(n19979) );
  NAND2_X1 U13788 ( .A1(n19976), .A2(n19979), .ZN(n10742) );
  NAND2_X1 U13789 ( .A1(n10729), .A2(n10747), .ZN(n10733) );
  XNOR2_X1 U13790 ( .A(n10753), .B(n10728), .ZN(n10746) );
  NAND2_X1 U13791 ( .A1(n10729), .A2(n10746), .ZN(n10730) );
  OR2_X1 U13792 ( .A1(n10759), .A2(n10730), .ZN(n10732) );
  INV_X1 U13793 ( .A(n10763), .ZN(n10731) );
  OAI21_X1 U13794 ( .B1(n10759), .B2(n10733), .A(n13514), .ZN(n10734) );
  NAND2_X1 U13795 ( .A1(n10734), .A2(n15803), .ZN(n10738) );
  NOR2_X1 U13796 ( .A1(n10735), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16380) );
  NAND2_X1 U13797 ( .A1(n16380), .A2(n11138), .ZN(n10737) );
  NOR2_X1 U13798 ( .A1(n15803), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n10736) );
  NAND2_X1 U13799 ( .A1(n10737), .A2(n10736), .ZN(n16401) );
  NAND2_X1 U13800 ( .A1(n10738), .A2(n16401), .ZN(n19977) );
  INV_X1 U13801 ( .A(n16383), .ZN(n10739) );
  NAND2_X1 U13802 ( .A1(n10739), .A2(n19997), .ZN(n10740) );
  NAND2_X1 U13803 ( .A1(n10742), .A2(n10741), .ZN(n13082) );
  NAND2_X1 U13804 ( .A1(n19994), .A2(n19997), .ZN(n10743) );
  NAND2_X1 U13805 ( .A1(n10743), .A2(n10749), .ZN(n10745) );
  AOI21_X1 U13806 ( .B1(n10745), .B2(n10744), .A(n10759), .ZN(n10757) );
  OAI21_X1 U13807 ( .B1(n19997), .B2(n10747), .A(n10746), .ZN(n10748) );
  OAI21_X1 U13808 ( .B1(n19997), .B2(n10749), .A(n10748), .ZN(n10750) );
  NAND2_X1 U13809 ( .A1(n10750), .A2(n16384), .ZN(n10755) );
  OAI21_X1 U13810 ( .B1(n10753), .B2(n10752), .A(n10751), .ZN(n10754) );
  NAND2_X1 U13811 ( .A1(n10755), .A2(n10754), .ZN(n10756) );
  AOI21_X1 U13812 ( .B1(n10757), .B2(n10756), .A(n10763), .ZN(n10758) );
  MUX2_X1 U13813 ( .A(n15700), .B(n10758), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n10762) );
  NAND2_X1 U13814 ( .A1(n10760), .A2(n10759), .ZN(n10761) );
  NAND2_X1 U13815 ( .A1(n16389), .A2(n19997), .ZN(n13771) );
  AOI21_X1 U13816 ( .B1(n10765), .B2(n16384), .A(n19364), .ZN(n10766) );
  NAND2_X1 U13817 ( .A1(n13771), .A2(n10766), .ZN(n10786) );
  NAND2_X1 U13818 ( .A1(n10768), .A2(n10218), .ZN(n10769) );
  NAND2_X1 U13819 ( .A1(n10767), .A2(n10769), .ZN(n10781) );
  NAND2_X1 U13820 ( .A1(n10771), .A2(n10770), .ZN(n10772) );
  NAND2_X1 U13821 ( .A1(n10772), .A2(n15558), .ZN(n10773) );
  NAND2_X1 U13822 ( .A1(n10773), .A2(n12726), .ZN(n11199) );
  NAND2_X1 U13823 ( .A1(n19348), .A2(n10774), .ZN(n11194) );
  INV_X1 U13824 ( .A(n15558), .ZN(n13447) );
  AOI21_X1 U13825 ( .B1(n11194), .B2(n16384), .A(n13447), .ZN(n10775) );
  OR2_X1 U13826 ( .A1(n10775), .A2(n10205), .ZN(n10776) );
  AND2_X1 U13827 ( .A1(n11199), .A2(n10776), .ZN(n10780) );
  AND2_X1 U13828 ( .A1(n10778), .A2(n10777), .ZN(n10779) );
  NAND3_X1 U13829 ( .A1(n10781), .A2(n10780), .A3(n10779), .ZN(n11195) );
  NAND2_X1 U13830 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19993) );
  INV_X1 U13831 ( .A(n19993), .ZN(n19864) );
  INV_X1 U13832 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19851) );
  INV_X1 U13833 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19872) );
  NOR2_X1 U13834 ( .A1(n19851), .A2(n19872), .ZN(n19863) );
  NOR2_X1 U13835 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19866) );
  NOR3_X1 U13836 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19863), .A3(n19866), 
        .ZN(n19995) );
  INV_X1 U13837 ( .A(n19995), .ZN(n19858) );
  NOR2_X1 U13838 ( .A1(n19864), .A2(n19858), .ZN(n13511) );
  AND3_X1 U13839 ( .A1(n16398), .A2(n13514), .A3(n13511), .ZN(n10783) );
  NOR2_X1 U13840 ( .A1(n11195), .A2(n10783), .ZN(n13767) );
  MUX2_X1 U13841 ( .A(n16398), .B(n10205), .S(n19348), .Z(n10784) );
  NAND3_X1 U13842 ( .A1(n10784), .A2(n13514), .A3(n19993), .ZN(n10785) );
  NAND3_X1 U13843 ( .A1(n10786), .A2(n13767), .A3(n10785), .ZN(n10789) );
  NAND2_X1 U13844 ( .A1(n10205), .A2(n13511), .ZN(n10787) );
  NOR2_X1 U13845 ( .A1(n13771), .A2(n10787), .ZN(n10788) );
  AND2_X1 U13846 ( .A1(n15803), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12730) );
  NAND2_X1 U13847 ( .A1(n13475), .A2(n16344), .ZN(n11240) );
  INV_X1 U13848 ( .A(n10793), .ZN(n10791) );
  NAND2_X1 U13849 ( .A1(n16355), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16354) );
  INV_X1 U13850 ( .A(n16354), .ZN(n10795) );
  XOR2_X1 U13851 ( .A(n10982), .B(n10794), .Z(n10796) );
  NAND2_X1 U13852 ( .A1(n10795), .A2(n10796), .ZN(n10797) );
  XNOR2_X1 U13853 ( .A(n10796), .B(n16354), .ZN(n13532) );
  NAND2_X1 U13854 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13532), .ZN(
        n13531) );
  NAND2_X1 U13855 ( .A1(n10797), .A2(n13531), .ZN(n10799) );
  XNOR2_X1 U13856 ( .A(n11221), .B(n10799), .ZN(n13675) );
  XNOR2_X1 U13857 ( .A(n10798), .B(n10989), .ZN(n13674) );
  NAND2_X1 U13858 ( .A1(n13675), .A2(n13674), .ZN(n13673) );
  NAND2_X1 U13859 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10799), .ZN(
        n10800) );
  NAND2_X1 U13860 ( .A1(n13673), .A2(n10800), .ZN(n10801) );
  INV_X1 U13861 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20944) );
  XNOR2_X1 U13862 ( .A(n10801), .B(n20944), .ZN(n13916) );
  NAND2_X1 U13863 ( .A1(n13917), .A2(n13916), .ZN(n10803) );
  NAND2_X1 U13864 ( .A1(n10801), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10802) );
  OAI21_X1 U13865 ( .B1(n19292), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n19294), .ZN(n10805) );
  NAND2_X1 U13866 ( .A1(n19292), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10804) );
  NAND2_X1 U13867 ( .A1(n10805), .A2(n10804), .ZN(n14136) );
  INV_X1 U13868 ( .A(n10806), .ZN(n10813) );
  INV_X1 U13869 ( .A(n14139), .ZN(n10810) );
  INV_X1 U13870 ( .A(n10808), .ZN(n10809) );
  NAND2_X1 U13871 ( .A1(n10810), .A2(n10809), .ZN(n10811) );
  NAND2_X1 U13872 ( .A1(n14246), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14245) );
  NAND2_X1 U13873 ( .A1(n10812), .A2(n14139), .ZN(n10814) );
  NAND2_X1 U13874 ( .A1(n10814), .A2(n10813), .ZN(n10815) );
  NAND2_X1 U13875 ( .A1(n10816), .A2(n11013), .ZN(n10817) );
  NAND2_X1 U13876 ( .A1(n10820), .A2(n10817), .ZN(n14265) );
  XNOR2_X1 U13877 ( .A(n10820), .B(n16324), .ZN(n15264) );
  NAND2_X1 U13878 ( .A1(n10819), .A2(n10818), .ZN(n15267) );
  INV_X1 U13879 ( .A(n10820), .ZN(n10821) );
  NAND2_X1 U13880 ( .A1(n10821), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10822) );
  NAND2_X1 U13881 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15478) );
  INV_X1 U13882 ( .A(n15478), .ZN(n10823) );
  AND2_X1 U13883 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n10823), .ZN(
        n15458) );
  AND2_X1 U13884 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10824) );
  NAND2_X1 U13885 ( .A1(n15458), .A2(n10824), .ZN(n16286) );
  INV_X1 U13886 ( .A(n16286), .ZN(n11213) );
  AND2_X1 U13887 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15433) );
  AND2_X1 U13888 ( .A1(n15433), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11226) );
  AND2_X1 U13889 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11227) );
  INV_X1 U13890 ( .A(n11227), .ZN(n15207) );
  OR2_X1 U13891 ( .A1(n15207), .A2(n21096), .ZN(n10825) );
  NOR2_X2 U13892 ( .A1(n15205), .A2(n10825), .ZN(n15180) );
  NAND2_X1 U13893 ( .A1(n15180), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15182) );
  NOR2_X2 U13894 ( .A1(n15182), .A2(n15342), .ZN(n14304) );
  NAND2_X1 U13895 ( .A1(n14304), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14305) );
  NOR2_X2 U13896 ( .A1(n14305), .A2(n15322), .ZN(n15159) );
  INV_X1 U13897 ( .A(n12626), .ZN(n15288) );
  XNOR2_X1 U13898 ( .A(n10826), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13481) );
  NAND2_X1 U13899 ( .A1(n11211), .A2(n19979), .ZN(n19343) );
  OR2_X1 U13900 ( .A1(n13481), .A2(n19343), .ZN(n11239) );
  INV_X1 U13901 ( .A(n10828), .ZN(n10829) );
  NOR2_X2 U13902 ( .A1(n11220), .A2(n10829), .ZN(n19338) );
  INV_X1 U13903 ( .A(n10896), .ZN(n10881) );
  OR2_X1 U13904 ( .A1(n10896), .A2(n10831), .ZN(n10838) );
  INV_X1 U13905 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10832) );
  OR2_X1 U13906 ( .A1(n10956), .A2(n10832), .ZN(n10834) );
  NAND2_X1 U13907 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10833) );
  OAI211_X1 U13908 ( .C1(n10951), .C2(n10835), .A(n10834), .B(n10833), .ZN(
        n10836) );
  INV_X1 U13909 ( .A(n10836), .ZN(n10837) );
  NAND2_X1 U13910 ( .A1(n10838), .A2(n10837), .ZN(n13688) );
  INV_X1 U13911 ( .A(n10841), .ZN(n10843) );
  AOI22_X1 U13912 ( .A1(n10909), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10846) );
  OAI21_X1 U13913 ( .B1(n10951), .B2(n20945), .A(n10846), .ZN(n10847) );
  AOI21_X1 U13914 ( .B1(n10881), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10847), .ZN(n13740) );
  INV_X1 U13915 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13854) );
  OR2_X1 U13916 ( .A1(n10896), .A2(n14254), .ZN(n10849) );
  AOI22_X1 U13917 ( .A1(n10909), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10848) );
  OAI211_X1 U13918 ( .C1(n13854), .C2(n10951), .A(n10849), .B(n10848), .ZN(
        n13849) );
  OR2_X1 U13919 ( .A1(n10896), .A2(n16337), .ZN(n10851) );
  AOI22_X1 U13920 ( .A1(n10909), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10850) );
  OAI211_X1 U13921 ( .C1(n10951), .C2(n13747), .A(n10851), .B(n10850), .ZN(
        n13746) );
  OR2_X1 U13922 ( .A1(n10896), .A2(n16324), .ZN(n10853) );
  AOI22_X1 U13923 ( .A1(n10909), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10852) );
  OAI211_X1 U13924 ( .C1(n10854), .C2(n10951), .A(n10853), .B(n10852), .ZN(
        n13889) );
  OR2_X1 U13925 ( .A1(n10896), .A2(n15493), .ZN(n10860) );
  INV_X1 U13926 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10857) );
  INV_X1 U13927 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15253) );
  OR2_X1 U13928 ( .A1(n10956), .A2(n15253), .ZN(n10856) );
  NAND2_X1 U13929 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10855) );
  OAI211_X1 U13930 ( .C1(n10951), .C2(n10857), .A(n10856), .B(n10855), .ZN(
        n10858) );
  INV_X1 U13931 ( .A(n10858), .ZN(n10859) );
  OR2_X1 U13932 ( .A1(n10896), .A2(n16269), .ZN(n10862) );
  AOI22_X1 U13933 ( .A1(n10909), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10861) );
  OAI211_X1 U13934 ( .C1(n13994), .C2(n10951), .A(n10862), .B(n10861), .ZN(
        n13989) );
  OR2_X1 U13935 ( .A1(n10896), .A2(n10612), .ZN(n10864) );
  AOI22_X1 U13936 ( .A1(n10909), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10863) );
  OAI211_X1 U13937 ( .C1(n13948), .C2(n10951), .A(n10864), .B(n10863), .ZN(
        n13946) );
  INV_X1 U13938 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13939 ( .A1(n10909), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10865) );
  OAI21_X1 U13940 ( .B1(n10951), .B2(n10866), .A(n10865), .ZN(n10867) );
  AOI21_X1 U13941 ( .B1(n10881), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10867), .ZN(n14062) );
  NAND2_X1 U13942 ( .A1(n10881), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10869) );
  AOI22_X1 U13943 ( .A1(n10909), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10868) );
  OAI211_X1 U13944 ( .C1(n10870), .C2(n10951), .A(n10869), .B(n10868), .ZN(
        n14026) );
  OR2_X1 U13945 ( .A1(n10896), .A2(n16251), .ZN(n10873) );
  AOI22_X1 U13946 ( .A1(n10909), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10872) );
  NAND2_X1 U13947 ( .A1(n10959), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10871) );
  INV_X1 U13948 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10877) );
  OR2_X1 U13949 ( .A1(n10896), .A2(n10874), .ZN(n10876) );
  AOI22_X1 U13950 ( .A1(n10909), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10875) );
  OAI211_X1 U13951 ( .C1(n10877), .C2(n10951), .A(n10876), .B(n10875), .ZN(
        n14186) );
  AOI22_X1 U13952 ( .A1(n10909), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10878) );
  OAI21_X1 U13953 ( .B1(n10951), .B2(n10879), .A(n10878), .ZN(n10880) );
  AOI21_X1 U13954 ( .B1(n10881), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10880), .ZN(n14209) );
  INV_X1 U13955 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10885) );
  OR2_X1 U13956 ( .A1(n10896), .A2(n10882), .ZN(n10884) );
  AOI22_X1 U13957 ( .A1(n10909), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10883) );
  OAI211_X1 U13958 ( .C1(n10885), .C2(n10951), .A(n10884), .B(n10883), .ZN(
        n14228) );
  OR2_X1 U13959 ( .A1(n10896), .A2(n15417), .ZN(n10892) );
  INV_X1 U13960 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10889) );
  INV_X1 U13961 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n10886) );
  OR2_X1 U13962 ( .A1(n10956), .A2(n10886), .ZN(n10888) );
  NAND2_X1 U13963 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10887) );
  OAI211_X1 U13964 ( .C1(n10951), .C2(n10889), .A(n10888), .B(n10887), .ZN(
        n10890) );
  INV_X1 U13965 ( .A(n10890), .ZN(n10891) );
  NAND2_X1 U13966 ( .A1(n10892), .A2(n10891), .ZN(n14274) );
  INV_X1 U13967 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10895) );
  OR2_X1 U13968 ( .A1(n10896), .A2(n20966), .ZN(n10894) );
  AOI22_X1 U13969 ( .A1(n10909), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10893) );
  OAI211_X1 U13970 ( .C1(n10895), .C2(n10951), .A(n10894), .B(n10893), .ZN(
        n15038) );
  INV_X1 U13971 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15035) );
  INV_X1 U13972 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15378) );
  OR2_X1 U13973 ( .A1(n10896), .A2(n15378), .ZN(n10898) );
  AOI22_X1 U13974 ( .A1(n10909), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10897) );
  OAI211_X1 U13975 ( .C1(n15035), .C2(n10951), .A(n10898), .B(n10897), .ZN(
        n15030) );
  OR2_X1 U13976 ( .A1(n10896), .A2(n21096), .ZN(n10901) );
  INV_X1 U13977 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19906) );
  INV_X1 U13978 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18941) );
  OAI22_X1 U13979 ( .A1(n10956), .A2(n19906), .B1(n15803), .B2(n18941), .ZN(
        n10899) );
  INV_X1 U13980 ( .A(n10899), .ZN(n10900) );
  OAI211_X1 U13981 ( .C1(n18942), .C2(n10951), .A(n10901), .B(n10900), .ZN(
        n15024) );
  OR2_X1 U13982 ( .A1(n10896), .A2(n15357), .ZN(n10908) );
  INV_X1 U13983 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10905) );
  INV_X1 U13984 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10902) );
  OR2_X1 U13985 ( .A1(n10956), .A2(n10902), .ZN(n10904) );
  NAND2_X1 U13986 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10903) );
  OAI211_X1 U13987 ( .C1(n10951), .C2(n10905), .A(n10904), .B(n10903), .ZN(
        n10906) );
  INV_X1 U13988 ( .A(n10906), .ZN(n10907) );
  INV_X1 U13989 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10912) );
  OR2_X1 U13990 ( .A1(n10896), .A2(n15342), .ZN(n10911) );
  AOI22_X1 U13991 ( .A1(n10909), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10910) );
  OAI211_X1 U13992 ( .C1(n10951), .C2(n10912), .A(n10911), .B(n10910), .ZN(
        n15012) );
  OR2_X1 U13993 ( .A1(n10896), .A2(n14308), .ZN(n10917) );
  INV_X1 U13994 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19911) );
  OR2_X1 U13995 ( .A1(n10956), .A2(n19911), .ZN(n10914) );
  NAND2_X1 U13996 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10913) );
  OAI211_X1 U13997 ( .C1(n10951), .C2(n9810), .A(n10914), .B(n10913), .ZN(
        n10915) );
  INV_X1 U13998 ( .A(n10915), .ZN(n10916) );
  OR2_X1 U13999 ( .A1(n10896), .A2(n15322), .ZN(n10922) );
  INV_X1 U14000 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14998) );
  INV_X1 U14001 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19913) );
  OR2_X1 U14002 ( .A1(n10956), .A2(n19913), .ZN(n10919) );
  NAND2_X1 U14003 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10918) );
  OAI211_X1 U14004 ( .C1(n10951), .C2(n14998), .A(n10919), .B(n10918), .ZN(
        n10920) );
  INV_X1 U14005 ( .A(n10920), .ZN(n10921) );
  NAND2_X1 U14006 ( .A1(n10922), .A2(n10921), .ZN(n14996) );
  NAND2_X1 U14007 ( .A1(n14309), .A2(n14996), .ZN(n14987) );
  INV_X1 U14008 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15323) );
  OR2_X1 U14009 ( .A1(n10896), .A2(n15323), .ZN(n10928) );
  INV_X1 U14010 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15162) );
  OR2_X1 U14011 ( .A1(n10956), .A2(n15162), .ZN(n10924) );
  NAND2_X1 U14012 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10923) );
  OAI211_X1 U14013 ( .C1(n10951), .C2(n10925), .A(n10924), .B(n10923), .ZN(
        n10926) );
  INV_X1 U14014 ( .A(n10926), .ZN(n10927) );
  AND2_X1 U14015 ( .A1(n10928), .A2(n10927), .ZN(n14988) );
  INV_X1 U14016 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15152) );
  OR2_X1 U14017 ( .A1(n10896), .A2(n15152), .ZN(n10934) );
  INV_X1 U14018 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10931) );
  INV_X1 U14019 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19918) );
  OR2_X1 U14020 ( .A1(n10956), .A2(n19918), .ZN(n10930) );
  NAND2_X1 U14021 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10929) );
  OAI211_X1 U14022 ( .C1(n10951), .C2(n10931), .A(n10930), .B(n10929), .ZN(
        n10932) );
  INV_X1 U14023 ( .A(n10932), .ZN(n10933) );
  AND2_X1 U14024 ( .A1(n10934), .A2(n10933), .ZN(n14978) );
  INV_X1 U14025 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15142) );
  OR2_X1 U14026 ( .A1(n10896), .A2(n15142), .ZN(n10940) );
  INV_X1 U14027 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19919) );
  OR2_X1 U14028 ( .A1(n10956), .A2(n19919), .ZN(n10936) );
  NAND2_X1 U14029 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10935) );
  OAI211_X1 U14030 ( .C1(n10951), .C2(n10937), .A(n10936), .B(n10935), .ZN(
        n10938) );
  INV_X1 U14031 ( .A(n10938), .ZN(n10939) );
  AND2_X1 U14032 ( .A1(n10940), .A2(n10939), .ZN(n14969) );
  INV_X1 U14033 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10941) );
  OR2_X1 U14034 ( .A1(n10896), .A2(n10941), .ZN(n10947) );
  INV_X1 U14035 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19921) );
  OR2_X1 U14036 ( .A1(n10956), .A2(n19921), .ZN(n10943) );
  NAND2_X1 U14037 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10942) );
  OAI211_X1 U14038 ( .C1(n10951), .C2(n10944), .A(n10943), .B(n10942), .ZN(
        n10945) );
  INV_X1 U14039 ( .A(n10945), .ZN(n10946) );
  NAND2_X1 U14040 ( .A1(n10947), .A2(n10946), .ZN(n12632) );
  OR2_X1 U14041 ( .A1(n10896), .A2(n15274), .ZN(n10954) );
  INV_X1 U14042 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19925) );
  OR2_X1 U14043 ( .A1(n10956), .A2(n19925), .ZN(n10949) );
  NAND2_X1 U14044 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10948) );
  OAI211_X1 U14045 ( .C1(n10951), .C2(n10950), .A(n10949), .B(n10948), .ZN(
        n10952) );
  INV_X1 U14046 ( .A(n10952), .ZN(n10953) );
  AND2_X1 U14047 ( .A1(n10954), .A2(n10953), .ZN(n12742) );
  INV_X1 U14048 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n10955) );
  INV_X1 U14049 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15803) );
  OAI22_X1 U14050 ( .A1(n10956), .A2(n10955), .B1(n15803), .B2(n9967), .ZN(
        n10958) );
  NOR2_X1 U14051 ( .A1(n10896), .A2(n9971), .ZN(n10957) );
  AOI211_X1 U14052 ( .C1(n10959), .C2(P2_EBX_REG_31__SCAN_IN), .A(n10958), .B(
        n10957), .ZN(n10960) );
  XNOR2_X1 U14053 ( .A(n10961), .B(n10960), .ZN(n16116) );
  INV_X1 U14054 ( .A(n16116), .ZN(n11238) );
  NOR2_X1 U14055 ( .A1(n15558), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14056 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n10965) );
  NAND2_X1 U14057 ( .A1(n11160), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U14058 ( .A1(n10965), .A2(n10964), .ZN(n15086) );
  AND2_X2 U14059 ( .A1(n19348), .A2(n9674), .ZN(n10967) );
  INV_X1 U14060 ( .A(n10966), .ZN(n11011) );
  INV_X1 U14061 ( .A(n10967), .ZN(n11012) );
  INV_X1 U14062 ( .A(n10969), .ZN(n13446) );
  NAND2_X1 U14063 ( .A1(n10978), .A2(n13446), .ZN(n10991) );
  OAI22_X1 U14064 ( .A1(n15558), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19973), 
        .B2(n19986), .ZN(n10970) );
  INV_X1 U14065 ( .A(n10970), .ZN(n10971) );
  AND2_X1 U14066 ( .A1(n10991), .A2(n10971), .ZN(n10972) );
  NAND2_X1 U14067 ( .A1(n11160), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U14068 ( .A1(n13447), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10974) );
  OAI211_X1 U14069 ( .C1(n19348), .C2(n16351), .A(n10974), .B(n19950), .ZN(
        n10975) );
  INV_X1 U14070 ( .A(n10975), .ZN(n10976) );
  AOI22_X1 U14071 ( .A1(n10978), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n10995), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n10980) );
  INV_X1 U14072 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19874) );
  NAND2_X1 U14073 ( .A1(n11160), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10979) );
  NAND2_X1 U14074 ( .A1(n10980), .A2(n10979), .ZN(n10988) );
  INV_X1 U14075 ( .A(n10988), .ZN(n10981) );
  OR2_X1 U14076 ( .A1(n10982), .A2(n11012), .ZN(n10986) );
  AND2_X1 U14077 ( .A1(n15558), .A2(n19950), .ZN(n10984) );
  NOR2_X1 U14078 ( .A1(n10498), .A2(n19950), .ZN(n10983) );
  AOI21_X1 U14079 ( .B1(n10969), .B2(n10984), .A(n10983), .ZN(n10985) );
  NAND2_X1 U14080 ( .A1(n10986), .A2(n10985), .ZN(n13606) );
  INV_X1 U14081 ( .A(n13606), .ZN(n10987) );
  NAND2_X1 U14082 ( .A1(n10967), .A2(n10989), .ZN(n10990) );
  OAI211_X1 U14083 ( .C1(n19986), .C2(n19957), .A(n10991), .B(n10990), .ZN(
        n10992) );
  AND3_X1 U14084 ( .A1(n13609), .A2(n10993), .A3(n10992), .ZN(n10994) );
  AOI22_X1 U14085 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U14086 ( .A1(n11160), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10996) );
  NAND2_X1 U14087 ( .A1(n10997), .A2(n10996), .ZN(n13666) );
  NAND2_X1 U14088 ( .A1(n11160), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14089 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11001) );
  AOI22_X1 U14090 ( .A1(n10967), .A2(n10999), .B1(n11187), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n11000) );
  NAND3_X1 U14091 ( .A1(n11002), .A2(n11001), .A3(n11000), .ZN(n13931) );
  NAND2_X1 U14092 ( .A1(n11160), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U14093 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11005) );
  NAND2_X1 U14094 ( .A1(n10967), .A2(n11003), .ZN(n11004) );
  AOI22_X1 U14095 ( .A1(n11160), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n10967), 
        .B2(n11007), .ZN(n11009) );
  AOI22_X1 U14096 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U14097 ( .A1(n11009), .A2(n11008), .ZN(n14142) );
  NAND2_X1 U14098 ( .A1(n14143), .A2(n14142), .ZN(n14141) );
  INV_X1 U14099 ( .A(n14141), .ZN(n11010) );
  AOI21_X1 U14100 ( .B1(n10967), .B2(n11011), .A(n11010), .ZN(n14250) );
  AOI222_X1 U14101 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n11160), .B1(n11184), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n11187), .ZN(n14249) );
  AOI22_X1 U14102 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U14103 ( .A1(n11160), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11014) );
  NAND2_X1 U14104 ( .A1(n11015), .A2(n11014), .ZN(n16340) );
  INV_X1 U14105 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11016) );
  OAI22_X1 U14106 ( .A1(n11130), .A2(n15590), .B1(n11138), .B2(n11016), .ZN(
        n11019) );
  INV_X1 U14107 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n19381) );
  OAI22_X1 U14108 ( .A1(n11137), .A2(n11017), .B1(n11132), .B2(n19381), .ZN(
        n11018) );
  NOR2_X1 U14109 ( .A1(n11019), .A2(n11018), .ZN(n11034) );
  INV_X1 U14110 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11020) );
  OAI22_X1 U14111 ( .A1(n11131), .A2(n11020), .B1(n11133), .B2(n12817), .ZN(
        n11023) );
  OAI22_X1 U14112 ( .A1(n11143), .A2(n15575), .B1(n11141), .B2(n11021), .ZN(
        n11022) );
  NOR2_X1 U14113 ( .A1(n11023), .A2(n11022), .ZN(n11033) );
  AOI22_X1 U14114 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12924), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14115 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11026) );
  OR2_X1 U14116 ( .A1(n11087), .A2(n14023), .ZN(n11025) );
  NAND2_X1 U14117 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11024) );
  NAND4_X1 U14118 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11031) );
  OAI22_X1 U14119 ( .A1(n12882), .A2(n11029), .B1(n13779), .B2(n11028), .ZN(
        n11030) );
  NOR2_X1 U14120 ( .A1(n11031), .A2(n11030), .ZN(n11032) );
  AOI22_X1 U14121 ( .A1(n11160), .A2(P2_REIP_REG_8__SCAN_IN), .B1(n10967), 
        .B2(n10090), .ZN(n11036) );
  AOI22_X1 U14122 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14123 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12914), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14124 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12911), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14125 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U14126 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11037) );
  NAND4_X1 U14127 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(
        n11049) );
  AOI22_X1 U14128 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11047) );
  NAND2_X1 U14129 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11042) );
  NAND2_X1 U14130 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11041) );
  OAI211_X1 U14131 ( .C1(n11087), .C2(n12949), .A(n11042), .B(n11041), .ZN(
        n11043) );
  INV_X1 U14132 ( .A(n11043), .ZN(n11046) );
  AOI22_X1 U14133 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U14134 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11044) );
  NAND4_X1 U14135 ( .A1(n11047), .A2(n11046), .A3(n11045), .A4(n11044), .ZN(
        n11048) );
  AOI22_X1 U14136 ( .A1(n11160), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n10967), 
        .B2(n13896), .ZN(n11051) );
  AOI22_X1 U14137 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11050) );
  NAND2_X1 U14138 ( .A1(n11051), .A2(n11050), .ZN(n15490) );
  NAND2_X1 U14139 ( .A1(n11160), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14140 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14141 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12912), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14142 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12914), .B1(
        n12916), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14143 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14144 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11052) );
  NAND4_X1 U14145 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11064) );
  AOI22_X1 U14146 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U14147 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11057) );
  NAND2_X1 U14148 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11056) );
  OAI211_X1 U14149 ( .C1(n11087), .C2(n12975), .A(n11057), .B(n11056), .ZN(
        n11058) );
  INV_X1 U14150 ( .A(n11058), .ZN(n11061) );
  AOI22_X1 U14151 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11060) );
  NAND2_X1 U14152 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11059) );
  NAND4_X1 U14153 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(
        n11063) );
  NAND2_X1 U14154 ( .A1(n10967), .A2(n13987), .ZN(n11065) );
  AOI22_X1 U14155 ( .A1(n11160), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11187), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14156 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12914), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14157 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12911), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14158 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14159 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11068) );
  NAND4_X1 U14160 ( .A1(n11071), .A2(n11070), .A3(n11069), .A4(n11068), .ZN(
        n11080) );
  AOI22_X1 U14161 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U14162 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11073) );
  NAND2_X1 U14163 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11072) );
  OAI211_X1 U14164 ( .C1(n11087), .C2(n13001), .A(n11073), .B(n11072), .ZN(
        n11074) );
  INV_X1 U14165 ( .A(n11074), .ZN(n11077) );
  AOI22_X1 U14166 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U14167 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11075) );
  NAND4_X1 U14168 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11079) );
  AOI22_X1 U14169 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n11184), .B1(
        n10967), .B2(n14064), .ZN(n11081) );
  NAND2_X1 U14170 ( .A1(n11082), .A2(n11081), .ZN(n15476) );
  AOI22_X1 U14171 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12916), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14172 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12911), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14173 ( .A1(n12914), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14174 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11083) );
  NAND4_X1 U14175 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11096) );
  AOI22_X1 U14176 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U14177 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14178 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11088) );
  OAI211_X1 U14179 ( .C1(n11087), .C2(n13023), .A(n11089), .B(n11088), .ZN(
        n11090) );
  INV_X1 U14180 ( .A(n11090), .ZN(n11093) );
  AOI22_X1 U14181 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12930), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U14182 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11091) );
  NAND4_X1 U14183 ( .A1(n11094), .A2(n11093), .A3(n11092), .A4(n11091), .ZN(
        n11095) );
  AOI22_X1 U14184 ( .A1(n11160), .A2(P2_REIP_REG_12__SCAN_IN), .B1(n10967), 
        .B2(n14063), .ZN(n11098) );
  AOI22_X1 U14185 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14186 ( .A1(n11160), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11184), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14187 ( .A1(n12914), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14188 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14189 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14190 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11099) );
  NAND4_X1 U14191 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n11111) );
  AOI22_X1 U14192 ( .A1(n12921), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12922), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U14193 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11104) );
  NAND2_X1 U14194 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11103) );
  OAI211_X1 U14195 ( .C1(n11087), .C2(n14032), .A(n11104), .B(n11103), .ZN(
        n11105) );
  INV_X1 U14196 ( .A(n11105), .ZN(n11108) );
  AOI22_X1 U14197 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11107) );
  NAND2_X1 U14198 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11106) );
  NAND4_X1 U14199 ( .A1(n11109), .A2(n11108), .A3(n11107), .A4(n11106), .ZN(
        n11110) );
  AOI22_X1 U14200 ( .A1(n10967), .A2(n14084), .B1(n11187), .B2(
        P2_EAX_REG_13__SCAN_IN), .ZN(n11112) );
  NAND2_X1 U14201 ( .A1(n11113), .A2(n11112), .ZN(n15457) );
  AOI22_X1 U14202 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12909), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14203 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12910), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14204 ( .A1(n12914), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14205 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12916), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11114) );
  NAND4_X1 U14206 ( .A1(n11117), .A2(n11116), .A3(n11115), .A4(n11114), .ZN(
        n11126) );
  AOI22_X1 U14207 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U14208 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11119) );
  NAND2_X1 U14209 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11118) );
  OAI211_X1 U14210 ( .C1(n11087), .C2(n13062), .A(n11119), .B(n11118), .ZN(
        n11120) );
  INV_X1 U14211 ( .A(n11120), .ZN(n11123) );
  AOI22_X1 U14212 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12930), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U14213 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11121) );
  NAND4_X1 U14214 ( .A1(n11124), .A2(n11123), .A3(n11122), .A4(n11121), .ZN(
        n11125) );
  AOI22_X1 U14215 ( .A1(n11160), .A2(P2_REIP_REG_14__SCAN_IN), .B1(n10967), 
        .B2(n14086), .ZN(n11128) );
  AOI22_X1 U14216 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14217 ( .A1(n11160), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11184), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11159) );
  OAI22_X1 U14218 ( .A1(n13427), .A2(n11131), .B1(n11130), .B2(n11129), .ZN(
        n11135) );
  INV_X1 U14219 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15564) );
  OAI22_X1 U14220 ( .A1(n11133), .A2(n12927), .B1(n11132), .B2(n15564), .ZN(
        n11134) );
  NOR2_X1 U14221 ( .A1(n11135), .A2(n11134), .ZN(n11156) );
  INV_X1 U14222 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11139) );
  OAI22_X1 U14223 ( .A1(n11139), .A2(n11138), .B1(n11137), .B2(n11136), .ZN(
        n11145) );
  OAI22_X1 U14224 ( .A1(n11143), .A2(n11142), .B1(n11141), .B2(n11140), .ZN(
        n11144) );
  NOR2_X1 U14225 ( .A1(n11145), .A2(n11144), .ZN(n11155) );
  AOI22_X1 U14226 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12923), .B1(
        n12924), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14227 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11148) );
  OR2_X1 U14228 ( .A1(n11087), .A2(n13424), .ZN(n11147) );
  NAND2_X1 U14229 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11146) );
  NAND4_X1 U14230 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11153) );
  OAI22_X1 U14231 ( .A1(n11151), .A2(n13779), .B1(n12882), .B2(n11150), .ZN(
        n11152) );
  NOR2_X1 U14232 ( .A1(n11153), .A2(n11152), .ZN(n11154) );
  INV_X1 U14233 ( .A(n14204), .ZN(n11157) );
  AOI22_X1 U14234 ( .A1(n10967), .A2(n11157), .B1(n11187), .B2(
        P2_EAX_REG_15__SCAN_IN), .ZN(n11158) );
  NAND2_X1 U14235 ( .A1(n11159), .A2(n11158), .ZN(n15445) );
  AOI222_X1 U14236 ( .A1(n11160), .A2(P2_REIP_REG_16__SCAN_IN), .B1(n11184), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n11187), .C2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U14237 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U14238 ( .A1(n11160), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14239 ( .A1(n11162), .A2(n11161), .ZN(n14196) );
  NAND2_X1 U14240 ( .A1(n11160), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14241 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14242 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11166) );
  NAND2_X1 U14243 ( .A1(n11160), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U14244 ( .A1(n11166), .A2(n11165), .ZN(n15106) );
  AOI22_X1 U14245 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11168) );
  NAND2_X1 U14246 ( .A1(n11160), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U14247 ( .A1(n11168), .A2(n11167), .ZN(n15379) );
  AND2_X2 U14248 ( .A1(n15105), .A2(n15379), .ZN(n15381) );
  AOI22_X1 U14249 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U14250 ( .A1(n11160), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11169) );
  NAND2_X1 U14251 ( .A1(n11170), .A2(n11169), .ZN(n15095) );
  AOI222_X1 U14252 ( .A1(n11160), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n11184), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n11187), .C2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15360) );
  NAND2_X1 U14253 ( .A1(n11160), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14254 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11171) );
  AND2_X1 U14255 ( .A1(n11172), .A2(n11171), .ZN(n14313) );
  AOI22_X1 U14256 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U14257 ( .A1(n11160), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U14258 ( .A1(n11174), .A2(n11173), .ZN(n15073) );
  NAND2_X1 U14259 ( .A1(n14312), .A2(n15073), .ZN(n15065) );
  NAND2_X1 U14260 ( .A1(n11160), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14261 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11175) );
  AND2_X1 U14262 ( .A1(n11176), .A2(n11175), .ZN(n15067) );
  INV_X1 U14263 ( .A(n15067), .ZN(n11177) );
  NAND2_X1 U14264 ( .A1(n11160), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14265 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11178) );
  AND2_X1 U14266 ( .A1(n11179), .A2(n11178), .ZN(n15052) );
  NAND2_X1 U14267 ( .A1(n11160), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14268 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n11180) );
  AND2_X1 U14269 ( .A1(n11181), .A2(n11180), .ZN(n15046) );
  AOI22_X1 U14270 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11183) );
  NAND2_X1 U14271 ( .A1(n11160), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U14272 ( .A1(n11183), .A2(n11182), .ZN(n12630) );
  AOI22_X1 U14273 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n11187), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U14274 ( .A1(n11160), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14275 ( .A1(n11186), .A2(n11185), .ZN(n12720) );
  NAND2_X1 U14276 ( .A1(n12629), .A2(n12720), .ZN(n12724) );
  AOI222_X1 U14277 ( .A1(n11160), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11184), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n11187), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U14278 ( .A1(n11189), .A2(n19997), .ZN(n11192) );
  NAND2_X1 U14279 ( .A1(n11191), .A2(n11190), .ZN(n13777) );
  NAND2_X1 U14280 ( .A1(n11192), .A2(n13777), .ZN(n11193) );
  NAND2_X1 U14281 ( .A1(n11211), .A2(n11193), .ZN(n19330) );
  NOR2_X2 U14282 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19938) );
  NAND2_X1 U14283 ( .A1(n19938), .A2(n15803), .ZN(n18919) );
  INV_X2 U14284 ( .A(n19091), .ZN(n19291) );
  NAND2_X1 U14285 ( .A1(n19291), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13476) );
  NAND2_X1 U14286 ( .A1(n12626), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11233) );
  INV_X1 U14287 ( .A(n11233), .ZN(n11216) );
  NAND2_X1 U14288 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15317) );
  NAND2_X1 U14289 ( .A1(n11211), .A2(n16385), .ZN(n15427) );
  AND2_X1 U14290 ( .A1(n9699), .A2(n11203), .ZN(n13444) );
  OAI22_X1 U14291 ( .A1(n11196), .A2(n19364), .B1(n16384), .B2(n10218), .ZN(
        n11197) );
  NOR2_X1 U14292 ( .A1(n13444), .A2(n11197), .ZN(n11208) );
  NAND2_X1 U14293 ( .A1(n11198), .A2(n19997), .ZN(n14168) );
  NAND2_X1 U14294 ( .A1(n14168), .A2(n11199), .ZN(n11201) );
  NAND2_X1 U14295 ( .A1(n11201), .A2(n11200), .ZN(n11207) );
  OAI21_X1 U14296 ( .B1(n11203), .B2(n11202), .A(n11196), .ZN(n11205) );
  NAND2_X1 U14297 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  OR2_X1 U14298 ( .A1(n14165), .A2(n11209), .ZN(n11210) );
  NAND2_X1 U14299 ( .A1(n11211), .A2(n11210), .ZN(n11219) );
  INV_X1 U14300 ( .A(n15427), .ZN(n11222) );
  NAND2_X1 U14301 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13683) );
  INV_X1 U14302 ( .A(n13683), .ZN(n13614) );
  NAND2_X1 U14303 ( .A1(n11221), .A2(n13683), .ZN(n11212) );
  OAI221_X1 U14304 ( .B1(n11222), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n11222), .C2(n13614), .A(n11212), .ZN(n13929) );
  NAND2_X1 U14305 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14144) );
  INV_X1 U14306 ( .A(n14144), .ZN(n11224) );
  NAND2_X1 U14307 ( .A1(n19336), .A2(n11224), .ZN(n14248) );
  NAND3_X1 U14308 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n16334), .ZN(n16287) );
  NAND2_X1 U14309 ( .A1(n11213), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11214) );
  NAND2_X1 U14310 ( .A1(n15442), .A2(n11226), .ZN(n15418) );
  NOR2_X1 U14311 ( .A1(n15400), .A2(n15207), .ZN(n15341) );
  INV_X1 U14312 ( .A(n15341), .ZN(n15373) );
  NOR3_X1 U14313 ( .A1(n21096), .A2(n15357), .A3(n15373), .ZN(n15343) );
  NAND2_X1 U14314 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15343), .ZN(
        n15316) );
  NAND2_X1 U14315 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15321), .ZN(
        n11215) );
  NOR2_X1 U14316 ( .A1(n15317), .A2(n11215), .ZN(n15289) );
  AND2_X1 U14317 ( .A1(n11216), .A2(n15289), .ZN(n15275) );
  NAND3_X1 U14318 ( .A1(n15275), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n9971), .ZN(n11217) );
  OAI211_X1 U14319 ( .C1(n16115), .C2(n19330), .A(n13476), .B(n11217), .ZN(
        n11218) );
  INV_X1 U14320 ( .A(n11218), .ZN(n11237) );
  INV_X1 U14321 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16337) );
  NOR2_X1 U14322 ( .A1(n16337), .A2(n16324), .ZN(n16326) );
  INV_X1 U14323 ( .A(n11219), .ZN(n15429) );
  AND2_X1 U14324 ( .A1(n11220), .A2(n19328), .ZN(n16348) );
  AOI21_X1 U14325 ( .B1(n15429), .B2(n13683), .A(n16348), .ZN(n13676) );
  NAND2_X1 U14326 ( .A1(n15429), .A2(n11221), .ZN(n13682) );
  NAND3_X1 U14327 ( .A1(n11222), .A2(n11221), .A3(n13683), .ZN(n13681) );
  AND2_X1 U14328 ( .A1(n13682), .A2(n13681), .ZN(n11223) );
  NAND2_X1 U14329 ( .A1(n11235), .A2(n20944), .ZN(n13928) );
  NAND2_X1 U14330 ( .A1(n14145), .A2(n11224), .ZN(n11225) );
  NAND2_X1 U14331 ( .A1(n15473), .A2(n11225), .ZN(n16321) );
  OAI221_X1 U14332 ( .B1(n16359), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        n16359), .C2(n16326), .A(n16321), .ZN(n15492) );
  NOR3_X1 U14333 ( .A1(n16251), .A2(n16286), .A3(n15492), .ZN(n15424) );
  NAND2_X1 U14334 ( .A1(n11226), .A2(n15424), .ZN(n15414) );
  NOR2_X1 U14335 ( .A1(n15417), .A2(n15414), .ZN(n15397) );
  NAND2_X1 U14336 ( .A1(n15397), .A2(n11227), .ZN(n11228) );
  NAND3_X1 U14337 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U14338 ( .A1(n11235), .A2(n11229), .ZN(n11230) );
  NAND2_X1 U14339 ( .A1(n11230), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U14340 ( .A1(n14311), .A2(n15473), .ZN(n15331) );
  OAI21_X1 U14341 ( .B1(n15322), .B2(n15323), .A(n15473), .ZN(n11232) );
  NAND2_X1 U14342 ( .A1(n11235), .A2(n11233), .ZN(n11234) );
  NAND2_X1 U14343 ( .A1(n15302), .A2(n11234), .ZN(n15282) );
  AOI21_X1 U14344 ( .B1(n15274), .B2(n11235), .A(n15282), .ZN(n11236) );
  NAND2_X4 U14345 ( .A1(n13957), .A2(n11248), .ZN(n12182) );
  AND2_X2 U14346 ( .A1(n13960), .A2(n14918), .ZN(n11466) );
  AOI22_X1 U14347 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14348 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11244) );
  INV_X4 U14349 ( .A(n9664), .ZN(n12227) );
  AND2_X2 U14350 ( .A1(n11249), .A2(n13707), .ZN(n11349) );
  AOI22_X1 U14351 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11242) );
  AND2_X2 U14352 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13954) );
  AND2_X2 U14353 ( .A1(n11246), .A2(n13954), .ZN(n12201) );
  NOR2_X2 U14354 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11247) );
  AND2_X4 U14355 ( .A1(n11247), .A2(n13954), .ZN(n11459) );
  AOI22_X1 U14356 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11253) );
  AND2_X4 U14357 ( .A1(n13707), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13952) );
  NAND2_X4 U14358 ( .A1(n13952), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12209) );
  INV_X1 U14359 ( .A(n12209), .ZN(n11350) );
  NAND2_X1 U14360 ( .A1(n11350), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11252) );
  AND2_X2 U14361 ( .A1(n11248), .A2(n11249), .ZN(n11488) );
  NAND2_X1 U14362 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11251) );
  NAND2_X1 U14363 ( .A1(n12240), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11250) );
  NAND4_X1 U14364 ( .A1(n11253), .A2(n11252), .A3(n11251), .A4(n11250), .ZN(
        n11259) );
  AND2_X4 U14365 ( .A1(n13952), .A2(n13956), .ZN(n11379) );
  INV_X1 U14366 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11257) );
  NAND2_X1 U14367 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11256) );
  NAND2_X1 U14368 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11255) );
  NOR2_X1 U14369 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  AND2_X2 U14370 ( .A1(n11261), .A2(n11260), .ZN(n11473) );
  AOI22_X1 U14371 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U14372 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11264) );
  NAND2_X1 U14373 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11263) );
  NAND2_X1 U14374 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11262) );
  NAND2_X1 U14375 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11269) );
  BUF_X4 U14376 ( .A(n11466), .Z(n12187) );
  NAND2_X1 U14377 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11268) );
  NAND2_X1 U14378 ( .A1(n11287), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11267) );
  NAND2_X1 U14379 ( .A1(n12227), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11266) );
  NAND2_X1 U14380 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11274) );
  NAND2_X1 U14381 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11273) );
  NAND2_X1 U14382 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11272) );
  NAND2_X1 U14383 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11271) );
  INV_X1 U14384 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U14385 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14386 ( .A1(n11349), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11275) );
  OAI211_X1 U14387 ( .C1(n12209), .C2(n12016), .A(n11276), .B(n11275), .ZN(
        n11277) );
  INV_X1 U14388 ( .A(n11277), .ZN(n11278) );
  NAND2_X1 U14389 ( .A1(n11474), .A2(n11541), .ZN(n11409) );
  NAND2_X1 U14390 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14391 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11284) );
  NAND2_X1 U14392 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11283) );
  BUF_X2 U14393 ( .A(n11340), .Z(n12065) );
  NAND2_X1 U14394 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11282) );
  AND4_X2 U14395 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n11303) );
  NAND2_X1 U14396 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11291) );
  NAND2_X1 U14397 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11290) );
  NAND2_X1 U14398 ( .A1(n11287), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11289) );
  NAND2_X1 U14399 ( .A1(n12227), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11288) );
  AND4_X2 U14400 ( .A1(n11291), .A2(n11290), .A3(n11289), .A4(n11288), .ZN(
        n11302) );
  AOI22_X1 U14401 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11295) );
  NAND2_X1 U14402 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11294) );
  NAND2_X1 U14403 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11293) );
  NAND2_X1 U14404 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11292) );
  INV_X1 U14405 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11298) );
  NAND2_X1 U14406 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11297) );
  NAND2_X1 U14407 ( .A1(n11349), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11296) );
  OAI211_X1 U14408 ( .C1(n12209), .C2(n11298), .A(n11297), .B(n11296), .ZN(
        n11299) );
  INV_X1 U14409 ( .A(n11299), .ZN(n11300) );
  NAND2_X1 U14410 ( .A1(n11422), .A2(n11541), .ZN(n12446) );
  NAND2_X1 U14411 ( .A1(n11409), .A2(n12446), .ZN(n11337) );
  AOI22_X1 U14412 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11307) );
  NAND2_X1 U14413 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11306) );
  NAND2_X1 U14414 ( .A1(n11287), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11305) );
  NAND2_X1 U14415 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14416 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14417 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U14418 ( .A1(n12227), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11308) );
  INV_X1 U14419 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11312) );
  NAND2_X1 U14420 ( .A1(n11340), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11315) );
  NAND2_X1 U14421 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11314) );
  NAND2_X1 U14422 ( .A1(n11349), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11313) );
  INV_X1 U14423 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12183) );
  NAND2_X1 U14424 ( .A1(n11466), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11318) );
  NAND2_X1 U14425 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11317) );
  OAI211_X1 U14426 ( .C1(n12209), .C2(n12183), .A(n11318), .B(n11317), .ZN(
        n11319) );
  INV_X1 U14427 ( .A(n11319), .ZN(n11320) );
  AOI22_X1 U14428 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12170), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14429 ( .A1(n11779), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12144), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14430 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14431 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14432 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11331) );
  NAND2_X1 U14433 ( .A1(n11350), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11330) );
  NAND2_X1 U14434 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14435 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11328) );
  AOI22_X1 U14436 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11334) );
  NAND2_X1 U14437 ( .A1(n9638), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14438 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11332) );
  AOI22_X1 U14439 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11344) );
  INV_X1 U14440 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12088) );
  INV_X1 U14441 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11338) );
  OAI22_X1 U14442 ( .A1(n12184), .A2(n12088), .B1(n12182), .B2(n11338), .ZN(
        n11339) );
  INV_X1 U14443 ( .A(n11339), .ZN(n11343) );
  AOI22_X1 U14444 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14445 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11341) );
  NAND4_X1 U14446 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .ZN(
        n11356) );
  NAND2_X1 U14447 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11348) );
  NAND2_X1 U14448 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11347) );
  NAND2_X1 U14449 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14450 ( .A1(n11459), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11345) );
  AND4_X1 U14451 ( .A1(n11348), .A2(n11347), .A3(n11346), .A4(n11345), .ZN(
        n11354) );
  AOI22_X1 U14452 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11353) );
  NAND2_X1 U14453 ( .A1(n11350), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14454 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11351) );
  NAND4_X1 U14455 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11355) );
  NAND2_X1 U14456 ( .A1(n13724), .A2(n12586), .ZN(n11359) );
  OAI22_X1 U14457 ( .A1(n12184), .A2(n11361), .B1(n12182), .B2(n11360), .ZN(
        n11362) );
  INV_X1 U14458 ( .A(n11362), .ZN(n11365) );
  NAND4_X1 U14459 ( .A1(n11366), .A2(n11365), .A3(n11364), .A4(n11363), .ZN(
        n11377) );
  AOI22_X1 U14460 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11375) );
  NAND2_X1 U14461 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11371) );
  NAND2_X1 U14462 ( .A1(n11367), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11370) );
  NAND2_X1 U14463 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11369) );
  NAND2_X1 U14464 ( .A1(n11459), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11368) );
  INV_X2 U14465 ( .A(n12209), .ZN(n11454) );
  NAND2_X1 U14466 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11373) );
  NAND2_X1 U14467 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11372) );
  NOR2_X1 U14468 ( .A1(n12586), .A2(n11412), .ZN(n11378) );
  AOI22_X1 U14469 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U14470 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11382) );
  NAND2_X1 U14471 ( .A1(n11488), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U14472 ( .A1(n12240), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11380) );
  INV_X1 U14473 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11384) );
  OAI22_X1 U14474 ( .A1(n12184), .A2(n11485), .B1(n12182), .B2(n11384), .ZN(
        n11388) );
  NAND2_X1 U14475 ( .A1(n12144), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11386) );
  NAND2_X1 U14476 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U14477 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  NOR2_X2 U14478 ( .A1(n11388), .A2(n11387), .ZN(n11398) );
  NAND2_X1 U14479 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11392) );
  NAND2_X1 U14480 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11391) );
  NAND2_X1 U14481 ( .A1(n11287), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11390) );
  NAND2_X1 U14482 ( .A1(n12227), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11389) );
  AND4_X2 U14483 ( .A1(n11392), .A2(n11391), .A3(n11390), .A4(n11389), .ZN(
        n11397) );
  NAND2_X1 U14484 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11394) );
  NAND2_X1 U14485 ( .A1(n11349), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11393) );
  OAI211_X1 U14486 ( .C1(n12209), .C2(n12063), .A(n11394), .B(n11393), .ZN(
        n11395) );
  INV_X1 U14487 ( .A(n11395), .ZN(n11396) );
  NAND4_X4 U14488 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n20275) );
  INV_X1 U14489 ( .A(n11402), .ZN(n11400) );
  AND2_X4 U14490 ( .A1(n11404), .A2(n20275), .ZN(n13573) );
  NAND2_X1 U14491 ( .A1(n12444), .A2(n13573), .ZN(n12320) );
  NAND2_X4 U14492 ( .A1(n13404), .A2(n11412), .ZN(n12566) );
  NAND2_X1 U14493 ( .A1(n12342), .A2(n20275), .ZN(n11426) );
  INV_X1 U14494 ( .A(n11405), .ZN(n11406) );
  NAND2_X1 U14495 ( .A1(n12523), .A2(n11406), .ZN(n12595) );
  NAND2_X1 U14496 ( .A1(n9631), .A2(n13870), .ZN(n11431) );
  AND2_X2 U14497 ( .A1(n20275), .A2(n20295), .ZN(n12403) );
  NAND2_X1 U14498 ( .A1(n11431), .A2(n11407), .ZN(n12452) );
  OR2_X2 U14499 ( .A1(n11408), .A2(n11404), .ZN(n11433) );
  AND3_X2 U14500 ( .A1(n12595), .A2(n12452), .A3(n11433), .ZN(n12590) );
  INV_X1 U14501 ( .A(n13870), .ZN(n11411) );
  INV_X1 U14502 ( .A(n11409), .ZN(n11410) );
  INV_X1 U14503 ( .A(n11413), .ZN(n13724) );
  NAND2_X1 U14504 ( .A1(n11412), .A2(n13724), .ZN(n12592) );
  OAI21_X1 U14505 ( .B1(n12586), .B2(n11426), .A(n12592), .ZN(n11424) );
  NAND3_X1 U14506 ( .A1(n20261), .A2(n20280), .A3(n13404), .ZN(n11439) );
  NAND2_X1 U14507 ( .A1(n11439), .A2(n14036), .ZN(n11414) );
  INV_X1 U14508 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20857) );
  NAND2_X1 U14509 ( .A1(n20008), .A2(n20857), .ZN(n20842) );
  NAND2_X1 U14510 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_1__SCAN_IN), 
        .ZN(n11416) );
  NAND2_X1 U14511 ( .A1(n20842), .A2(n11416), .ZN(n12442) );
  NAND2_X1 U14512 ( .A1(n16108), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15779) );
  INV_X1 U14513 ( .A(n15779), .ZN(n11419) );
  NAND2_X1 U14514 ( .A1(n16097), .A2(n9758), .ZN(n12641) );
  MUX2_X1 U14515 ( .A(n11419), .B(n12641), .S(n20701), .Z(n11420) );
  NAND2_X1 U14516 ( .A1(n11421), .A2(n11420), .ZN(n11496) );
  OR2_X1 U14517 ( .A1(n11439), .A2(n11422), .ZN(n12591) );
  NAND2_X1 U14518 ( .A1(n16097), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20013) );
  INV_X1 U14519 ( .A(n20013), .ZN(n11423) );
  AND3_X1 U14520 ( .A1(n12591), .A2(n11423), .A3(n14036), .ZN(n11430) );
  INV_X1 U14521 ( .A(n11424), .ZN(n13702) );
  NAND2_X1 U14522 ( .A1(n11425), .A2(n15770), .ZN(n11429) );
  AND2_X1 U14523 ( .A1(n14033), .A2(n12555), .ZN(n13568) );
  NAND2_X1 U14524 ( .A1(n13568), .A2(n11427), .ZN(n11428) );
  NAND3_X1 U14525 ( .A1(n11431), .A2(n20275), .A3(n14922), .ZN(n11432) );
  NAND3_X1 U14526 ( .A1(n11434), .A2(n11433), .A3(n11432), .ZN(n11497) );
  INV_X1 U14527 ( .A(n11500), .ZN(n11443) );
  NAND2_X1 U14528 ( .A1(n20779), .A2(n20701), .ZN(n20662) );
  NAND2_X1 U14529 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20633) );
  NAND2_X1 U14530 ( .A1(n20662), .A2(n20633), .ZN(n20591) );
  NAND2_X1 U14531 ( .A1(n15779), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11444) );
  OAI21_X1 U14532 ( .B1(n12641), .B2(n20591), .A(n11444), .ZN(n11436) );
  INV_X1 U14533 ( .A(n11436), .ZN(n11437) );
  INV_X1 U14534 ( .A(n11438), .ZN(n11442) );
  OR2_X1 U14535 ( .A1(n11439), .A2(n20275), .ZN(n12319) );
  NOR2_X1 U14536 ( .A1(n12319), .A2(n20295), .ZN(n13700) );
  INV_X1 U14537 ( .A(n12446), .ZN(n11540) );
  NAND2_X1 U14538 ( .A1(n13700), .A2(n11540), .ZN(n12582) );
  NAND2_X1 U14539 ( .A1(n11440), .A2(n12582), .ZN(n11441) );
  AND2_X1 U14540 ( .A1(n11444), .A2(n11435), .ZN(n11445) );
  NAND2_X1 U14541 ( .A1(n11478), .A2(n11447), .ZN(n11452) );
  INV_X1 U14542 ( .A(n12641), .ZN(n11576) );
  XNOR2_X1 U14543 ( .A(n20633), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20269) );
  NAND2_X1 U14544 ( .A1(n11576), .A2(n20269), .ZN(n11450) );
  NAND2_X1 U14545 ( .A1(n15779), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11449) );
  NAND2_X1 U14547 ( .A1(n11453), .A2(n13970), .ZN(n13697) );
  INV_X1 U14548 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U14549 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11456) );
  NAND2_X1 U14550 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11455) );
  OAI211_X1 U14551 ( .C1(n12232), .C2(n11457), .A(n11456), .B(n11455), .ZN(
        n11458) );
  INV_X1 U14552 ( .A(n11458), .ZN(n11463) );
  INV_X1 U14553 ( .A(n12201), .ZN(n12033) );
  INV_X2 U14554 ( .A(n12033), .ZN(n12228) );
  AOI22_X1 U14555 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11462) );
  INV_X1 U14556 ( .A(n11488), .ZN(n12035) );
  AOI22_X1 U14557 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11461) );
  NAND2_X1 U14558 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11460) );
  NAND4_X1 U14559 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11472) );
  AOI22_X1 U14560 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11470) );
  INV_X1 U14561 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11464) );
  OAI22_X1 U14562 ( .A1(n12184), .A2(n11464), .B1(n12182), .B2(n12088), .ZN(
        n11465) );
  INV_X1 U14563 ( .A(n11465), .ZN(n11469) );
  AOI22_X1 U14564 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14565 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11467) );
  NAND4_X1 U14566 ( .A1(n11470), .A2(n11469), .A3(n11468), .A4(n11467), .ZN(
        n11471) );
  INV_X1 U14567 ( .A(n11579), .ZN(n11476) );
  AOI22_X1 U14568 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11476), .B2(n11475), .ZN(n11477) );
  NAND2_X1 U14569 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11482) );
  AOI22_X1 U14570 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14571 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U14572 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11479) );
  NAND4_X1 U14573 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11487) );
  NAND2_X1 U14574 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11484) );
  NAND2_X1 U14575 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11483) );
  OAI211_X1 U14576 ( .C1(n11485), .C2(n12182), .A(n11484), .B(n11483), .ZN(
        n11486) );
  NOR2_X1 U14577 ( .A1(n11487), .A2(n11486), .ZN(n11494) );
  AOI22_X1 U14578 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11492) );
  INV_X2 U14579 ( .A(n12035), .ZN(n12149) );
  AOI22_X1 U14580 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14581 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14582 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11489) );
  AND4_X1 U14583 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(
        n11493) );
  NAND2_X1 U14584 ( .A1(n11494), .A2(n11493), .ZN(n12345) );
  NAND2_X1 U14585 ( .A1(n11531), .A2(n12345), .ZN(n11495) );
  INV_X1 U14586 ( .A(n11496), .ZN(n11499) );
  INV_X1 U14587 ( .A(n11497), .ZN(n11498) );
  NAND2_X1 U14588 ( .A1(n11499), .A2(n11498), .ZN(n11501) );
  AOI22_X1 U14589 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14590 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14591 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12240), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14592 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11502) );
  AND4_X1 U14593 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11515) );
  AOI22_X1 U14594 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11509) );
  NAND2_X1 U14595 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14596 ( .A1(n12119), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14597 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11506) );
  NAND4_X1 U14598 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11513) );
  INV_X1 U14599 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U14600 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11511) );
  INV_X1 U14601 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12031) );
  OR2_X1 U14602 ( .A1(n12184), .A2(n12031), .ZN(n11510) );
  OAI211_X1 U14603 ( .C1(n12232), .C2(n11549), .A(n11511), .B(n11510), .ZN(
        n11512) );
  NOR2_X1 U14604 ( .A1(n11513), .A2(n11512), .ZN(n11514) );
  INV_X1 U14605 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U14606 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U14607 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11516) );
  OAI211_X1 U14608 ( .C1(n12232), .C2(n11699), .A(n11517), .B(n11516), .ZN(
        n11518) );
  INV_X1 U14609 ( .A(n11518), .ZN(n11522) );
  AOI22_X1 U14610 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14611 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12240), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U14612 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11519) );
  NAND4_X1 U14613 ( .A1(n11522), .A2(n11521), .A3(n11520), .A4(n11519), .ZN(
        n11530) );
  AOI22_X1 U14614 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11528) );
  INV_X1 U14615 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11523) );
  INV_X1 U14616 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n21093) );
  OAI22_X1 U14617 ( .A1(n12184), .A2(n11523), .B1(n12182), .B2(n21093), .ZN(
        n11524) );
  INV_X1 U14618 ( .A(n11524), .ZN(n11527) );
  AOI22_X1 U14619 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14620 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11525) );
  NAND4_X1 U14621 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11529) );
  XNOR2_X1 U14622 ( .A(n12351), .B(n12407), .ZN(n11532) );
  NAND2_X1 U14623 ( .A1(n11532), .A2(n11531), .ZN(n11552) );
  INV_X1 U14624 ( .A(n12345), .ZN(n12341) );
  NAND2_X1 U14625 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11533) );
  INV_X1 U14626 ( .A(n11534), .ZN(n11535) );
  NAND2_X1 U14627 ( .A1(n11540), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11605) );
  XNOR2_X1 U14628 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20082) );
  INV_X2 U14629 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20780) );
  AOI21_X1 U14630 ( .B1(n12225), .B2(n20082), .A(n12258), .ZN(n11543) );
  NAND2_X1 U14631 ( .A1(n11602), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11542) );
  OAI211_X1 U14632 ( .C1(n11605), .C2(n9848), .A(n11543), .B(n11542), .ZN(
        n11544) );
  INV_X1 U14633 ( .A(n11544), .ZN(n11545) );
  NAND2_X1 U14634 ( .A1(n12258), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11571) );
  NAND2_X1 U14635 ( .A1(n11546), .A2(n11571), .ZN(n13790) );
  INV_X1 U14636 ( .A(n12302), .ZN(n11698) );
  AOI21_X1 U14637 ( .B1(n20290), .B2(n12407), .A(n9758), .ZN(n11548) );
  INV_X1 U14638 ( .A(n12351), .ZN(n12346) );
  NAND2_X1 U14639 ( .A1(n20261), .A2(n12346), .ZN(n11547) );
  OAI211_X1 U14640 ( .C1(n11698), .C2(n11549), .A(n11548), .B(n11547), .ZN(
        n11551) );
  NAND2_X1 U14641 ( .A1(n11550), .A2(n11551), .ZN(n11555) );
  INV_X1 U14642 ( .A(n11551), .ZN(n11553) );
  NAND2_X1 U14643 ( .A1(n11555), .A2(n11554), .ZN(n12353) );
  OR2_X1 U14644 ( .A1(n11556), .A2(n11771), .ZN(n11560) );
  AOI22_X1 U14645 ( .A1(n11602), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20780), .ZN(n11558) );
  INV_X1 U14646 ( .A(n11605), .ZN(n11631) );
  NAND2_X1 U14647 ( .A1(n11631), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11557) );
  AND2_X1 U14648 ( .A1(n11558), .A2(n11557), .ZN(n11559) );
  NAND2_X1 U14649 ( .A1(n11560), .A2(n11559), .ZN(n13658) );
  NAND2_X1 U14650 ( .A1(n13659), .A2(n13658), .ZN(n13657) );
  INV_X1 U14651 ( .A(n13658), .ZN(n11562) );
  INV_X1 U14652 ( .A(n12225), .ZN(n11561) );
  NAND2_X1 U14653 ( .A1(n11562), .A2(n12225), .ZN(n11563) );
  NAND2_X1 U14654 ( .A1(n13657), .A2(n11563), .ZN(n13867) );
  OR2_X1 U14655 ( .A1(n20338), .A2(n11771), .ZN(n11568) );
  AOI22_X1 U14656 ( .A1(n11602), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20780), .ZN(n11566) );
  NAND2_X1 U14657 ( .A1(n11631), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11565) );
  AND2_X1 U14658 ( .A1(n11566), .A2(n11565), .ZN(n11567) );
  NAND2_X1 U14659 ( .A1(n11568), .A2(n11567), .ZN(n13866) );
  NAND2_X1 U14660 ( .A1(n13867), .A2(n13866), .ZN(n13865) );
  INV_X1 U14661 ( .A(n13865), .ZN(n11569) );
  NAND2_X1 U14662 ( .A1(n11570), .A2(n11569), .ZN(n13788) );
  NAND2_X1 U14663 ( .A1(n11572), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11578) );
  INV_X1 U14664 ( .A(n20633), .ZN(n20375) );
  NAND2_X1 U14665 ( .A1(n20590), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20470) );
  INV_X1 U14666 ( .A(n20470), .ZN(n11573) );
  NAND2_X1 U14667 ( .A1(n20375), .A2(n11573), .ZN(n20507) );
  NAND2_X1 U14668 ( .A1(n20507), .A2(n20590), .ZN(n11575) );
  NAND2_X1 U14669 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20778) );
  INV_X1 U14670 ( .A(n20778), .ZN(n11574) );
  NAND2_X1 U14671 ( .A1(n20375), .A2(n11574), .ZN(n20775) );
  AND2_X1 U14672 ( .A1(n11575), .A2(n20775), .ZN(n20538) );
  AOI22_X1 U14673 ( .A1(n20538), .A2(n11576), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15779), .ZN(n11577) );
  INV_X1 U14674 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U14675 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11581) );
  NAND2_X1 U14676 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11580) );
  OAI211_X1 U14677 ( .C1(n12232), .C2(n11582), .A(n11581), .B(n11580), .ZN(
        n11583) );
  INV_X1 U14678 ( .A(n11583), .ZN(n11587) );
  AOI22_X1 U14679 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14680 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11585) );
  NAND2_X1 U14681 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11584) );
  NAND4_X1 U14682 ( .A1(n11587), .A2(n11586), .A3(n11585), .A4(n11584), .ZN(
        n11596) );
  AOI22_X1 U14683 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11594) );
  INV_X1 U14684 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11589) );
  INV_X1 U14685 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11588) );
  OAI22_X1 U14686 ( .A1(n12184), .A2(n11589), .B1(n12182), .B2(n11588), .ZN(
        n11590) );
  INV_X1 U14687 ( .A(n11590), .ZN(n11593) );
  AOI22_X1 U14688 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14689 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11591) );
  NAND4_X1 U14690 ( .A1(n11594), .A2(n11593), .A3(n11592), .A4(n11591), .ZN(
        n11595) );
  AOI22_X1 U14691 ( .A1(n12277), .A2(n12378), .B1(n12302), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14692 ( .A1(n20260), .A2(n11857), .ZN(n11608) );
  INV_X1 U14693 ( .A(n11561), .ZN(n12654) );
  INV_X1 U14694 ( .A(n11599), .ZN(n11601) );
  INV_X1 U14695 ( .A(n11633), .ZN(n11600) );
  OAI21_X1 U14696 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11601), .A(
        n11600), .ZN(n14046) );
  AOI22_X1 U14697 ( .A1(n12654), .A2(n14046), .B1(n12258), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U14698 ( .A1(n12259), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11603) );
  OAI211_X1 U14699 ( .C1(n11605), .C2(n13956), .A(n11604), .B(n11603), .ZN(
        n11606) );
  INV_X1 U14700 ( .A(n11606), .ZN(n11607) );
  NAND2_X1 U14701 ( .A1(n11608), .A2(n11607), .ZN(n13875) );
  NAND2_X1 U14702 ( .A1(n13876), .A2(n13875), .ZN(n13874) );
  INV_X1 U14703 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11613) );
  NAND2_X1 U14704 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11612) );
  NAND2_X1 U14705 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11611) );
  OAI211_X1 U14706 ( .C1(n12232), .C2(n11613), .A(n11612), .B(n11611), .ZN(
        n11614) );
  INV_X1 U14707 ( .A(n11614), .ZN(n11618) );
  AOI22_X1 U14708 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14709 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12149), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14710 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11615) );
  NAND4_X1 U14711 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11626) );
  AOI22_X1 U14712 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12239), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11624) );
  INV_X1 U14713 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11619) );
  INV_X1 U14714 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12142) );
  OAI22_X1 U14715 ( .A1(n12184), .A2(n11619), .B1(n12182), .B2(n12142), .ZN(
        n11620) );
  INV_X1 U14716 ( .A(n11620), .ZN(n11623) );
  AOI22_X1 U14717 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9627), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14718 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14719 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11625) );
  AOI22_X1 U14720 ( .A1(n12277), .A2(n12377), .B1(n12302), .B2(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14721 ( .A1(n11629), .A2(n11628), .ZN(n11630) );
  AND2_X1 U14722 ( .A1(n11662), .A2(n11630), .ZN(n12368) );
  NAND2_X1 U14723 ( .A1(n11631), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11636) );
  INV_X1 U14724 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20066) );
  AOI21_X1 U14725 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20066), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11632) );
  AOI21_X1 U14726 ( .B1(n12259), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11632), .ZN(
        n11635) );
  OAI21_X1 U14727 ( .B1(n11633), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11665), .ZN(n20192) );
  NOR2_X1 U14728 ( .A1(n20192), .A2(n11561), .ZN(n11634) );
  AOI21_X1 U14729 ( .B1(n11636), .B2(n11635), .A(n11634), .ZN(n11637) );
  NAND2_X1 U14730 ( .A1(n11639), .A2(n11638), .ZN(n13906) );
  INV_X1 U14731 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11642) );
  NAND2_X1 U14732 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11641) );
  NAND2_X1 U14733 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11640) );
  OAI211_X1 U14734 ( .C1(n12232), .C2(n11642), .A(n11641), .B(n11640), .ZN(
        n11643) );
  INV_X1 U14735 ( .A(n11643), .ZN(n11647) );
  AOI22_X1 U14736 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14737 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11645) );
  NAND2_X1 U14738 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11644) );
  NAND4_X1 U14739 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11656) );
  AOI22_X1 U14740 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11654) );
  INV_X1 U14741 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11649) );
  INV_X1 U14742 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11648) );
  OAI22_X1 U14743 ( .A1(n12184), .A2(n11649), .B1(n12182), .B2(n11648), .ZN(
        n11650) );
  INV_X1 U14744 ( .A(n11650), .ZN(n11653) );
  AOI22_X1 U14745 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14746 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14747 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11655) );
  NAND2_X1 U14748 ( .A1(n12277), .A2(n12388), .ZN(n11658) );
  NAND2_X1 U14749 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11657) );
  NAND2_X1 U14750 ( .A1(n11658), .A2(n11657), .ZN(n11660) );
  INV_X1 U14751 ( .A(n11660), .ZN(n11661) );
  NAND2_X1 U14752 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  NAND2_X1 U14753 ( .A1(n11694), .A2(n11663), .ZN(n12376) );
  INV_X1 U14754 ( .A(n12376), .ZN(n11664) );
  NAND2_X1 U14755 ( .A1(n11664), .A2(n11857), .ZN(n11671) );
  INV_X1 U14756 ( .A(n12258), .ZN(n11901) );
  NAND2_X1 U14757 ( .A1(n11665), .A2(n11668), .ZN(n11666) );
  INV_X1 U14758 ( .A(n11688), .ZN(n11689) );
  NAND2_X1 U14759 ( .A1(n11666), .A2(n11689), .ZN(n20063) );
  NAND2_X1 U14760 ( .A1(n20063), .A2(n12225), .ZN(n11667) );
  OAI21_X1 U14761 ( .B1(n11901), .B2(n11668), .A(n11667), .ZN(n11669) );
  AOI21_X1 U14762 ( .B1(n12259), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11669), .ZN(
        n11670) );
  INV_X1 U14763 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14069) );
  INV_X1 U14764 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14765 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11673) );
  NAND2_X1 U14766 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11672) );
  OAI211_X1 U14767 ( .C1(n12232), .C2(n11674), .A(n11673), .B(n11672), .ZN(
        n11675) );
  INV_X1 U14768 ( .A(n11675), .ZN(n11679) );
  AOI22_X1 U14769 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14770 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11677) );
  NAND2_X1 U14771 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11676) );
  NAND4_X1 U14772 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11687) );
  AOI22_X1 U14773 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11685) );
  INV_X1 U14774 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11680) );
  INV_X1 U14775 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12204) );
  OAI22_X1 U14776 ( .A1(n12184), .A2(n11680), .B1(n12182), .B2(n12204), .ZN(
        n11681) );
  INV_X1 U14777 ( .A(n11681), .ZN(n11684) );
  AOI22_X1 U14778 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14779 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11682) );
  NAND4_X1 U14780 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11686) );
  AOI22_X1 U14781 ( .A1(n12277), .A2(n12397), .B1(n12302), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11695) );
  NAND2_X1 U14782 ( .A1(n11694), .A2(n11695), .ZN(n12386) );
  NAND2_X1 U14783 ( .A1(n12386), .A2(n11857), .ZN(n11693) );
  INV_X1 U14784 ( .A(n11701), .ZN(n11703) );
  INV_X1 U14785 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11690) );
  NAND2_X1 U14786 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  NAND2_X1 U14787 ( .A1(n11703), .A2(n11691), .ZN(n20054) );
  AOI22_X1 U14788 ( .A1(n20054), .A2(n12225), .B1(n12258), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U14789 ( .A1(n13907), .A2(n14068), .ZN(n14003) );
  INV_X1 U14790 ( .A(n14003), .ZN(n11710) );
  NAND2_X1 U14791 ( .A1(n12277), .A2(n12407), .ZN(n11697) );
  OAI21_X1 U14792 ( .B1(n11699), .B2(n11698), .A(n11697), .ZN(n11700) );
  INV_X1 U14793 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11707) );
  INV_X1 U14794 ( .A(n11730), .ZN(n11705) );
  INV_X1 U14795 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11702) );
  NAND2_X1 U14796 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  NAND2_X1 U14797 ( .A1(n11705), .A2(n11704), .ZN(n20044) );
  AOI22_X1 U14798 ( .A1(n20044), .A2(n12225), .B1(n12258), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11706) );
  OAI21_X1 U14799 ( .B1(n12220), .B2(n11707), .A(n11706), .ZN(n11708) );
  NAND2_X1 U14800 ( .A1(n11710), .A2(n11709), .ZN(n14001) );
  INV_X1 U14801 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11711) );
  OAI22_X1 U14802 ( .A1(n12184), .A2(n11711), .B1(n12182), .B2(n12031), .ZN(
        n11712) );
  INV_X1 U14803 ( .A(n11712), .ZN(n11716) );
  AOI22_X1 U14804 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14805 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14806 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U14807 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n11726) );
  INV_X1 U14808 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14809 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11718) );
  NAND2_X1 U14810 ( .A1(n12234), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11717) );
  OAI211_X1 U14811 ( .C1(n12232), .C2(n11719), .A(n11718), .B(n11717), .ZN(
        n11720) );
  INV_X1 U14812 ( .A(n11720), .ZN(n11724) );
  AOI22_X1 U14813 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11723) );
  INV_X1 U14814 ( .A(n12018), .ZN(n12241) );
  AOI22_X1 U14815 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U14816 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11721) );
  NAND4_X1 U14817 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n11725) );
  OAI21_X1 U14818 ( .B1(n11726), .B2(n11725), .A(n11857), .ZN(n11729) );
  NAND2_X1 U14819 ( .A1(n12259), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11728) );
  XNOR2_X1 U14820 ( .A(n11730), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14239) );
  AOI22_X1 U14821 ( .A1(n14239), .A2(n12225), .B1(n12258), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11727) );
  XNOR2_X1 U14822 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11768), .ZN(
        n14774) );
  INV_X1 U14823 ( .A(n14774), .ZN(n11752) );
  AOI22_X1 U14824 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11737) );
  INV_X1 U14825 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11732) );
  INV_X1 U14826 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11731) );
  OAI22_X1 U14827 ( .A1(n12184), .A2(n11732), .B1(n12182), .B2(n11731), .ZN(
        n11733) );
  INV_X1 U14828 ( .A(n11733), .ZN(n11736) );
  AOI22_X1 U14829 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14830 ( .A1(n12119), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14831 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11747) );
  INV_X1 U14832 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11740) );
  NAND2_X1 U14833 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14834 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11738) );
  OAI211_X1 U14835 ( .C1(n12232), .C2(n11740), .A(n11739), .B(n11738), .ZN(
        n11741) );
  INV_X1 U14836 ( .A(n11741), .ZN(n11745) );
  AOI22_X1 U14837 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14838 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11743) );
  NAND2_X1 U14839 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11742) );
  NAND4_X1 U14840 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11746) );
  OAI21_X1 U14841 ( .B1(n11747), .B2(n11746), .A(n11857), .ZN(n11750) );
  NAND2_X1 U14842 ( .A1(n12259), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11749) );
  NAND2_X1 U14843 ( .A1(n12258), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11748) );
  NAND3_X1 U14844 ( .A1(n11750), .A2(n11749), .A3(n11748), .ZN(n11751) );
  AOI21_X1 U14845 ( .B1(n11752), .B2(n12654), .A(n11751), .ZN(n14158) );
  AND2_X2 U14846 ( .A1(n14075), .A2(n14160), .ZN(n14159) );
  INV_X1 U14847 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U14848 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11755) );
  INV_X1 U14849 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11753) );
  OR2_X1 U14850 ( .A1(n12184), .A2(n11753), .ZN(n11754) );
  OAI211_X1 U14851 ( .C1(n12232), .C2(n11756), .A(n11755), .B(n11754), .ZN(
        n11757) );
  INV_X1 U14852 ( .A(n11757), .ZN(n11761) );
  AOI22_X1 U14853 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14854 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11759) );
  NAND2_X1 U14855 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11758) );
  NAND4_X1 U14856 ( .A1(n11761), .A2(n11760), .A3(n11759), .A4(n11758), .ZN(
        n11767) );
  AOI22_X1 U14857 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U14858 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14859 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14860 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11762) );
  NAND4_X1 U14861 ( .A1(n11765), .A2(n11764), .A3(n11763), .A4(n11762), .ZN(
        n11766) );
  NOR2_X1 U14862 ( .A1(n11767), .A2(n11766), .ZN(n11772) );
  XNOR2_X1 U14863 ( .A(n11773), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14767) );
  NAND2_X1 U14864 ( .A1(n14767), .A2(n12225), .ZN(n11770) );
  AOI22_X1 U14865 ( .A1(n12259), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12258), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11769) );
  OAI211_X1 U14866 ( .C1(n11772), .C2(n11771), .A(n11770), .B(n11769), .ZN(
        n14212) );
  INV_X1 U14867 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11776) );
  OAI21_X1 U14868 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11774), .A(
        n11813), .ZN(n15950) );
  NAND2_X1 U14869 ( .A1(n15950), .A2(n12654), .ZN(n11775) );
  OAI21_X1 U14870 ( .B1(n11776), .B2(n11901), .A(n11775), .ZN(n11777) );
  AOI21_X1 U14871 ( .B1(n12259), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11777), .ZN(
        n14471) );
  AOI22_X1 U14872 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14873 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14874 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14875 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11780) );
  AND4_X1 U14876 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11790) );
  AOI22_X1 U14877 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11980), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14878 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14879 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11785) );
  NAND2_X1 U14880 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11784) );
  AND3_X1 U14881 ( .A1(n11786), .A2(n11785), .A3(n11784), .ZN(n11788) );
  NAND2_X1 U14882 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11787) );
  NAND4_X1 U14883 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11791) );
  NAND2_X1 U14884 ( .A1(n11857), .A2(n11791), .ZN(n14644) );
  INV_X1 U14885 ( .A(n14644), .ZN(n11792) );
  XNOR2_X1 U14886 ( .A(n11829), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14756) );
  NAND2_X1 U14887 ( .A1(n14756), .A2(n12225), .ZN(n11812) );
  INV_X1 U14888 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U14889 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14890 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14891 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14892 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11795) );
  AND4_X1 U14893 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11806) );
  AOI22_X1 U14894 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U14895 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11802) );
  AOI22_X1 U14896 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U14897 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11800) );
  NAND2_X1 U14898 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11799) );
  AND4_X1 U14899 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11804) );
  NAND2_X1 U14900 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11803) );
  NAND4_X1 U14901 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n11807) );
  NAND2_X1 U14902 ( .A1(n11857), .A2(n11807), .ZN(n11809) );
  NAND2_X1 U14903 ( .A1(n12258), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11808) );
  OAI211_X1 U14904 ( .C1(n12220), .C2(n14640), .A(n11809), .B(n11808), .ZN(
        n11810) );
  INV_X1 U14905 ( .A(n11810), .ZN(n11811) );
  NAND2_X1 U14906 ( .A1(n11812), .A2(n11811), .ZN(n14473) );
  INV_X1 U14907 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14642) );
  XNOR2_X1 U14908 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11813), .ZN(
        n15939) );
  OAI22_X1 U14909 ( .A1(n15939), .A2(n11561), .B1(n11901), .B2(n11793), .ZN(
        n11814) );
  INV_X1 U14910 ( .A(n11814), .ZN(n11828) );
  AOI22_X1 U14911 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U14912 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12239), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U14913 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14914 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12242), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11815) );
  AND4_X1 U14915 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11825) );
  AOI22_X1 U14916 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14917 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12149), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14918 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U14919 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11819) );
  AND3_X1 U14920 ( .A1(n11821), .A2(n11820), .A3(n11819), .ZN(n11823) );
  NAND2_X1 U14921 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11822) );
  NAND4_X1 U14922 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11826) );
  NAND2_X1 U14923 ( .A1(n11857), .A2(n11826), .ZN(n11827) );
  OAI211_X1 U14924 ( .C1(n12220), .C2(n14642), .A(n11828), .B(n11827), .ZN(
        n14563) );
  INV_X1 U14925 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14639) );
  AOI21_X1 U14926 ( .B1(n21078), .B2(n11830), .A(n11883), .ZN(n15933) );
  OR2_X1 U14927 ( .A1(n15933), .A2(n11561), .ZN(n11844) );
  AOI22_X1 U14928 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14929 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14930 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14931 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11831) );
  AND4_X1 U14932 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11841) );
  AOI22_X1 U14933 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14934 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14935 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11836) );
  NAND2_X1 U14936 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11835) );
  AND3_X1 U14937 ( .A1(n11837), .A2(n11836), .A3(n11835), .ZN(n11839) );
  NAND2_X1 U14938 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11838) );
  NAND4_X1 U14939 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n11842) );
  AOI22_X1 U14940 ( .A1(n11857), .A2(n11842), .B1(n12258), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11843) );
  OAI211_X1 U14941 ( .C1(n12220), .C2(n14639), .A(n11844), .B(n11843), .ZN(
        n14554) );
  NAND2_X1 U14942 ( .A1(n14474), .A2(n14554), .ZN(n14455) );
  INV_X1 U14943 ( .A(n14455), .ZN(n11865) );
  XNOR2_X1 U14944 ( .A(n11883), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14744) );
  AOI22_X1 U14945 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14946 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14947 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14948 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U14949 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11859) );
  INV_X1 U14950 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11851) );
  NAND2_X1 U14951 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11850) );
  NAND2_X1 U14952 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11849) );
  OAI211_X1 U14953 ( .C1(n12232), .C2(n11851), .A(n11850), .B(n11849), .ZN(
        n11852) );
  INV_X1 U14954 ( .A(n11852), .ZN(n11856) );
  AOI22_X1 U14955 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14956 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11854) );
  NAND2_X1 U14957 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11853) );
  NAND4_X1 U14958 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11858) );
  OAI21_X1 U14959 ( .B1(n11859), .B2(n11858), .A(n11857), .ZN(n11862) );
  NAND2_X1 U14960 ( .A1(n12259), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U14961 ( .A1(n12258), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11860) );
  NAND3_X1 U14962 ( .A1(n11862), .A2(n11861), .A3(n11860), .ZN(n11863) );
  AOI21_X1 U14963 ( .B1(n14744), .B2(n12654), .A(n11863), .ZN(n14459) );
  INV_X1 U14964 ( .A(n14459), .ZN(n11864) );
  NAND2_X1 U14965 ( .A1(n11865), .A2(n11864), .ZN(n14457) );
  INV_X1 U14966 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12032) );
  NAND2_X1 U14967 ( .A1(n11287), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U14968 ( .A1(n12119), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11866) );
  OAI211_X1 U14969 ( .C1(n12232), .C2(n12032), .A(n11867), .B(n11866), .ZN(
        n11868) );
  INV_X1 U14970 ( .A(n11868), .ZN(n11872) );
  AOI22_X1 U14971 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14972 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11980), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U14973 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11869) );
  NAND4_X1 U14974 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11878) );
  AOI22_X1 U14975 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14976 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14977 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14978 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11873) );
  NAND4_X1 U14979 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11877) );
  NOR2_X1 U14980 ( .A1(n11878), .A2(n11877), .ZN(n11882) );
  INV_X1 U14981 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20418) );
  OAI21_X1 U14982 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20418), .A(
        n20780), .ZN(n11879) );
  INV_X1 U14983 ( .A(n11879), .ZN(n11880) );
  AOI21_X1 U14984 ( .B1(n12259), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11880), .ZN(
        n11881) );
  OAI21_X1 U14985 ( .B1(n12255), .B2(n11882), .A(n11881), .ZN(n11886) );
  OAI21_X1 U14986 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11884), .A(
        n11923), .ZN(n15928) );
  OR2_X1 U14987 ( .A1(n11561), .A2(n15928), .ZN(n11885) );
  NAND2_X1 U14988 ( .A1(n11886), .A2(n11885), .ZN(n14547) );
  INV_X1 U14989 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11889) );
  NAND2_X1 U14990 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U14991 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11887) );
  OAI211_X1 U14992 ( .C1(n12209), .C2(n11889), .A(n11888), .B(n11887), .ZN(
        n11890) );
  INV_X1 U14993 ( .A(n11890), .ZN(n11894) );
  AOI22_X1 U14994 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14995 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11892) );
  NAND2_X1 U14996 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11891) );
  NAND4_X1 U14997 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11900) );
  AOI22_X1 U14998 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U14999 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15000 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U15001 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11895) );
  NAND4_X1 U15002 ( .A1(n11898), .A2(n11897), .A3(n11896), .A4(n11895), .ZN(
        n11899) );
  NOR2_X1 U15003 ( .A1(n11900), .A2(n11899), .ZN(n11904) );
  XNOR2_X1 U15004 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11923), .ZN(
        n14735) );
  INV_X1 U15005 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14731) );
  OAI22_X1 U15006 ( .A1(n11561), .A2(n14735), .B1(n11901), .B2(n14731), .ZN(
        n11902) );
  AOI21_X1 U15007 ( .B1(n12259), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11902), .ZN(
        n11903) );
  OAI21_X1 U15008 ( .B1(n12255), .B2(n11904), .A(n11903), .ZN(n14446) );
  AND2_X2 U15009 ( .A1(n14444), .A2(n14446), .ZN(n14445) );
  INV_X1 U15010 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U15011 ( .A1(n12234), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11906) );
  NAND2_X1 U15012 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11905) );
  OAI211_X1 U15013 ( .C1(n12232), .C2(n11907), .A(n11906), .B(n11905), .ZN(
        n11908) );
  INV_X1 U15014 ( .A(n11908), .ZN(n11912) );
  AOI22_X1 U15015 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15016 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11910) );
  NAND2_X1 U15017 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11909) );
  NAND4_X1 U15018 ( .A1(n11912), .A2(n11911), .A3(n11910), .A4(n11909), .ZN(
        n11918) );
  AOI22_X1 U15019 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U15020 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15021 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15022 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U15023 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11917) );
  NOR2_X1 U15024 ( .A1(n11918), .A2(n11917), .ZN(n11922) );
  NAND2_X1 U15025 ( .A1(n20780), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11919) );
  NAND2_X1 U15026 ( .A1(n11561), .A2(n11919), .ZN(n11920) );
  AOI21_X1 U15027 ( .B1(n12259), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11920), .ZN(
        n11921) );
  OAI21_X1 U15028 ( .B1(n12255), .B2(n11922), .A(n11921), .ZN(n11926) );
  OAI21_X1 U15029 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11924), .A(
        n11966), .ZN(n15921) );
  OR2_X1 U15030 ( .A1(n11561), .A2(n15921), .ZN(n11925) );
  INV_X1 U15031 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11927) );
  OR2_X1 U15032 ( .A1(n11928), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U15033 ( .A1(n11929), .A2(n12012), .ZN(n15907) );
  INV_X1 U15034 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11932) );
  NAND2_X1 U15035 ( .A1(n12119), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U15036 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11930) );
  OAI211_X1 U15037 ( .C1(n12232), .C2(n11932), .A(n11931), .B(n11930), .ZN(
        n11933) );
  INV_X1 U15038 ( .A(n11933), .ZN(n11937) );
  AOI22_X1 U15039 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U15040 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12239), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U15041 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11934) );
  NAND4_X1 U15042 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n11943) );
  AOI22_X1 U15043 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11980), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15044 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15045 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12241), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15046 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12242), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11938) );
  NAND4_X1 U15047 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11942) );
  NOR2_X1 U15048 ( .A1(n11943), .A2(n11942), .ZN(n11946) );
  OAI21_X1 U15049 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20418), .A(
        n20780), .ZN(n11945) );
  NAND2_X1 U15050 ( .A1(n12259), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n11944) );
  OAI211_X1 U15051 ( .C1(n12255), .C2(n11946), .A(n11945), .B(n11944), .ZN(
        n11947) );
  OAI21_X1 U15052 ( .B1(n15907), .B2(n11561), .A(n11947), .ZN(n14525) );
  INV_X1 U15053 ( .A(n14525), .ZN(n11970) );
  AOI22_X1 U15054 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U15055 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15056 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15057 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11948) );
  NAND4_X1 U15058 ( .A1(n11951), .A2(n11950), .A3(n11949), .A4(n11948), .ZN(
        n11961) );
  AOI22_X1 U15059 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U15060 ( .A1(n11287), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11955) );
  NAND2_X1 U15061 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11954) );
  NAND2_X1 U15062 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11953) );
  NAND2_X1 U15063 ( .A1(n11459), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11952) );
  AND4_X1 U15064 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11958) );
  NAND2_X1 U15065 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11957) );
  NAND2_X1 U15066 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11956) );
  NAND4_X1 U15067 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  NOR2_X1 U15068 ( .A1(n11961), .A2(n11960), .ZN(n11965) );
  NAND2_X1 U15069 ( .A1(n20780), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11962) );
  NAND2_X1 U15070 ( .A1(n11561), .A2(n11962), .ZN(n11963) );
  AOI21_X1 U15071 ( .B1(n12259), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11963), .ZN(
        n11964) );
  OAI21_X1 U15072 ( .B1(n12255), .B2(n11965), .A(n11964), .ZN(n11968) );
  XNOR2_X1 U15073 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n11966), .ZN(
        n14719) );
  NAND2_X1 U15074 ( .A1(n12654), .A2(n14719), .ZN(n11967) );
  NAND2_X1 U15075 ( .A1(n11968), .A2(n11967), .ZN(n14526) );
  INV_X1 U15076 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11974) );
  NAND2_X1 U15077 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11973) );
  NAND2_X1 U15078 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11972) );
  OAI211_X1 U15079 ( .C1(n12209), .C2(n11974), .A(n11973), .B(n11972), .ZN(
        n11975) );
  INV_X1 U15080 ( .A(n11975), .ZN(n11979) );
  AOI22_X1 U15081 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15082 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11977) );
  NAND2_X1 U15083 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11976) );
  NAND4_X1 U15084 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11986) );
  AOI22_X1 U15085 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15086 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11980), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15087 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15088 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11981) );
  NAND4_X1 U15089 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11985) );
  NOR2_X1 U15090 ( .A1(n11986), .A2(n11985), .ZN(n11990) );
  NAND2_X1 U15091 ( .A1(n20780), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11987) );
  NAND2_X1 U15092 ( .A1(n11561), .A2(n11987), .ZN(n11988) );
  AOI21_X1 U15093 ( .B1(n12259), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11988), .ZN(
        n11989) );
  OAI21_X1 U15094 ( .B1(n12255), .B2(n11990), .A(n11989), .ZN(n11992) );
  XNOR2_X1 U15095 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12012), .ZN(
        n15902) );
  NAND2_X1 U15096 ( .A1(n12654), .A2(n15902), .ZN(n11991) );
  AOI22_X1 U15097 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12239), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15098 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15099 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15100 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11993) );
  NAND4_X1 U15101 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n12006) );
  AOI22_X1 U15102 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12004) );
  NAND2_X1 U15103 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12000) );
  NAND2_X1 U15104 ( .A1(n12240), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11999) );
  NAND2_X1 U15105 ( .A1(n9638), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11998) );
  NAND2_X1 U15106 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11997) );
  AND4_X1 U15107 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12003) );
  NAND2_X1 U15108 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12002) );
  NAND2_X1 U15109 ( .A1(n11454), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12001) );
  NAND4_X1 U15110 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12005) );
  NOR2_X1 U15111 ( .A1(n12006), .A2(n12005), .ZN(n12010) );
  OAI21_X1 U15112 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20418), .A(
        n20780), .ZN(n12007) );
  INV_X1 U15113 ( .A(n12007), .ZN(n12008) );
  AOI21_X1 U15114 ( .B1(n12259), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12008), .ZN(
        n12009) );
  OAI21_X1 U15115 ( .B1(n12255), .B2(n12010), .A(n12009), .ZN(n12015) );
  INV_X1 U15116 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12011) );
  OAI21_X1 U15117 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12013), .A(
        n12076), .ZN(n15901) );
  OR2_X1 U15118 ( .A1(n11561), .A2(n15901), .ZN(n12014) );
  INV_X1 U15119 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12017) );
  OAI22_X1 U15120 ( .A1(n12018), .A2(n12017), .B1(n9664), .B2(n12016), .ZN(
        n12019) );
  AOI21_X1 U15121 ( .B1(n11454), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12019), .ZN(n12023) );
  AOI22_X1 U15122 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12228), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15123 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12021) );
  NAND2_X1 U15124 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12020) );
  NAND4_X1 U15125 ( .A1(n12023), .A2(n12022), .A3(n12021), .A4(n12020), .ZN(
        n12029) );
  AOI22_X1 U15126 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12210), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15127 ( .A1(n11980), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15128 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15129 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12024) );
  NAND4_X1 U15130 ( .A1(n12027), .A2(n12026), .A3(n12025), .A4(n12024), .ZN(
        n12028) );
  NOR2_X1 U15131 ( .A1(n12029), .A2(n12028), .ZN(n12052) );
  INV_X1 U15132 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12040) );
  INV_X1 U15133 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12030) );
  OAI22_X1 U15134 ( .A1(n9628), .A2(n12031), .B1(n12184), .B2(n12030), .ZN(
        n12037) );
  INV_X1 U15135 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12034) );
  OAI22_X1 U15136 ( .A1(n12035), .A2(n12034), .B1(n12033), .B2(n12032), .ZN(
        n12036) );
  AOI211_X1 U15137 ( .C1(n12175), .C2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n12037), .B(n12036), .ZN(n12039) );
  AOI22_X1 U15138 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12038) );
  OAI211_X1 U15139 ( .C1(n12209), .C2(n12040), .A(n12039), .B(n12038), .ZN(
        n12046) );
  AOI22_X1 U15140 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12239), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15141 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15142 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15143 ( .A1(n12148), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12041) );
  NAND4_X1 U15144 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12045) );
  NOR2_X1 U15145 ( .A1(n12046), .A2(n12045), .ZN(n12053) );
  XOR2_X1 U15146 ( .A(n12052), .B(n12053), .Z(n12047) );
  INV_X1 U15147 ( .A(n12255), .ZN(n12222) );
  NAND2_X1 U15148 ( .A1(n12047), .A2(n12222), .ZN(n12051) );
  INV_X1 U15149 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15829) );
  OAI21_X1 U15150 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15829), .A(n11561), 
        .ZN(n12048) );
  AOI21_X1 U15151 ( .B1(n12259), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12048), .ZN(
        n12050) );
  XNOR2_X1 U15152 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12076), .ZN(
        n15822) );
  AOI21_X1 U15153 ( .B1(n12051), .B2(n12050), .A(n12049), .ZN(n14504) );
  NOR2_X1 U15154 ( .A1(n12053), .A2(n12052), .ZN(n12085) );
  INV_X1 U15155 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U15156 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12055) );
  NAND2_X1 U15157 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12054) );
  OAI211_X1 U15158 ( .C1(n12232), .C2(n12056), .A(n12055), .B(n12054), .ZN(
        n12057) );
  INV_X1 U15159 ( .A(n12057), .ZN(n12061) );
  AOI22_X1 U15160 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15161 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12148), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12059) );
  NAND2_X1 U15162 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12058) );
  NAND4_X1 U15163 ( .A1(n12061), .A2(n12060), .A3(n12059), .A4(n12058), .ZN(
        n12071) );
  AOI22_X1 U15164 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12241), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12069) );
  INV_X1 U15165 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12062) );
  OAI22_X1 U15166 ( .A1(n12184), .A2(n12063), .B1(n12182), .B2(n12062), .ZN(
        n12064) );
  INV_X1 U15167 ( .A(n12064), .ZN(n12068) );
  AOI22_X1 U15168 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12067) );
  INV_X1 U15169 ( .A(n9664), .ZN(n12119) );
  AOI22_X1 U15170 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U15171 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12070) );
  OR2_X1 U15172 ( .A1(n12071), .A2(n12070), .ZN(n12084) );
  INV_X1 U15173 ( .A(n12084), .ZN(n12072) );
  XNOR2_X1 U15174 ( .A(n12085), .B(n12072), .ZN(n12075) );
  INV_X1 U15175 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U15176 ( .A1(n20780), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12073) );
  OAI211_X1 U15177 ( .C1(n12220), .C2(n14595), .A(n11561), .B(n12073), .ZN(
        n12074) );
  AOI21_X1 U15178 ( .B1(n12075), .B2(n12222), .A(n12074), .ZN(n12083) );
  INV_X1 U15179 ( .A(n12078), .ZN(n12080) );
  INV_X1 U15180 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12079) );
  NAND2_X1 U15181 ( .A1(n12080), .A2(n12079), .ZN(n12081) );
  NAND2_X1 U15182 ( .A1(n12130), .A2(n12081), .ZN(n15821) );
  NOR2_X1 U15183 ( .A1(n15821), .A2(n11561), .ZN(n12082) );
  NAND2_X1 U15184 ( .A1(n12085), .A2(n12084), .ZN(n12106) );
  INV_X1 U15185 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15186 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15187 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12086) );
  OAI211_X1 U15188 ( .C1(n12238), .C2(n12088), .A(n12087), .B(n12086), .ZN(
        n12089) );
  INV_X1 U15189 ( .A(n12089), .ZN(n12091) );
  AOI22_X1 U15190 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12090) );
  OAI211_X1 U15191 ( .C1(n12209), .C2(n12092), .A(n12091), .B(n12090), .ZN(
        n12098) );
  AOI22_X1 U15192 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15193 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15194 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12240), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15195 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12093) );
  NAND4_X1 U15196 ( .A1(n12096), .A2(n12095), .A3(n12094), .A4(n12093), .ZN(
        n12097) );
  NOR2_X1 U15197 ( .A1(n12098), .A2(n12097), .ZN(n12107) );
  XOR2_X1 U15198 ( .A(n12106), .B(n12107), .Z(n12099) );
  NAND2_X1 U15199 ( .A1(n12099), .A2(n12222), .ZN(n12102) );
  INV_X1 U15200 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14696) );
  AOI21_X1 U15201 ( .B1(n14696), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12100) );
  AOI21_X1 U15202 ( .B1(n12259), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12100), .ZN(
        n12101) );
  NAND2_X1 U15203 ( .A1(n12102), .A2(n12101), .ZN(n12104) );
  XNOR2_X1 U15204 ( .A(n12130), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14694) );
  NAND2_X1 U15205 ( .A1(n14694), .A2(n12225), .ZN(n12103) );
  NAND2_X1 U15206 ( .A1(n12104), .A2(n12103), .ZN(n14408) );
  NOR2_X1 U15207 ( .A1(n12107), .A2(n12106), .ZN(n12139) );
  INV_X1 U15208 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12110) );
  NAND2_X1 U15209 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12109) );
  NAND2_X1 U15210 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12108) );
  OAI211_X1 U15211 ( .C1(n12232), .C2(n12110), .A(n12109), .B(n12108), .ZN(
        n12111) );
  INV_X1 U15212 ( .A(n12111), .ZN(n12115) );
  AOI22_X1 U15213 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15214 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12240), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12113) );
  NAND2_X1 U15215 ( .A1(n11379), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12112) );
  NAND4_X1 U15216 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12125) );
  AOI22_X1 U15217 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12123) );
  INV_X1 U15218 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12117) );
  INV_X1 U15219 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12116) );
  OAI22_X1 U15220 ( .A1(n12117), .A2(n12182), .B1(n12184), .B2(n12116), .ZN(
        n12118) );
  INV_X1 U15221 ( .A(n12118), .ZN(n12122) );
  AOI22_X1 U15222 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15223 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12119), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15224 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12124) );
  OR2_X1 U15225 ( .A1(n12125), .A2(n12124), .ZN(n12138) );
  INV_X1 U15226 ( .A(n12138), .ZN(n12126) );
  XNOR2_X1 U15227 ( .A(n12139), .B(n12126), .ZN(n12127) );
  NAND2_X1 U15228 ( .A1(n12127), .A2(n12222), .ZN(n12137) );
  NAND2_X1 U15229 ( .A1(n20780), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12128) );
  NAND2_X1 U15230 ( .A1(n11561), .A2(n12128), .ZN(n12129) );
  AOI21_X1 U15231 ( .B1(n12259), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12129), .ZN(
        n12136) );
  INV_X1 U15232 ( .A(n12131), .ZN(n12133) );
  INV_X1 U15233 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U15234 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  NAND2_X1 U15235 ( .A1(n12162), .A2(n12134), .ZN(n14681) );
  NOR2_X1 U15236 ( .A1(n14681), .A2(n11561), .ZN(n12135) );
  AOI21_X1 U15237 ( .B1(n12137), .B2(n12136), .A(n12135), .ZN(n14393) );
  NAND2_X1 U15238 ( .A1(n12139), .A2(n12138), .ZN(n12168) );
  INV_X1 U15239 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15240 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15241 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12228), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12140) );
  OAI211_X1 U15242 ( .C1(n12238), .C2(n12142), .A(n12141), .B(n12140), .ZN(
        n12143) );
  INV_X1 U15243 ( .A(n12143), .ZN(n12146) );
  AOI22_X1 U15244 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9627), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12145) );
  OAI211_X1 U15245 ( .C1(n12147), .C2(n12232), .A(n12146), .B(n12145), .ZN(
        n12155) );
  AOI22_X1 U15246 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12239), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15247 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12148), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15248 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12242), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15249 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15250 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12154) );
  NOR2_X1 U15251 ( .A1(n12155), .A2(n12154), .ZN(n12169) );
  XOR2_X1 U15252 ( .A(n12168), .B(n12169), .Z(n12156) );
  NAND2_X1 U15253 ( .A1(n12156), .A2(n12222), .ZN(n12161) );
  NAND2_X1 U15254 ( .A1(n20780), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12157) );
  NAND2_X1 U15255 ( .A1(n11561), .A2(n12157), .ZN(n12158) );
  AOI21_X1 U15256 ( .B1(n12259), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12158), .ZN(
        n12160) );
  XNOR2_X1 U15257 ( .A(n12162), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14678) );
  AOI21_X1 U15258 ( .B1(n12161), .B2(n12160), .A(n12159), .ZN(n14379) );
  INV_X1 U15259 ( .A(n12162), .ZN(n12163) );
  INV_X1 U15260 ( .A(n12164), .ZN(n12166) );
  INV_X1 U15261 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12165) );
  NAND2_X1 U15262 ( .A1(n12166), .A2(n12165), .ZN(n12167) );
  NAND2_X1 U15263 ( .A1(n12226), .A2(n12167), .ZN(n14667) );
  NOR2_X1 U15264 ( .A1(n12169), .A2(n12168), .ZN(n12199) );
  INV_X1 U15265 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12173) );
  NAND2_X1 U15266 ( .A1(n12170), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12172) );
  NAND2_X1 U15267 ( .A1(n12211), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12171) );
  OAI211_X1 U15268 ( .C1(n12232), .C2(n12173), .A(n12172), .B(n12171), .ZN(
        n12174) );
  INV_X1 U15269 ( .A(n12174), .ZN(n12179) );
  AOI22_X1 U15270 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11459), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12178) );
  INV_X1 U15271 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n21087) );
  AOI22_X1 U15272 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12240), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12177) );
  NAND2_X1 U15273 ( .A1(n12175), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12176) );
  NAND4_X1 U15274 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n12193) );
  AOI22_X1 U15275 ( .A1(n12239), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11287), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12191) );
  INV_X1 U15276 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12181) );
  OAI22_X1 U15277 ( .A1(n12184), .A2(n12183), .B1(n12182), .B2(n12181), .ZN(
        n12185) );
  INV_X1 U15278 ( .A(n12185), .ZN(n12190) );
  AOI22_X1 U15279 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15280 ( .A1(n12187), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15281 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12192) );
  OR2_X1 U15282 ( .A1(n12193), .A2(n12192), .ZN(n12198) );
  XNOR2_X1 U15283 ( .A(n12199), .B(n12198), .ZN(n12196) );
  AOI21_X1 U15284 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20780), .A(
        n12654), .ZN(n12195) );
  NAND2_X1 U15285 ( .A1(n12259), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12194) );
  OAI211_X1 U15286 ( .C1(n12196), .C2(n12255), .A(n12195), .B(n12194), .ZN(
        n12197) );
  OAI21_X1 U15287 ( .B1(n11561), .B2(n14667), .A(n12197), .ZN(n14367) );
  XNOR2_X1 U15288 ( .A(n12226), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14335) );
  NAND2_X1 U15289 ( .A1(n12199), .A2(n12198), .ZN(n12249) );
  INV_X1 U15290 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15291 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12239), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15292 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12202) );
  OAI211_X1 U15293 ( .C1(n12238), .C2(n12204), .A(n12203), .B(n12202), .ZN(
        n12205) );
  INV_X1 U15294 ( .A(n12205), .ZN(n12207) );
  AOI22_X1 U15295 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12242), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12206) );
  OAI211_X1 U15296 ( .C1(n12209), .C2(n12208), .A(n12207), .B(n12206), .ZN(
        n12218) );
  AOI22_X1 U15297 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15298 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12240), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15299 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15300 ( .A1(n12212), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12211), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12213) );
  NAND4_X1 U15301 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12217) );
  NOR2_X1 U15302 ( .A1(n12218), .A2(n12217), .ZN(n12250) );
  XOR2_X1 U15303 ( .A(n12249), .B(n12250), .Z(n12223) );
  INV_X1 U15304 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14343) );
  NOR2_X1 U15305 ( .A1(n20418), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12219) );
  OAI22_X1 U15306 ( .A1(n12220), .A2(n14343), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12219), .ZN(n12221) );
  AOI21_X1 U15307 ( .B1(n12223), .B2(n12222), .A(n12221), .ZN(n12224) );
  AOI21_X1 U15308 ( .B1(n12225), .B2(n14335), .A(n12224), .ZN(n13472) );
  INV_X1 U15309 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14332) );
  INV_X1 U15310 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12644) );
  XNOR2_X1 U15311 ( .A(n12645), .B(n12644), .ZN(n14656) );
  INV_X1 U15312 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15313 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12227), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15314 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9638), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12229) );
  OAI211_X1 U15315 ( .C1(n12232), .C2(n12231), .A(n12230), .B(n12229), .ZN(
        n12233) );
  INV_X1 U15316 ( .A(n12233), .ZN(n12237) );
  AOI22_X1 U15317 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12234), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12236) );
  OAI211_X1 U15318 ( .C1(n12238), .C2(n21093), .A(n12237), .B(n12236), .ZN(
        n12248) );
  AOI22_X1 U15319 ( .A1(n12200), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12239), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15320 ( .A1(n12210), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12186), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15321 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12240), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15322 ( .A1(n12242), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11349), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12243) );
  NAND4_X1 U15323 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12247) );
  NOR2_X1 U15324 ( .A1(n12248), .A2(n12247), .ZN(n12252) );
  NOR2_X1 U15325 ( .A1(n12250), .A2(n12249), .ZN(n12251) );
  XOR2_X1 U15326 ( .A(n12252), .B(n12251), .Z(n12256) );
  AOI21_X1 U15327 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20780), .A(
        n12654), .ZN(n12254) );
  NAND2_X1 U15328 ( .A1(n12259), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12253) );
  OAI211_X1 U15329 ( .C1(n12256), .C2(n12255), .A(n12254), .B(n12253), .ZN(
        n12257) );
  OAI21_X1 U15330 ( .B1(n11561), .B2(n14656), .A(n12257), .ZN(n13402) );
  AOI22_X1 U15331 ( .A1(n12259), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12258), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12260) );
  XNOR2_X1 U15332 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U15333 ( .A1(n12286), .A2(n12285), .ZN(n12284) );
  NAND2_X1 U15334 ( .A1(n20779), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12261) );
  NAND2_X1 U15335 ( .A1(n20537), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12265) );
  NAND2_X1 U15336 ( .A1(n11241), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12262) );
  NAND2_X1 U15337 ( .A1(n12265), .A2(n12262), .ZN(n12272) );
  INV_X1 U15338 ( .A(n12272), .ZN(n12263) );
  XNOR2_X1 U15339 ( .A(n13956), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12271) );
  AOI222_X1 U15340 ( .A1(n12266), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12266), .B2(n16100), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n16100), .ZN(n12315) );
  AND2_X1 U15341 ( .A1(n12315), .A2(n12277), .ZN(n12305) );
  NOR2_X1 U15342 ( .A1(n9758), .A2(n20295), .ZN(n12288) );
  INV_X1 U15343 ( .A(n12288), .ZN(n12268) );
  NAND3_X1 U15344 ( .A1(n12287), .A2(n20275), .A3(n12268), .ZN(n12301) );
  AOI21_X1 U15345 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n12310) );
  NAND2_X1 U15346 ( .A1(n12273), .A2(n12272), .ZN(n12275) );
  NAND2_X1 U15347 ( .A1(n12275), .A2(n12274), .ZN(n12312) );
  INV_X1 U15348 ( .A(n12312), .ZN(n12276) );
  INV_X1 U15349 ( .A(n12296), .ZN(n12300) );
  NAND2_X1 U15350 ( .A1(n13621), .A2(n20295), .ZN(n12278) );
  INV_X1 U15351 ( .A(n12295), .ZN(n12299) );
  INV_X1 U15352 ( .A(n12286), .ZN(n12279) );
  OAI21_X1 U15353 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20701), .A(
        n12279), .ZN(n12281) );
  INV_X1 U15354 ( .A(n12281), .ZN(n12280) );
  OAI21_X1 U15355 ( .B1(n20261), .B2(n12586), .A(n12280), .ZN(n12283) );
  NAND2_X1 U15356 ( .A1(n12302), .A2(n12403), .ZN(n12304) );
  OAI21_X1 U15357 ( .B1(n12287), .B2(n12281), .A(n12304), .ZN(n12282) );
  OAI21_X1 U15358 ( .B1(n12283), .B2(n12295), .A(n12282), .ZN(n12290) );
  INV_X1 U15359 ( .A(n12290), .ZN(n12294) );
  OAI21_X1 U15360 ( .B1(n12286), .B2(n12285), .A(n12284), .ZN(n12313) );
  NOR2_X1 U15361 ( .A1(n12287), .A2(n13621), .ZN(n12289) );
  AOI211_X1 U15362 ( .C1(n12302), .C2(n12313), .A(n12289), .B(n12288), .ZN(
        n12291) );
  INV_X1 U15363 ( .A(n12291), .ZN(n12293) );
  AOI22_X1 U15364 ( .A1(n12291), .A2(n12290), .B1(n12301), .B2(n12313), .ZN(
        n12292) );
  AOI21_X1 U15365 ( .B1(n12294), .B2(n12293), .A(n12292), .ZN(n12298) );
  AOI211_X1 U15366 ( .C1(n12302), .C2(n12312), .A(n12296), .B(n12295), .ZN(
        n12297) );
  INV_X1 U15367 ( .A(n12306), .ZN(n12307) );
  NAND2_X1 U15368 ( .A1(n14922), .A2(n20261), .ZN(n12309) );
  NAND2_X1 U15369 ( .A1(n12309), .A2(n11405), .ZN(n12457) );
  NOR2_X1 U15370 ( .A1(n12457), .A2(n14033), .ZN(n13705) );
  INV_X1 U15371 ( .A(n12310), .ZN(n12311) );
  NOR3_X1 U15372 ( .A1(n12313), .A2(n12312), .A3(n12311), .ZN(n12316) );
  OAI21_X1 U15373 ( .B1(n12316), .B2(n12315), .A(n12314), .ZN(n13574) );
  NAND2_X1 U15374 ( .A1(n13574), .A2(n13580), .ZN(n13570) );
  AND2_X1 U15375 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20850) );
  INV_X1 U15376 ( .A(n20850), .ZN(n15768) );
  NAND2_X1 U15377 ( .A1(n13621), .A2(n15768), .ZN(n12317) );
  NOR2_X1 U15378 ( .A1(n13570), .A2(n12317), .ZN(n12318) );
  AOI21_X1 U15379 ( .B1(n15774), .B2(n13705), .A(n12318), .ZN(n13730) );
  INV_X1 U15380 ( .A(n12319), .ZN(n13711) );
  INV_X1 U15381 ( .A(n11541), .ZN(n13412) );
  AND4_X1 U15382 ( .A1(n14340), .A2(n20290), .A3(n13412), .A4(n11422), .ZN(
        n13405) );
  NAND2_X1 U15383 ( .A1(n13711), .A2(n13405), .ZN(n12322) );
  NAND2_X1 U15384 ( .A1(n15774), .A2(n15768), .ZN(n13723) );
  OR2_X1 U15385 ( .A1(n13723), .A2(n12320), .ZN(n12321) );
  NAND3_X1 U15386 ( .A1(n13730), .A2(n12322), .A3(n12321), .ZN(n12323) );
  NOR2_X1 U15387 ( .A1(n15779), .A2(n9758), .ZN(n13407) );
  INV_X2 U15388 ( .A(n13869), .ZN(n14637) );
  AND2_X1 U15389 ( .A1(n14637), .A2(n13412), .ZN(n12324) );
  NOR4_X1 U15390 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12328) );
  NOR4_X1 U15391 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12327) );
  NOR4_X1 U15392 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12326) );
  NOR4_X1 U15393 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12325) );
  AND4_X1 U15394 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12333) );
  NOR4_X1 U15395 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12331) );
  NOR4_X1 U15396 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12330) );
  NOR4_X1 U15397 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12329) );
  INV_X1 U15398 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20858) );
  AND4_X1 U15399 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n20858), .ZN(
        n12332) );
  NAND2_X1 U15400 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  AOI22_X1 U15401 ( .A1(n14633), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n13869), .ZN(n12335) );
  INV_X1 U15402 ( .A(n12335), .ZN(n12338) );
  INV_X1 U15403 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16481) );
  NOR2_X1 U15404 ( .A1(n14628), .A2(n16481), .ZN(n12337) );
  NAND2_X1 U15405 ( .A1(n12340), .A2(n12339), .ZN(P1_U2873) );
  OR2_X1 U15406 ( .A1(n12351), .A2(n12341), .ZN(n12361) );
  XNOR2_X1 U15407 ( .A(n12361), .B(n12360), .ZN(n12343) );
  AND2_X1 U15408 ( .A1(n20261), .A2(n12342), .ZN(n12350) );
  AOI21_X1 U15409 ( .B1(n12343), .B2(n15770), .A(n12350), .ZN(n12344) );
  OAI21_X1 U15410 ( .B1(n13980), .B2(n12375), .A(n12344), .ZN(n13786) );
  OAI211_X1 U15411 ( .C1(n12346), .C2(n12345), .A(n12361), .B(n15770), .ZN(
        n12347) );
  AND3_X1 U15412 ( .A1(n12347), .A2(n11405), .A3(n20295), .ZN(n12348) );
  AOI21_X1 U15413 ( .B1(n12351), .B2(n15770), .A(n12350), .ZN(n12352) );
  NAND2_X1 U15414 ( .A1(n13662), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12354) );
  INV_X1 U15415 ( .A(n12354), .ZN(n12356) );
  NAND2_X1 U15416 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  INV_X1 U15417 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20238) );
  XNOR2_X1 U15418 ( .A(n12358), .B(n20238), .ZN(n13787) );
  NAND2_X1 U15419 ( .A1(n12358), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12359) );
  INV_X1 U15420 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20220) );
  NAND2_X1 U15421 ( .A1(n20260), .A2(n12403), .ZN(n12365) );
  NAND2_X1 U15422 ( .A1(n12361), .A2(n12360), .ZN(n12380) );
  INV_X1 U15423 ( .A(n12378), .ZN(n12362) );
  XNOR2_X1 U15424 ( .A(n12380), .B(n12362), .ZN(n12363) );
  NAND2_X1 U15425 ( .A1(n12363), .A2(n15770), .ZN(n12364) );
  NAND2_X1 U15426 ( .A1(n12365), .A2(n12364), .ZN(n13910) );
  NAND2_X1 U15427 ( .A1(n12368), .A2(n12403), .ZN(n12372) );
  NAND2_X1 U15428 ( .A1(n12380), .A2(n12378), .ZN(n12369) );
  XNOR2_X1 U15429 ( .A(n12369), .B(n12377), .ZN(n12370) );
  NAND2_X1 U15430 ( .A1(n12370), .A2(n15770), .ZN(n12371) );
  NAND2_X1 U15431 ( .A1(n12372), .A2(n12371), .ZN(n12373) );
  INV_X1 U15432 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20213) );
  XNOR2_X1 U15433 ( .A(n12373), .B(n20213), .ZN(n20185) );
  NAND2_X1 U15434 ( .A1(n12373), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12374) );
  OR2_X1 U15435 ( .A1(n12376), .A2(n12375), .ZN(n12383) );
  AND2_X1 U15436 ( .A1(n12378), .A2(n12377), .ZN(n12379) );
  NAND2_X1 U15437 ( .A1(n12380), .A2(n12379), .ZN(n12387) );
  XNOR2_X1 U15438 ( .A(n12387), .B(n12388), .ZN(n12381) );
  NAND2_X1 U15439 ( .A1(n12381), .A2(n15770), .ZN(n12382) );
  NAND2_X1 U15440 ( .A1(n12383), .A2(n12382), .ZN(n12384) );
  INV_X1 U15441 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16093) );
  XNOR2_X1 U15442 ( .A(n12384), .B(n16093), .ZN(n15963) );
  NAND2_X1 U15443 ( .A1(n15964), .A2(n15963), .ZN(n15962) );
  NAND2_X1 U15444 ( .A1(n12384), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12385) );
  NAND2_X1 U15445 ( .A1(n15962), .A2(n12385), .ZN(n15959) );
  NAND3_X1 U15446 ( .A1(n12406), .A2(n12386), .A3(n12403), .ZN(n12392) );
  INV_X1 U15447 ( .A(n12387), .ZN(n12389) );
  NAND2_X1 U15448 ( .A1(n12389), .A2(n12388), .ZN(n12396) );
  XNOR2_X1 U15449 ( .A(n12396), .B(n12397), .ZN(n12390) );
  NAND2_X1 U15450 ( .A1(n12390), .A2(n15770), .ZN(n12391) );
  NAND2_X1 U15451 ( .A1(n12392), .A2(n12391), .ZN(n15957) );
  OR2_X1 U15452 ( .A1(n15957), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12393) );
  NAND2_X1 U15453 ( .A1(n15957), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12394) );
  NAND2_X1 U15454 ( .A1(n12395), .A2(n12403), .ZN(n12401) );
  INV_X1 U15455 ( .A(n12396), .ZN(n12398) );
  NAND2_X1 U15456 ( .A1(n12398), .A2(n12397), .ZN(n12410) );
  XNOR2_X1 U15457 ( .A(n12410), .B(n12407), .ZN(n12399) );
  NAND2_X1 U15458 ( .A1(n12399), .A2(n15770), .ZN(n12400) );
  NAND2_X1 U15459 ( .A1(n12401), .A2(n12400), .ZN(n12402) );
  OR2_X1 U15460 ( .A1(n12402), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15952) );
  NAND2_X1 U15461 ( .A1(n12402), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15951) );
  NAND2_X1 U15462 ( .A1(n12403), .A2(n12407), .ZN(n12404) );
  INV_X1 U15463 ( .A(n12407), .ZN(n12409) );
  INV_X1 U15464 ( .A(n15770), .ZN(n12408) );
  OR3_X1 U15465 ( .A1(n12410), .A2(n12409), .A3(n12408), .ZN(n12411) );
  NAND2_X1 U15466 ( .A1(n12419), .A2(n12411), .ZN(n14236) );
  OR2_X1 U15467 ( .A1(n14236), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12412) );
  NAND2_X1 U15468 ( .A1(n14236), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12413) );
  INV_X1 U15469 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16060) );
  NOR2_X1 U15470 ( .A1(n14761), .A2(n16060), .ZN(n12415) );
  NAND2_X1 U15471 ( .A1(n14862), .A2(n16060), .ZN(n12416) );
  INV_X1 U15472 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12613) );
  INV_X1 U15473 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16014) );
  OR2_X1 U15474 ( .A1(n12419), .A2(n16014), .ZN(n12417) );
  INV_X1 U15475 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12601) );
  AND2_X1 U15476 ( .A1(n12422), .A2(n14741), .ZN(n14727) );
  NAND2_X1 U15477 ( .A1(n12419), .A2(n12613), .ZN(n12418) );
  NAND2_X1 U15478 ( .A1(n14859), .A2(n12418), .ZN(n14855) );
  NAND2_X1 U15479 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14749) );
  OAI21_X1 U15480 ( .B1(n16014), .B2(n14749), .A(n14761), .ZN(n12420) );
  INV_X1 U15481 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12503) );
  NAND2_X1 U15482 ( .A1(n12419), .A2(n12503), .ZN(n14857) );
  NAND2_X1 U15483 ( .A1(n12420), .A2(n14857), .ZN(n12421) );
  XNOR2_X1 U15484 ( .A(n14862), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15926) );
  NAND2_X1 U15485 ( .A1(n14862), .A2(n12601), .ZN(n14740) );
  NAND2_X1 U15486 ( .A1(n15926), .A2(n14740), .ZN(n15924) );
  AOI21_X1 U15487 ( .B1(n14727), .B2(n14739), .A(n15924), .ZN(n14725) );
  NAND2_X1 U15488 ( .A1(n14725), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12426) );
  INV_X1 U15489 ( .A(n12422), .ZN(n12424) );
  NOR2_X1 U15490 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14750) );
  AND2_X1 U15491 ( .A1(n14750), .A2(n12503), .ZN(n12423) );
  NOR2_X1 U15492 ( .A1(n14761), .A2(n12423), .ZN(n14724) );
  INV_X1 U15493 ( .A(n14741), .ZN(n15922) );
  NOR2_X1 U15494 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12427) );
  INV_X1 U15495 ( .A(n12428), .ZN(n12429) );
  XNOR2_X1 U15496 ( .A(n14862), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15915) );
  NAND2_X1 U15497 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15797) );
  INV_X1 U15498 ( .A(n15797), .ZN(n12616) );
  NAND2_X1 U15499 ( .A1(n15895), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12433) );
  INV_X1 U15500 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14716) );
  INV_X1 U15501 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15994) );
  INV_X1 U15502 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15980) );
  NAND2_X1 U15503 ( .A1(n15980), .A2(n15800), .ZN(n12430) );
  INV_X1 U15504 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14702) );
  INV_X1 U15505 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14822) );
  NAND2_X1 U15506 ( .A1(n14702), .A2(n14822), .ZN(n12432) );
  INV_X1 U15507 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14660) );
  NOR2_X1 U15508 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14797) );
  INV_X1 U15509 ( .A(n14797), .ZN(n12434) );
  NOR2_X1 U15510 ( .A1(n12436), .A2(n12434), .ZN(n12435) );
  AND2_X1 U15511 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14823) );
  AND2_X1 U15512 ( .A1(n14823), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12607) );
  NAND2_X1 U15513 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12606) );
  INV_X1 U15514 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14788) );
  NAND2_X1 U15515 ( .A1(n15943), .A2(n14788), .ZN(n14650) );
  NOR2_X1 U15516 ( .A1(n14650), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12439) );
  NAND2_X1 U15517 ( .A1(n14761), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13468) );
  INV_X1 U15518 ( .A(n13468), .ZN(n12437) );
  AOI22_X1 U15519 ( .A1(n13469), .A2(n12439), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14649), .ZN(n12441) );
  OR2_X1 U15520 ( .A1(n12442), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15791) );
  AOI21_X1 U15521 ( .B1(n20275), .B2(n15791), .A(n20850), .ZN(n12443) );
  NAND2_X1 U15522 ( .A1(n13574), .A2(n12443), .ZN(n12449) );
  NAND2_X1 U15523 ( .A1(n13621), .A2(n15791), .ZN(n12663) );
  AND2_X1 U15524 ( .A1(n12663), .A2(n15768), .ZN(n12445) );
  NAND2_X1 U15525 ( .A1(n12444), .A2(n12445), .ZN(n15769) );
  NAND3_X1 U15526 ( .A1(n15769), .A2(n11404), .A3(n12446), .ZN(n12447) );
  NAND2_X1 U15527 ( .A1(n15774), .A2(n12447), .ZN(n12448) );
  MUX2_X1 U15528 ( .A(n12449), .B(n12448), .S(n20280), .Z(n12456) );
  NOR2_X1 U15529 ( .A1(n14922), .A2(n13621), .ZN(n12597) );
  INV_X1 U15530 ( .A(n12597), .ZN(n12450) );
  OR2_X1 U15531 ( .A1(n13870), .A2(n11474), .ZN(n12451) );
  NAND2_X1 U15532 ( .A1(n10097), .A2(n12451), .ZN(n12585) );
  NOR2_X1 U15533 ( .A1(n12457), .A2(n12585), .ZN(n12453) );
  OAI21_X1 U15534 ( .B1(n13580), .B2(n12453), .A(n12452), .ZN(n13726) );
  INV_X1 U15535 ( .A(n13726), .ZN(n12454) );
  INV_X1 U15536 ( .A(n13407), .ZN(n20010) );
  INV_X1 U15537 ( .A(n12598), .ZN(n12461) );
  NOR2_X1 U15538 ( .A1(n12585), .A2(n12586), .ZN(n12639) );
  INV_X1 U15539 ( .A(n14033), .ZN(n13569) );
  OR2_X1 U15540 ( .A1(n12639), .A2(n13569), .ZN(n12458) );
  INV_X1 U15541 ( .A(n12457), .ZN(n12638) );
  NAND2_X1 U15542 ( .A1(n12458), .A2(n12638), .ZN(n13576) );
  OAI211_X1 U15543 ( .C1(n20290), .C2(n12582), .A(n11438), .B(n13576), .ZN(
        n12459) );
  INV_X1 U15544 ( .A(n12459), .ZN(n12460) );
  INV_X1 U15545 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20254) );
  INV_X1 U15546 ( .A(n12566), .ZN(n12462) );
  OAI21_X1 U15547 ( .B1(n12534), .B2(n20254), .A(n12533), .ZN(n12463) );
  INV_X1 U15548 ( .A(n12463), .ZN(n12465) );
  MUX2_X1 U15549 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12464) );
  NAND2_X1 U15550 ( .A1(n12465), .A2(n12464), .ZN(n12468) );
  NAND2_X1 U15551 ( .A1(n12566), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12467) );
  INV_X1 U15552 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13904) );
  NAND2_X1 U15553 ( .A1(n12555), .A2(n13904), .ZN(n12466) );
  NAND2_X1 U15554 ( .A1(n12467), .A2(n12466), .ZN(n13901) );
  XNOR2_X1 U15555 ( .A(n12468), .B(n13901), .ZN(n20089) );
  INV_X1 U15556 ( .A(n12468), .ZN(n12469) );
  AOI21_X1 U15557 ( .B1(n20089), .B2(n13573), .A(n12469), .ZN(n13858) );
  OAI21_X1 U15558 ( .B1(n12534), .B2(n20238), .A(n12533), .ZN(n12470) );
  INV_X1 U15559 ( .A(n12470), .ZN(n12472) );
  MUX2_X1 U15560 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12471) );
  NAND2_X1 U15561 ( .A1(n12472), .A2(n12471), .ZN(n13857) );
  INV_X1 U15562 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12473) );
  NAND2_X1 U15563 ( .A1(n12553), .A2(n12473), .ZN(n12477) );
  NAND2_X1 U15564 ( .A1(n13573), .A2(n12473), .ZN(n12475) );
  NAND2_X1 U15565 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12474) );
  NAND3_X1 U15566 ( .A1(n12475), .A2(n12474), .A3(n12566), .ZN(n12476) );
  AND2_X1 U15567 ( .A1(n12477), .A2(n12476), .ZN(n13886) );
  MUX2_X1 U15568 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12479) );
  NAND2_X1 U15569 ( .A1(n12568), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12478) );
  INV_X1 U15570 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20115) );
  NAND2_X1 U15571 ( .A1(n13573), .A2(n20115), .ZN(n12483) );
  NAND2_X1 U15572 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12482) );
  NAND3_X1 U15573 ( .A1(n12483), .A2(n12482), .A3(n12566), .ZN(n12484) );
  OAI21_X1 U15574 ( .B1(n12564), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12484), .ZN(
        n16086) );
  INV_X1 U15575 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16080) );
  OAI21_X1 U15576 ( .B1(n12534), .B2(n16080), .A(n12533), .ZN(n12485) );
  INV_X1 U15577 ( .A(n12485), .ZN(n12487) );
  MUX2_X1 U15578 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12486) );
  NAND2_X1 U15579 ( .A1(n12487), .A2(n12486), .ZN(n14071) );
  INV_X1 U15580 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20035) );
  NAND2_X1 U15581 ( .A1(n12553), .A2(n20035), .ZN(n12491) );
  NAND2_X1 U15582 ( .A1(n13573), .A2(n20035), .ZN(n12489) );
  NAND2_X1 U15583 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12488) );
  NAND3_X1 U15584 ( .A1(n12489), .A2(n12488), .A3(n12566), .ZN(n12490) );
  AND2_X1 U15585 ( .A1(n12491), .A2(n12490), .ZN(n14005) );
  MUX2_X1 U15586 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12493) );
  NAND2_X1 U15587 ( .A1(n12568), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12492) );
  INV_X1 U15588 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U15589 ( .A1(n13573), .A2(n14178), .ZN(n12495) );
  NAND2_X1 U15590 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12494) );
  NAND3_X1 U15591 ( .A1(n12495), .A2(n12494), .A3(n12566), .ZN(n12496) );
  OAI21_X1 U15592 ( .B1(n12564), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12496), .ZN(
        n14163) );
  MUX2_X1 U15593 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12498) );
  NAND2_X1 U15594 ( .A1(n12568), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12497) );
  INV_X1 U15595 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15893) );
  NAND2_X1 U15596 ( .A1(n12553), .A2(n15893), .ZN(n12502) );
  NAND2_X1 U15597 ( .A1(n13573), .A2(n15893), .ZN(n12500) );
  NAND2_X1 U15598 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12499) );
  NAND3_X1 U15599 ( .A1(n12500), .A2(n12499), .A3(n12566), .ZN(n12501) );
  OAI21_X1 U15600 ( .B1(n12534), .B2(n12503), .A(n12533), .ZN(n12504) );
  INV_X1 U15601 ( .A(n12504), .ZN(n12506) );
  MUX2_X1 U15602 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12505) );
  NAND2_X1 U15603 ( .A1(n12506), .A2(n12505), .ZN(n14565) );
  INV_X1 U15604 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14559) );
  NAND2_X1 U15605 ( .A1(n12553), .A2(n14559), .ZN(n12510) );
  NAND2_X1 U15606 ( .A1(n13573), .A2(n14559), .ZN(n12508) );
  NAND2_X1 U15607 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12507) );
  NAND3_X1 U15608 ( .A1(n12508), .A2(n12507), .A3(n12566), .ZN(n12509) );
  AND2_X1 U15609 ( .A1(n12510), .A2(n12509), .ZN(n14477) );
  NAND2_X1 U15610 ( .A1(n14565), .A2(n14477), .ZN(n12511) );
  OAI21_X1 U15611 ( .B1(n12534), .B2(n16014), .A(n12533), .ZN(n12512) );
  INV_X1 U15612 ( .A(n12512), .ZN(n12514) );
  MUX2_X1 U15613 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12513) );
  NAND2_X1 U15614 ( .A1(n12514), .A2(n12513), .ZN(n14555) );
  INV_X1 U15615 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14550) );
  NAND2_X1 U15616 ( .A1(n12553), .A2(n14550), .ZN(n12518) );
  NAND2_X1 U15617 ( .A1(n13573), .A2(n14550), .ZN(n12516) );
  NAND2_X1 U15618 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12515) );
  NAND3_X1 U15619 ( .A1(n12516), .A2(n12515), .A3(n12566), .ZN(n12517) );
  AND2_X1 U15620 ( .A1(n12518), .A2(n12517), .ZN(n14462) );
  NAND2_X1 U15621 ( .A1(n14555), .A2(n14462), .ZN(n12519) );
  INV_X1 U15622 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16015) );
  OAI21_X1 U15623 ( .B1(n12534), .B2(n16015), .A(n12533), .ZN(n12520) );
  INV_X1 U15624 ( .A(n12520), .ZN(n12522) );
  MUX2_X1 U15625 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12521) );
  NAND2_X1 U15626 ( .A1(n12522), .A2(n12521), .ZN(n14543) );
  OR2_X1 U15627 ( .A1(n12524), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12526) );
  NAND2_X1 U15628 ( .A1(n12584), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n12525) );
  OAI211_X1 U15629 ( .C1(n12564), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12526), .B(
        n12525), .ZN(n12527) );
  INV_X1 U15630 ( .A(n12527), .ZN(n14447) );
  MUX2_X1 U15631 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12529) );
  NAND2_X1 U15632 ( .A1(n12568), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12528) );
  AND3_X1 U15633 ( .A1(n12529), .A2(n12533), .A3(n12528), .ZN(n14535) );
  INV_X1 U15634 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14529) );
  NAND2_X1 U15635 ( .A1(n13573), .A2(n14529), .ZN(n12531) );
  NAND2_X1 U15636 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12530) );
  NAND3_X1 U15637 ( .A1(n12531), .A2(n12530), .A3(n12566), .ZN(n12532) );
  OAI21_X1 U15638 ( .B1(n12564), .B2(P1_EBX_REG_19__SCAN_IN), .A(n12532), .ZN(
        n14434) );
  OAI21_X1 U15639 ( .B1(n12534), .B2(n15800), .A(n12533), .ZN(n12535) );
  INV_X1 U15640 ( .A(n12535), .ZN(n12537) );
  MUX2_X1 U15641 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12536) );
  NAND2_X1 U15642 ( .A1(n12537), .A2(n12536), .ZN(n14521) );
  INV_X1 U15643 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n12538) );
  NAND2_X1 U15644 ( .A1(n12553), .A2(n12538), .ZN(n12542) );
  NAND2_X1 U15645 ( .A1(n13573), .A2(n12538), .ZN(n12540) );
  NAND2_X1 U15646 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12539) );
  NAND3_X1 U15647 ( .A1(n12540), .A2(n12539), .A3(n12566), .ZN(n12541) );
  AND2_X1 U15648 ( .A1(n12542), .A2(n12541), .ZN(n14424) );
  INV_X1 U15649 ( .A(n12567), .ZN(n12543) );
  INV_X1 U15650 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15833) );
  NAND2_X1 U15651 ( .A1(n12543), .A2(n15833), .ZN(n12547) );
  INV_X1 U15652 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15979) );
  NAND2_X1 U15653 ( .A1(n12566), .A2(n15979), .ZN(n12545) );
  NAND2_X1 U15654 ( .A1(n13573), .A2(n15833), .ZN(n12544) );
  NAND3_X1 U15655 ( .A1(n12545), .A2(n12555), .A3(n12544), .ZN(n12546) );
  AND2_X1 U15656 ( .A1(n12547), .A2(n12546), .ZN(n14514) );
  INV_X1 U15657 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14508) );
  NAND2_X1 U15658 ( .A1(n13573), .A2(n14508), .ZN(n12549) );
  NAND2_X1 U15659 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12548) );
  NAND3_X1 U15660 ( .A1(n12549), .A2(n12548), .A3(n12566), .ZN(n12550) );
  OAI21_X1 U15661 ( .B1(n12564), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12550), .ZN(
        n14505) );
  MUX2_X1 U15662 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12552) );
  NAND2_X1 U15663 ( .A1(n12568), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12551) );
  AND2_X1 U15664 ( .A1(n12552), .A2(n12551), .ZN(n14500) );
  INV_X1 U15665 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n12554) );
  NAND2_X1 U15666 ( .A1(n12553), .A2(n12554), .ZN(n12559) );
  NAND2_X1 U15667 ( .A1(n13573), .A2(n12554), .ZN(n12557) );
  NAND2_X1 U15668 ( .A1(n12555), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12556) );
  NAND3_X1 U15669 ( .A1(n12557), .A2(n12556), .A3(n12566), .ZN(n12558) );
  AND2_X1 U15670 ( .A1(n12559), .A2(n12558), .ZN(n14415) );
  MUX2_X1 U15671 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12561) );
  NAND2_X1 U15672 ( .A1(n12568), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12560) );
  NAND2_X1 U15673 ( .A1(n12561), .A2(n12560), .ZN(n14400) );
  OR2_X1 U15674 ( .A1(n12524), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12563) );
  NAND2_X1 U15675 ( .A1(n12584), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n12562) );
  OAI211_X1 U15676 ( .C1(n12564), .C2(P1_EBX_REG_27__SCAN_IN), .A(n12563), .B(
        n12562), .ZN(n12565) );
  INV_X1 U15677 ( .A(n12565), .ZN(n14387) );
  MUX2_X1 U15678 ( .A(n12567), .B(n12566), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12570) );
  NAND2_X1 U15679 ( .A1(n12568), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12569) );
  AND2_X1 U15680 ( .A1(n12570), .A2(n12569), .ZN(n14370) );
  OR2_X1 U15681 ( .A1(n12524), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12571) );
  INV_X1 U15682 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14347) );
  NAND2_X1 U15683 ( .A1(n13573), .A2(n14347), .ZN(n12572) );
  NAND2_X1 U15684 ( .A1(n12571), .A2(n12572), .ZN(n13409) );
  MUX2_X1 U15685 ( .A(n13409), .B(n12572), .S(n12584), .Z(n14329) );
  NAND2_X1 U15686 ( .A1(n12524), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12575) );
  NAND2_X1 U15687 ( .A1(n12573), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12574) );
  NAND2_X1 U15688 ( .A1(n12575), .A2(n12574), .ZN(n13410) );
  AOI22_X1 U15689 ( .A1(n12524), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n12573), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12578) );
  INV_X1 U15690 ( .A(n12578), .ZN(n12579) );
  OR2_X1 U15691 ( .A1(n13575), .A2(n20275), .ZN(n13626) );
  OAI21_X1 U15692 ( .B1(n12582), .B2(n11474), .A(n13626), .ZN(n12583) );
  NAND2_X1 U15693 ( .A1(n12585), .A2(n12584), .ZN(n12588) );
  INV_X1 U15694 ( .A(n14036), .ZN(n12587) );
  NAND2_X1 U15695 ( .A1(n12587), .A2(n12586), .ZN(n12594) );
  AND2_X1 U15696 ( .A1(n12588), .A2(n12594), .ZN(n12589) );
  AND2_X1 U15697 ( .A1(n12590), .A2(n12589), .ZN(n13704) );
  NAND3_X1 U15698 ( .A1(n13704), .A2(n12592), .A3(n12591), .ZN(n12593) );
  INV_X1 U15699 ( .A(n14823), .ZN(n12605) );
  AND2_X1 U15700 ( .A1(n13580), .A2(n20275), .ZN(n15750) );
  AND2_X1 U15701 ( .A1(n12595), .A2(n12594), .ZN(n12596) );
  NAND2_X1 U15702 ( .A1(n12597), .A2(n12596), .ZN(n13403) );
  INV_X1 U15703 ( .A(n13403), .ZN(n13706) );
  INV_X1 U15704 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20223) );
  NAND2_X1 U15705 ( .A1(n14902), .A2(n20223), .ZN(n12599) );
  OR2_X1 U15706 ( .A1(n12598), .A2(n20209), .ZN(n20253) );
  NAND2_X1 U15707 ( .A1(n20242), .A2(n16044), .ZN(n16066) );
  INV_X1 U15708 ( .A(n20226), .ZN(n14889) );
  NAND2_X1 U15709 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16045) );
  NAND2_X1 U15710 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20210) );
  NOR2_X1 U15711 ( .A1(n16093), .A2(n20210), .ZN(n14865) );
  INV_X1 U15712 ( .A(n14865), .ZN(n12600) );
  INV_X1 U15713 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16072) );
  INV_X1 U15714 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16078) );
  NOR3_X1 U15715 ( .A1(n16072), .A2(n16078), .A3(n16080), .ZN(n16046) );
  NAND3_X1 U15716 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16046), .ZN(n14886) );
  NOR3_X1 U15717 ( .A1(n16045), .A2(n12600), .A3(n14886), .ZN(n14888) );
  NAND3_X1 U15718 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n14888), .ZN(n16028) );
  NOR2_X1 U15719 ( .A1(n12601), .A2(n16015), .ZN(n16011) );
  NAND3_X1 U15720 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n16011), .ZN(n16001) );
  NOR2_X1 U15721 ( .A1(n16001), .A2(n15994), .ZN(n12617) );
  NAND2_X1 U15722 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12617), .ZN(
        n14849) );
  NOR2_X1 U15723 ( .A1(n16028), .A2(n14849), .ZN(n14850) );
  NAND2_X1 U15724 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12611) );
  OAI21_X1 U15725 ( .B1(n20223), .B2(n20254), .A(n20238), .ZN(n20228) );
  NAND2_X1 U15726 ( .A1(n14865), .A2(n20228), .ZN(n16061) );
  OR3_X1 U15727 ( .A1(n14886), .A2(n12611), .A3(n16061), .ZN(n14869) );
  OAI21_X1 U15728 ( .B1(n14849), .B2(n14869), .A(n20206), .ZN(n12602) );
  OAI211_X1 U15729 ( .C1(n14889), .C2(n14850), .A(n16044), .B(n12602), .ZN(
        n15988) );
  NAND2_X1 U15730 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15981) );
  INV_X1 U15731 ( .A(n15981), .ZN(n12603) );
  NAND2_X1 U15732 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n12603), .ZN(
        n12604) );
  INV_X1 U15733 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14782) );
  INV_X1 U15734 ( .A(n12606), .ZN(n14798) );
  NAND2_X1 U15735 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12609) );
  INV_X1 U15736 ( .A(n12607), .ZN(n14818) );
  AOI22_X1 U15737 ( .A1(n20206), .A2(n14702), .B1(n15798), .B2(n14818), .ZN(
        n12608) );
  NAND2_X1 U15738 ( .A1(n12610), .A2(n12608), .ZN(n14833) );
  AOI21_X1 U15739 ( .B1(n16013), .B2(n12609), .A(n14833), .ZN(n14803) );
  OAI21_X1 U15740 ( .B1(n20242), .B2(n14798), .A(n14803), .ZN(n14793) );
  AOI211_X1 U15741 ( .C1(n16013), .C2(n14788), .A(n14782), .B(n14793), .ZN(
        n14780) );
  AOI211_X1 U15742 ( .C1(n12610), .C2(n20242), .A(n12440), .B(n14780), .ZN(
        n12620) );
  INV_X1 U15743 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20909) );
  NOR2_X1 U15744 ( .A1(n20244), .A2(n20909), .ZN(n12647) );
  NOR2_X1 U15745 ( .A1(n12613), .A2(n12611), .ZN(n14879) );
  NAND2_X1 U15746 ( .A1(n14888), .A2(n14879), .ZN(n14871) );
  INV_X1 U15747 ( .A(n14871), .ZN(n12612) );
  NAND2_X1 U15748 ( .A1(n20222), .A2(n12612), .ZN(n12615) );
  NAND2_X1 U15749 ( .A1(n12615), .A2(n12614), .ZN(n16002) );
  AND4_X1 U15750 ( .A1(n12617), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n12616), .A4(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12618) );
  NOR3_X1 U15751 ( .A1(n14836), .A2(n14818), .A3(n14660), .ZN(n14808) );
  NAND3_X1 U15752 ( .A1(n14808), .A2(n14798), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14781) );
  NOR3_X1 U15753 ( .A1(n14781), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14782), .ZN(n12619) );
  NOR2_X1 U15754 ( .A1(n12621), .A2(n15117), .ZN(n12623) );
  XOR2_X1 U15755 ( .A(n12623), .B(n12622), .Z(n13094) );
  OAI21_X1 U15756 ( .B1(n12624), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12625), .ZN(n13083) );
  NOR2_X1 U15757 ( .A1(n13083), .A2(n19343), .ZN(n12628) );
  INV_X1 U15758 ( .A(n15289), .ZN(n15303) );
  OAI21_X1 U15759 ( .B1(n12626), .B2(n15303), .A(n15302), .ZN(n15295) );
  NOR2_X1 U15760 ( .A1(n15045), .A2(n12630), .ZN(n12631) );
  INV_X1 U15761 ( .A(n16124), .ZN(n14353) );
  NAND2_X1 U15762 ( .A1(n14353), .A2(n16350), .ZN(n12636) );
  OAI21_X1 U15763 ( .B1(n14970), .B2(n12632), .A(n12743), .ZN(n16125) );
  NOR3_X1 U15764 ( .A1(n15303), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15288), .ZN(n12633) );
  NOR2_X1 U15765 ( .A1(n19328), .A2(n19921), .ZN(n13089) );
  OAI211_X1 U15766 ( .C1(n13094), .C2(n19331), .A(n12637), .B(n10069), .ZN(
        P2_U3017) );
  NAND2_X1 U15767 ( .A1(n12640), .A2(n20200), .ZN(n12651) );
  AND3_X1 U15768 ( .A1(n9758), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16104) );
  NOR2_X2 U15769 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20791) );
  NAND2_X1 U15770 ( .A1(n20782), .A2(n12641), .ZN(n20936) );
  AND2_X1 U15771 ( .A1(n20936), .A2(n9758), .ZN(n12642) );
  NOR2_X1 U15772 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20780), .ZN(n20938) );
  AOI21_X1 U15773 ( .B1(n20418), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n20938), 
        .ZN(n13660) );
  INV_X1 U15774 ( .A(n13660), .ZN(n12643) );
  NOR2_X1 U15775 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  XNOR2_X1 U15776 ( .A(n12646), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14043) );
  AOI21_X1 U15777 ( .B1(n20194), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12647), .ZN(n12648) );
  OAI21_X1 U15778 ( .B1(n20193), .B2(n14043), .A(n12648), .ZN(n12649) );
  AOI21_X1 U15779 ( .B1(n12658), .B2(n20189), .A(n12649), .ZN(n12650) );
  NAND2_X1 U15780 ( .A1(n12651), .A2(n12650), .ZN(P1_U2968) );
  INV_X1 U15781 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20671) );
  NOR3_X1 U15782 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n20671), .ZN(n15775) );
  INV_X1 U15783 ( .A(n13570), .ZN(n12652) );
  NAND2_X1 U15784 ( .A1(n12652), .A2(n13407), .ZN(n13525) );
  AND2_X1 U15785 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n9758), .ZN(n12653) );
  NAND2_X1 U15786 ( .A1(n12654), .A2(n12653), .ZN(n12655) );
  NOR2_X1 U15787 ( .A1(n14043), .A2(n16108), .ZN(n12657) );
  NAND2_X1 U15788 ( .A1(n12658), .A2(n20052), .ZN(n12680) );
  INV_X1 U15789 ( .A(n12669), .ZN(n12661) );
  NAND2_X1 U15790 ( .A1(n20275), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12667) );
  NOR2_X1 U15791 ( .A1(n20850), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12662) );
  NOR2_X1 U15792 ( .A1(n12667), .A2(n12662), .ZN(n12660) );
  NAND2_X1 U15793 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12672) );
  INV_X1 U15794 ( .A(n12672), .ZN(n12666) );
  NAND2_X1 U15795 ( .A1(n12663), .A2(n12662), .ZN(n12670) );
  NAND2_X1 U15796 ( .A1(n20092), .A2(n20071), .ZN(n20100) );
  INV_X1 U15797 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20897) );
  INV_X1 U15798 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20867) );
  INV_X1 U15799 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20862) );
  NAND3_X1 U15800 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20070) );
  NOR2_X1 U15801 ( .A1(n20862), .A2(n20070), .ZN(n20072) );
  NAND3_X1 U15802 ( .A1(n20072), .A2(P1_REIP_REG_6__SCAN_IN), .A3(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20032) );
  NOR2_X1 U15803 ( .A1(n20867), .A2(n20032), .ZN(n14177) );
  NAND2_X1 U15804 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14177), .ZN(n14100) );
  NAND2_X1 U15805 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14433) );
  NAND4_X1 U15806 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14431) );
  NAND3_X1 U15807 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14437) );
  NOR2_X1 U15808 ( .A1(n14431), .A2(n14437), .ZN(n14436) );
  NAND4_X1 U15809 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14436), .A3(
        P1_REIP_REG_20__SCAN_IN), .A4(P1_REIP_REG_19__SCAN_IN), .ZN(n12664) );
  NOR2_X1 U15810 ( .A1(n14433), .A2(n12664), .ZN(n14421) );
  NAND4_X1 U15811 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14421), .A3(
        P1_REIP_REG_22__SCAN_IN), .A4(P1_REIP_REG_21__SCAN_IN), .ZN(n14410) );
  NOR2_X1 U15812 ( .A1(n14100), .A2(n14410), .ZN(n15813) );
  NAND2_X1 U15813 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15813), .ZN(n14409) );
  NOR2_X1 U15814 ( .A1(n20897), .A2(n14409), .ZN(n14394) );
  AND2_X1 U15815 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n14394), .ZN(n14381) );
  AND2_X1 U15816 ( .A1(n20092), .A2(n14381), .ZN(n14380) );
  NAND3_X1 U15817 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .A3(n14380), .ZN(n12665) );
  NAND2_X1 U15818 ( .A1(n20100), .A2(n12665), .ZN(n14371) );
  OAI21_X1 U15819 ( .B1(n12666), .B2(n20071), .A(n14371), .ZN(n14362) );
  INV_X1 U15820 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12675) );
  INV_X1 U15821 ( .A(n12667), .ZN(n12668) );
  NOR2_X1 U15822 ( .A1(n12669), .A2(n12668), .ZN(n12671) );
  AND3_X1 U15823 ( .A1(n20090), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14381), 
        .ZN(n14373) );
  NAND2_X1 U15824 ( .A1(n14373), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14358) );
  NOR3_X1 U15825 ( .A1(n14358), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n12672), 
        .ZN(n12673) );
  AOI21_X1 U15826 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(n20103), .A(n12673), .ZN(
        n12674) );
  OAI21_X1 U15827 ( .B1(n20102), .B2(n12675), .A(n12674), .ZN(n12676) );
  AOI21_X1 U15828 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(n14362), .A(n12676), 
        .ZN(n12677) );
  NAND2_X1 U15829 ( .A1(n12680), .A2(n12679), .ZN(P1_U2809) );
  NAND2_X1 U15830 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12683), .ZN(
        n12684) );
  INV_X1 U15831 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16256) );
  INV_X1 U15832 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19008) );
  INV_X1 U15833 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18985) );
  INV_X1 U15834 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18963) );
  INV_X1 U15835 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16224) );
  INV_X1 U15836 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12705) );
  INV_X1 U15837 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12709) );
  INV_X1 U15838 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15143) );
  XNOR2_X1 U15839 ( .A(n12713), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16118) );
  AOI21_X1 U15840 ( .B1(n16256), .B2(n12692), .A(n12681), .ZN(n19020) );
  AOI21_X1 U15841 ( .B1(n15244), .B2(n12690), .A(n12682), .ZN(n19041) );
  AOI21_X1 U15842 ( .B1(n16284), .B2(n12688), .A(n12691), .ZN(n19064) );
  AOI21_X1 U15843 ( .B1(n15268), .B2(n12687), .A(n12689), .ZN(n19081) );
  AOI21_X1 U15844 ( .B1(n19104), .B2(n12685), .A(n9651), .ZN(n19109) );
  AOI21_X1 U15845 ( .B1(n19301), .B2(n12684), .A(n12686), .ZN(n19289) );
  AOI21_X1 U15846 ( .B1(n19311), .B2(n14953), .A(n12683), .ZN(n14122) );
  AOI22_X1 U15847 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13085), .ZN(n14961) );
  AOI22_X1 U15848 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14953), .B2(n13085), .ZN(
        n14960) );
  NAND2_X1 U15849 ( .A1(n14961), .A2(n14960), .ZN(n14959) );
  NOR2_X1 U15850 ( .A1(n14122), .A2(n14959), .ZN(n14939) );
  OAI21_X1 U15851 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12683), .A(
        n12684), .ZN(n14940) );
  NAND2_X1 U15852 ( .A1(n14939), .A2(n14940), .ZN(n19132) );
  NOR2_X1 U15853 ( .A1(n19289), .A2(n19132), .ZN(n19117) );
  OAI21_X1 U15854 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12686), .A(
        n12685), .ZN(n19119) );
  NAND2_X1 U15855 ( .A1(n19117), .A2(n19119), .ZN(n19107) );
  NOR2_X1 U15856 ( .A1(n19109), .A2(n19107), .ZN(n19094) );
  OAI21_X1 U15857 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n9651), .A(
        n12687), .ZN(n19095) );
  NAND2_X1 U15858 ( .A1(n19094), .A2(n19095), .ZN(n19079) );
  NOR2_X1 U15859 ( .A1(n19081), .A2(n19079), .ZN(n19069) );
  OAI21_X1 U15860 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n12689), .A(
        n12688), .ZN(n19071) );
  NAND2_X1 U15861 ( .A1(n19069), .A2(n19071), .ZN(n19062) );
  NOR2_X1 U15862 ( .A1(n19064), .A2(n19062), .ZN(n19049) );
  OAI21_X1 U15863 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12691), .A(
        n12690), .ZN(n19051) );
  NAND2_X1 U15864 ( .A1(n19049), .A2(n19051), .ZN(n19039) );
  NOR2_X1 U15865 ( .A1(n19041), .A2(n19039), .ZN(n19030) );
  OAI21_X1 U15866 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n12682), .A(
        n12692), .ZN(n19032) );
  NAND2_X1 U15867 ( .A1(n19030), .A2(n19032), .ZN(n19018) );
  NOR2_X1 U15868 ( .A1(n19020), .A2(n19018), .ZN(n19010) );
  AOI21_X1 U15869 ( .B1(n19008), .B2(n12694), .A(n12693), .ZN(n16237) );
  INV_X1 U15870 ( .A(n16237), .ZN(n19012) );
  NAND2_X1 U15871 ( .A1(n19010), .A2(n19012), .ZN(n18996) );
  OAI21_X1 U15872 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12693), .A(
        n12696), .ZN(n18998) );
  INV_X1 U15873 ( .A(n18998), .ZN(n12695) );
  AOI21_X1 U15874 ( .B1(n18985), .B2(n12696), .A(n12698), .ZN(n12697) );
  INV_X1 U15875 ( .A(n12697), .ZN(n18992) );
  NAND2_X1 U15876 ( .A1(n18991), .A2(n18992), .ZN(n18990) );
  NAND2_X1 U15877 ( .A1(n9704), .A2(n18990), .ZN(n18979) );
  OAI21_X1 U15878 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12698), .A(
        n12699), .ZN(n18980) );
  NAND2_X1 U15879 ( .A1(n18979), .A2(n18980), .ZN(n18978) );
  NAND2_X1 U15880 ( .A1(n18978), .A2(n9704), .ZN(n18968) );
  AOI21_X1 U15881 ( .B1(n18963), .B2(n12699), .A(n12700), .ZN(n16226) );
  INV_X1 U15882 ( .A(n16226), .ZN(n18969) );
  OAI21_X1 U15883 ( .B1(n12700), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n9718), .ZN(n18957) );
  AOI21_X1 U15884 ( .B1(n18941), .B2(n9718), .A(n12701), .ZN(n15202) );
  INV_X1 U15885 ( .A(n15202), .ZN(n18948) );
  NAND2_X1 U15886 ( .A1(n18946), .A2(n9704), .ZN(n15740) );
  OAI21_X1 U15887 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12701), .A(
        n12702), .ZN(n15741) );
  NAND2_X1 U15888 ( .A1(n15740), .A2(n15741), .ZN(n15739) );
  NAND2_X1 U15889 ( .A1(n15739), .A2(n9704), .ZN(n16190) );
  AOI21_X1 U15890 ( .B1(n16224), .B2(n12702), .A(n12703), .ZN(n16216) );
  INV_X1 U15891 ( .A(n16216), .ZN(n16191) );
  OAI21_X1 U15892 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12703), .A(
        n12704), .ZN(n16183) );
  AOI21_X1 U15893 ( .B1(n12704), .B2(n12705), .A(n9716), .ZN(n15174) );
  INV_X1 U15894 ( .A(n15174), .ZN(n16171) );
  NAND2_X1 U15895 ( .A1(n16169), .A2(n9704), .ZN(n16159) );
  OR2_X1 U15896 ( .A1(n9716), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12706) );
  NAND2_X1 U15897 ( .A1(n12708), .A2(n12706), .ZN(n16160) );
  NAND2_X1 U15898 ( .A1(n16159), .A2(n16160), .ZN(n16158) );
  NAND2_X1 U15899 ( .A1(n16158), .A2(n9704), .ZN(n16149) );
  INV_X1 U15900 ( .A(n12710), .ZN(n12707) );
  AOI21_X1 U15901 ( .B1(n12709), .B2(n12708), .A(n12707), .ZN(n15151) );
  INV_X1 U15902 ( .A(n15151), .ZN(n16150) );
  NAND2_X1 U15903 ( .A1(n16148), .A2(n9704), .ZN(n16138) );
  AND2_X1 U15904 ( .A1(n12710), .A2(n15143), .ZN(n12711) );
  OR2_X1 U15905 ( .A1(n12711), .A2(n12712), .ZN(n16139) );
  NAND2_X1 U15906 ( .A1(n16138), .A2(n16139), .ZN(n16137) );
  NAND2_X1 U15907 ( .A1(n16137), .A2(n9704), .ZN(n16128) );
  INV_X1 U15908 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12715) );
  INV_X1 U15909 ( .A(n12712), .ZN(n12714) );
  AOI21_X1 U15910 ( .B1(n12715), .B2(n12714), .A(n12713), .ZN(n13092) );
  INV_X1 U15911 ( .A(n13092), .ZN(n16129) );
  NAND2_X1 U15912 ( .A1(n9704), .A2(n16127), .ZN(n16117) );
  INV_X1 U15913 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n18922) );
  NAND4_X1 U15914 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19777), .A3(n13085), 
        .A4(n18922), .ZN(n19847) );
  AOI21_X1 U15915 ( .B1(n16118), .B2(n16117), .A(n19847), .ZN(n12719) );
  INV_X1 U15916 ( .A(n16117), .ZN(n12717) );
  INV_X1 U15917 ( .A(n16118), .ZN(n12716) );
  NAND2_X1 U15918 ( .A1(n12719), .A2(n12718), .ZN(n12749) );
  INV_X1 U15919 ( .A(n12629), .ZN(n12722) );
  INV_X1 U15920 ( .A(n12720), .ZN(n12721) );
  NAND2_X1 U15921 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  NAND2_X1 U15922 ( .A1(n13514), .A2(n19843), .ZN(n12728) );
  INV_X1 U15923 ( .A(n12728), .ZN(n12725) );
  AND2_X1 U15924 ( .A1(n11189), .A2(n12725), .ZN(n18920) );
  INV_X1 U15925 ( .A(n13511), .ZN(n13769) );
  NOR2_X1 U15926 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13769), .ZN(n12734) );
  AND2_X1 U15927 ( .A1(n12726), .A2(n12734), .ZN(n16397) );
  NOR2_X1 U15928 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19864), .ZN(n12744) );
  INV_X1 U15929 ( .A(n12744), .ZN(n12735) );
  AND2_X1 U15930 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12735), .ZN(n12729) );
  NOR2_X1 U15931 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19950), .ZN(n19721) );
  NAND2_X1 U15932 ( .A1(n12730), .A2(n19721), .ZN(n16408) );
  NAND3_X1 U15933 ( .A1(n19328), .A2(n16408), .A3(n19847), .ZN(n12731) );
  OAI22_X1 U15934 ( .A1(n12732), .A2(n19149), .B1(n19925), .B2(n19142), .ZN(
        n12741) );
  INV_X1 U15935 ( .A(n13510), .ZN(n12733) );
  NOR2_X1 U15936 ( .A1(n13549), .A2(n12734), .ZN(n16114) );
  INV_X1 U15937 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12736) );
  NAND2_X1 U15938 ( .A1(n12736), .A2(n12735), .ZN(n12737) );
  NOR2_X1 U15939 ( .A1(n13510), .A2(n12737), .ZN(n12738) );
  NAND2_X1 U15940 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19142), .ZN(n19139) );
  AOI22_X1 U15941 ( .A1(n19146), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19127), .ZN(n12739) );
  INV_X1 U15942 ( .A(n12739), .ZN(n12740) );
  AOI211_X1 U15943 ( .C1(n15278), .C2(n19098), .A(n12741), .B(n12740), .ZN(
        n12747) );
  XNOR2_X1 U15944 ( .A(n12743), .B(n12742), .ZN(n15124) );
  INV_X1 U15945 ( .A(n15124), .ZN(n12745) );
  NAND2_X1 U15946 ( .A1(n12749), .A2(n12748), .ZN(P2_U2825) );
  NAND2_X1 U15947 ( .A1(n12750), .A2(n12768), .ZN(n12756) );
  NAND2_X1 U15948 ( .A1(n10184), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12751) );
  NOR2_X1 U15949 ( .A1(n12752), .A2(n19957), .ZN(n19719) );
  INV_X1 U15950 ( .A(n19833), .ZN(n12754) );
  INV_X1 U15951 ( .A(n19537), .ZN(n16367) );
  OAI21_X1 U15952 ( .B1(n16367), .B2(n19957), .A(n12752), .ZN(n12753) );
  AND3_X1 U15953 ( .A1(n12754), .A2(n19938), .A3(n12753), .ZN(n19683) );
  AOI21_X1 U15954 ( .B1(n12770), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19683), .ZN(n12755) );
  NOR2_X1 U15955 ( .A1(n13031), .A2(n12758), .ZN(n12759) );
  NAND2_X1 U15956 ( .A1(n12779), .A2(n12759), .ZN(n13736) );
  NAND2_X1 U15957 ( .A1(n12770), .A2(n15516), .ZN(n12762) );
  NAND2_X1 U15958 ( .A1(n10498), .A2(n19973), .ZN(n19684) );
  INV_X1 U15959 ( .A(n19684), .ZN(n12761) );
  NOR2_X1 U15960 ( .A1(n19537), .A2(n12761), .ZN(n19463) );
  NAND2_X1 U15961 ( .A1(n19463), .A2(n19938), .ZN(n19632) );
  NAND2_X1 U15962 ( .A1(n12762), .A2(n19632), .ZN(n12763) );
  INV_X1 U15963 ( .A(n12768), .ZN(n13088) );
  AOI22_X1 U15964 ( .A1(n12770), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19938), .B2(n19973), .ZN(n12764) );
  NAND2_X1 U15965 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12765) );
  NAND2_X1 U15966 ( .A1(n13861), .A2(n13860), .ZN(n12767) );
  INV_X1 U15967 ( .A(n13597), .ZN(n14173) );
  NAND2_X1 U15968 ( .A1(n14173), .A2(n12765), .ZN(n12766) );
  NAND2_X1 U15969 ( .A1(n12767), .A2(n12766), .ZN(n13755) );
  NAND2_X1 U15970 ( .A1(n12769), .A2(n12768), .ZN(n12772) );
  XNOR2_X1 U15971 ( .A(n19537), .B(n19957), .ZN(n19464) );
  AOI22_X1 U15972 ( .A1(n12770), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19938), .B2(n19464), .ZN(n12771) );
  NAND2_X1 U15973 ( .A1(n12772), .A2(n12771), .ZN(n12775) );
  NOR2_X1 U15974 ( .A1(n13031), .A2(n12773), .ZN(n12774) );
  OR2_X1 U15975 ( .A1(n12775), .A2(n12774), .ZN(n12776) );
  NAND2_X1 U15976 ( .A1(n12777), .A2(n12776), .ZN(n13757) );
  OR2_X2 U15977 ( .A1(n13755), .A2(n13757), .ZN(n12778) );
  NAND2_X1 U15978 ( .A1(n13691), .A2(n13692), .ZN(n13693) );
  NOR2_X1 U15979 ( .A1(n13031), .A2(n12780), .ZN(n13734) );
  NAND2_X1 U15980 ( .A1(n13896), .A2(n13987), .ZN(n12781) );
  AND2_X1 U15981 ( .A1(n14084), .A2(n14086), .ZN(n12783) );
  INV_X1 U15982 ( .A(n12930), .ZN(n12871) );
  INV_X1 U15983 ( .A(n12929), .ZN(n12870) );
  OAI22_X1 U15984 ( .A1(n19501), .A2(n12871), .B1(n12870), .B2(n12784), .ZN(
        n12785) );
  AOI21_X1 U15985 ( .B1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12913), .A(
        n12785), .ZN(n12787) );
  AOI22_X1 U15986 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12924), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12786) );
  OAI211_X1 U15987 ( .C1(n12788), .C2(n11087), .A(n12787), .B(n12786), .ZN(
        n12796) );
  AOI22_X1 U15988 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12914), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15989 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12912), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U15990 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U15991 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12789) );
  NAND4_X1 U15992 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n12795) );
  OAI22_X1 U15993 ( .A1(n12793), .A2(n13779), .B1(n12882), .B2(n19756), .ZN(
        n12794) );
  NOR3_X1 U15994 ( .A1(n12796), .A2(n12795), .A3(n12794), .ZN(n14278) );
  AOI22_X1 U15995 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12914), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U15996 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12911), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U15997 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U15998 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12797) );
  NAND4_X1 U15999 ( .A1(n12800), .A2(n12799), .A3(n12798), .A4(n12797), .ZN(
        n12810) );
  AOI22_X1 U16000 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12808) );
  NAND2_X1 U16001 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12802) );
  NAND2_X1 U16002 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12801) );
  OAI211_X1 U16003 ( .C1(n11087), .C2(n12803), .A(n12802), .B(n12801), .ZN(
        n12804) );
  INV_X1 U16004 ( .A(n12804), .ZN(n12807) );
  AOI22_X1 U16005 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U16006 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12805) );
  NAND4_X1 U16007 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n12809) );
  OR2_X1 U16008 ( .A1(n12810), .A2(n12809), .ZN(n14194) );
  AOI22_X1 U16009 ( .A1(n12914), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16010 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16011 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U16012 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12811) );
  NAND4_X1 U16013 ( .A1(n12814), .A2(n12813), .A3(n12812), .A4(n12811), .ZN(
        n12824) );
  AOI22_X1 U16014 ( .A1(n12921), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12922), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12822) );
  NAND2_X1 U16015 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12816) );
  NAND2_X1 U16016 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12815) );
  OAI211_X1 U16017 ( .C1(n11087), .C2(n12817), .A(n12816), .B(n12815), .ZN(
        n12818) );
  INV_X1 U16018 ( .A(n12818), .ZN(n12821) );
  AOI22_X1 U16019 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U16020 ( .A1(n12913), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12819) );
  NAND4_X1 U16021 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n12823) );
  NOR2_X1 U16022 ( .A1(n12824), .A2(n12823), .ZN(n14207) );
  INV_X1 U16023 ( .A(n14207), .ZN(n14191) );
  NAND2_X1 U16024 ( .A1(n14194), .A2(n14191), .ZN(n12825) );
  INV_X1 U16025 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12993) );
  INV_X1 U16026 ( .A(n12923), .ZN(n12856) );
  INV_X1 U16027 ( .A(n12924), .ZN(n12855) );
  INV_X1 U16028 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12827) );
  OAI22_X1 U16029 ( .A1(n12993), .A2(n12856), .B1(n12855), .B2(n12827), .ZN(
        n12831) );
  INV_X1 U16030 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12829) );
  INV_X1 U16031 ( .A(n12913), .ZN(n12859) );
  AOI22_X1 U16032 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12828) );
  OAI21_X1 U16033 ( .B1(n12829), .B2(n12859), .A(n12828), .ZN(n12830) );
  AOI211_X1 U16034 ( .C1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .C2(n10458), .A(
        n12831), .B(n12830), .ZN(n12838) );
  AOI22_X1 U16035 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U16036 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12914), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16037 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12911), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16038 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U16039 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12832) );
  AND4_X1 U16040 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12836) );
  NAND3_X1 U16041 ( .A1(n12838), .A2(n12837), .A3(n12836), .ZN(n15037) );
  OAI22_X1 U16042 ( .A1(n12840), .A2(n12871), .B1(n12870), .B2(n12839), .ZN(
        n12841) );
  AOI21_X1 U16043 ( .B1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12913), .A(
        n12841), .ZN(n12843) );
  AOI22_X1 U16044 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12924), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12842) );
  OAI211_X1 U16045 ( .C1(n12844), .C2(n11087), .A(n12843), .B(n12842), .ZN(
        n12853) );
  AOI22_X1 U16046 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12914), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U16047 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12912), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U16048 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U16049 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12845) );
  NAND4_X1 U16050 ( .A1(n12848), .A2(n12847), .A3(n12846), .A4(n12845), .ZN(
        n12852) );
  OAI22_X1 U16051 ( .A1(n12850), .A2(n13779), .B1(n12882), .B2(n12849), .ZN(
        n12851) );
  NOR3_X1 U16052 ( .A1(n12853), .A2(n12852), .A3(n12851), .ZN(n15028) );
  OAI22_X1 U16053 ( .A1(n12856), .A2(n13038), .B1(n12855), .B2(n12854), .ZN(
        n12861) );
  AOI22_X1 U16054 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12857) );
  OAI21_X1 U16055 ( .B1(n12859), .B2(n12858), .A(n12857), .ZN(n12860) );
  AOI211_X1 U16056 ( .C1(n10458), .C2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n12861), .B(n12860), .ZN(n12868) );
  AOI22_X1 U16057 ( .A1(n12921), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12922), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U16058 ( .A1(n12914), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U16059 ( .A1(n12911), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12912), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16060 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U16061 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12862) );
  AND4_X1 U16062 ( .A1(n12865), .A2(n12864), .A3(n12863), .A4(n12862), .ZN(
        n12866) );
  NAND3_X1 U16063 ( .A1(n12868), .A2(n12867), .A3(n12866), .ZN(n15023) );
  NAND2_X1 U16064 ( .A1(n15022), .A2(n15023), .ZN(n15015) );
  OAI22_X1 U16065 ( .A1(n12872), .A2(n12871), .B1(n12870), .B2(n12869), .ZN(
        n12873) );
  AOI21_X1 U16066 ( .B1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12913), .A(
        n12873), .ZN(n12875) );
  AOI22_X1 U16067 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12924), .B1(
        n12923), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12874) );
  OAI211_X1 U16068 ( .C1(n12876), .C2(n11087), .A(n12875), .B(n12874), .ZN(
        n12886) );
  AOI22_X1 U16069 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12914), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U16070 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12912), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16071 ( .A1(n12916), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12931), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U16072 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12910), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12877) );
  NAND4_X1 U16073 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n12885) );
  OAI22_X1 U16074 ( .A1(n12883), .A2(n13779), .B1(n12882), .B2(n12881), .ZN(
        n12884) );
  NOR3_X1 U16075 ( .A1(n12886), .A2(n12885), .A3(n12884), .ZN(n15018) );
  AOI22_X1 U16076 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16077 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13419), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12898) );
  INV_X1 U16078 ( .A(n12888), .ZN(n13432) );
  AOI22_X1 U16079 ( .A1(n13432), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12897) );
  INV_X1 U16080 ( .A(n10339), .ZN(n15514) );
  NAND2_X1 U16081 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12894) );
  INV_X1 U16082 ( .A(n12890), .ZN(n12893) );
  INV_X1 U16083 ( .A(n12891), .ZN(n12892) );
  AND2_X1 U16084 ( .A1(n12893), .A2(n12892), .ZN(n13060) );
  OAI211_X1 U16085 ( .C1(n15514), .C2(n14023), .A(n12894), .B(n13060), .ZN(
        n12895) );
  INV_X1 U16086 ( .A(n12895), .ZN(n12896) );
  NAND4_X1 U16087 ( .A1(n12899), .A2(n12898), .A3(n12897), .A4(n12896), .ZN(
        n12908) );
  AOI22_X1 U16088 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U16089 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16090 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12904) );
  INV_X1 U16091 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12901) );
  NAND2_X1 U16092 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12900) );
  INV_X1 U16093 ( .A(n13060), .ZN(n13425) );
  OAI211_X1 U16094 ( .C1(n15514), .C2(n12901), .A(n12900), .B(n13425), .ZN(
        n12902) );
  INV_X1 U16095 ( .A(n12902), .ZN(n12903) );
  NAND4_X1 U16096 ( .A1(n12906), .A2(n12905), .A3(n12904), .A4(n12903), .ZN(
        n12907) );
  AND2_X1 U16097 ( .A1(n12908), .A2(n12907), .ZN(n12960) );
  NAND2_X1 U16098 ( .A1(n19997), .A2(n12960), .ZN(n12938) );
  AOI22_X1 U16099 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12910), .B1(
        n12909), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16100 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12912), .B1(
        n12911), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16101 ( .A1(n12914), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12913), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16102 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12916), .B1(
        n12915), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12917) );
  NAND4_X1 U16103 ( .A1(n12920), .A2(n12919), .A3(n12918), .A4(n12917), .ZN(
        n12937) );
  AOI22_X1 U16104 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12922), .B1(
        n12921), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U16105 ( .A1(n12923), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12926) );
  NAND2_X1 U16106 ( .A1(n12924), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12925) );
  OAI211_X1 U16107 ( .C1(n11087), .C2(n12927), .A(n12926), .B(n12925), .ZN(
        n12928) );
  INV_X1 U16108 ( .A(n12928), .ZN(n12934) );
  AOI22_X1 U16109 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12930), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12933) );
  NAND2_X1 U16110 ( .A1(n12931), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12932) );
  NAND4_X1 U16111 ( .A1(n12935), .A2(n12934), .A3(n12933), .A4(n12932), .ZN(
        n12936) );
  OR2_X1 U16112 ( .A1(n12937), .A2(n12936), .ZN(n12957) );
  XNOR2_X1 U16113 ( .A(n12938), .B(n12957), .ZN(n12963) );
  NAND2_X1 U16114 ( .A1(n19348), .A2(n12960), .ZN(n15008) );
  AOI22_X1 U16116 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16117 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U16118 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U16119 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12941) );
  OAI211_X1 U16120 ( .C1(n15514), .C2(n12942), .A(n12941), .B(n13425), .ZN(
        n12943) );
  INV_X1 U16121 ( .A(n12943), .ZN(n12944) );
  NAND4_X1 U16122 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        n12956) );
  AOI22_X1 U16123 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U16124 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U16125 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12952) );
  NAND2_X1 U16126 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12948) );
  OAI211_X1 U16127 ( .C1(n15514), .C2(n12949), .A(n12948), .B(n13060), .ZN(
        n12950) );
  INV_X1 U16128 ( .A(n12950), .ZN(n12951) );
  NAND4_X1 U16129 ( .A1(n12954), .A2(n12953), .A3(n12952), .A4(n12951), .ZN(
        n12955) );
  NAND2_X1 U16130 ( .A1(n12956), .A2(n12955), .ZN(n12964) );
  NAND2_X1 U16131 ( .A1(n12957), .A2(n12960), .ZN(n12965) );
  XOR2_X1 U16132 ( .A(n12964), .B(n12965), .Z(n12958) );
  NAND2_X1 U16133 ( .A1(n12958), .A2(n12983), .ZN(n15002) );
  INV_X1 U16134 ( .A(n12964), .ZN(n12959) );
  NAND2_X1 U16135 ( .A1(n19348), .A2(n12959), .ZN(n15003) );
  INV_X1 U16136 ( .A(n12960), .ZN(n12961) );
  NOR2_X1 U16137 ( .A1(n15003), .A2(n12961), .ZN(n12962) );
  NOR2_X2 U16138 ( .A1(n15001), .A2(n10093), .ZN(n12988) );
  NOR2_X1 U16139 ( .A1(n12965), .A2(n12964), .ZN(n12984) );
  AOI22_X1 U16140 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16141 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16142 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12970) );
  INV_X1 U16143 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U16144 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12966) );
  OAI211_X1 U16145 ( .C1(n15514), .C2(n12967), .A(n12966), .B(n13425), .ZN(
        n12968) );
  INV_X1 U16146 ( .A(n12968), .ZN(n12969) );
  NAND4_X1 U16147 ( .A1(n12972), .A2(n12971), .A3(n12970), .A4(n12969), .ZN(
        n12982) );
  AOI22_X1 U16148 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U16149 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16150 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12978) );
  NAND2_X1 U16151 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12974) );
  OAI211_X1 U16152 ( .C1(n15514), .C2(n12975), .A(n12974), .B(n13060), .ZN(
        n12976) );
  INV_X1 U16153 ( .A(n12976), .ZN(n12977) );
  NAND4_X1 U16154 ( .A1(n12980), .A2(n12979), .A3(n12978), .A4(n12977), .ZN(
        n12981) );
  AND2_X1 U16155 ( .A1(n12982), .A2(n12981), .ZN(n12986) );
  NAND2_X1 U16156 ( .A1(n12984), .A2(n12986), .ZN(n13009) );
  OAI211_X1 U16157 ( .C1(n12984), .C2(n12986), .A(n13009), .B(n12983), .ZN(
        n12989) );
  INV_X1 U16158 ( .A(n12989), .ZN(n12985) );
  XNOR2_X1 U16159 ( .A(n12988), .B(n12985), .ZN(n14993) );
  INV_X1 U16160 ( .A(n12986), .ZN(n12987) );
  NOR2_X1 U16161 ( .A1(n19997), .A2(n12987), .ZN(n14995) );
  NAND2_X1 U16162 ( .A1(n14993), .A2(n14995), .ZN(n14994) );
  AOI22_X1 U16164 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16165 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16166 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U16167 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12992) );
  OAI211_X1 U16168 ( .C1(n15514), .C2(n12993), .A(n12992), .B(n13425), .ZN(
        n12994) );
  INV_X1 U16169 ( .A(n12994), .ZN(n12995) );
  NAND4_X1 U16170 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n13008) );
  AOI22_X1 U16171 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16172 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U16173 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13004) );
  NAND2_X1 U16174 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13000) );
  OAI211_X1 U16175 ( .C1(n15514), .C2(n13001), .A(n13000), .B(n13060), .ZN(
        n13002) );
  INV_X1 U16176 ( .A(n13002), .ZN(n13003) );
  NAND4_X1 U16177 ( .A1(n13006), .A2(n13005), .A3(n13004), .A4(n13003), .ZN(
        n13007) );
  NAND2_X1 U16178 ( .A1(n13008), .A2(n13007), .ZN(n13011) );
  AOI21_X1 U16179 ( .B1(n13009), .B2(n13011), .A(n13031), .ZN(n13010) );
  NAND2_X1 U16180 ( .A1(n13010), .A2(n13032), .ZN(n13013) );
  NOR2_X1 U16181 ( .A1(n19997), .A2(n13011), .ZN(n14985) );
  NAND2_X1 U16182 ( .A1(n14983), .A2(n14985), .ZN(n14984) );
  INV_X1 U16183 ( .A(n13012), .ZN(n13014) );
  NAND2_X1 U16184 ( .A1(n14984), .A2(n10065), .ZN(n13034) );
  AOI22_X1 U16185 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16186 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U16187 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13019) );
  INV_X1 U16188 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U16189 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13015) );
  OAI211_X1 U16190 ( .C1(n15514), .C2(n13016), .A(n13015), .B(n13425), .ZN(
        n13017) );
  INV_X1 U16191 ( .A(n13017), .ZN(n13018) );
  NAND4_X1 U16192 ( .A1(n13021), .A2(n13020), .A3(n13019), .A4(n13018), .ZN(
        n13030) );
  AOI22_X1 U16193 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U16194 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U16195 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U16196 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13022) );
  OAI211_X1 U16197 ( .C1(n15514), .C2(n13023), .A(n13022), .B(n13060), .ZN(
        n13024) );
  INV_X1 U16198 ( .A(n13024), .ZN(n13025) );
  NAND4_X1 U16199 ( .A1(n13028), .A2(n13027), .A3(n13026), .A4(n13025), .ZN(
        n13029) );
  NAND2_X1 U16200 ( .A1(n13030), .A2(n13029), .ZN(n13035) );
  NOR2_X1 U16201 ( .A1(n13032), .A2(n13035), .ZN(n13052) );
  AOI211_X1 U16202 ( .C1(n13035), .C2(n13032), .A(n13031), .B(n13052), .ZN(
        n13033) );
  INV_X1 U16203 ( .A(n13035), .ZN(n13036) );
  NAND2_X1 U16204 ( .A1(n19348), .A2(n13036), .ZN(n14975) );
  AOI22_X1 U16205 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16206 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16207 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U16208 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13037) );
  OAI211_X1 U16209 ( .C1(n15514), .C2(n13038), .A(n13037), .B(n13425), .ZN(
        n13039) );
  INV_X1 U16210 ( .A(n13039), .ZN(n13040) );
  NAND4_X1 U16211 ( .A1(n13043), .A2(n13042), .A3(n13041), .A4(n13040), .ZN(
        n13051) );
  AOI22_X1 U16212 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U16213 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U16214 ( .A1(n13431), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13047) );
  NAND2_X1 U16215 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13044) );
  OAI211_X1 U16216 ( .C1(n15514), .C2(n14032), .A(n13044), .B(n13060), .ZN(
        n13045) );
  INV_X1 U16217 ( .A(n13045), .ZN(n13046) );
  NAND4_X1 U16218 ( .A1(n13049), .A2(n13048), .A3(n13047), .A4(n13046), .ZN(
        n13050) );
  AND2_X1 U16219 ( .A1(n13051), .A2(n13050), .ZN(n14967) );
  INV_X1 U16220 ( .A(n13052), .ZN(n14965) );
  NAND2_X1 U16221 ( .A1(n19997), .A2(n14967), .ZN(n13053) );
  NOR2_X1 U16222 ( .A1(n14965), .A2(n13053), .ZN(n13071) );
  AOI22_X1 U16223 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16224 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16225 ( .A1(n12991), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13057) );
  NAND2_X1 U16226 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13054) );
  OAI211_X1 U16227 ( .C1(n10545), .C2(n15514), .A(n13054), .B(n13425), .ZN(
        n13055) );
  INV_X1 U16228 ( .A(n13055), .ZN(n13056) );
  NAND4_X1 U16229 ( .A1(n13059), .A2(n13058), .A3(n13057), .A4(n13056), .ZN(
        n13069) );
  AOI22_X1 U16230 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U16231 ( .A1(n12991), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16232 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U16233 ( .A1(n9636), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13061) );
  OAI211_X1 U16234 ( .C1(n15514), .C2(n13062), .A(n13061), .B(n13060), .ZN(
        n13063) );
  INV_X1 U16235 ( .A(n13063), .ZN(n13064) );
  NAND4_X1 U16236 ( .A1(n13067), .A2(n13066), .A3(n13065), .A4(n13064), .ZN(
        n13068) );
  AND2_X1 U16237 ( .A1(n13069), .A2(n13068), .ZN(n13070) );
  NAND2_X1 U16238 ( .A1(n13071), .A2(n13070), .ZN(n13416) );
  OAI21_X1 U16239 ( .B1(n13071), .B2(n13070), .A(n13416), .ZN(n13072) );
  INV_X1 U16240 ( .A(n13418), .ZN(n13076) );
  NAND2_X1 U16241 ( .A1(n13073), .A2(n13072), .ZN(n14348) );
  OR2_X1 U16242 ( .A1(n16389), .A2(n13777), .ZN(n13768) );
  INV_X1 U16243 ( .A(n11209), .ZN(n13074) );
  NAND2_X1 U16244 ( .A1(n13768), .A2(n13074), .ZN(n13075) );
  NAND2_X1 U16245 ( .A1(n15036), .A2(n15558), .ZN(n15044) );
  NAND2_X1 U16246 ( .A1(n15042), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13077) );
  INV_X1 U16247 ( .A(n19843), .ZN(n13775) );
  NOR2_X1 U16248 ( .A1(n16384), .A2(n13775), .ZN(n13081) );
  OR2_X1 U16249 ( .A1(n13515), .A2(n19997), .ZN(n19323) );
  INV_X1 U16250 ( .A(n13515), .ZN(n13084) );
  NAND2_X1 U16251 ( .A1(n15803), .A2(n19950), .ZN(n15697) );
  INV_X1 U16252 ( .A(n15697), .ZN(n19940) );
  OR2_X1 U16253 ( .A1(n19938), .A2(n19940), .ZN(n19969) );
  NAND2_X1 U16254 ( .A1(n19969), .A2(n13085), .ZN(n13086) );
  NAND2_X2 U16255 ( .A1(n13515), .A2(n13086), .ZN(n19312) );
  NAND2_X1 U16256 ( .A1(n18922), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13087) );
  NAND2_X1 U16257 ( .A1(n13088), .A2(n13087), .ZN(n19314) );
  AND2_X1 U16258 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19958) );
  INV_X1 U16259 ( .A(n19312), .ZN(n19313) );
  AOI21_X1 U16260 ( .B1(n19313), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n13089), .ZN(n13090) );
  OAI21_X1 U16261 ( .B1(n16125), .B2(n19305), .A(n13090), .ZN(n13091) );
  NAND2_X2 U16262 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18865), .ZN(
        n13104) );
  AOI22_X1 U16263 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13097) );
  OAI21_X1 U16264 ( .B1(n17058), .B2(n21086), .A(n13097), .ZN(n13114) );
  INV_X1 U16265 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16979) );
  OR3_X2 U16266 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n13103), .ZN(n13131) );
  AOI22_X1 U16267 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13112) );
  NOR4_X2 U16268 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n18879), .ZN(n13138) );
  INV_X1 U16269 ( .A(n13138), .ZN(n13098) );
  INV_X1 U16270 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13102) );
  NOR2_X4 U16271 ( .A1(n18856), .A2(n13100), .ZN(n16984) );
  AOI22_X1 U16272 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13101) );
  OAI21_X1 U16273 ( .B1(n17229), .B2(n13102), .A(n13101), .ZN(n13110) );
  INV_X1 U16274 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17274) );
  NOR2_X2 U16275 ( .A1(n13105), .A2(n13104), .ZN(n17251) );
  AOI22_X1 U16276 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13108) );
  INV_X4 U16277 ( .A(n16912), .ZN(n17254) );
  AOI22_X1 U16278 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13107) );
  OAI211_X1 U16279 ( .C1(n17250), .C2(n17274), .A(n13108), .B(n13107), .ZN(
        n13109) );
  AOI211_X1 U16280 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n13110), .B(n13109), .ZN(n13111) );
  OAI211_X1 U16281 ( .C1(n13126), .C2(n16979), .A(n13112), .B(n13111), .ZN(
        n13113) );
  INV_X1 U16282 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U16283 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13115) );
  OAI21_X1 U16284 ( .B1(n17199), .B2(n17174), .A(n13115), .ZN(n13125) );
  INV_X1 U16285 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15608) );
  AOI22_X1 U16286 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13123) );
  INV_X1 U16287 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16288 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U16289 ( .B1(n17229), .B2(n13117), .A(n13116), .ZN(n13121) );
  INV_X1 U16290 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U16291 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16292 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13118) );
  OAI211_X1 U16293 ( .C1(n17250), .C2(n17280), .A(n13119), .B(n13118), .ZN(
        n13120) );
  AOI211_X1 U16294 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n13121), .B(n13120), .ZN(n13122) );
  OAI211_X1 U16295 ( .C1(n17226), .C2(n15608), .A(n13123), .B(n13122), .ZN(
        n13124) );
  INV_X1 U16296 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U16297 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16298 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13127) );
  OAI211_X1 U16299 ( .C1(n9629), .C2(n17239), .A(n13128), .B(n13127), .ZN(
        n13129) );
  AOI22_X1 U16300 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13137) );
  INV_X2 U16301 ( .A(n17229), .ZN(n13171) );
  AOI22_X1 U16302 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13195), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U16303 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U16304 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13133) );
  NAND2_X1 U16305 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13132) );
  INV_X1 U16306 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U16307 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13138), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13139) );
  OAI21_X1 U16308 ( .B1(n17250), .B2(n17289), .A(n13139), .ZN(n13145) );
  INV_X1 U16309 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n21126) );
  AOI22_X1 U16310 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13140), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13143) );
  AOI22_X1 U16311 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13142) );
  OAI211_X1 U16312 ( .C1(n17229), .C2(n21126), .A(n13143), .B(n13142), .ZN(
        n13144) );
  AOI211_X1 U16313 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n13145), .B(n13144), .ZN(n13154) );
  AOI22_X1 U16314 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13146) );
  INV_X1 U16315 ( .A(n13146), .ZN(n13149) );
  INV_X1 U16316 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U16317 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13150) );
  OAI21_X1 U16318 ( .B1(n17058), .B2(n17218), .A(n13150), .ZN(n13151) );
  INV_X1 U16319 ( .A(n13151), .ZN(n13152) );
  INV_X1 U16320 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U16321 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13167) );
  INV_X1 U16322 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U16323 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16324 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13157) );
  OAI211_X1 U16325 ( .C1(n17250), .C2(n17283), .A(n13158), .B(n13157), .ZN(
        n13165) );
  AOI22_X1 U16326 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U16327 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U16328 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13171), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13161) );
  INV_X1 U16329 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13159) );
  NAND4_X1 U16330 ( .A1(n13163), .A2(n13162), .A3(n13161), .A4(n13160), .ZN(
        n13164) );
  NAND2_X1 U16331 ( .A1(n13208), .A2(n17432), .ZN(n13212) );
  INV_X1 U16332 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16333 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U16334 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13196), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U16335 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13169) );
  OAI211_X1 U16336 ( .C1(n17250), .C2(n17277), .A(n13170), .B(n13169), .ZN(
        n13177) );
  AOI22_X1 U16337 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16338 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U16339 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U16340 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13172) );
  NAND4_X1 U16341 ( .A1(n13175), .A2(n13174), .A3(n13173), .A4(n13172), .ZN(
        n13176) );
  AOI211_X1 U16342 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n13177), .B(n13176), .ZN(n13178) );
  INV_X1 U16343 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21077) );
  AOI22_X1 U16344 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13190) );
  INV_X1 U16345 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U16346 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U16347 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13181) );
  OAI211_X1 U16348 ( .C1(n17250), .C2(n17270), .A(n13182), .B(n13181), .ZN(
        n13188) );
  AOI22_X1 U16349 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13196), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13186) );
  AOI22_X1 U16350 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U16351 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13184) );
  NAND2_X1 U16352 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13183) );
  NAND4_X1 U16353 ( .A1(n13186), .A2(n13185), .A3(n13184), .A4(n13183), .ZN(
        n13187) );
  AOI211_X1 U16354 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n13188), .B(n13187), .ZN(n13189) );
  OAI211_X1 U16355 ( .C1(n21077), .C2(n15640), .A(n13190), .B(n13189), .ZN(
        n16464) );
  NAND2_X1 U16356 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17937) );
  INV_X1 U16357 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18154) );
  XNOR2_X1 U16358 ( .A(n13192), .B(n17422), .ZN(n17869) );
  INV_X1 U16359 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18227) );
  NOR2_X1 U16360 ( .A1(n18227), .A2(n13193), .ZN(n13207) );
  INV_X1 U16361 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18861) );
  NOR2_X1 U16362 ( .A1(n13363), .A2(n18861), .ZN(n13206) );
  AOI22_X1 U16363 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16364 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U16365 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13195), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13197) );
  OAI211_X1 U16366 ( .C1(n17250), .C2(n17119), .A(n13198), .B(n13197), .ZN(
        n13204) );
  AOI22_X1 U16367 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13202) );
  AOI22_X1 U16368 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13201) );
  AOI22_X1 U16369 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13200) );
  NAND2_X1 U16370 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13199) );
  NAND4_X1 U16371 ( .A1(n13202), .A2(n13201), .A3(n13200), .A4(n13199), .ZN(
        n13203) );
  NOR2_X1 U16372 ( .A1(n13206), .A2(n17917), .ZN(n17906) );
  XOR2_X1 U16373 ( .A(n13208), .B(n17432), .Z(n13209) );
  XNOR2_X1 U16374 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13209), .ZN(
        n17897) );
  NOR2_X1 U16375 ( .A1(n17898), .A2(n17897), .ZN(n17896) );
  INV_X1 U16376 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18202) );
  NAND2_X1 U16377 ( .A1(n13211), .A2(n18202), .ZN(n13213) );
  XNOR2_X1 U16378 ( .A(n13212), .B(n17428), .ZN(n17883) );
  XNOR2_X1 U16379 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13214), .ZN(
        n17859) );
  OAI21_X1 U16380 ( .B1(n16466), .B2(n16464), .A(n17834), .ZN(n13216) );
  INV_X1 U16381 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18160) );
  INV_X1 U16382 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18086) );
  INV_X1 U16383 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17814) );
  NOR2_X1 U16384 ( .A1(n18148), .A2(n17814), .ZN(n18123) );
  NAND2_X1 U16385 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18123), .ZN(
        n18096) );
  INV_X1 U16386 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17779) );
  NOR3_X1 U16387 ( .A1(n18086), .A2(n18096), .A3(n17779), .ZN(n17747) );
  NAND2_X1 U16388 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17747), .ZN(
        n13393) );
  INV_X1 U16389 ( .A(n13393), .ZN(n18057) );
  NAND2_X1 U16390 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18057), .ZN(
        n18045) );
  INV_X1 U16391 ( .A(n18045), .ZN(n17992) );
  NAND2_X1 U16392 ( .A1(n13354), .A2(n17992), .ZN(n13221) );
  NAND2_X1 U16393 ( .A1(n13221), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13220) );
  INV_X1 U16394 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18059) );
  NOR3_X1 U16395 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17746) );
  NOR2_X1 U16396 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17757) );
  INV_X1 U16397 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18072) );
  NAND4_X1 U16398 ( .A1(n17746), .A2(n17757), .A3(n18086), .A4(n18072), .ZN(
        n13218) );
  OAI21_X1 U16399 ( .B1(n17744), .B2(n13218), .A(n17834), .ZN(n13222) );
  INV_X1 U16400 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21117) );
  NAND2_X1 U16401 ( .A1(n13222), .A2(n13221), .ZN(n17727) );
  NAND2_X1 U16402 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17712) );
  INV_X1 U16403 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21089) );
  INV_X1 U16404 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17664) );
  NAND2_X1 U16405 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17672) );
  NOR3_X1 U16406 ( .A1(n21089), .A2(n17664), .A3(n17672), .ZN(n18002) );
  NAND2_X1 U16407 ( .A1(n18002), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17974) );
  NOR2_X1 U16408 ( .A1(n17712), .A2(n17974), .ZN(n17993) );
  INV_X1 U16409 ( .A(n17993), .ZN(n13356) );
  INV_X1 U16410 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17986) );
  NOR2_X1 U16411 ( .A1(n13356), .A2(n17986), .ZN(n17623) );
  NAND2_X1 U16412 ( .A1(n17727), .A2(n17623), .ZN(n13224) );
  INV_X1 U16413 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18028) );
  NAND2_X1 U16414 ( .A1(n17709), .A2(n18028), .ZN(n13223) );
  NOR2_X1 U16415 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13223), .ZN(
        n17663) );
  NAND2_X1 U16416 ( .A1(n17663), .A2(n17664), .ZN(n17655) );
  NOR2_X2 U16417 ( .A1(n17616), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17615) );
  INV_X1 U16418 ( .A(n17974), .ZN(n17958) );
  INV_X1 U16419 ( .A(n17712), .ZN(n18039) );
  NAND2_X1 U16420 ( .A1(n18039), .A2(n17727), .ZN(n17662) );
  NOR2_X1 U16421 ( .A1(n17607), .A2(n17834), .ZN(n13226) );
  INV_X1 U16422 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17949) );
  OR2_X1 U16423 ( .A1(n17745), .A2(n17615), .ZN(n17606) );
  INV_X1 U16424 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17944) );
  NOR3_X2 U16425 ( .A1(n17580), .A2(n17745), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15722) );
  INV_X1 U16426 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16425) );
  NAND2_X1 U16427 ( .A1(n15722), .A2(n16425), .ZN(n15784) );
  NAND2_X1 U16428 ( .A1(n17745), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16462) );
  INV_X1 U16429 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16444) );
  AOI21_X1 U16430 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n17834), .ZN(n13227) );
  NOR2_X1 U16431 ( .A1(n15783), .A2(n16444), .ZN(n13230) );
  NAND2_X1 U16432 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16444), .ZN(
        n16442) );
  OAI22_X1 U16433 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17834), .B1(
        n15784), .B2(n16442), .ZN(n13228) );
  NOR2_X1 U16434 ( .A1(n13230), .A2(n13229), .ZN(n13231) );
  AOI21_X1 U16435 ( .B1(n13232), .B2(n10068), .A(n13231), .ZN(n16452) );
  INV_X1 U16436 ( .A(n16464), .ZN(n17416) );
  OAI22_X1 U16437 ( .A1(n18865), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18255), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U16438 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18714), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18873), .ZN(n13344) );
  OAI21_X1 U16439 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18865), .A(
        n13234), .ZN(n13235) );
  OAI22_X1 U16440 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13235), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21095), .ZN(n13241) );
  NOR2_X1 U16441 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21095), .ZN(
        n13236) );
  NAND2_X1 U16442 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13235), .ZN(
        n13240) );
  AOI22_X1 U16443 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13241), .B1(
        n13236), .B2(n13240), .ZN(n13244) );
  AOI21_X1 U16444 ( .B1(n18879), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n13343), .ZN(n13347) );
  AND2_X1 U16445 ( .A1(n13344), .A2(n13347), .ZN(n13243) );
  OAI21_X1 U16446 ( .B1(n13239), .B2(n13238), .A(n13244), .ZN(n13237) );
  INV_X1 U16447 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14293) );
  AND2_X1 U16448 ( .A1(n13240), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13242) );
  OAI22_X1 U16449 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14293), .B1(
        n13242), .B2(n13241), .ZN(n13345) );
  AOI22_X1 U16450 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13245) );
  OAI21_X1 U16451 ( .B1(n13131), .B2(n17291), .A(n13245), .ZN(n13255) );
  AOI22_X1 U16452 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16453 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16454 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13246) );
  OAI22_X1 U16455 ( .A1(n17229), .A2(n17102), .B1(n9629), .B2(n17101), .ZN(
        n13252) );
  AOI22_X1 U16456 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13250) );
  NAND3_X1 U16457 ( .A1(n13250), .A2(n13249), .A3(n10080), .ZN(n13251) );
  AOI211_X4 U16458 ( .C1(n13196), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n13255), .B(n13254), .ZN(n18892) );
  AOI22_X1 U16459 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13256) );
  OAI21_X1 U16460 ( .B1(n13131), .B2(n17119), .A(n13256), .ZN(n13265) );
  AOI22_X1 U16461 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13263) );
  OAI21_X1 U16462 ( .B1(n17250), .B2(n21110), .A(n13257), .ZN(n13261) );
  INV_X1 U16463 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U16464 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13259) );
  AOI22_X1 U16465 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13258) );
  OAI211_X1 U16466 ( .C1(n17229), .C2(n17126), .A(n13259), .B(n13258), .ZN(
        n13260) );
  AOI211_X1 U16467 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n13261), .B(n13260), .ZN(n13262) );
  OAI211_X1 U16468 ( .C1(n17058), .C2(n17122), .A(n13263), .B(n13262), .ZN(
        n13264) );
  NAND2_X1 U16469 ( .A1(n18892), .A2(n18262), .ZN(n13335) );
  NAND2_X1 U16470 ( .A1(n13352), .A2(n13335), .ZN(n18912) );
  INV_X1 U16471 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17172) );
  AOI22_X1 U16472 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13266) );
  OAI21_X1 U16473 ( .B1(n17208), .B2(n17172), .A(n13266), .ZN(n13275) );
  INV_X1 U16474 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U16475 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13273) );
  INV_X1 U16476 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15601) );
  INV_X1 U16477 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17181) );
  OAI22_X1 U16478 ( .A1(n17264), .A2(n15601), .B1(n17250), .B2(n17181), .ZN(
        n13271) );
  AOI22_X1 U16479 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13269) );
  AOI22_X1 U16480 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U16481 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13267) );
  NAND3_X1 U16482 ( .A1(n13269), .A2(n13268), .A3(n13267), .ZN(n13270) );
  AOI211_X1 U16483 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n13271), .B(n13270), .ZN(n13272) );
  OAI211_X1 U16484 ( .C1(n17058), .C2(n17060), .A(n13273), .B(n13272), .ZN(
        n13274) );
  AOI22_X1 U16485 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13285) );
  INV_X1 U16486 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U16487 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U16488 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13276) );
  OAI211_X1 U16489 ( .C1(n17250), .C2(n17155), .A(n13277), .B(n13276), .ZN(
        n13283) );
  AOI22_X1 U16490 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16491 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U16492 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13279) );
  NAND2_X1 U16493 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13278) );
  NAND4_X1 U16494 ( .A1(n13281), .A2(n13280), .A3(n13279), .A4(n13278), .ZN(
        n13282) );
  AOI211_X1 U16495 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n13283), .B(n13282), .ZN(n13284) );
  AOI22_X1 U16496 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U16497 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U16498 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13293) );
  OAI22_X1 U16499 ( .A1(n13131), .A2(n17277), .B1(n17264), .B2(n21120), .ZN(
        n13291) );
  AOI22_X1 U16500 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U16501 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13288) );
  AOI22_X1 U16502 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13287) );
  NAND2_X1 U16503 ( .A1(n17236), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13286) );
  NAND4_X1 U16504 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13290) );
  AOI211_X1 U16505 ( .C1(n9635), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n13291), .B(n13290), .ZN(n13292) );
  NAND4_X1 U16506 ( .A1(n13295), .A2(n13294), .A3(n13293), .A4(n13292), .ZN(
        n17300) );
  NOR2_X1 U16507 ( .A1(n18289), .A2(n17300), .ZN(n13326) );
  AOI22_X1 U16508 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16509 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16510 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13303) );
  INV_X1 U16511 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20947) );
  OAI22_X1 U16512 ( .A1(n17264), .A2(n17218), .B1(n13156), .B2(n20947), .ZN(
        n13301) );
  AOI22_X1 U16513 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13299) );
  AOI22_X1 U16514 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13298) );
  AOI22_X1 U16515 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U16516 ( .A1(n17215), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13296) );
  NAND4_X1 U16517 ( .A1(n13299), .A2(n13298), .A3(n13297), .A4(n13296), .ZN(
        n13300) );
  INV_X1 U16518 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U16519 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U16520 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17230), .ZN(n13306) );
  OAI211_X1 U16521 ( .C1(n17250), .C2(n17137), .A(n13307), .B(n13306), .ZN(
        n13313) );
  AOI22_X1 U16522 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17254), .ZN(n13311) );
  AOI22_X1 U16523 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n13141), .ZN(n13310) );
  AOI22_X1 U16524 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17253), .ZN(n13309) );
  NAND2_X1 U16525 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n16984), .ZN(
        n13308) );
  NAND4_X1 U16526 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13312) );
  AOI22_X1 U16527 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U16528 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U16529 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13323) );
  INV_X1 U16530 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17198) );
  INV_X1 U16531 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n21072) );
  OAI22_X1 U16532 ( .A1(n17058), .A2(n17198), .B1(n17264), .B2(n21072), .ZN(
        n13321) );
  AOI22_X1 U16533 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U16534 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U16535 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U16536 ( .A1(n17236), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13316) );
  NAND4_X1 U16537 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13320) );
  NAND2_X1 U16538 ( .A1(n17340), .A2(n13337), .ZN(n13339) );
  NAND2_X1 U16539 ( .A1(n18700), .A2(n13353), .ZN(n14288) );
  NAND2_X1 U16540 ( .A1(n13326), .A2(n18699), .ZN(n15592) );
  NAND3_X2 U16541 ( .A1(n18285), .A2(n13353), .A3(n18262), .ZN(n17512) );
  INV_X1 U16542 ( .A(n13337), .ZN(n18277) );
  INV_X1 U16543 ( .A(n18281), .ZN(n15591) );
  INV_X1 U16544 ( .A(n13349), .ZN(n18273) );
  OAI211_X1 U16545 ( .C1(n18285), .C2(n15591), .A(n18273), .B(n13352), .ZN(
        n13328) );
  NAND2_X1 U16546 ( .A1(n18289), .A2(n17300), .ZN(n18708) );
  AOI21_X1 U16547 ( .B1(n17340), .B2(n18708), .A(n13335), .ZN(n14283) );
  AOI211_X1 U16548 ( .C1(n13337), .C2(n13336), .A(n14284), .B(n14283), .ZN(
        n13341) );
  INV_X1 U16549 ( .A(n13489), .ZN(n13340) );
  NAND3_X1 U16550 ( .A1(n18268), .A2(n13340), .A3(n13339), .ZN(n13342) );
  NAND2_X2 U16551 ( .A1(n18129), .A2(n17934), .ZN(n18156) );
  NOR2_X4 U16552 ( .A1(n18268), .A2(n18156), .ZN(n15702) );
  XOR2_X1 U16553 ( .A(n13344), .B(n13343), .Z(n13346) );
  AOI21_X1 U16554 ( .B1(n13346), .B2(n13348), .A(n13345), .ZN(n18695) );
  AOI21_X1 U16555 ( .B1(n13348), .B2(n13347), .A(n16576), .ZN(n18696) );
  NOR2_X1 U16556 ( .A1(n18892), .A2(n13349), .ZN(n15704) );
  NAND2_X1 U16557 ( .A1(n15704), .A2(n13350), .ZN(n15708) );
  NAND3_X1 U16558 ( .A1(n13353), .A2(n13352), .A3(n13351), .ZN(n14285) );
  NAND2_X1 U16559 ( .A1(n18859), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18754) );
  NOR2_X1 U16560 ( .A1(n18754), .A2(n18910), .ZN(n18902) );
  NOR2_X4 U16561 ( .A1(n16579), .A2(n18892), .ZN(n17920) );
  INV_X2 U16562 ( .A(n17920), .ZN(n17931) );
  NAND2_X1 U16563 ( .A1(n16452), .A2(n17829), .ZN(n13400) );
  INV_X1 U16564 ( .A(n17744), .ZN(n13355) );
  NAND2_X1 U16565 ( .A1(n18164), .A2(n17834), .ZN(n17833) );
  INV_X1 U16566 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17796) );
  NOR2_X1 U16567 ( .A1(n18096), .A2(n17796), .ZN(n18106) );
  NAND2_X1 U16568 ( .A1(n18106), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18067) );
  NAND2_X1 U16569 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17962) );
  OR2_X1 U16570 ( .A1(n17962), .A2(n17937), .ZN(n16460) );
  OR2_X1 U16571 ( .A1(n13356), .A2(n16460), .ZN(n15711) );
  NAND2_X1 U16572 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16436) );
  NOR2_X1 U16573 ( .A1(n16436), .A2(n16425), .ZN(n15782) );
  INV_X1 U16574 ( .A(n15782), .ZN(n16445) );
  NAND2_X1 U16575 ( .A1(n16437), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13357) );
  XNOR2_X1 U16576 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13357), .ZN(
        n16453) );
  NOR2_X4 U16577 ( .A1(n16464), .A2(n17931), .ZN(n17842) );
  NAND2_X1 U16578 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18251) );
  NAND2_X1 U16579 ( .A1(n18850), .A2(n18251), .ZN(n18901) );
  INV_X1 U16580 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18893) );
  NOR2_X1 U16581 ( .A1(n18859), .A2(n18893), .ZN(n17886) );
  NOR2_X4 U16582 ( .A1(n18859), .A2(n17868), .ZN(n17789) );
  NAND4_X1 U16583 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16773) );
  NAND2_X1 U16584 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17731) );
  NAND2_X1 U16585 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17695) );
  NAND2_X1 U16586 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17649) );
  NAND2_X1 U16587 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17611) );
  NAND2_X1 U16588 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17575) );
  NAND2_X1 U16589 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n13359), .ZN(
        n13360) );
  INV_X1 U16590 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17923) );
  NAND2_X1 U16591 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16426), .ZN(
        n13358) );
  XOR2_X2 U16592 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13358), .Z(
        n16884) );
  INV_X1 U16593 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18833) );
  NOR2_X1 U16594 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18911) );
  INV_X1 U16595 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18898) );
  NOR2_X1 U16596 ( .A1(n18833), .A2(n18229), .ZN(n16449) );
  NOR2_X1 U16597 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18910), .ZN(n17646) );
  NAND2_X1 U16598 ( .A1(n18859), .A2(n18910), .ZN(n18897) );
  AOI21_X1 U16599 ( .B1(n18251), .B2(n18897), .A(n18874), .ZN(n18261) );
  NOR3_X1 U16600 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18893), .ZN(n18604) );
  INV_X2 U16601 ( .A(n18363), .ZN(n18636) );
  OR2_X1 U16602 ( .A1(n13360), .A2(n17769), .ZN(n16415) );
  INV_X1 U16603 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16606) );
  XOR2_X1 U16604 ( .A(n16606), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n13361) );
  NOR2_X1 U16605 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17715), .ZN(
        n16428) );
  INV_X1 U16606 ( .A(n13359), .ZN(n16431) );
  NOR2_X1 U16607 ( .A1(n16431), .A2(n17923), .ZN(n16595) );
  INV_X1 U16608 ( .A(n17646), .ZN(n17928) );
  NAND2_X1 U16609 ( .A1(n18636), .A2(n13360), .ZN(n16432) );
  OAI211_X1 U16610 ( .C1(n16595), .C2(n17928), .A(n16432), .B(n17927), .ZN(
        n16435) );
  NOR2_X1 U16611 ( .A1(n16428), .A2(n16435), .ZN(n16414) );
  OAI22_X1 U16612 ( .A1(n16415), .A2(n13361), .B1(n16414), .B2(n16606), .ZN(
        n13362) );
  AOI211_X1 U16613 ( .C1(n17789), .C2(n13498), .A(n16449), .B(n13362), .ZN(
        n13397) );
  NAND2_X1 U16614 ( .A1(n13363), .A2(n17926), .ZN(n13366) );
  NAND2_X1 U16615 ( .A1(n10083), .A2(n13366), .ZN(n13365) );
  NAND2_X1 U16616 ( .A1(n17432), .A2(n13365), .ZN(n13375) );
  NOR2_X1 U16617 ( .A1(n17428), .A2(n13375), .ZN(n13364) );
  NAND2_X1 U16618 ( .A1(n13364), .A2(n17422), .ZN(n13381) );
  NOR2_X1 U16619 ( .A1(n17419), .A2(n13381), .ZN(n13385) );
  NAND2_X1 U16620 ( .A1(n13385), .A2(n16464), .ZN(n13386) );
  XOR2_X1 U16621 ( .A(n17422), .B(n13364), .Z(n13379) );
  INV_X1 U16622 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18192) );
  XNOR2_X1 U16623 ( .A(n17432), .B(n13365), .ZN(n13373) );
  NOR2_X1 U16624 ( .A1(n18192), .A2(n13373), .ZN(n13374) );
  XOR2_X1 U16625 ( .A(n10083), .B(n13366), .Z(n13367) );
  NOR2_X1 U16626 ( .A1(n13367), .A2(n18227), .ZN(n13372) );
  XNOR2_X1 U16627 ( .A(n18227), .B(n13367), .ZN(n17908) );
  INV_X1 U16628 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18876) );
  NOR2_X1 U16629 ( .A1(n17448), .A2(n18876), .ZN(n13370) );
  INV_X1 U16630 ( .A(n17926), .ZN(n13369) );
  NAND3_X1 U16631 ( .A1(n13369), .A2(n17448), .A3(n18876), .ZN(n13368) );
  OAI221_X1 U16632 ( .B1(n13370), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n13369), .C2(n17448), .A(n13368), .ZN(n17907) );
  NOR2_X1 U16633 ( .A1(n17908), .A2(n17907), .ZN(n13371) );
  NOR2_X1 U16634 ( .A1(n13372), .A2(n13371), .ZN(n17895) );
  XNOR2_X1 U16635 ( .A(n18192), .B(n13373), .ZN(n17894) );
  NOR2_X1 U16636 ( .A1(n17895), .A2(n17894), .ZN(n17893) );
  NOR2_X1 U16637 ( .A1(n13374), .A2(n17893), .ZN(n13376) );
  XNOR2_X1 U16638 ( .A(n17428), .B(n13375), .ZN(n13377) );
  NOR2_X1 U16639 ( .A1(n13376), .A2(n13377), .ZN(n13378) );
  XNOR2_X1 U16640 ( .A(n13377), .B(n13376), .ZN(n17881) );
  NOR2_X1 U16641 ( .A1(n18202), .A2(n17881), .ZN(n17880) );
  NOR2_X1 U16642 ( .A1(n13378), .A2(n17880), .ZN(n17874) );
  XNOR2_X1 U16643 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13379), .ZN(
        n17873) );
  XNOR2_X1 U16644 ( .A(n17419), .B(n13381), .ZN(n13383) );
  NOR2_X1 U16645 ( .A1(n13382), .A2(n13383), .ZN(n13384) );
  INV_X1 U16646 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18155) );
  XNOR2_X1 U16647 ( .A(n13383), .B(n13382), .ZN(n17862) );
  NOR2_X1 U16648 ( .A1(n13384), .A2(n17861), .ZN(n13387) );
  XOR2_X1 U16649 ( .A(n17416), .B(n13385), .Z(n13388) );
  NAND2_X1 U16650 ( .A1(n13387), .A2(n13388), .ZN(n17851) );
  NAND2_X1 U16651 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17851), .ZN(
        n13390) );
  NOR2_X1 U16652 ( .A1(n13386), .A2(n13390), .ZN(n13392) );
  INV_X1 U16653 ( .A(n13386), .ZN(n13391) );
  OR2_X1 U16654 ( .A1(n13388), .A2(n13387), .ZN(n17852) );
  OAI21_X1 U16655 ( .B1(n13391), .B2(n13390), .A(n17852), .ZN(n13389) );
  AOI21_X1 U16656 ( .B1(n13391), .B2(n13390), .A(n13389), .ZN(n17841) );
  NOR2_X2 U16657 ( .A1(n18117), .A2(n13393), .ZN(n18076) );
  NAND3_X1 U16658 ( .A1(n15782), .A2(n17940), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13394) );
  XOR2_X1 U16659 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13394), .Z(
        n16457) );
  INV_X1 U16660 ( .A(n16457), .ZN(n13395) );
  NOR2_X4 U16661 ( .A1(n18268), .A2(n16579), .ZN(n17916) );
  NAND2_X1 U16662 ( .A1(n13400), .A2(n13399), .ZN(P3_U2799) );
  INV_X1 U16663 ( .A(n14658), .ZN(n14574) );
  NAND4_X1 U16664 ( .A1(n13405), .A2(n20280), .A3(n13404), .A4(n13573), .ZN(
        n13406) );
  NAND2_X1 U16665 ( .A1(n13727), .A2(n13406), .ZN(n13408) );
  OAI22_X1 U16666 ( .A1(n14330), .A2(n12555), .B1(n14368), .B2(n13409), .ZN(
        n13411) );
  XNOR2_X1 U16667 ( .A(n13411), .B(n13410), .ZN(n14778) );
  INV_X1 U16668 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13413) );
  OAI22_X1 U16669 ( .A1(n14778), .A2(n14557), .B1(n13413), .B2(n20116), .ZN(
        n13414) );
  INV_X1 U16670 ( .A(n13414), .ZN(n13415) );
  INV_X1 U16671 ( .A(n13416), .ZN(n13417) );
  AOI22_X1 U16672 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U16673 ( .A1(n13419), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13420) );
  NAND2_X1 U16674 ( .A1(n13421), .A2(n13420), .ZN(n13439) );
  AOI22_X1 U16675 ( .A1(n12991), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10343), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13423) );
  AOI21_X1 U16676 ( .B1(n9636), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n13425), .ZN(n13422) );
  OAI211_X1 U16677 ( .C1(n15514), .C2(n13424), .A(n13423), .B(n13422), .ZN(
        n13438) );
  OAI21_X1 U16678 ( .B1(n10126), .B2(n13426), .A(n13425), .ZN(n13430) );
  OAI22_X1 U16679 ( .A1(n13428), .A2(n19377), .B1(n12889), .B2(n13427), .ZN(
        n13429) );
  AOI211_X1 U16680 ( .C1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n10339), .A(
        n13430), .B(n13429), .ZN(n13436) );
  AOI22_X1 U16681 ( .A1(n12999), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13431), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U16682 ( .A1(n13433), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13432), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13434) );
  NAND3_X1 U16683 ( .A1(n13436), .A2(n13435), .A3(n13434), .ZN(n13437) );
  OAI21_X1 U16684 ( .B1(n13439), .B2(n13438), .A(n13437), .ZN(n13440) );
  XNOR2_X1 U16685 ( .A(n13441), .B(n13440), .ZN(n14327) );
  NAND2_X1 U16686 ( .A1(n16385), .A2(n16389), .ZN(n13443) );
  AND2_X1 U16687 ( .A1(n11196), .A2(n19993), .ZN(n13512) );
  NAND3_X1 U16688 ( .A1(n11189), .A2(n13514), .A3(n13512), .ZN(n13442) );
  NAND2_X1 U16689 ( .A1(n13443), .A2(n13442), .ZN(n13766) );
  NAND2_X1 U16690 ( .A1(n19187), .A2(n13448), .ZN(n16196) );
  NOR4_X1 U16691 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n13452) );
  NOR4_X1 U16692 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13451) );
  NOR4_X1 U16693 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13450) );
  NOR4_X1 U16694 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13449) );
  NAND4_X1 U16695 ( .A1(n13452), .A2(n13451), .A3(n13450), .A4(n13449), .ZN(
        n13457) );
  NOR4_X1 U16696 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13455) );
  NOR4_X1 U16697 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13454) );
  NOR4_X1 U16698 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13453) );
  INV_X1 U16699 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19876) );
  NAND4_X1 U16700 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n19876), .ZN(
        n13456) );
  OAI21_X1 U16701 ( .B1(n13457), .B2(n13456), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13458) );
  INV_X2 U16702 ( .A(n19167), .ZN(n19166) );
  NAND2_X1 U16703 ( .A1(n19166), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13460) );
  INV_X1 U16704 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14569) );
  OR2_X1 U16705 ( .A1(n19166), .A2(n14569), .ZN(n13459) );
  NAND2_X1 U16706 ( .A1(n13460), .A2(n13459), .ZN(n19170) );
  INV_X1 U16707 ( .A(n19170), .ZN(n13462) );
  INV_X1 U16708 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13461) );
  OAI22_X1 U16709 ( .A1(n16196), .A2(n13462), .B1(n19187), .B2(n13461), .ZN(
        n13463) );
  AOI21_X1 U16710 ( .B1(n15278), .B2(n19206), .A(n13463), .ZN(n13466) );
  AND2_X1 U16711 ( .A1(n10184), .A2(n15558), .ZN(n13464) );
  NAND2_X1 U16712 ( .A1(n19187), .A2(n13464), .ZN(n13593) );
  AOI22_X1 U16713 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19160), .B1(n19159), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n13465) );
  OAI21_X1 U16714 ( .B1(n14327), .B2(n19210), .A(n13467), .ZN(P2_U2889) );
  NAND2_X1 U16715 ( .A1(n20209), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14790) );
  OAI21_X1 U16716 ( .B1(n15913), .B2(n14332), .A(n14790), .ZN(n13470) );
  AOI21_X1 U16717 ( .B1(n20199), .B2(n14335), .A(n13470), .ZN(n13474) );
  NAND2_X1 U16718 ( .A1(n13475), .A2(n19318), .ZN(n13482) );
  OAI21_X1 U16719 ( .B1(n19312), .B2(n9967), .A(n13476), .ZN(n13477) );
  INV_X1 U16720 ( .A(n13477), .ZN(n13478) );
  NOR2_X1 U16721 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13484) );
  NOR4_X1 U16722 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13483) );
  NAND4_X1 U16723 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13484), .A4(n13483), .ZN(n13487) );
  NOR2_X1 U16724 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13487), .ZN(n16557)
         );
  INV_X1 U16725 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20929) );
  NOR3_X1 U16726 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20929), .ZN(n13486) );
  NOR4_X1 U16727 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13485) );
  NAND4_X1 U16728 ( .A1(n20256), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13486), .A4(
        n13485), .ZN(U214) );
  NOR2_X1 U16729 ( .A1(n19166), .A2(n13487), .ZN(n16480) );
  NAND2_X1 U16730 ( .A1(n16480), .A2(U214), .ZN(U212) );
  NOR3_X1 U16731 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16928) );
  INV_X1 U16732 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16919) );
  NAND2_X1 U16733 ( .A1(n16928), .A2(n16919), .ZN(n16918) );
  NOR2_X1 U16734 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16918), .ZN(n16900) );
  INV_X1 U16735 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U16736 ( .A1(n16900), .A2(n15596), .ZN(n16886) );
  INV_X1 U16737 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16864) );
  NAND2_X1 U16738 ( .A1(n16871), .A2(n16864), .ZN(n16862) );
  INV_X1 U16739 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16844) );
  NAND2_X1 U16740 ( .A1(n16847), .A2(n16844), .ZN(n16843) );
  INV_X1 U16741 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16819) );
  NAND2_X1 U16742 ( .A1(n16820), .A2(n16819), .ZN(n16811) );
  INV_X1 U16743 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17150) );
  NAND2_X1 U16744 ( .A1(n16797), .A2(n17150), .ZN(n16792) );
  INV_X1 U16745 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16765) );
  NAND2_X1 U16746 ( .A1(n16770), .A2(n16765), .ZN(n16763) );
  INV_X1 U16747 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17114) );
  NAND2_X1 U16748 ( .A1(n16749), .A2(n17114), .ZN(n16743) );
  INV_X1 U16749 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16721) );
  NAND2_X1 U16750 ( .A1(n16728), .A2(n16721), .ZN(n16720) );
  INV_X1 U16751 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16696) );
  NAND2_X1 U16752 ( .A1(n16704), .A2(n16696), .ZN(n16695) );
  NOR2_X1 U16753 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16695), .ZN(n16683) );
  INV_X1 U16754 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16679) );
  NAND2_X1 U16755 ( .A1(n16683), .A2(n16679), .ZN(n16678) );
  NOR2_X1 U16756 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16678), .ZN(n16650) );
  INV_X1 U16757 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21056) );
  NAND2_X1 U16758 ( .A1(n16650), .A2(n21056), .ZN(n13491) );
  NOR2_X1 U16759 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n13491), .ZN(n16646) );
  NAND2_X1 U16760 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18904) );
  NAND2_X1 U16761 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18268), .ZN(n13490) );
  AOI211_X4 U16762 ( .C1(n18893), .C2(n18904), .A(n13503), .B(n13490), .ZN(
        n16955) );
  AOI211_X1 U16763 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n13491), .A(n16646), .B(
        n16954), .ZN(n13509) );
  INV_X1 U16764 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18824) );
  INV_X1 U16765 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18820) );
  NAND2_X1 U16766 ( .A1(n18768), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18908) );
  INV_X2 U16767 ( .A(n18908), .ZN(n18843) );
  NAND2_X1 U16768 ( .A1(n18843), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18836) );
  OAI211_X1 U16769 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18768), .B(n18830), .ZN(n18891) );
  INV_X1 U16770 ( .A(n18904), .ZN(n18895) );
  AOI211_X1 U16771 ( .C1(n18891), .C2(n18892), .A(n18895), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n13504) );
  INV_X1 U16772 ( .A(n13504), .ZN(n18745) );
  INV_X1 U16773 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18818) );
  INV_X1 U16774 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18800) );
  INV_X1 U16775 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18796) );
  INV_X1 U16776 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18792) );
  INV_X1 U16777 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18788) );
  INV_X1 U16778 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18784) );
  INV_X1 U16779 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18780) );
  NAND2_X1 U16780 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16926) );
  NOR2_X1 U16781 ( .A1(n18780), .A2(n16926), .ZN(n16901) );
  NAND2_X1 U16782 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16901), .ZN(n16890) );
  NOR2_X1 U16783 ( .A1(n18784), .A2(n16890), .ZN(n16867) );
  NAND2_X1 U16784 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16867), .ZN(n16861) );
  NOR2_X1 U16785 ( .A1(n18788), .A2(n16861), .ZN(n16850) );
  NAND2_X1 U16786 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16850), .ZN(n16832) );
  NOR2_X1 U16787 ( .A1(n18792), .A2(n16832), .ZN(n16821) );
  NAND2_X1 U16788 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16821), .ZN(n16808) );
  NOR2_X1 U16789 ( .A1(n18796), .A2(n16808), .ZN(n16800) );
  NAND2_X1 U16790 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16800), .ZN(n16785) );
  NOR2_X1 U16791 ( .A1(n18800), .A2(n16785), .ZN(n16776) );
  NAND2_X1 U16792 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16776), .ZN(n16775) );
  NAND2_X1 U16793 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16755) );
  NOR2_X1 U16794 ( .A1(n16775), .A2(n16755), .ZN(n16738) );
  NAND2_X1 U16795 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16738), .ZN(n16736) );
  NAND2_X1 U16796 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16719) );
  NOR2_X1 U16797 ( .A1(n16736), .A2(n16719), .ZN(n16707) );
  NAND2_X1 U16798 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16707), .ZN(n16671) );
  NAND2_X1 U16799 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16682) );
  NOR3_X1 U16800 ( .A1(n18818), .A2(n16671), .A3(n16682), .ZN(n13492) );
  NAND2_X1 U16801 ( .A1(n16925), .A2(n13492), .ZN(n16670) );
  NOR2_X1 U16802 ( .A1(n18820), .A2(n16670), .ZN(n16658) );
  NAND2_X1 U16803 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16658), .ZN(n16593) );
  INV_X1 U16804 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18822) );
  INV_X1 U16805 ( .A(n18913), .ZN(n18900) );
  NAND3_X1 U16806 ( .A1(n18898), .A2(n18910), .A3(n18893), .ZN(n18759) );
  NOR2_X2 U16807 ( .A1(n18859), .A2(n18759), .ZN(n16935) );
  NOR2_X1 U16808 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18850), .ZN(n18752) );
  INV_X1 U16809 ( .A(n18752), .ZN(n18600) );
  OR2_X1 U16810 ( .A1(n18754), .A2(n18600), .ZN(n18749) );
  AND2_X1 U16811 ( .A1(n16958), .A2(n13492), .ZN(n16661) );
  NAND2_X1 U16812 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16661), .ZN(n16653) );
  NOR2_X1 U16813 ( .A1(n18822), .A2(n16653), .ZN(n13493) );
  NAND2_X1 U16814 ( .A1(n16948), .A2(n16958), .ZN(n16957) );
  INV_X1 U16815 ( .A(n16957), .ZN(n16662) );
  AOI21_X1 U16816 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n13493), .A(n16662), 
        .ZN(n16643) );
  INV_X1 U16817 ( .A(n16643), .ZN(n13494) );
  AOI21_X1 U16818 ( .B1(n18824), .B2(n16593), .A(n13494), .ZN(n13508) );
  NOR2_X1 U16819 ( .A1(n17610), .A2(n17923), .ZN(n13500) );
  INV_X1 U16820 ( .A(n13500), .ZN(n13496) );
  NOR2_X1 U16821 ( .A1(n17611), .A2(n13496), .ZN(n17561) );
  INV_X1 U16822 ( .A(n17561), .ZN(n13495) );
  NOR2_X1 U16823 ( .A1(n9844), .A2(n13495), .ZN(n16598) );
  AOI21_X1 U16824 ( .B1(n9844), .B2(n13495), .A(n16598), .ZN(n17591) );
  INV_X1 U16825 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17621) );
  AOI22_X1 U16826 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13500), .B1(
        n13496), .B2(n17621), .ZN(n17617) );
  INV_X1 U16827 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17651) );
  NAND2_X1 U16828 ( .A1(n17678), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17645) );
  NOR2_X1 U16829 ( .A1(n9836), .A2(n17645), .ZN(n13499) );
  NAND2_X1 U16830 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13499), .ZN(
        n13497) );
  AOI22_X1 U16831 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17638), .B1(
        n17651), .B2(n13497), .ZN(n17653) );
  NAND2_X1 U16832 ( .A1(n17716), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16746) );
  NOR2_X1 U16833 ( .A1(n9840), .A2(n16746), .ZN(n17693) );
  NAND2_X1 U16834 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17693), .ZN(
        n16725) );
  NOR2_X1 U16835 ( .A1(n17730), .A2(n17923), .ZN(n17729) );
  NAND2_X1 U16836 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17729), .ZN(
        n16759) );
  INV_X1 U16837 ( .A(n16759), .ZN(n16747) );
  INV_X1 U16838 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16946) );
  NAND2_X1 U16839 ( .A1(n16747), .A2(n16946), .ZN(n16750) );
  OAI21_X1 U16840 ( .B1(n16725), .B2(n16750), .A(n13498), .ZN(n16715) );
  OAI21_X1 U16841 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16884), .A(
        n16715), .ZN(n16703) );
  AOI21_X1 U16842 ( .B1(n9836), .B2(n17645), .A(n13499), .ZN(n17681) );
  NOR2_X1 U16843 ( .A1(n16702), .A2(n16884), .ZN(n16692) );
  INV_X1 U16844 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17668) );
  XNOR2_X1 U16845 ( .A(n17668), .B(n13499), .ZN(n17671) );
  NOR2_X1 U16846 ( .A1(n16691), .A2(n16884), .ZN(n16685) );
  NAND2_X1 U16847 ( .A1(n17638), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17602) );
  AOI21_X1 U16848 ( .B1(n9843), .B2(n17602), .A(n13500), .ZN(n17632) );
  NOR2_X1 U16849 ( .A1(n17617), .A2(n16665), .ZN(n16664) );
  NOR2_X1 U16850 ( .A1(n16664), .A2(n16884), .ZN(n16652) );
  INV_X1 U16851 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16655) );
  NAND2_X1 U16852 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13500), .ZN(
        n13501) );
  AOI21_X1 U16853 ( .B1(n16655), .B2(n13501), .A(n17561), .ZN(n17603) );
  AOI211_X1 U16854 ( .C1(n17591), .C2(n13502), .A(n16596), .B(n18757), .ZN(
        n13507) );
  AOI211_X4 U16855 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18268), .A(n13504), .B(
        n13503), .ZN(n16956) );
  INV_X1 U16856 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n13505) );
  OAI22_X1 U16857 ( .A1(n9844), .A2(n16944), .B1(n16947), .B2(n13505), .ZN(
        n13506) );
  OR4_X1 U16858 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13506), .ZN(
        P3_U2645) );
  OR2_X1 U16859 ( .A1(n10767), .A2(n13775), .ZN(n13550) );
  INV_X1 U16860 ( .A(n13514), .ZN(n16386) );
  NOR2_X1 U16861 ( .A1(n13550), .A2(n16386), .ZN(n19141) );
  INV_X1 U16862 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20007) );
  OAI211_X1 U16863 ( .C1(n19141), .C2(n20007), .A(n18919), .B(n13510), .ZN(
        P2_U2814) );
  NOR2_X1 U16864 ( .A1(n13512), .A2(n13511), .ZN(n13513) );
  AND3_X1 U16865 ( .A1(n11189), .A2(n13514), .A3(n13513), .ZN(n16379) );
  OR2_X1 U16866 ( .A1(n16379), .A2(n13775), .ZN(n19984) );
  INV_X1 U16867 ( .A(n19984), .ZN(n13517) );
  INV_X1 U16868 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13516) );
  OAI21_X1 U16869 ( .B1(n13517), .B2(n13516), .A(n13515), .ZN(P2_U2819) );
  INV_X1 U16870 ( .A(n11196), .ZN(n13520) );
  INV_X1 U16871 ( .A(n18920), .ZN(n19991) );
  INV_X1 U16872 ( .A(n18919), .ZN(n13518) );
  OAI21_X1 U16873 ( .B1(n13518), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19991), 
        .ZN(n13519) );
  OAI21_X1 U16874 ( .B1(n13520), .B2(n19991), .A(n13519), .ZN(P2_U3612) );
  INV_X1 U16875 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13590) );
  NAND2_X2 U16876 ( .A1(n13521), .A2(n19993), .ZN(n19287) );
  NOR2_X1 U16877 ( .A1(n13540), .A2(n19284), .ZN(n13523) );
  NAND2_X1 U16878 ( .A1(n13523), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13522) );
  INV_X1 U16879 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16513) );
  INV_X1 U16880 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U16881 ( .A1(n19167), .A2(n16513), .B1(n17541), .B2(n19166), .ZN(
        n19183) );
  NAND2_X1 U16882 ( .A1(n13540), .A2(n19183), .ZN(n13543) );
  OAI211_X1 U16883 ( .C1(n13590), .C2(n13549), .A(n13522), .B(n13543), .ZN(
        P2_U2960) );
  INV_X1 U16884 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13524) );
  INV_X1 U16885 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13559) );
  INV_X1 U16886 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16529) );
  INV_X1 U16887 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18263) );
  AOI22_X1 U16888 ( .A1(n19167), .A2(n16529), .B1(n18263), .B2(n19166), .ZN(
        n19157) );
  INV_X1 U16889 ( .A(n19157), .ZN(n19265) );
  OAI222_X1 U16890 ( .A1(n13524), .A2(n13542), .B1(n13549), .B2(n13559), .C1(
        n19287), .C2(n19265), .ZN(P2_U2952) );
  AND2_X1 U16891 ( .A1(n20791), .A2(n16108), .ZN(n13566) );
  AOI21_X1 U16892 ( .B1(n13525), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13566), 
        .ZN(n13526) );
  NAND2_X1 U16893 ( .A1(n13620), .A2(n13526), .ZN(P1_U2801) );
  INV_X1 U16894 ( .A(n13527), .ZN(n15506) );
  NAND2_X1 U16895 ( .A1(n13529), .A2(n13528), .ZN(n13530) );
  XNOR2_X1 U16896 ( .A(n13530), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13617) );
  NOR2_X1 U16897 ( .A1(n19091), .A2(n19874), .ZN(n13610) );
  OAI21_X1 U16898 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13532), .A(
        n13531), .ZN(n13613) );
  NOR2_X1 U16899 ( .A1(n19323), .A2(n13613), .ZN(n13533) );
  AOI211_X1 U16900 ( .C1(n19313), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13610), .B(n13533), .ZN(n13534) );
  OAI21_X1 U16901 ( .B1(n19304), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13534), .ZN(n13535) );
  AOI21_X1 U16902 ( .B1(n19318), .B2(n13617), .A(n13535), .ZN(n13536) );
  OAI21_X1 U16903 ( .B1(n15506), .B2(n19305), .A(n13536), .ZN(P2_U3013) );
  INV_X1 U16904 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19229) );
  NAND2_X1 U16905 ( .A1(n19285), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U16906 ( .A1(n19166), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13538) );
  INV_X1 U16907 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16510) );
  OR2_X1 U16908 ( .A1(n19166), .A2(n16510), .ZN(n13537) );
  NAND2_X1 U16909 ( .A1(n13538), .A2(n13537), .ZN(n19178) );
  NAND2_X1 U16910 ( .A1(n13540), .A2(n19178), .ZN(n13547) );
  OAI211_X1 U16911 ( .C1(n19229), .C2(n13549), .A(n13539), .B(n13547), .ZN(
        P2_U2977) );
  NAND2_X1 U16912 ( .A1(n19285), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13541) );
  NAND2_X1 U16913 ( .A1(n13540), .A2(n19170), .ZN(n13545) );
  OAI211_X1 U16914 ( .C1(n13461), .C2(n13549), .A(n13541), .B(n13545), .ZN(
        P2_U2966) );
  INV_X1 U16915 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19233) );
  NAND2_X1 U16916 ( .A1(n19285), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13544) );
  OAI211_X1 U16917 ( .C1(n19233), .C2(n13549), .A(n13544), .B(n13543), .ZN(
        P2_U2975) );
  INV_X1 U16918 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19221) );
  NAND2_X1 U16919 ( .A1(n19285), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13546) );
  OAI211_X1 U16920 ( .C1(n19221), .C2(n13549), .A(n13546), .B(n13545), .ZN(
        P2_U2981) );
  INV_X1 U16921 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13565) );
  NAND2_X1 U16922 ( .A1(n19285), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13548) );
  OAI211_X1 U16923 ( .C1(n13565), .C2(n13549), .A(n13548), .B(n13547), .ZN(
        P2_U2962) );
  INV_X1 U16924 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14351) );
  OAI21_X1 U16925 ( .B1(n13771), .B2(n13550), .A(n13549), .ZN(n13551) );
  INV_X1 U16926 ( .A(n19249), .ZN(n13553) );
  NAND2_X1 U16927 ( .A1(n13553), .A2(n13552), .ZN(n13592) );
  NAND2_X1 U16928 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n16402) );
  OR2_X1 U16929 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16402), .ZN(n19217) );
  AND2_X2 U16930 ( .A1(n19249), .A2(n19217), .ZN(n19247) );
  AOI22_X1 U16931 ( .A1(n9637), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13554) );
  OAI21_X1 U16932 ( .B1(n14351), .B2(n13592), .A(n13554), .ZN(P2_U2922) );
  INV_X1 U16933 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13556) );
  AOI22_X1 U16934 ( .A1(n9637), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U16935 ( .B1(n13556), .B2(n13592), .A(n13555), .ZN(P2_U2929) );
  INV_X1 U16936 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15047) );
  AOI22_X1 U16937 ( .A1(n9637), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13557) );
  OAI21_X1 U16938 ( .B1(n15047), .B2(n13592), .A(n13557), .ZN(P2_U2923) );
  AOI22_X1 U16939 ( .A1(n9637), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13558) );
  OAI21_X1 U16940 ( .B1(n13559), .B2(n13592), .A(n13558), .ZN(P2_U2935) );
  INV_X1 U16941 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U16942 ( .A1(n9637), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13560) );
  OAI21_X1 U16943 ( .B1(n13561), .B2(n13592), .A(n13560), .ZN(P2_U2933) );
  INV_X1 U16944 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15108) );
  AOI22_X1 U16945 ( .A1(n9637), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13562) );
  OAI21_X1 U16946 ( .B1(n15108), .B2(n13592), .A(n13562), .ZN(P2_U2932) );
  INV_X1 U16947 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U16948 ( .A1(n9637), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13563) );
  OAI21_X1 U16949 ( .B1(n15097), .B2(n13592), .A(n13563), .ZN(P2_U2930) );
  AOI22_X1 U16950 ( .A1(n9637), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13564) );
  OAI21_X1 U16951 ( .B1(n13565), .B2(n13592), .A(n13564), .ZN(P2_U2925) );
  INV_X1 U16952 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15078) );
  INV_X1 U16953 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n20949) );
  INV_X1 U16954 ( .A(n19247), .ZN(n19216) );
  INV_X1 U16955 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16556) );
  OAI222_X1 U16956 ( .A1(n13592), .A2(n15078), .B1(n19217), .B2(n20949), .C1(
        n19216), .C2(n16556), .ZN(P2_U2926) );
  OAI21_X1 U16957 ( .B1(n13566), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n14035), 
        .ZN(n13567) );
  OAI21_X1 U16958 ( .B1(n13568), .B2(n14035), .A(n13567), .ZN(P1_U3487) );
  OR2_X1 U16959 ( .A1(n15774), .A2(n13569), .ZN(n13572) );
  NAND2_X1 U16960 ( .A1(n13570), .A2(n13575), .ZN(n13571) );
  NAND2_X1 U16961 ( .A1(n13572), .A2(n13571), .ZN(n20011) );
  INV_X1 U16962 ( .A(n15791), .ZN(n13627) );
  NOR2_X1 U16963 ( .A1(n13573), .A2(n13627), .ZN(n13721) );
  AOI21_X1 U16964 ( .B1(n13721), .B2(n14033), .A(n20850), .ZN(n20930) );
  NOR2_X1 U16965 ( .A1(n20011), .A2(n20930), .ZN(n15761) );
  OR2_X1 U16966 ( .A1(n15761), .A2(n20010), .ZN(n13581) );
  INV_X1 U16967 ( .A(n13581), .ZN(n20018) );
  INV_X1 U16968 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13583) );
  INV_X1 U16969 ( .A(n13574), .ZN(n13579) );
  NAND2_X1 U16970 ( .A1(n13576), .A2(n13575), .ZN(n13577) );
  MUX2_X1 U16971 ( .A(n13577), .B(n13706), .S(n15774), .Z(n13578) );
  AOI21_X1 U16972 ( .B1(n13580), .B2(n13579), .A(n13578), .ZN(n15763) );
  OR2_X1 U16973 ( .A1(n15763), .A2(n13581), .ZN(n13582) );
  OAI21_X1 U16974 ( .B1(n20018), .B2(n13583), .A(n13582), .ZN(P1_U3484) );
  AOI22_X1 U16975 ( .A1(n9637), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13584) );
  OAI21_X1 U16976 ( .B1(n13461), .B2(n13592), .A(n13584), .ZN(P2_U2921) );
  INV_X1 U16977 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14198) );
  AOI22_X1 U16978 ( .A1(n9637), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13585) );
  OAI21_X1 U16979 ( .B1(n14198), .B2(n13592), .A(n13585), .ZN(P2_U2934) );
  INV_X1 U16980 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U16981 ( .A1(n9637), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13586) );
  OAI21_X1 U16982 ( .B1(n15058), .B2(n13592), .A(n13586), .ZN(P2_U2924) );
  INV_X1 U16983 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U16984 ( .A1(n9637), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13587) );
  OAI21_X1 U16985 ( .B1(n13588), .B2(n13592), .A(n13587), .ZN(P2_U2931) );
  AOI22_X1 U16986 ( .A1(n9637), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13589) );
  OAI21_X1 U16987 ( .B1(n13590), .B2(n13592), .A(n13589), .ZN(P2_U2927) );
  INV_X1 U16988 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15089) );
  AOI22_X1 U16989 ( .A1(n9637), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U16990 ( .B1(n15089), .B2(n13592), .A(n13591), .ZN(P2_U2928) );
  NAND2_X1 U16991 ( .A1(n16196), .A2(n13593), .ZN(n19189) );
  AND2_X1 U16992 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19950), .ZN(n13594) );
  OAI211_X1 U16993 ( .C1(n19348), .C2(n19346), .A(n15543), .B(n13594), .ZN(
        n13595) );
  INV_X1 U16994 ( .A(n13595), .ZN(n13596) );
  INV_X1 U16995 ( .A(n13598), .ZN(n13599) );
  OAI21_X1 U16996 ( .B1(n13601), .B2(n13600), .A(n13599), .ZN(n19143) );
  INV_X1 U16997 ( .A(n19143), .ZN(n16349) );
  NOR2_X1 U16998 ( .A1(n14110), .A2(n19143), .ZN(n19209) );
  INV_X1 U16999 ( .A(n19209), .ZN(n13602) );
  OAI211_X1 U17000 ( .C1(n19970), .C2(n16349), .A(n13602), .B(n19191), .ZN(
        n13604) );
  AOI22_X1 U17001 ( .A1(n19206), .A2(n16349), .B1(n19205), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13603) );
  OAI211_X1 U17002 ( .C1(n19214), .C2(n19265), .A(n13604), .B(n13603), .ZN(
        P2_U2919) );
  INV_X1 U17003 ( .A(n13605), .ZN(n13607) );
  NAND2_X1 U17004 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  NAND2_X1 U17005 ( .A1(n13609), .A2(n13608), .ZN(n19965) );
  NAND2_X1 U17006 ( .A1(n16350), .A2(n19965), .ZN(n13612) );
  AOI21_X1 U17007 ( .B1(n16348), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13610), .ZN(n13611) );
  OAI211_X1 U17008 ( .C1(n13613), .C2(n19343), .A(n13612), .B(n13611), .ZN(
        n13616) );
  AOI211_X1 U17009 ( .C1(n15508), .C2(n16351), .A(n13614), .B(n16359), .ZN(
        n13615) );
  AOI211_X1 U17010 ( .C1(n13617), .C2(n16344), .A(n13616), .B(n13615), .ZN(
        n13618) );
  OAI21_X1 U17011 ( .B1(n15506), .B2(n16341), .A(n13618), .ZN(P2_U3045) );
  NOR2_X1 U17012 ( .A1(n15770), .A2(n15768), .ZN(n13619) );
  OR2_X1 U17013 ( .A1(n20151), .A2(n20275), .ZN(n13794) );
  INV_X1 U17014 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13625) );
  OR2_X1 U17015 ( .A1(n20151), .A2(n13621), .ZN(n13795) );
  INV_X1 U17016 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13622) );
  NOR2_X1 U17017 ( .A1(n20257), .A2(n13622), .ZN(n13623) );
  AOI21_X1 U17018 ( .B1(DATAI_15_), .B2(n20257), .A(n13623), .ZN(n14636) );
  INV_X1 U17019 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13624) );
  OAI222_X1 U17020 ( .A1(n13794), .A2(n13625), .B1(n13795), .B2(n14636), .C1(
        n13624), .C2(n13824), .ZN(P1_U2967) );
  INV_X1 U17021 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13632) );
  INV_X1 U17022 ( .A(n13626), .ZN(n13628) );
  OAI21_X1 U17023 ( .B1(n15750), .B2(n13628), .A(n13627), .ZN(n13720) );
  INV_X1 U17024 ( .A(n13720), .ZN(n13629) );
  NAND2_X1 U17025 ( .A1(n20121), .A2(n11412), .ZN(n13656) );
  NAND2_X1 U17026 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16106) );
  NOR2_X1 U17027 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16106), .ZN(n20120) );
  INV_X2 U17028 ( .A(n20123), .ZN(n20138) );
  AOI22_X1 U17029 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13631) );
  OAI21_X1 U17030 ( .B1(n13632), .B2(n13656), .A(n13631), .ZN(P1_U2906) );
  INV_X1 U17031 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U17032 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13633) );
  OAI21_X1 U17033 ( .B1(n13634), .B2(n13656), .A(n13633), .ZN(P1_U2910) );
  INV_X1 U17034 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U17035 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13635) );
  OAI21_X1 U17036 ( .B1(n13636), .B2(n13656), .A(n13635), .ZN(P1_U2919) );
  INV_X1 U17037 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13638) );
  AOI22_X1 U17038 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13637) );
  OAI21_X1 U17039 ( .B1(n13638), .B2(n13656), .A(n13637), .ZN(P1_U2908) );
  INV_X1 U17040 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U17041 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13639) );
  OAI21_X1 U17042 ( .B1(n13640), .B2(n13656), .A(n13639), .ZN(P1_U2909) );
  INV_X1 U17043 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14629) );
  AOI22_X1 U17044 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13641) );
  OAI21_X1 U17045 ( .B1(n14629), .B2(n13656), .A(n13641), .ZN(P1_U2920) );
  AOI22_X1 U17046 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13642) );
  OAI21_X1 U17047 ( .B1(n14343), .B2(n13656), .A(n13642), .ZN(P1_U2907) );
  INV_X1 U17048 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13644) );
  AOI22_X1 U17049 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13643) );
  OAI21_X1 U17050 ( .B1(n13644), .B2(n13656), .A(n13643), .ZN(P1_U2917) );
  INV_X1 U17051 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U17052 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13645) );
  OAI21_X1 U17053 ( .B1(n13646), .B2(n13656), .A(n13645), .ZN(P1_U2913) );
  INV_X1 U17054 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U17055 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13647) );
  OAI21_X1 U17056 ( .B1(n14604), .B2(n13656), .A(n13647), .ZN(P1_U2914) );
  INV_X1 U17057 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13649) );
  AOI22_X1 U17058 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13648) );
  OAI21_X1 U17059 ( .B1(n13649), .B2(n13656), .A(n13648), .ZN(P1_U2911) );
  AOI22_X1 U17060 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13650) );
  OAI21_X1 U17061 ( .B1(n14595), .B2(n13656), .A(n13650), .ZN(P1_U2912) );
  INV_X1 U17062 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13652) );
  AOI22_X1 U17063 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13651) );
  OAI21_X1 U17064 ( .B1(n13652), .B2(n13656), .A(n13651), .ZN(P1_U2918) );
  INV_X1 U17065 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U17066 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13653) );
  OAI21_X1 U17067 ( .B1(n13654), .B2(n13656), .A(n13653), .ZN(P1_U2915) );
  INV_X1 U17068 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14612) );
  AOI22_X1 U17069 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20120), .B1(n20138), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13655) );
  OAI21_X1 U17070 ( .B1(n14612), .B2(n13656), .A(n13655), .ZN(P1_U2916) );
  OAI21_X1 U17071 ( .B1(n13659), .B2(n13658), .A(n13657), .ZN(n20108) );
  NAND2_X1 U17072 ( .A1(n13660), .A2(n15913), .ZN(n13664) );
  INV_X1 U17073 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13661) );
  NOR2_X1 U17074 ( .A1(n20244), .A2(n13661), .ZN(n14901) );
  OAI21_X1 U17075 ( .B1(n13662), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12354), .ZN(n14897) );
  NOR2_X1 U17076 ( .A1(n14897), .A2(n20016), .ZN(n13663) );
  AOI211_X1 U17077 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13664), .A(
        n14901), .B(n13663), .ZN(n13665) );
  OAI21_X1 U17078 ( .B1(n20258), .B2(n20108), .A(n13665), .ZN(P1_U2999) );
  NAND2_X1 U17079 ( .A1(n13667), .A2(n13666), .ZN(n13669) );
  AND2_X1 U17080 ( .A1(n13669), .A2(n9922), .ZN(n19951) );
  AOI21_X1 U17081 ( .B1(n13672), .B2(n13671), .A(n13670), .ZN(n19308) );
  NAND2_X1 U17082 ( .A1(n19308), .A2(n16344), .ZN(n13680) );
  OAI21_X1 U17083 ( .B1(n13675), .B2(n13674), .A(n13673), .ZN(n19302) );
  INV_X1 U17084 ( .A(n19302), .ZN(n13678) );
  OAI21_X1 U17085 ( .B1(n15427), .B2(n13683), .A(n13676), .ZN(n13677) );
  AOI22_X1 U17086 ( .A1(n16329), .A2(n13678), .B1(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13677), .ZN(n13679) );
  OAI211_X1 U17087 ( .C1(n19951), .C2(n19330), .A(n13680), .B(n13679), .ZN(
        n13685) );
  NAND2_X1 U17088 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19291), .ZN(n19309) );
  OAI211_X1 U17089 ( .C1(n13683), .C2(n13682), .A(n13681), .B(n19309), .ZN(
        n13684) );
  AOI211_X1 U17090 ( .C1(n19338), .C2(n14127), .A(n13685), .B(n13684), .ZN(
        n13686) );
  INV_X1 U17091 ( .A(n13686), .ZN(P2_U3044) );
  XOR2_X1 U17092 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13846), .Z(n13690)
         );
  INV_X1 U17093 ( .A(n13850), .ZN(n13687) );
  OAI21_X1 U17094 ( .B1(n13739), .B2(n13688), .A(n13687), .ZN(n19120) );
  MUX2_X1 U17095 ( .A(n19120), .B(n10835), .S(n15042), .Z(n13689) );
  OAI21_X1 U17096 ( .B1(n13690), .B2(n15044), .A(n13689), .ZN(P2_U2882) );
  NOR2_X1 U17097 ( .A1(n15036), .A2(n10281), .ZN(n13695) );
  AOI21_X1 U17098 ( .B1(n14948), .B2(n15036), .A(n13695), .ZN(n13696) );
  OAI21_X1 U17099 ( .B1(n14104), .B2(n15044), .A(n13696), .ZN(P2_U2884) );
  INV_X1 U17100 ( .A(n15750), .ZN(n13716) );
  XNOR2_X1 U17101 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13715) );
  INV_X1 U17102 ( .A(n13698), .ZN(n20265) );
  INV_X1 U17103 ( .A(n12444), .ZN(n13719) );
  INV_X1 U17104 ( .A(n13700), .ZN(n13701) );
  AND4_X1 U17105 ( .A1(n13699), .A2(n13702), .A3(n13719), .A4(n13701), .ZN(
        n13703) );
  NAND2_X1 U17106 ( .A1(n13704), .A2(n13703), .ZN(n14924) );
  NAND2_X1 U17107 ( .A1(n20265), .A2(n14924), .ZN(n13714) );
  OR2_X1 U17108 ( .A1(n13706), .A2(n13705), .ZN(n13958) );
  INV_X1 U17109 ( .A(n13952), .ZN(n13709) );
  INV_X1 U17110 ( .A(n13707), .ZN(n14919) );
  NAND2_X1 U17111 ( .A1(n14919), .A2(n11241), .ZN(n13708) );
  NAND2_X1 U17112 ( .A1(n13709), .A2(n13708), .ZN(n13717) );
  INV_X1 U17113 ( .A(n14922), .ZN(n13710) );
  NAND2_X1 U17114 ( .A1(n13711), .A2(n13710), .ZN(n13963) );
  NOR2_X1 U17115 ( .A1(n13963), .A2(n13717), .ZN(n13712) );
  AOI21_X1 U17116 ( .B1(n13958), .B2(n13717), .A(n13712), .ZN(n13713) );
  OAI211_X1 U17117 ( .C1(n13716), .C2(n13715), .A(n13714), .B(n13713), .ZN(
        n13951) );
  AOI22_X1 U17118 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20254), .B2(n12440), .ZN(
        n14926) );
  NOR2_X1 U17119 ( .A1(n16108), .A2(n20223), .ZN(n14928) );
  INV_X1 U17120 ( .A(n13717), .ZN(n13718) );
  AOI222_X1 U17121 ( .A1(n13951), .A2(n16097), .B1(n14926), .B2(n14928), .C1(
        n14930), .C2(n13718), .ZN(n13732) );
  AND2_X1 U17122 ( .A1(n13720), .A2(n13719), .ZN(n13722) );
  OR3_X1 U17123 ( .A1(n13723), .A2(n13722), .A3(n13721), .ZN(n13729) );
  NOR2_X1 U17124 ( .A1(n14036), .A2(n13724), .ZN(n13725) );
  NOR2_X1 U17125 ( .A1(n13726), .A2(n13725), .ZN(n13728) );
  NAND4_X1 U17126 ( .A1(n13730), .A2(n13729), .A3(n13728), .A4(n13727), .ZN(
        n13973) );
  INV_X1 U17127 ( .A(n13973), .ZN(n15747) );
  OR2_X1 U17128 ( .A1(n9758), .A2(n16106), .ZN(n16111) );
  INV_X1 U17129 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20017) );
  OAI22_X1 U17130 ( .A1(n15747), .A2(n20010), .B1(n16111), .B2(n20017), .ZN(
        n16096) );
  AOI21_X1 U17131 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n9758), .A(n16096), 
        .ZN(n14932) );
  NAND2_X1 U17132 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14932), .ZN(
        n13731) );
  OAI21_X1 U17133 ( .B1(n13732), .B2(n14932), .A(n13731), .ZN(P1_U3472) );
  NAND2_X1 U17134 ( .A1(n10184), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13733) );
  NAND2_X1 U17135 ( .A1(n13693), .A2(n13733), .ZN(n13738) );
  INV_X1 U17136 ( .A(n13734), .ZN(n13735) );
  NAND2_X1 U17137 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  OAI21_X1 U17138 ( .B1(n13738), .B2(n13737), .A(n13846), .ZN(n19131) );
  AOI21_X1 U17139 ( .B1(n13741), .B2(n13740), .A(n13739), .ZN(n19339) );
  NOR2_X1 U17140 ( .A1(n15036), .A2(n20945), .ZN(n13742) );
  AOI21_X1 U17141 ( .B1(n19339), .B2(n15036), .A(n13742), .ZN(n13743) );
  OAI21_X1 U17142 ( .B1(n19131), .B2(n15044), .A(n13743), .ZN(P2_U2883) );
  XNOR2_X1 U17143 ( .A(n13744), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13749) );
  OAI21_X1 U17144 ( .B1(n13745), .B2(n13746), .A(n9706), .ZN(n19102) );
  MUX2_X1 U17145 ( .A(n19102), .B(n13747), .S(n15042), .Z(n13748) );
  OAI21_X1 U17146 ( .B1(n13749), .B2(n15044), .A(n13748), .ZN(P2_U2880) );
  INV_X1 U17147 ( .A(n14924), .ZN(n13750) );
  OAI22_X1 U17148 ( .A1(n11556), .A2(n13750), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14922), .ZN(n15749) );
  INV_X1 U17149 ( .A(n14930), .ZN(n14934) );
  OAI22_X1 U17150 ( .A1(n14934), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n16108), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13751) );
  AOI21_X1 U17151 ( .B1(n16097), .B2(n15749), .A(n13751), .ZN(n13754) );
  AOI21_X1 U17152 ( .B1(n15750), .B2(n16097), .A(n14932), .ZN(n13753) );
  OAI22_X1 U17153 ( .A1(n13754), .A2(n14932), .B1(n13753), .B2(n13752), .ZN(
        P1_U3474) );
  MUX2_X1 U17154 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n14127), .S(n15036), .Z(
        n13758) );
  AOI21_X1 U17155 ( .B1(n19955), .B2(n15029), .A(n13758), .ZN(n13759) );
  INV_X1 U17156 ( .A(n13759), .ZN(P2_U2885) );
  INV_X1 U17157 ( .A(n13760), .ZN(n13761) );
  NOR2_X1 U17158 ( .A1(n13761), .A2(n11209), .ZN(n15519) );
  CLKBUF_X1 U17159 ( .A(n13762), .Z(n15503) );
  AND2_X1 U17160 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15516), .ZN(
        n13778) );
  INV_X1 U17161 ( .A(n13778), .ZN(n13763) );
  NAND2_X1 U17162 ( .A1(n15503), .A2(n13763), .ZN(n13765) );
  INV_X1 U17163 ( .A(n10330), .ZN(n13764) );
  NAND2_X1 U17164 ( .A1(n13764), .A2(n16364), .ZN(n15513) );
  OAI211_X1 U17165 ( .C1(n15519), .C2(n10339), .A(n13765), .B(n15513), .ZN(
        n16360) );
  NOR2_X1 U17166 ( .A1(n13085), .A2(n16402), .ZN(n16411) );
  INV_X1 U17167 ( .A(n13766), .ZN(n13774) );
  AND2_X1 U17168 ( .A1(n13768), .A2(n13767), .ZN(n13773) );
  OR2_X1 U17169 ( .A1(n10767), .A2(n13769), .ZN(n13770) );
  OR2_X1 U17170 ( .A1(n13771), .A2(n13770), .ZN(n13772) );
  OAI22_X1 U17171 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19950), .B1(n16392), 
        .B2(n13775), .ZN(n13776) );
  AOI21_X1 U17172 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16411), .A(n13776), .ZN(
        n15696) );
  AOI21_X1 U17173 ( .B1(n19940), .B2(n16360), .A(n15696), .ZN(n13784) );
  INV_X1 U17174 ( .A(n16404), .ZN(n15525) );
  INV_X1 U17175 ( .A(n13777), .ZN(n16387) );
  OR2_X1 U17176 ( .A1(n16385), .A2(n16387), .ZN(n15522) );
  AOI22_X1 U17177 ( .A1(n15522), .A2(n15513), .B1(n13778), .B2(n15503), .ZN(
        n13780) );
  OAI21_X1 U17178 ( .B1(n13780), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13779), .ZN(n13781) );
  AOI21_X1 U17179 ( .B1(n14948), .B2(n14165), .A(n13781), .ZN(n16362) );
  INV_X1 U17180 ( .A(n16362), .ZN(n13782) );
  AOI22_X1 U17181 ( .A1(n19947), .A2(n15525), .B1(n19940), .B2(n13782), .ZN(
        n13783) );
  OAI22_X1 U17182 ( .A1(n13784), .A2(n10138), .B1(n15696), .B2(n13783), .ZN(
        P2_U3596) );
  OAI21_X1 U17183 ( .B1(n13787), .B2(n13786), .A(n13785), .ZN(n20231) );
  INV_X1 U17184 ( .A(n13788), .ZN(n13789) );
  AOI21_X1 U17185 ( .B1(n13790), .B2(n13865), .A(n13789), .ZN(n20084) );
  AOI22_X1 U17186 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13791) );
  OAI21_X1 U17187 ( .B1(n20193), .B2(n20082), .A(n13791), .ZN(n13792) );
  AOI21_X1 U17188 ( .B1(n20084), .B2(n20189), .A(n13792), .ZN(n13793) );
  OAI21_X1 U17189 ( .B1(n20016), .B2(n20231), .A(n13793), .ZN(P1_U2997) );
  AOI22_X1 U17190 ( .A1(n20181), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20176), .ZN(n13799) );
  NAND2_X1 U17191 ( .A1(n20257), .A2(DATAI_1_), .ZN(n13797) );
  NAND2_X1 U17192 ( .A1(n20256), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13796) );
  AND2_X1 U17193 ( .A1(n13797), .A2(n13796), .ZN(n20277) );
  INV_X1 U17194 ( .A(n20277), .ZN(n13798) );
  NAND2_X1 U17195 ( .A1(n20166), .A2(n13798), .ZN(n13827) );
  NAND2_X1 U17196 ( .A1(n13799), .A2(n13827), .ZN(P1_U2938) );
  AOI22_X1 U17197 ( .A1(n20181), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20176), .ZN(n13803) );
  NAND2_X1 U17198 ( .A1(n20257), .A2(DATAI_5_), .ZN(n13801) );
  NAND2_X1 U17199 ( .A1(n20256), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13800) );
  AND2_X1 U17200 ( .A1(n13801), .A2(n13800), .ZN(n20297) );
  INV_X1 U17201 ( .A(n20297), .ZN(n13802) );
  NAND2_X1 U17202 ( .A1(n20166), .A2(n13802), .ZN(n13829) );
  NAND2_X1 U17203 ( .A1(n13803), .A2(n13829), .ZN(P1_U2942) );
  AOI22_X1 U17204 ( .A1(n20181), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20176), .ZN(n13807) );
  NAND2_X1 U17205 ( .A1(n20257), .A2(DATAI_7_), .ZN(n13805) );
  NAND2_X1 U17206 ( .A1(n20256), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13804) );
  AND2_X1 U17207 ( .A1(n13805), .A2(n13804), .ZN(n20309) );
  INV_X1 U17208 ( .A(n20309), .ZN(n13806) );
  NAND2_X1 U17209 ( .A1(n20166), .A2(n13806), .ZN(n13837) );
  NAND2_X1 U17210 ( .A1(n13807), .A2(n13837), .ZN(P1_U2959) );
  AOI22_X1 U17211 ( .A1(n20181), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20176), .ZN(n13811) );
  NAND2_X1 U17212 ( .A1(n20257), .A2(DATAI_3_), .ZN(n13809) );
  NAND2_X1 U17213 ( .A1(n20256), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13808) );
  AND2_X1 U17214 ( .A1(n13809), .A2(n13808), .ZN(n20286) );
  INV_X1 U17215 ( .A(n20286), .ZN(n13810) );
  NAND2_X1 U17216 ( .A1(n20166), .A2(n13810), .ZN(n13825) );
  NAND2_X1 U17217 ( .A1(n13811), .A2(n13825), .ZN(P1_U2940) );
  AOI22_X1 U17218 ( .A1(n20181), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20176), .ZN(n13815) );
  NAND2_X1 U17219 ( .A1(n20257), .A2(DATAI_4_), .ZN(n13813) );
  NAND2_X1 U17220 ( .A1(n20256), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13812) );
  AND2_X1 U17221 ( .A1(n13813), .A2(n13812), .ZN(n20292) );
  INV_X1 U17222 ( .A(n20292), .ZN(n13814) );
  NAND2_X1 U17223 ( .A1(n20166), .A2(n13814), .ZN(n13841) );
  NAND2_X1 U17224 ( .A1(n13815), .A2(n13841), .ZN(P1_U2941) );
  AOI22_X1 U17225 ( .A1(n20181), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20176), .ZN(n13819) );
  NAND2_X1 U17226 ( .A1(n20257), .A2(DATAI_0_), .ZN(n13817) );
  NAND2_X1 U17227 ( .A1(n20256), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13816) );
  AND2_X1 U17228 ( .A1(n13817), .A2(n13816), .ZN(n20267) );
  INV_X1 U17229 ( .A(n20267), .ZN(n13818) );
  NAND2_X1 U17230 ( .A1(n20166), .A2(n13818), .ZN(n13843) );
  NAND2_X1 U17231 ( .A1(n13819), .A2(n13843), .ZN(P1_U2937) );
  AOI22_X1 U17232 ( .A1(n20181), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20176), .ZN(n13823) );
  NAND2_X1 U17233 ( .A1(n20257), .A2(DATAI_2_), .ZN(n13821) );
  NAND2_X1 U17234 ( .A1(n20256), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13820) );
  AND2_X1 U17235 ( .A1(n13821), .A2(n13820), .ZN(n20282) );
  INV_X1 U17236 ( .A(n20282), .ZN(n13822) );
  NAND2_X1 U17237 ( .A1(n20166), .A2(n13822), .ZN(n13835) );
  NAND2_X1 U17238 ( .A1(n13823), .A2(n13835), .ZN(P1_U2939) );
  INV_X1 U17239 ( .A(n13824), .ZN(n20176) );
  AOI22_X1 U17240 ( .A1(n20181), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20176), .ZN(n13826) );
  NAND2_X1 U17241 ( .A1(n13826), .A2(n13825), .ZN(P1_U2955) );
  AOI22_X1 U17242 ( .A1(n20181), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20176), .ZN(n13828) );
  NAND2_X1 U17243 ( .A1(n13828), .A2(n13827), .ZN(P1_U2953) );
  AOI22_X1 U17244 ( .A1(n20181), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20176), .ZN(n13830) );
  NAND2_X1 U17245 ( .A1(n13830), .A2(n13829), .ZN(P1_U2957) );
  AOI22_X1 U17246 ( .A1(n20181), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20176), .ZN(n13834) );
  NAND2_X1 U17247 ( .A1(n20257), .A2(DATAI_6_), .ZN(n13832) );
  NAND2_X1 U17248 ( .A1(n20256), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13831) );
  AND2_X1 U17249 ( .A1(n13832), .A2(n13831), .ZN(n20301) );
  INV_X1 U17250 ( .A(n20301), .ZN(n13833) );
  NAND2_X1 U17251 ( .A1(n20166), .A2(n13833), .ZN(n13839) );
  NAND2_X1 U17252 ( .A1(n13834), .A2(n13839), .ZN(P1_U2958) );
  AOI22_X1 U17253 ( .A1(n20181), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20176), .ZN(n13836) );
  NAND2_X1 U17254 ( .A1(n13836), .A2(n13835), .ZN(P1_U2954) );
  AOI22_X1 U17255 ( .A1(n20181), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20176), .ZN(n13838) );
  NAND2_X1 U17256 ( .A1(n13838), .A2(n13837), .ZN(P1_U2944) );
  AOI22_X1 U17257 ( .A1(n20181), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20176), .ZN(n13840) );
  NAND2_X1 U17258 ( .A1(n13840), .A2(n13839), .ZN(P1_U2943) );
  AOI22_X1 U17259 ( .A1(n20181), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20176), .ZN(n13842) );
  NAND2_X1 U17260 ( .A1(n13842), .A2(n13841), .ZN(P1_U2956) );
  AOI22_X1 U17261 ( .A1(n20181), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20176), .ZN(n13844) );
  NAND2_X1 U17262 ( .A1(n13844), .A2(n13843), .ZN(P1_U2952) );
  NOR2_X1 U17263 ( .A1(n13846), .A2(n13845), .ZN(n13848) );
  INV_X1 U17264 ( .A(n13744), .ZN(n13847) );
  OAI211_X1 U17265 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13848), .A(
        n13847), .B(n15029), .ZN(n13853) );
  NOR2_X1 U17266 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  NOR2_X1 U17267 ( .A1(n13745), .A2(n13851), .ZN(n19111) );
  NAND2_X1 U17268 ( .A1(n19111), .A2(n15036), .ZN(n13852) );
  OAI211_X1 U17269 ( .C1(n15036), .C2(n13854), .A(n13853), .B(n13852), .ZN(
        P2_U2881) );
  INV_X1 U17270 ( .A(n20084), .ZN(n13873) );
  INV_X1 U17271 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13859) );
  INV_X1 U17272 ( .A(n13855), .ZN(n13856) );
  OAI21_X1 U17273 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n20227) );
  OAI222_X1 U17274 ( .A1(n13873), .A2(n14568), .B1(n20116), .B2(n13859), .C1(
        n20227), .C2(n14557), .ZN(P1_U2870) );
  MUX2_X1 U17275 ( .A(n10494), .B(n15506), .S(n15036), .Z(n13862) );
  OAI21_X1 U17276 ( .B1(n19960), .B2(n15044), .A(n13862), .ZN(P2_U2886) );
  MUX2_X1 U17277 ( .A(n14166), .B(n13863), .S(n15042), .Z(n13864) );
  OAI21_X1 U17278 ( .B1(n14110), .B2(n15044), .A(n13864), .ZN(P2_U2887) );
  XNOR2_X1 U17279 ( .A(n20089), .B(n12573), .ZN(n20245) );
  INV_X1 U17280 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13868) );
  OAI21_X1 U17281 ( .B1(n13867), .B2(n13866), .A(n13865), .ZN(n20203) );
  OAI222_X1 U17282 ( .A1(n20245), .A2(n14557), .B1(n20116), .B2(n13868), .C1(
        n20203), .C2(n14568), .ZN(P1_U2871) );
  NAND2_X1 U17283 ( .A1(n13870), .A2(n11541), .ZN(n13871) );
  INV_X1 U17284 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20137) );
  INV_X1 U17285 ( .A(n13871), .ZN(n13872) );
  OAI222_X1 U17286 ( .A1(n14647), .A2(n13873), .B1(n14637), .B2(n20137), .C1(
        n14645), .C2(n20282), .ZN(P1_U2902) );
  OAI21_X1 U17287 ( .B1(n13876), .B2(n13875), .A(n13874), .ZN(n14050) );
  INV_X1 U17288 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20135) );
  OAI222_X1 U17289 ( .A1(n14647), .A2(n14050), .B1(n14637), .B2(n20135), .C1(
        n14645), .C2(n20286), .ZN(P1_U2901) );
  INV_X1 U17290 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20144) );
  OAI222_X1 U17291 ( .A1(n14647), .A2(n20108), .B1(n14637), .B2(n20144), .C1(
        n14645), .C2(n20267), .ZN(P1_U2904) );
  INV_X1 U17292 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20140) );
  OAI222_X1 U17293 ( .A1(n14647), .A2(n20203), .B1(n14637), .B2(n20140), .C1(
        n14645), .C2(n20277), .ZN(P1_U2903) );
  XOR2_X1 U17294 ( .A(n19951), .B(n19955), .Z(n13881) );
  OR2_X1 U17295 ( .A1(n19963), .A2(n19965), .ZN(n13878) );
  NAND2_X1 U17296 ( .A1(n19963), .A2(n19965), .ZN(n13877) );
  NAND2_X1 U17297 ( .A1(n13878), .A2(n13877), .ZN(n19208) );
  NOR2_X1 U17298 ( .A1(n19208), .A2(n19209), .ZN(n19207) );
  INV_X1 U17299 ( .A(n13878), .ZN(n13879) );
  NOR2_X1 U17300 ( .A1(n19207), .A2(n13879), .ZN(n13880) );
  NOR2_X1 U17301 ( .A1(n13881), .A2(n13880), .ZN(n14051) );
  AOI21_X1 U17302 ( .B1(n13881), .B2(n13880), .A(n14051), .ZN(n13885) );
  INV_X1 U17303 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16522) );
  INV_X1 U17304 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18271) );
  AOI22_X1 U17305 ( .A1(n19167), .A2(n16522), .B1(n18271), .B2(n19166), .ZN(
        n19252) );
  AOI22_X1 U17306 ( .A1(n19189), .A2(n19252), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19205), .ZN(n13884) );
  INV_X1 U17307 ( .A(n19951), .ZN(n13882) );
  NAND2_X1 U17308 ( .A1(n13882), .A2(n19206), .ZN(n13883) );
  OAI211_X1 U17309 ( .C1(n13885), .C2(n19210), .A(n13884), .B(n13883), .ZN(
        P2_U2917) );
  OR2_X1 U17310 ( .A1(n13855), .A2(n13886), .ZN(n13887) );
  AND2_X1 U17311 ( .A1(n13942), .A2(n13887), .ZN(n20214) );
  INV_X1 U17312 ( .A(n20116), .ZN(n14566) );
  AOI22_X1 U17313 ( .A1(n20111), .A2(n20214), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14566), .ZN(n13888) );
  OAI21_X1 U17314 ( .B1(n14050), .B2(n14542), .A(n13888), .ZN(P1_U2869) );
  INV_X1 U17315 ( .A(n13889), .ZN(n13890) );
  NAND2_X1 U17316 ( .A1(n9706), .A2(n13890), .ZN(n13891) );
  AND2_X1 U17317 ( .A1(n13891), .A2(n13897), .ZN(n19085) );
  INV_X1 U17318 ( .A(n19085), .ZN(n15270) );
  OAI211_X1 U17319 ( .C1(n9717), .C2(n10090), .A(n15029), .B(n13893), .ZN(
        n13895) );
  NAND2_X1 U17320 ( .A1(n15042), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13894) );
  OAI211_X1 U17321 ( .C1(n15270), .C2(n15042), .A(n13895), .B(n13894), .ZN(
        P2_U2879) );
  INV_X1 U17322 ( .A(n13896), .ZN(n13985) );
  XNOR2_X1 U17323 ( .A(n13893), .B(n13985), .ZN(n13900) );
  AOI21_X1 U17324 ( .B1(n13898), .B2(n13897), .A(n9705), .ZN(n15494) );
  INV_X1 U17325 ( .A(n15494), .ZN(n19074) );
  MUX2_X1 U17326 ( .A(n10857), .B(n19074), .S(n15036), .Z(n13899) );
  OAI21_X1 U17327 ( .B1(n13900), .B2(n15044), .A(n13899), .ZN(P2_U2878) );
  OR2_X1 U17328 ( .A1(n12524), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13902) );
  AND2_X1 U17329 ( .A1(n13902), .A2(n13901), .ZN(n20098) );
  INV_X1 U17330 ( .A(n20098), .ZN(n13903) );
  OAI222_X1 U17331 ( .A1(n20108), .A2(n14568), .B1(n13904), .B2(n20116), .C1(
        n13903), .C2(n14557), .ZN(P1_U2872) );
  AND2_X1 U17332 ( .A1(n13906), .A2(n13905), .ZN(n13908) );
  OR2_X1 U17333 ( .A1(n13908), .A2(n13907), .ZN(n15966) );
  INV_X1 U17334 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20131) );
  OAI222_X1 U17335 ( .A1(n14647), .A2(n15966), .B1(n14637), .B2(n20131), .C1(
        n14645), .C2(n20297), .ZN(P1_U2899) );
  OAI21_X1 U17336 ( .B1(n13911), .B2(n13910), .A(n13909), .ZN(n20215) );
  INV_X1 U17337 ( .A(n14050), .ZN(n13914) );
  AOI22_X1 U17338 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13912) );
  OAI21_X1 U17339 ( .B1(n20193), .B2(n14046), .A(n13912), .ZN(n13913) );
  AOI21_X1 U17340 ( .B1(n13914), .B2(n20189), .A(n13913), .ZN(n13915) );
  OAI21_X1 U17341 ( .B1(n20215), .B2(n20016), .A(n13915), .ZN(P1_U2996) );
  XOR2_X1 U17342 ( .A(n13917), .B(n13916), .Z(n13939) );
  OAI21_X1 U17343 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14943), .A(
        n13918), .ZN(n13920) );
  XNOR2_X1 U17344 ( .A(n13920), .B(n13919), .ZN(n13936) );
  INV_X1 U17345 ( .A(n14940), .ZN(n13923) );
  INV_X1 U17346 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14945) );
  OAI22_X1 U17347 ( .A1(n19312), .A2(n14945), .B1(n13921), .B2(n19091), .ZN(
        n13922) );
  AOI21_X1 U17348 ( .B1(n19290), .B2(n13923), .A(n13922), .ZN(n13925) );
  NAND2_X1 U17349 ( .A1(n14948), .A2(n19319), .ZN(n13924) );
  OAI211_X1 U17350 ( .C1(n13936), .C2(n19297), .A(n13925), .B(n13924), .ZN(
        n13926) );
  AOI21_X1 U17351 ( .B1(n13939), .B2(n16265), .A(n13926), .ZN(n13927) );
  INV_X1 U17352 ( .A(n13927), .ZN(P2_U3011) );
  NOR2_X1 U17353 ( .A1(n13929), .A2(n13928), .ZN(n13938) );
  INV_X1 U17354 ( .A(n13930), .ZN(n13933) );
  XNOR2_X1 U17355 ( .A(n13931), .B(n9657), .ZN(n19198) );
  INV_X1 U17356 ( .A(n19198), .ZN(n19945) );
  OAI22_X1 U17357 ( .A1(n19330), .A2(n19945), .B1(n13921), .B2(n19091), .ZN(
        n13932) );
  AOI21_X1 U17358 ( .B1(n13933), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13932), .ZN(n13935) );
  NAND2_X1 U17359 ( .A1(n14948), .A2(n19338), .ZN(n13934) );
  OAI211_X1 U17360 ( .C1(n13936), .C2(n19331), .A(n13935), .B(n13934), .ZN(
        n13937) );
  AOI211_X1 U17361 ( .C1(n13939), .C2(n16329), .A(n13938), .B(n13937), .ZN(
        n13940) );
  INV_X1 U17362 ( .A(n13940), .ZN(P2_U3043) );
  NAND2_X1 U17363 ( .A1(n13942), .A2(n13941), .ZN(n13943) );
  AND2_X1 U17364 ( .A1(n16087), .A2(n13943), .ZN(n20208) );
  INV_X1 U17365 ( .A(n20208), .ZN(n20065) );
  INV_X1 U17366 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21105) );
  XOR2_X1 U17367 ( .A(n13874), .B(n13944), .Z(n20188) );
  INV_X1 U17368 ( .A(n20188), .ZN(n14000) );
  OAI222_X1 U17369 ( .A1(n14557), .A2(n20065), .B1(n20116), .B2(n21105), .C1(
        n14568), .C2(n14000), .ZN(P1_U2868) );
  XNOR2_X1 U17370 ( .A(n13945), .B(n14064), .ZN(n13950) );
  OR2_X1 U17371 ( .A1(n13991), .A2(n13946), .ZN(n13947) );
  NAND2_X1 U17372 ( .A1(n13947), .A2(n14061), .ZN(n19054) );
  MUX2_X1 U17373 ( .A(n19054), .B(n13948), .S(n15042), .Z(n13949) );
  OAI21_X1 U17374 ( .B1(n13950), .B2(n15044), .A(n13949), .ZN(P2_U2876) );
  NOR2_X1 U17375 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16108), .ZN(n13966) );
  MUX2_X1 U17376 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13951), .S(
        n13973), .Z(n15746) );
  AOI22_X1 U17377 ( .A1(n13966), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16108), .B2(n15746), .ZN(n13968) );
  NOR2_X1 U17378 ( .A1(n13952), .A2(n13956), .ZN(n13953) );
  NOR2_X1 U17379 ( .A1(n12175), .A2(n13953), .ZN(n14935) );
  XNOR2_X1 U17380 ( .A(n13954), .B(n13956), .ZN(n13955) );
  NAND2_X1 U17381 ( .A1(n15750), .A2(n13955), .ZN(n13962) );
  MUX2_X1 U17382 ( .A(n13957), .B(n13956), .S(n13707), .Z(n13959) );
  OAI21_X1 U17383 ( .B1(n13960), .B2(n13959), .A(n13958), .ZN(n13961) );
  OAI211_X1 U17384 ( .C1(n14935), .C2(n13963), .A(n13962), .B(n13961), .ZN(
        n13964) );
  AOI21_X1 U17385 ( .B1(n20536), .B2(n14924), .A(n13964), .ZN(n14937) );
  INV_X1 U17386 ( .A(n14937), .ZN(n13965) );
  MUX2_X1 U17387 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13965), .S(
        n13973), .Z(n15758) );
  AOI22_X1 U17388 ( .A1(n13966), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n15758), .B2(n16108), .ZN(n13967) );
  NOR2_X1 U17389 ( .A1(n13968), .A2(n13967), .ZN(n15767) );
  INV_X1 U17390 ( .A(n15767), .ZN(n13969) );
  NOR2_X1 U17391 ( .A1(n13969), .A2(n14918), .ZN(n13995) );
  INV_X1 U17392 ( .A(n20415), .ZN(n20668) );
  NOR2_X1 U17393 ( .A1(n13970), .A2(n20668), .ZN(n13971) );
  XOR2_X1 U17394 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n13971), .Z(
        n20069) );
  INV_X1 U17395 ( .A(n13699), .ZN(n13972) );
  NAND2_X1 U17396 ( .A1(n20069), .A2(n13972), .ZN(n16095) );
  NAND2_X1 U17397 ( .A1(n13973), .A2(n16108), .ZN(n13974) );
  INV_X1 U17398 ( .A(n13974), .ZN(n13977) );
  NAND2_X1 U17399 ( .A1(n13974), .A2(n16100), .ZN(n13975) );
  OAI21_X1 U17400 ( .B1(n16108), .B2(n20017), .A(n13975), .ZN(n13976) );
  AOI21_X1 U17401 ( .B1(n16095), .B2(n13977), .A(n13976), .ZN(n15766) );
  INV_X1 U17402 ( .A(n16111), .ZN(n13978) );
  AOI21_X1 U17403 ( .B1(n16108), .B2(n20780), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n20931) );
  NAND2_X1 U17404 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20671), .ZN(n13996) );
  INV_X1 U17405 ( .A(n20338), .ZN(n14911) );
  NAND2_X1 U17406 ( .A1(n20791), .A2(n20418), .ZN(n20666) );
  NOR3_X1 U17407 ( .A1(n20338), .A2(n20782), .A3(n20418), .ZN(n13981) );
  MUX2_X1 U17408 ( .A(n20787), .B(n13981), .S(n13980), .Z(n13982) );
  AOI21_X1 U17409 ( .B1(n13996), .B2(n20265), .A(n13982), .ZN(n13984) );
  NAND2_X1 U17410 ( .A1(n20255), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13983) );
  OAI21_X1 U17411 ( .B1(n20255), .B2(n13984), .A(n13983), .ZN(P1_U3476) );
  NOR2_X1 U17412 ( .A1(n13893), .A2(n13985), .ZN(n13988) );
  INV_X1 U17413 ( .A(n13945), .ZN(n13986) );
  OAI211_X1 U17414 ( .C1(n13988), .C2(n13987), .A(n13986), .B(n15029), .ZN(
        n13993) );
  NOR2_X1 U17415 ( .A1(n9705), .A2(n13989), .ZN(n13990) );
  OR2_X1 U17416 ( .A1(n13991), .A2(n13990), .ZN(n19068) );
  INV_X1 U17417 ( .A(n19068), .ZN(n16281) );
  NAND2_X1 U17418 ( .A1(n16281), .A2(n15036), .ZN(n13992) );
  OAI211_X1 U17419 ( .C1(n15036), .C2(n13994), .A(n13993), .B(n13992), .ZN(
        P2_U2877) );
  INV_X1 U17420 ( .A(n20255), .ZN(n13999) );
  NOR3_X1 U17421 ( .A1(n13995), .A2(n15766), .A3(n16106), .ZN(n15773) );
  INV_X1 U17422 ( .A(n13996), .ZN(n14913) );
  OAI22_X1 U17423 ( .A1(n12353), .A2(n20782), .B1(n11556), .B2(n14913), .ZN(
        n13997) );
  OAI21_X1 U17424 ( .B1(n15773), .B2(n13997), .A(n13999), .ZN(n13998) );
  OAI21_X1 U17425 ( .B1(n13999), .B2(n20701), .A(n13998), .ZN(P1_U3478) );
  INV_X1 U17426 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20133) );
  OAI222_X1 U17427 ( .A1(n14645), .A2(n20292), .B1(n14647), .B2(n14000), .C1(
        n14637), .C2(n20133), .ZN(P1_U2900) );
  NAND2_X1 U17428 ( .A1(n14003), .A2(n14002), .ZN(n14004) );
  AND2_X1 U17429 ( .A1(n14001), .A2(n14004), .ZN(n20041) );
  INV_X1 U17430 ( .A(n20041), .ZN(n14024) );
  OR2_X1 U17431 ( .A1(n9719), .A2(n14005), .ZN(n14006) );
  AND2_X1 U17432 ( .A1(n14078), .A2(n14006), .ZN(n20037) );
  AOI22_X1 U17433 ( .A1(n20037), .A2(n20111), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14566), .ZN(n14007) );
  OAI21_X1 U17434 ( .B1(n14024), .B2(n14568), .A(n14007), .ZN(P1_U2865) );
  NAND2_X1 U17435 ( .A1(n19947), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19722) );
  NAND2_X1 U17436 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19957), .ZN(
        n19633) );
  INV_X1 U17437 ( .A(n19633), .ZN(n14008) );
  NAND2_X1 U17438 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n14008), .ZN(
        n14018) );
  OAI21_X1 U17439 ( .B1(n19722), .B2(n19939), .A(n14018), .ZN(n14016) );
  NAND2_X1 U17440 ( .A1(n19537), .A2(n14008), .ZN(n14009) );
  INV_X1 U17441 ( .A(n14009), .ZN(n19675) );
  AND2_X1 U17442 ( .A1(n14009), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14010) );
  NAND2_X1 U17443 ( .A1(n14011), .A2(n14010), .ZN(n14020) );
  AOI21_X1 U17444 ( .B1(n19777), .B2(n15803), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19992) );
  NAND2_X1 U17445 ( .A1(n19992), .A2(n16402), .ZN(n14012) );
  OAI211_X1 U17446 ( .C1(n19950), .C2(n19675), .A(n14020), .B(n19788), .ZN(
        n14014) );
  INV_X1 U17447 ( .A(n14014), .ZN(n14015) );
  INV_X1 U17448 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16503) );
  INV_X1 U17449 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18265) );
  OAI22_X1 U17450 ( .A1(n16503), .A2(n19368), .B1(n18265), .B2(n19366), .ZN(
        n19790) );
  NAND2_X1 U17451 ( .A1(n19682), .A2(n19430), .ZN(n19671) );
  AOI22_X1 U17452 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19361), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19362), .ZN(n19793) );
  AOI22_X1 U17453 ( .A1(n19707), .A2(n19790), .B1(n19677), .B2(n19695), .ZN(
        n14022) );
  NOR2_X2 U17454 ( .A1(n19265), .A2(n19601), .ZN(n19782) );
  OAI21_X1 U17455 ( .B1(n14018), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19777), 
        .ZN(n14019) );
  AND2_X1 U17456 ( .A1(n14020), .A2(n14019), .ZN(n19676) );
  NAND2_X1 U17457 ( .A1(n19996), .A2(n19352), .ZN(n15582) );
  AOI22_X1 U17458 ( .A1(n19782), .A2(n19676), .B1(n19781), .B2(n19675), .ZN(
        n14021) );
  OAI211_X1 U17459 ( .C1(n19674), .C2(n14023), .A(n14022), .B(n14021), .ZN(
        P2_U3136) );
  OAI222_X1 U17460 ( .A1(n14647), .A2(n14024), .B1(n14637), .B2(n11707), .C1(
        n14645), .C2(n20309), .ZN(P1_U2897) );
  XNOR2_X1 U17461 ( .A(n14025), .B(n14084), .ZN(n14028) );
  OAI21_X1 U17462 ( .B1(n14026), .B2(n14060), .A(n14088), .ZN(n19033) );
  MUX2_X1 U17463 ( .A(n10870), .B(n19033), .S(n15036), .Z(n14027) );
  OAI21_X1 U17464 ( .B1(n14028), .B2(n15044), .A(n14027), .ZN(P2_U2874) );
  INV_X1 U17465 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16485) );
  INV_X1 U17466 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17310) );
  OAI22_X2 U17467 ( .A1(n16485), .A2(n19368), .B1(n17310), .B2(n19366), .ZN(
        n19763) );
  AOI22_X1 U17468 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19361), .ZN(n19710) );
  INV_X1 U17469 ( .A(n19710), .ZN(n19822) );
  AOI22_X1 U17470 ( .A1(n19677), .A2(n19763), .B1(n19707), .B2(n19822), .ZN(
        n14031) );
  AOI22_X1 U17471 ( .A1(n19167), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19166), .ZN(n19271) );
  NOR2_X2 U17472 ( .A1(n19271), .A2(n19601), .ZN(n19821) );
  AOI22_X1 U17473 ( .A1(n19676), .A2(n19821), .B1(n19675), .B2(n19820), .ZN(
        n14030) );
  OAI211_X1 U17474 ( .C1(n19674), .C2(n14032), .A(n14031), .B(n14030), .ZN(
        P2_U3141) );
  NOR2_X1 U17475 ( .A1(n14033), .A2(n14035), .ZN(n14034) );
  NOR2_X1 U17476 ( .A1(n20052), .A2(n14034), .ZN(n20109) );
  OAI21_X1 U17477 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20071), .A(n20092), .ZN(
        n20077) );
  INV_X1 U17478 ( .A(n20536), .ZN(n14914) );
  NOR2_X1 U17479 ( .A1(n14036), .A2(n14035), .ZN(n20104) );
  INV_X1 U17480 ( .A(n20104), .ZN(n14042) );
  INV_X1 U17481 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20243) );
  NOR2_X1 U17482 ( .A1(n20071), .A2(n20243), .ZN(n20079) );
  INV_X1 U17483 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14038) );
  INV_X1 U17484 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20078) );
  AND2_X1 U17485 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n14037) );
  AOI21_X1 U17486 ( .B1(n14038), .B2(n20078), .A(n14037), .ZN(n14039) );
  AOI22_X1 U17487 ( .A1(n20079), .A2(n14039), .B1(n20103), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14041) );
  NAND2_X1 U17488 ( .A1(n20214), .A2(n20099), .ZN(n14040) );
  OAI211_X1 U17489 ( .C1(n14914), .C2(n14042), .A(n14041), .B(n14040), .ZN(
        n14048) );
  AND2_X1 U17490 ( .A1(n14043), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14044) );
  OAI22_X1 U17491 ( .A1(n14046), .A2(n20101), .B1(n20102), .B2(n14045), .ZN(
        n14047) );
  AOI211_X1 U17492 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n20077), .A(n14048), .B(
        n14047), .ZN(n14049) );
  OAI21_X1 U17493 ( .B1(n20109), .B2(n14050), .A(n14049), .ZN(P1_U2837) );
  INV_X1 U17494 ( .A(n19955), .ZN(n14052) );
  AOI21_X1 U17495 ( .B1(n19951), .B2(n14052), .A(n14051), .ZN(n19200) );
  XNOR2_X1 U17496 ( .A(n19947), .B(n19198), .ZN(n19201) );
  NOR2_X1 U17497 ( .A1(n19200), .A2(n19201), .ZN(n19199) );
  NOR2_X1 U17498 ( .A1(n19947), .A2(n19198), .ZN(n14055) );
  XNOR2_X1 U17499 ( .A(n14054), .B(n14053), .ZN(n19329) );
  OAI21_X1 U17500 ( .B1(n19199), .B2(n14055), .A(n19329), .ZN(n19193) );
  XOR2_X1 U17501 ( .A(n19131), .B(n19193), .Z(n14059) );
  INV_X1 U17502 ( .A(n19329), .ZN(n14056) );
  AOI22_X1 U17503 ( .A1(n19206), .A2(n14056), .B1(n19205), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n14058) );
  INV_X1 U17504 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16519) );
  INV_X1 U17505 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18280) );
  AOI22_X1 U17506 ( .A1(n19167), .A2(n16519), .B1(n18280), .B2(n19166), .ZN(
        n19255) );
  NAND2_X1 U17507 ( .A1(n19189), .A2(n19255), .ZN(n14057) );
  OAI211_X1 U17508 ( .C1(n14059), .C2(n19210), .A(n14058), .B(n14057), .ZN(
        P2_U2915) );
  AOI21_X1 U17509 ( .B1(n14062), .B2(n14061), .A(n14060), .ZN(n19045) );
  INV_X1 U17510 ( .A(n19045), .ZN(n15243) );
  AOI21_X1 U17511 ( .B1(n13945), .B2(n14064), .A(n14063), .ZN(n14065) );
  OR3_X1 U17512 ( .A1(n14025), .A2(n14065), .A3(n15044), .ZN(n14067) );
  NAND2_X1 U17513 ( .A1(n15042), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14066) );
  OAI211_X1 U17514 ( .C1(n15243), .C2(n15042), .A(n14067), .B(n14066), .ZN(
        P2_U2875) );
  XOR2_X1 U17515 ( .A(n13907), .B(n14068), .Z(n20051) );
  INV_X1 U17516 ( .A(n20051), .ZN(n14073) );
  OAI222_X1 U17517 ( .A1(n14645), .A2(n20301), .B1(n14647), .B2(n14073), .C1(
        n14069), .C2(n14637), .ZN(P1_U2898) );
  NOR2_X1 U17518 ( .A1(n14070), .A2(n14071), .ZN(n14072) );
  OR2_X1 U17519 ( .A1(n9719), .A2(n14072), .ZN(n20047) );
  INV_X1 U17520 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14074) );
  OAI222_X1 U17521 ( .A1(n20047), .A2(n14557), .B1(n14074), .B2(n20116), .C1(
        n14568), .C2(n14073), .ZN(P1_U2866) );
  NAND2_X1 U17522 ( .A1(n14001), .A2(n14076), .ZN(n14077) );
  AND2_X1 U17523 ( .A1(n14157), .A2(n14077), .ZN(n14241) );
  INV_X1 U17524 ( .A(n14241), .ZN(n14083) );
  INV_X1 U17525 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14097) );
  INV_X1 U17526 ( .A(n14078), .ZN(n14079) );
  OAI21_X1 U17527 ( .B1(n14079), .B2(n10084), .A(n14162), .ZN(n16068) );
  OAI222_X1 U17528 ( .A1(n14083), .A2(n14568), .B1(n20116), .B2(n14097), .C1(
        n16068), .C2(n14557), .ZN(P1_U2864) );
  INV_X1 U17529 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14082) );
  NAND2_X1 U17530 ( .A1(n20257), .A2(DATAI_8_), .ZN(n14081) );
  NAND2_X1 U17531 ( .A1(n20256), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14080) );
  AND2_X1 U17532 ( .A1(n14081), .A2(n14080), .ZN(n20145) );
  OAI222_X1 U17533 ( .A1(n14083), .A2(n14647), .B1(n14082), .B2(n14637), .C1(
        n14645), .C2(n20145), .ZN(P1_U2896) );
  AND2_X1 U17534 ( .A1(n14025), .A2(n14084), .ZN(n14087) );
  OAI211_X1 U17535 ( .C1(n14087), .C2(n14086), .A(n15029), .B(n14085), .ZN(
        n14093) );
  NAND2_X1 U17536 ( .A1(n14089), .A2(n14088), .ZN(n14091) );
  INV_X1 U17537 ( .A(n14185), .ZN(n14090) );
  AND2_X1 U17538 ( .A1(n14091), .A2(n14090), .ZN(n19024) );
  NAND2_X1 U17539 ( .A1(n19024), .A2(n15036), .ZN(n14092) );
  OAI211_X1 U17540 ( .C1(n15036), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        P2_U2873) );
  INV_X1 U17541 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14095) );
  NAND3_X1 U17542 ( .A1(n20090), .A2(n14177), .A3(n14095), .ZN(n14096) );
  OAI211_X1 U17543 ( .C1(n20034), .C2(n14097), .A(n20244), .B(n14096), .ZN(
        n14098) );
  AOI21_X1 U17544 ( .B1(n20095), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n14098), .ZN(n14099) );
  OAI21_X1 U17545 ( .B1(n20101), .B2(n14239), .A(n14099), .ZN(n14102) );
  INV_X1 U17546 ( .A(n20092), .ZN(n20033) );
  NAND2_X1 U17547 ( .A1(n20100), .A2(n14423), .ZN(n14182) );
  OAI22_X1 U17548 ( .A1(n20088), .A2(n16068), .B1(n14095), .B2(n14182), .ZN(
        n14101) );
  AOI211_X1 U17549 ( .C1(n14241), .C2(n20052), .A(n14102), .B(n14101), .ZN(
        n14103) );
  INV_X1 U17550 ( .A(n14103), .ZN(P1_U2832) );
  NAND2_X1 U17551 ( .A1(n14104), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19542) );
  OAI21_X1 U17552 ( .B1(n19542), .B2(n15577), .A(n19938), .ZN(n14118) );
  NOR2_X1 U17553 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19957), .ZN(
        n19536) );
  NAND2_X1 U17554 ( .A1(n19536), .A2(n10498), .ZN(n14117) );
  INV_X1 U17555 ( .A(n14117), .ZN(n14105) );
  OR2_X1 U17556 ( .A1(n14118), .A2(n14105), .ZN(n14109) );
  NAND2_X1 U17557 ( .A1(n14114), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14106) );
  NAND2_X1 U17558 ( .A1(n14106), .A2(n19950), .ZN(n14107) );
  NOR2_X1 U17559 ( .A1(n19973), .A2(n14117), .ZN(n19510) );
  INV_X1 U17560 ( .A(n19510), .ZN(n14112) );
  AOI21_X1 U17561 ( .B1(n14107), .B2(n14112), .A(n19601), .ZN(n14108) );
  INV_X1 U17562 ( .A(n19548), .ZN(n14111) );
  INV_X1 U17563 ( .A(n19790), .ZN(n19698) );
  OAI22_X1 U17564 ( .A1(n19520), .A2(n19698), .B1(n15582), .B2(n14112), .ZN(
        n14113) );
  AOI21_X1 U17565 ( .B1(n19695), .B2(n19511), .A(n14113), .ZN(n14120) );
  INV_X1 U17566 ( .A(n14114), .ZN(n14115) );
  OAI21_X1 U17567 ( .B1(n14115), .B2(n19510), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14116) );
  OAI21_X1 U17568 ( .B1(n14118), .B2(n14117), .A(n14116), .ZN(n19512) );
  NAND2_X1 U17569 ( .A1(n19512), .A2(n19782), .ZN(n14119) );
  OAI211_X1 U17570 ( .C1(n19515), .C2(n14121), .A(n14120), .B(n14119), .ZN(
        P2_U3088) );
  INV_X1 U17571 ( .A(n14122), .ZN(n19303) );
  NAND2_X1 U17572 ( .A1(n9704), .A2(n14959), .ZN(n14123) );
  XOR2_X1 U17573 ( .A(n19303), .B(n14123), .Z(n14132) );
  INV_X1 U17574 ( .A(n19847), .ZN(n19123) );
  OAI22_X1 U17575 ( .A1(n10267), .A2(n19142), .B1(n14124), .B2(n19149), .ZN(
        n14126) );
  OAI22_X1 U17576 ( .A1(n19951), .A2(n19144), .B1(n19311), .B2(n19139), .ZN(
        n14125) );
  AOI211_X1 U17577 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n19146), .A(n14126), .B(
        n14125), .ZN(n14130) );
  NAND2_X1 U17578 ( .A1(n19955), .A2(n19141), .ZN(n14129) );
  NAND2_X1 U17579 ( .A1(n14127), .A2(n19151), .ZN(n14128) );
  NAND3_X1 U17580 ( .A1(n14130), .A2(n14129), .A3(n14128), .ZN(n14131) );
  AOI21_X1 U17581 ( .B1(n14132), .B2(n19123), .A(n14131), .ZN(n14133) );
  INV_X1 U17582 ( .A(n14133), .ZN(P2_U2853) );
  XNOR2_X1 U17583 ( .A(n14134), .B(n14135), .ZN(n14156) );
  INV_X1 U17584 ( .A(n10812), .ZN(n14140) );
  AOI21_X1 U17585 ( .B1(n14139), .B2(n14137), .A(n14136), .ZN(n14138) );
  AOI21_X1 U17586 ( .B1(n14140), .B2(n14139), .A(n14138), .ZN(n14154) );
  OAI21_X1 U17587 ( .B1(n14143), .B2(n14142), .A(n14141), .ZN(n19196) );
  OAI211_X1 U17588 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n19336), .B(n14144), .ZN(n14148) );
  INV_X1 U17589 ( .A(n14145), .ZN(n19337) );
  NAND2_X1 U17590 ( .A1(n19291), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n14151) );
  OAI21_X1 U17591 ( .B1(n16341), .B2(n19120), .A(n14151), .ZN(n14146) );
  AOI21_X1 U17592 ( .B1(n19337), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n14146), .ZN(n14147) );
  OAI211_X1 U17593 ( .C1(n19196), .C2(n19330), .A(n14148), .B(n14147), .ZN(
        n14149) );
  AOI21_X1 U17594 ( .B1(n14154), .B2(n16329), .A(n14149), .ZN(n14150) );
  OAI21_X1 U17595 ( .B1(n19331), .B2(n14156), .A(n14150), .ZN(P2_U3041) );
  OAI22_X1 U17596 ( .A1(n9975), .A2(n19312), .B1(n19304), .B2(n19119), .ZN(
        n14153) );
  OAI21_X1 U17597 ( .B1(n19305), .B2(n19120), .A(n14151), .ZN(n14152) );
  AOI211_X1 U17598 ( .C1(n14154), .C2(n16265), .A(n14153), .B(n14152), .ZN(
        n14155) );
  OAI21_X1 U17599 ( .B1(n19297), .B2(n14156), .A(n14155), .ZN(P2_U3009) );
  INV_X1 U17600 ( .A(n14158), .ZN(n14160) );
  INV_X1 U17601 ( .A(n14159), .ZN(n14213) );
  OAI21_X1 U17602 ( .B1(n14075), .B2(n14160), .A(n14213), .ZN(n14777) );
  INV_X1 U17603 ( .A(n14216), .ZN(n14161) );
  AOI21_X1 U17604 ( .B1(n14163), .B2(n14162), .A(n14161), .ZN(n16054) );
  AOI22_X1 U17605 ( .A1(n16054), .A2(n20111), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14566), .ZN(n14164) );
  OAI21_X1 U17606 ( .B1(n14777), .B2(n14568), .A(n14164), .ZN(P1_U2863) );
  INV_X1 U17607 ( .A(n14165), .ZN(n15524) );
  OR2_X1 U17608 ( .A1(n14166), .A2(n15524), .ZN(n14171) );
  INV_X1 U17609 ( .A(n15503), .ZN(n15518) );
  AND2_X1 U17610 ( .A1(n14168), .A2(n14167), .ZN(n15501) );
  MUX2_X1 U17611 ( .A(n15518), .B(n15501), .S(n14169), .Z(n14170) );
  NAND2_X1 U17612 ( .A1(n14171), .A2(n14170), .ZN(n16366) );
  INV_X1 U17613 ( .A(n14961), .ZN(n14172) );
  AOI22_X1 U17614 ( .A1(n9963), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n14172), .B2(n9704), .ZN(n15509) );
  AOI222_X1 U17615 ( .A1(n16366), .A2(n19940), .B1(n14173), .B2(n15525), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15509), .ZN(n14176) );
  NAND2_X1 U17616 ( .A1(n15696), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14175) );
  OAI21_X1 U17617 ( .B1(n14176), .B2(n15696), .A(n14175), .ZN(P2_U3601) );
  NAND3_X1 U17618 ( .A1(n20090), .A2(P1_REIP_REG_8__SCAN_IN), .A3(n14177), 
        .ZN(n14432) );
  INV_X1 U17619 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20870) );
  OAI22_X1 U17620 ( .A1(n20102), .A2(n14179), .B1(n14178), .B2(n20034), .ZN(
        n14180) );
  AOI211_X1 U17621 ( .C1(n16054), .C2(n20099), .A(n20209), .B(n14180), .ZN(
        n14181) );
  OAI221_X1 U17622 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n14432), .C1(n20870), 
        .C2(n14182), .A(n14181), .ZN(n14183) );
  AOI21_X1 U17623 ( .B1(n14774), .B2(n15877), .A(n14183), .ZN(n14184) );
  OAI21_X1 U17624 ( .B1(n15859), .B2(n14777), .A(n14184), .ZN(P1_U2831) );
  XNOR2_X1 U17625 ( .A(n14085), .B(n14204), .ZN(n14188) );
  OAI21_X1 U17626 ( .B1(n14186), .B2(n14185), .A(n14208), .ZN(n19013) );
  MUX2_X1 U17627 ( .A(n10877), .B(n19013), .S(n15036), .Z(n14187) );
  OAI21_X1 U17628 ( .B1(n14188), .B2(n15044), .A(n14187), .ZN(P2_U2872) );
  INV_X1 U17629 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14190) );
  INV_X1 U17630 ( .A(DATAI_9_), .ZN(n14189) );
  INV_X1 U17631 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n15075) );
  MUX2_X1 U17632 ( .A(n14189), .B(n15075), .S(n20256), .Z(n20148) );
  OAI222_X1 U17633 ( .A1(n14777), .A2(n14647), .B1(n14190), .B2(n14637), .C1(
        n14645), .C2(n20148), .ZN(P1_U2895) );
  NOR2_X1 U17634 ( .A1(n14085), .A2(n14204), .ZN(n14192) );
  AND2_X1 U17635 ( .A1(n14192), .A2(n14191), .ZN(n14205) );
  OR2_X1 U17636 ( .A1(n14085), .A2(n14193), .ZN(n14277) );
  OAI21_X1 U17637 ( .B1(n14205), .B2(n14194), .A(n14277), .ZN(n14234) );
  OR2_X1 U17638 ( .A1(n14196), .A2(n14195), .ZN(n14197) );
  AND2_X1 U17639 ( .A1(n14197), .A2(n15412), .ZN(n18989) );
  AOI22_X1 U17640 ( .A1(n19167), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19166), .ZN(n19349) );
  OAI22_X1 U17641 ( .A1(n16196), .A2(n19349), .B1(n19187), .B2(n14198), .ZN(
        n14202) );
  INV_X1 U17642 ( .A(n19160), .ZN(n15112) );
  INV_X1 U17643 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14200) );
  INV_X1 U17644 ( .A(n19159), .ZN(n15110) );
  INV_X1 U17645 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14199) );
  OAI22_X1 U17646 ( .A1(n15112), .A2(n14200), .B1(n15110), .B2(n14199), .ZN(
        n14201) );
  AOI211_X1 U17647 ( .C1(n19206), .C2(n18989), .A(n14202), .B(n14201), .ZN(
        n14203) );
  OAI21_X1 U17648 ( .B1(n14234), .B2(n19210), .A(n14203), .ZN(P2_U2902) );
  OR2_X1 U17649 ( .A1(n14085), .A2(n14204), .ZN(n14206) );
  AOI21_X1 U17650 ( .B1(n14207), .B2(n14206), .A(n14205), .ZN(n19162) );
  NAND2_X1 U17651 ( .A1(n19162), .A2(n15029), .ZN(n14211) );
  AOI21_X1 U17652 ( .B1(n14209), .B2(n14208), .A(n14229), .ZN(n19003) );
  NAND2_X1 U17653 ( .A1(n19003), .A2(n15036), .ZN(n14210) );
  OAI211_X1 U17654 ( .C1(n15036), .C2(n10879), .A(n14211), .B(n14210), .ZN(
        P2_U2871) );
  INV_X1 U17655 ( .A(n14212), .ZN(n14214) );
  AOI21_X1 U17656 ( .B1(n14214), .B2(n14213), .A(n9642), .ZN(n14769) );
  INV_X1 U17657 ( .A(n14769), .ZN(n14227) );
  NOR2_X1 U17658 ( .A1(n14433), .A2(n14423), .ZN(n14487) );
  NOR2_X1 U17659 ( .A1(n14486), .A2(n14487), .ZN(n15885) );
  NOR2_X1 U17660 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14432), .ZN(n14215) );
  AOI22_X1 U17661 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15885), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n14215), .ZN(n14222) );
  INV_X1 U17662 ( .A(n14767), .ZN(n14220) );
  AOI21_X1 U17663 ( .B1(n14217), .B2(n14216), .A(n15884), .ZN(n16049) );
  INV_X1 U17664 ( .A(n16049), .ZN(n14223) );
  AOI22_X1 U17665 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n20103), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20095), .ZN(n14218) );
  OAI21_X1 U17666 ( .B1(n20088), .B2(n14223), .A(n14218), .ZN(n14219) );
  AOI211_X1 U17667 ( .C1(n15877), .C2(n14220), .A(n20209), .B(n14219), .ZN(
        n14221) );
  OAI211_X1 U17668 ( .C1(n14227), .C2(n15859), .A(n14222), .B(n14221), .ZN(
        P1_U2830) );
  INV_X1 U17669 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14224) );
  OAI222_X1 U17670 ( .A1(n14227), .A2(n14568), .B1(n20116), .B2(n14224), .C1(
        n14223), .C2(n14557), .ZN(P1_U2862) );
  INV_X1 U17671 ( .A(DATAI_10_), .ZN(n14225) );
  MUX2_X1 U17672 ( .A(n14225), .B(n16510), .S(n20256), .Z(n20152) );
  INV_X1 U17673 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14226) );
  OAI222_X1 U17674 ( .A1(n14647), .A2(n14227), .B1(n14645), .B2(n20152), .C1(
        n14226), .C2(n14637), .ZN(P1_U2894) );
  NAND2_X1 U17675 ( .A1(n15042), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14233) );
  INV_X1 U17676 ( .A(n14228), .ZN(n14231) );
  INV_X1 U17677 ( .A(n14229), .ZN(n14230) );
  AOI21_X1 U17678 ( .B1(n14231), .B2(n14230), .A(n14273), .ZN(n18988) );
  NAND2_X1 U17679 ( .A1(n18988), .A2(n15036), .ZN(n14232) );
  OAI211_X1 U17680 ( .C1(n14234), .C2(n15044), .A(n14233), .B(n14232), .ZN(
        P2_U2870) );
  XOR2_X1 U17681 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14236), .Z(
        n14237) );
  XNOR2_X1 U17682 ( .A(n14235), .B(n14237), .ZN(n16067) );
  AOI22_X1 U17683 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14238) );
  OAI21_X1 U17684 ( .B1(n20193), .B2(n14239), .A(n14238), .ZN(n14240) );
  AOI21_X1 U17685 ( .B1(n14241), .B2(n20189), .A(n14240), .ZN(n14242) );
  OAI21_X1 U17686 ( .B1(n16067), .B2(n20016), .A(n14242), .ZN(P1_U2991) );
  XNOR2_X1 U17687 ( .A(n14243), .B(n14244), .ZN(n14263) );
  OAI21_X1 U17688 ( .B1(n14246), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14245), .ZN(n14247) );
  INV_X1 U17689 ( .A(n14247), .ZN(n14261) );
  NOR2_X1 U17690 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14248), .ZN(
        n16323) );
  XNOR2_X1 U17691 ( .A(n14250), .B(n14249), .ZN(n19188) );
  INV_X1 U17692 ( .A(n19188), .ZN(n14251) );
  NAND2_X1 U17693 ( .A1(n14251), .A2(n16350), .ZN(n14253) );
  AOI22_X1 U17694 ( .A1(n19111), .A2(n19338), .B1(n19291), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n14252) );
  OAI211_X1 U17695 ( .C1(n14254), .C2(n16321), .A(n14253), .B(n14252), .ZN(
        n14255) );
  AOI211_X1 U17696 ( .C1(n14261), .C2(n16329), .A(n16323), .B(n14255), .ZN(
        n14256) );
  OAI21_X1 U17697 ( .B1(n19331), .B2(n14263), .A(n14256), .ZN(P2_U3040) );
  INV_X1 U17698 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19880) );
  OAI22_X1 U17699 ( .A1(n19104), .A2(n19312), .B1(n19880), .B2(n19328), .ZN(
        n14260) );
  INV_X1 U17700 ( .A(n19111), .ZN(n14258) );
  INV_X1 U17701 ( .A(n19109), .ZN(n14257) );
  OAI22_X1 U17702 ( .A1(n14258), .A2(n19305), .B1(n19304), .B2(n14257), .ZN(
        n14259) );
  AOI211_X1 U17703 ( .C1(n14261), .C2(n16265), .A(n14260), .B(n14259), .ZN(
        n14262) );
  OAI21_X1 U17704 ( .B1(n19297), .B2(n14263), .A(n14262), .ZN(P2_U3008) );
  XOR2_X1 U17705 ( .A(n16337), .B(n14265), .Z(n14266) );
  XNOR2_X1 U17706 ( .A(n14264), .B(n14266), .ZN(n16347) );
  NAND2_X1 U17707 ( .A1(n15259), .A2(n15257), .ZN(n14268) );
  XNOR2_X1 U17708 ( .A(n14267), .B(n14268), .ZN(n16345) );
  INV_X1 U17709 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19882) );
  OAI22_X1 U17710 ( .A1(n19882), .A2(n19328), .B1(n19304), .B2(n19095), .ZN(
        n14270) );
  OAI22_X1 U17711 ( .A1(n19102), .A2(n19305), .B1(n19312), .B2(n9976), .ZN(
        n14269) );
  AOI211_X1 U17712 ( .C1(n16345), .C2(n19318), .A(n14270), .B(n14269), .ZN(
        n14271) );
  OAI21_X1 U17713 ( .B1(n16347), .B2(n19323), .A(n14271), .ZN(P2_U3007) );
  NOR2_X1 U17714 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  NOR2_X1 U17715 ( .A1(n14272), .A2(n14275), .ZN(n18977) );
  INV_X1 U17716 ( .A(n18977), .ZN(n14281) );
  AOI21_X1 U17717 ( .B1(n14278), .B2(n14277), .A(n14276), .ZN(n16212) );
  NAND2_X1 U17718 ( .A1(n16212), .A2(n15029), .ZN(n14280) );
  NAND2_X1 U17719 ( .A1(n15042), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14279) );
  OAI211_X1 U17720 ( .C1(n14281), .C2(n15042), .A(n14280), .B(n14279), .ZN(
        P2_U2869) );
  INV_X1 U17721 ( .A(n18911), .ZN(n18851) );
  OAI21_X1 U17722 ( .B1(n14282), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n14287), .ZN(n18739) );
  NOR2_X1 U17723 ( .A1(n18851), .A2(n18739), .ZN(n14292) );
  AOI211_X1 U17724 ( .C1(n16578), .C2(n14285), .A(n14284), .B(n14283), .ZN(
        n15706) );
  OR2_X1 U17725 ( .A1(n18268), .A2(n17512), .ZN(n18746) );
  NOR2_X1 U17726 ( .A1(n18895), .A2(n16576), .ZN(n15807) );
  INV_X1 U17727 ( .A(n18692), .ZN(n14289) );
  AOI221_X1 U17728 ( .B1(n17449), .B2(n15807), .C1(n15806), .C2(n15807), .A(
        n15593), .ZN(n14290) );
  NAND2_X1 U17729 ( .A1(n15706), .A2(n14290), .ZN(n18732) );
  NAND2_X1 U17730 ( .A1(n18898), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18260) );
  INV_X1 U17731 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18253) );
  NAND3_X1 U17732 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18848)
         );
  OR2_X1 U17733 ( .A1(n18253), .A2(n18848), .ZN(n14291) );
  OAI211_X1 U17734 ( .C1(n18750), .C2(n18742), .A(n18260), .B(n14291), .ZN(
        n18877) );
  MUX2_X1 U17735 ( .A(n14292), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18880), .Z(P3_U3284) );
  NAND3_X1 U17736 ( .A1(n17264), .A2(n14294), .A3(n14293), .ZN(n18252) );
  NOR2_X1 U17737 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18252), .ZN(n14295) );
  OAI21_X1 U17738 ( .B1(n14295), .B2(n18848), .A(n18362), .ZN(n18259) );
  INV_X1 U17739 ( .A(n18259), .ZN(n14296) );
  NOR2_X1 U17740 ( .A1(n17886), .A2(n18901), .ZN(n15693) );
  AOI21_X1 U17741 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15693), .ZN(n15694) );
  NOR2_X1 U17742 ( .A1(n14296), .A2(n15694), .ZN(n14298) );
  NAND2_X1 U17743 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18713), .ZN(n18430) );
  NAND2_X1 U17744 ( .A1(n18430), .A2(n18259), .ZN(n15692) );
  OR2_X1 U17745 ( .A1(n18604), .A2(n15692), .ZN(n14297) );
  MUX2_X1 U17746 ( .A(n14298), .B(n14297), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17747 ( .A(n14299), .ZN(n14300) );
  NOR2_X1 U17748 ( .A1(n14301), .A2(n14300), .ZN(n14302) );
  XNOR2_X1 U17749 ( .A(n14303), .B(n14302), .ZN(n14324) );
  INV_X1 U17750 ( .A(n14304), .ZN(n14307) );
  INV_X1 U17751 ( .A(n15171), .ZN(n14306) );
  AOI21_X1 U17752 ( .B1(n14308), .B2(n14307), .A(n14306), .ZN(n14319) );
  AOI21_X1 U17753 ( .B1(n14310), .B2(n15011), .A(n14309), .ZN(n16176) );
  INV_X1 U17754 ( .A(n16176), .ZN(n14316) );
  OAI21_X1 U17755 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15321), .A(
        n14311), .ZN(n14315) );
  AOI21_X1 U17756 ( .B1(n14313), .B2(n15088), .A(n14312), .ZN(n16197) );
  NOR2_X1 U17757 ( .A1(n19091), .A2(n19911), .ZN(n14321) );
  AOI21_X1 U17758 ( .B1(n16350), .B2(n16197), .A(n14321), .ZN(n14314) );
  OAI211_X1 U17759 ( .C1(n16341), .C2(n14316), .A(n14315), .B(n14314), .ZN(
        n14317) );
  AOI21_X1 U17760 ( .B1(n14319), .B2(n16329), .A(n14317), .ZN(n14318) );
  OAI21_X1 U17761 ( .B1(n14324), .B2(n19331), .A(n14318), .ZN(P2_U3022) );
  NAND2_X1 U17762 ( .A1(n14319), .A2(n16265), .ZN(n14323) );
  OAI22_X1 U17763 ( .A1(n9979), .A2(n19312), .B1(n19304), .B2(n16183), .ZN(
        n14320) );
  AOI211_X1 U17764 ( .C1(n16176), .C2(n19319), .A(n14321), .B(n14320), .ZN(
        n14322) );
  OAI211_X1 U17765 ( .C1(n14324), .C2(n19297), .A(n14323), .B(n14322), .ZN(
        P2_U2990) );
  NOR2_X1 U17766 ( .A1(n15124), .A2(n15042), .ZN(n14325) );
  AOI21_X1 U17767 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15042), .A(n14325), .ZN(
        n14326) );
  OAI21_X1 U17768 ( .B1(n14327), .B2(n15044), .A(n14326), .ZN(P2_U2857) );
  AND2_X1 U17769 ( .A1(n14368), .A2(n14329), .ZN(n14331) );
  INV_X1 U17770 ( .A(n14791), .ZN(n14338) );
  INV_X1 U17771 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20905) );
  OAI22_X1 U17772 ( .A1(n14358), .A2(P1_REIP_REG_29__SCAN_IN), .B1(n14347), 
        .B2(n20034), .ZN(n14334) );
  NOR2_X1 U17773 ( .A1(n20102), .A2(n14332), .ZN(n14333) );
  AOI211_X1 U17774 ( .C1(n15877), .C2(n14335), .A(n14334), .B(n14333), .ZN(
        n14336) );
  OAI21_X1 U17775 ( .B1(n20905), .B2(n14371), .A(n14336), .ZN(n14337) );
  AOI21_X1 U17776 ( .B1(n14338), .B2(n20099), .A(n14337), .ZN(n14339) );
  OAI21_X1 U17777 ( .B1(n14328), .B2(n15859), .A(n14339), .ZN(P1_U2811) );
  AND2_X1 U17778 ( .A1(n14340), .A2(n11541), .ZN(n14341) );
  NAND2_X1 U17779 ( .A1(n14637), .A2(n14341), .ZN(n14630) );
  INV_X1 U17780 ( .A(DATAI_13_), .ZN(n14342) );
  INV_X1 U17781 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14349) );
  MUX2_X1 U17782 ( .A(n14342), .B(n14349), .S(n20256), .Z(n20161) );
  OAI22_X1 U17783 ( .A1(n14630), .A2(n20161), .B1(n14637), .B2(n14343), .ZN(
        n14344) );
  AOI21_X1 U17784 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14625), .A(n14344), .ZN(
        n14346) );
  NAND2_X1 U17785 ( .A1(n14633), .A2(DATAI_29_), .ZN(n14345) );
  OAI211_X1 U17786 ( .C1(n14328), .C2(n14647), .A(n14346), .B(n14345), .ZN(
        P1_U2875) );
  OAI222_X1 U17787 ( .A1(n14542), .A2(n14328), .B1(n14347), .B2(n20116), .C1(
        n14791), .C2(n14557), .ZN(P1_U2843) );
  NAND2_X1 U17788 ( .A1(n14348), .A2(n19191), .ZN(n14356) );
  NOR2_X1 U17789 ( .A1(n19166), .A2(n14349), .ZN(n14350) );
  AOI21_X1 U17790 ( .B1(n19166), .B2(BUF2_REG_13__SCAN_IN), .A(n14350), .ZN(
        n19283) );
  OAI22_X1 U17791 ( .A1(n16196), .A2(n19283), .B1(n19187), .B2(n14351), .ZN(
        n14352) );
  AOI21_X1 U17792 ( .B1(n14353), .B2(n19206), .A(n14352), .ZN(n14355) );
  AOI22_X1 U17793 ( .A1(n19160), .A2(BUF1_REG_29__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14354) );
  OAI211_X1 U17794 ( .C1(n13418), .C2(n14356), .A(n14355), .B(n14354), .ZN(
        P2_U2890) );
  NAND2_X1 U17795 ( .A1(n14658), .A2(n20052), .ZN(n14364) );
  INV_X1 U17796 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14357) );
  OAI21_X1 U17797 ( .B1(n14358), .B2(n20905), .A(n14357), .ZN(n14361) );
  AOI22_X1 U17798 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n20103), .ZN(n14359) );
  OAI21_X1 U17799 ( .B1(n20101), .B2(n14656), .A(n14359), .ZN(n14360) );
  AOI21_X1 U17800 ( .B1(n14362), .B2(n14361), .A(n14360), .ZN(n14363) );
  OAI211_X1 U17801 ( .C1(n20088), .C2(n14778), .A(n14364), .B(n14363), .ZN(
        P1_U2810) );
  AOI21_X1 U17802 ( .B1(n14365), .B2(n14367), .A(n14366), .ZN(n14669) );
  INV_X1 U17803 ( .A(n14669), .ZN(n14580) );
  INV_X1 U17804 ( .A(n14368), .ZN(n14369) );
  AOI21_X1 U17805 ( .B1(n14370), .B2(n14386), .A(n14369), .ZN(n14802) );
  INV_X1 U17806 ( .A(n14371), .ZN(n14372) );
  OAI21_X1 U17807 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14373), .A(n14372), 
        .ZN(n14375) );
  AOI22_X1 U17808 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20103), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n14374) );
  OAI211_X1 U17809 ( .C1(n20101), .C2(n14667), .A(n14375), .B(n14374), .ZN(
        n14376) );
  AOI21_X1 U17810 ( .B1(n14802), .B2(n20099), .A(n14376), .ZN(n14377) );
  OAI21_X1 U17811 ( .B1(n14580), .B2(n15859), .A(n14377), .ZN(P1_U2812) );
  NOR2_X1 U17812 ( .A1(n14486), .A2(n14380), .ZN(n14404) );
  INV_X1 U17813 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14674) );
  INV_X1 U17814 ( .A(n14381), .ZN(n14382) );
  NOR3_X1 U17815 ( .A1(n20071), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14382), 
        .ZN(n14383) );
  AOI21_X1 U17816 ( .B1(n20103), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14383), .ZN(
        n14385) );
  NAND2_X1 U17817 ( .A1(n15877), .A2(n14678), .ZN(n14384) );
  OAI211_X1 U17818 ( .C1(n20102), .C2(n14674), .A(n14385), .B(n14384), .ZN(
        n14389) );
  OAI21_X1 U17819 ( .B1(n14398), .B2(n14387), .A(n14386), .ZN(n14811) );
  NOR2_X1 U17820 ( .A1(n14811), .A2(n20088), .ZN(n14388) );
  AOI211_X1 U17821 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14404), .A(n14389), 
        .B(n14388), .ZN(n14390) );
  OAI21_X1 U17822 ( .B1(n14675), .B2(n15859), .A(n14390), .ZN(P1_U2813) );
  INV_X1 U17823 ( .A(n14378), .ZN(n14392) );
  OAI21_X1 U17824 ( .B1(n14393), .B2(n14391), .A(n14392), .ZN(n14688) );
  INV_X1 U17825 ( .A(n14394), .ZN(n14395) );
  INV_X1 U17826 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14680) );
  OAI21_X1 U17827 ( .B1(n14395), .B2(n20071), .A(n14680), .ZN(n14403) );
  AOI22_X1 U17828 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20103), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n14396) );
  OAI21_X1 U17829 ( .B1(n20101), .B2(n14681), .A(n14396), .ZN(n14402) );
  INV_X1 U17830 ( .A(n14398), .ZN(n14399) );
  OAI21_X1 U17831 ( .B1(n14397), .B2(n14400), .A(n14399), .ZN(n14817) );
  NOR2_X1 U17832 ( .A1(n14817), .A2(n20088), .ZN(n14401) );
  AOI211_X1 U17833 ( .C1(n14404), .C2(n14403), .A(n14402), .B(n14401), .ZN(
        n14405) );
  OAI21_X1 U17834 ( .B1(n14688), .B2(n15859), .A(n14405), .ZN(P1_U2814) );
  INV_X1 U17835 ( .A(n14406), .ZN(n14407) );
  AOI21_X1 U17836 ( .B1(n14408), .B2(n14407), .A(n14391), .ZN(n14698) );
  INV_X1 U17837 ( .A(n14698), .ZN(n14594) );
  NOR2_X1 U17838 ( .A1(n20071), .A2(n14409), .ZN(n14418) );
  OAI21_X1 U17839 ( .B1(n14423), .B2(n14410), .A(n20100), .ZN(n15823) );
  OAI21_X1 U17840 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20071), .A(n15823), 
        .ZN(n14411) );
  AOI22_X1 U17841 ( .A1(n20103), .A2(P1_EBX_REG_25__SCAN_IN), .B1(n14411), 
        .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U17842 ( .A1(n15877), .A2(n14694), .ZN(n14412) );
  OAI211_X1 U17843 ( .C1(n20102), .C2(n14696), .A(n14413), .B(n14412), .ZN(
        n14417) );
  INV_X1 U17844 ( .A(n14397), .ZN(n14414) );
  OAI21_X1 U17845 ( .B1(n14415), .B2(n14499), .A(n14414), .ZN(n14831) );
  NOR2_X1 U17846 ( .A1(n14831), .A2(n20088), .ZN(n14416) );
  AOI211_X1 U17847 ( .C1(n14418), .C2(n20897), .A(n14417), .B(n14416), .ZN(
        n14419) );
  OAI21_X1 U17848 ( .B1(n14594), .B2(n15859), .A(n14419), .ZN(P1_U2815) );
  XNOR2_X1 U17849 ( .A(n9956), .B(n14512), .ZN(n15903) );
  INV_X1 U17850 ( .A(n15903), .ZN(n14611) );
  INV_X1 U17851 ( .A(n14421), .ZN(n14422) );
  NOR2_X1 U17852 ( .A1(n14422), .A2(n14432), .ZN(n15830) );
  INV_X1 U17853 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20890) );
  OAI21_X1 U17854 ( .B1(n14423), .B2(n14422), .A(n20100), .ZN(n15840) );
  OR2_X1 U17855 ( .A1(n14524), .A2(n14424), .ZN(n14425) );
  AND2_X1 U17856 ( .A1(n14515), .A2(n14425), .ZN(n14846) );
  AOI22_X1 U17857 ( .A1(n14846), .A2(n20099), .B1(n20095), .B2(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17858 ( .A1(n15877), .A2(n15902), .B1(n20103), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n14426) );
  OAI211_X1 U17859 ( .C1(n20890), .C2(n15840), .A(n14427), .B(n14426), .ZN(
        n14428) );
  AOI21_X1 U17860 ( .B1(n15830), .B2(n20890), .A(n14428), .ZN(n14429) );
  OAI21_X1 U17861 ( .B1(n14611), .B2(n15859), .A(n14429), .ZN(P1_U2819) );
  XNOR2_X1 U17862 ( .A(n14430), .B(n14526), .ZN(n14722) );
  INV_X1 U17863 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20884) );
  INV_X1 U17864 ( .A(n14431), .ZN(n14461) );
  NAND2_X1 U17865 ( .A1(n14461), .A2(n15888), .ZN(n14460) );
  NOR3_X1 U17866 ( .A1(n20884), .A2(n14437), .A3(n14460), .ZN(n15839) );
  INV_X1 U17867 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20887) );
  AND2_X1 U17868 ( .A1(n14538), .A2(n14434), .ZN(n14435) );
  NOR2_X1 U17869 ( .A1(n14522), .A2(n14435), .ZN(n15989) );
  AOI21_X1 U17870 ( .B1(n14487), .B2(n14436), .A(n14486), .ZN(n15853) );
  NOR3_X1 U17871 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14437), .A3(n14460), 
        .ZN(n15851) );
  OAI21_X1 U17872 ( .B1(n15853), .B2(n15851), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14438) );
  OAI211_X1 U17873 ( .C1(n20034), .C2(n14529), .A(n14438), .B(n20244), .ZN(
        n14439) );
  AOI21_X1 U17874 ( .B1(n15989), .B2(n20099), .A(n14439), .ZN(n14441) );
  NAND2_X1 U17875 ( .A1(n15877), .A2(n14719), .ZN(n14440) );
  OAI211_X1 U17876 ( .C1(n20102), .C2(n11927), .A(n14441), .B(n14440), .ZN(
        n14442) );
  AOI21_X1 U17877 ( .B1(n15839), .B2(n20887), .A(n14442), .ZN(n14443) );
  OAI21_X1 U17878 ( .B1(n14722), .B2(n15859), .A(n14443), .ZN(P1_U2821) );
  INV_X1 U17879 ( .A(n14445), .ZN(n14534) );
  OAI21_X1 U17880 ( .B1(n14444), .B2(n14446), .A(n14534), .ZN(n14732) );
  NAND2_X1 U17881 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15862) );
  INV_X1 U17882 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20883) );
  OAI21_X1 U17883 ( .B1(n15862), .B2(n14460), .A(n20883), .ZN(n14453) );
  OR2_X1 U17884 ( .A1(n14546), .A2(n14447), .ZN(n14448) );
  AND2_X1 U17885 ( .A1(n14536), .A2(n14448), .ZN(n16005) );
  INV_X1 U17886 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14541) );
  OAI21_X1 U17887 ( .B1(n20034), .B2(n14541), .A(n20244), .ZN(n14449) );
  AOI21_X1 U17888 ( .B1(n16005), .B2(n20099), .A(n14449), .ZN(n14451) );
  NAND2_X1 U17889 ( .A1(n15877), .A2(n14735), .ZN(n14450) );
  OAI211_X1 U17890 ( .C1(n20102), .C2(n14731), .A(n14451), .B(n14450), .ZN(
        n14452) );
  AOI21_X1 U17891 ( .B1(n14453), .B2(n15853), .A(n14452), .ZN(n14454) );
  OAI21_X1 U17892 ( .B1(n14732), .B2(n15859), .A(n14454), .ZN(P1_U2823) );
  INV_X1 U17893 ( .A(n14457), .ZN(n14458) );
  AOI21_X1 U17894 ( .B1(n14459), .B2(n14456), .A(n14458), .ZN(n14746) );
  INV_X1 U17895 ( .A(n14746), .ZN(n14638) );
  INV_X1 U17896 ( .A(n14460), .ZN(n15863) );
  INV_X1 U17897 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20880) );
  AOI21_X1 U17898 ( .B1(n14487), .B2(n14461), .A(n14486), .ZN(n15869) );
  NAND2_X1 U17899 ( .A1(n15869), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14468) );
  INV_X1 U17900 ( .A(n14556), .ZN(n14463) );
  AOI21_X1 U17901 ( .B1(n14463), .B2(n14555), .A(n14462), .ZN(n14464) );
  OR2_X1 U17902 ( .A1(n14464), .A2(n14544), .ZN(n14551) );
  INV_X1 U17903 ( .A(n14551), .ZN(n16023) );
  NAND2_X1 U17904 ( .A1(n16023), .A2(n20099), .ZN(n14465) );
  OAI211_X1 U17905 ( .C1(n14550), .C2(n20034), .A(n14465), .B(n20244), .ZN(
        n14466) );
  AOI21_X1 U17906 ( .B1(n20095), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n14466), .ZN(n14467) );
  OAI211_X1 U17907 ( .C1(n20101), .C2(n14744), .A(n14468), .B(n14467), .ZN(
        n14469) );
  AOI21_X1 U17908 ( .B1(n15863), .B2(n20880), .A(n14469), .ZN(n14470) );
  OAI21_X1 U17909 ( .B1(n14638), .B2(n15859), .A(n14470), .ZN(P1_U2825) );
  OAI21_X1 U17910 ( .B1(n9642), .B2(n11778), .A(n14472), .ZN(n14643) );
  OAI21_X1 U17911 ( .B1(n14643), .B2(n14644), .A(n14472), .ZN(n14564) );
  NAND2_X1 U17912 ( .A1(n14564), .A2(n14563), .ZN(n14562) );
  INV_X1 U17913 ( .A(n14473), .ZN(n14475) );
  AOI21_X1 U17914 ( .B1(n14562), .B2(n14475), .A(n14474), .ZN(n14758) );
  INV_X1 U17915 ( .A(n14758), .ZN(n14641) );
  NAND2_X1 U17916 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15868) );
  NOR2_X1 U17917 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15868), .ZN(n14485) );
  INV_X1 U17918 ( .A(n14565), .ZN(n14479) );
  INV_X1 U17919 ( .A(n14477), .ZN(n14478) );
  OAI21_X1 U17920 ( .B1(n14476), .B2(n14479), .A(n14478), .ZN(n14480) );
  AND2_X1 U17921 ( .A1(n14480), .A2(n14556), .ZN(n16031) );
  OAI21_X1 U17922 ( .B1(n20034), .B2(n14559), .A(n20244), .ZN(n14481) );
  AOI21_X1 U17923 ( .B1(n16031), .B2(n20099), .A(n14481), .ZN(n14483) );
  NAND2_X1 U17924 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14482) );
  OAI211_X1 U17925 ( .C1(n20101), .C2(n14756), .A(n14483), .B(n14482), .ZN(
        n14484) );
  AOI21_X1 U17926 ( .B1(n15888), .B2(n14485), .A(n14484), .ZN(n14490) );
  INV_X1 U17927 ( .A(n15868), .ZN(n14488) );
  AOI21_X1 U17928 ( .B1(n14488), .B2(n14487), .A(n14486), .ZN(n15878) );
  NAND2_X1 U17929 ( .A1(n15878), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n14489) );
  OAI211_X1 U17930 ( .C1(n14641), .C2(n15859), .A(n14490), .B(n14489), .ZN(
        P1_U2827) );
  INV_X1 U17931 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14491) );
  OAI22_X1 U17932 ( .A1(n12659), .A2(n14557), .B1(n20116), .B2(n14491), .ZN(
        P1_U2841) );
  AOI22_X1 U17933 ( .A1(n14802), .A2(n20111), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14566), .ZN(n14492) );
  OAI21_X1 U17934 ( .B1(n14580), .B2(n14542), .A(n14492), .ZN(P1_U2844) );
  INV_X1 U17935 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14493) );
  OAI222_X1 U17936 ( .A1(n14542), .A2(n14675), .B1(n14493), .B2(n20116), .C1(
        n14811), .C2(n14557), .ZN(P1_U2845) );
  INV_X1 U17937 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14494) );
  OAI222_X1 U17938 ( .A1(n14542), .A2(n14688), .B1(n14494), .B2(n20116), .C1(
        n14817), .C2(n14557), .ZN(P1_U2846) );
  INV_X1 U17939 ( .A(n14831), .ZN(n14495) );
  AOI22_X1 U17940 ( .A1(n14495), .A2(n20111), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14566), .ZN(n14496) );
  OAI21_X1 U17941 ( .B1(n14594), .B2(n14542), .A(n14496), .ZN(P1_U2847) );
  AOI21_X1 U17942 ( .B1(n14498), .B2(n14503), .A(n14406), .ZN(n15819) );
  INV_X1 U17943 ( .A(n15819), .ZN(n14600) );
  INV_X1 U17944 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14501) );
  AOI21_X1 U17945 ( .B1(n14500), .B2(n14507), .A(n14499), .ZN(n14839) );
  INV_X1 U17946 ( .A(n14839), .ZN(n15817) );
  OAI222_X1 U17947 ( .A1(n14542), .A2(n14600), .B1(n14501), .B2(n20116), .C1(
        n15817), .C2(n14557), .ZN(P1_U2848) );
  OAI21_X1 U17948 ( .B1(n14502), .B2(n14504), .A(n14503), .ZN(n15825) );
  NAND2_X1 U17949 ( .A1(n14517), .A2(n14505), .ZN(n14506) );
  AND2_X1 U17950 ( .A1(n14507), .A2(n14506), .ZN(n15972) );
  NOR2_X1 U17951 ( .A1(n20116), .A2(n14508), .ZN(n14509) );
  AOI21_X1 U17952 ( .B1(n15972), .B2(n20111), .A(n14509), .ZN(n14510) );
  OAI21_X1 U17953 ( .B1(n15825), .B2(n14542), .A(n14510), .ZN(P1_U2849) );
  AOI21_X1 U17954 ( .B1(n14420), .B2(n14512), .A(n14511), .ZN(n14513) );
  OR2_X1 U17955 ( .A1(n14513), .A2(n14502), .ZN(n15894) );
  NAND2_X1 U17956 ( .A1(n14515), .A2(n14514), .ZN(n14516) );
  NAND2_X1 U17957 ( .A1(n14517), .A2(n14516), .ZN(n15987) );
  OAI22_X1 U17958 ( .A1(n15987), .A2(n14557), .B1(n15833), .B2(n20116), .ZN(
        n14518) );
  INV_X1 U17959 ( .A(n14518), .ZN(n14519) );
  OAI21_X1 U17960 ( .B1(n15894), .B2(n14568), .A(n14519), .ZN(P1_U2850) );
  AOI22_X1 U17961 ( .A1(n14846), .A2(n20111), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14566), .ZN(n14520) );
  OAI21_X1 U17962 ( .B1(n14611), .B2(n14542), .A(n14520), .ZN(P1_U2851) );
  NOR2_X1 U17963 ( .A1(n14522), .A2(n14521), .ZN(n14523) );
  OR2_X1 U17964 ( .A1(n14524), .A2(n14523), .ZN(n15848) );
  INV_X1 U17965 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14528) );
  OAI21_X1 U17966 ( .B1(n14430), .B2(n14526), .A(n14525), .ZN(n14527) );
  AND2_X1 U17967 ( .A1(n14527), .A2(n9956), .ZN(n15846) );
  OAI222_X1 U17968 ( .A1(n15848), .A2(n14557), .B1(n20116), .B2(n14528), .C1(
        n15908), .C2(n14568), .ZN(P1_U2852) );
  NOR2_X1 U17969 ( .A1(n20116), .A2(n14529), .ZN(n14530) );
  AOI21_X1 U17970 ( .B1(n15989), .B2(n20111), .A(n14530), .ZN(n14531) );
  OAI21_X1 U17971 ( .B1(n14722), .B2(n14542), .A(n14531), .ZN(P1_U2853) );
  INV_X1 U17972 ( .A(n14430), .ZN(n14533) );
  AOI21_X1 U17973 ( .B1(n9955), .B2(n14534), .A(n14533), .ZN(n15918) );
  INV_X1 U17974 ( .A(n15918), .ZN(n14623) );
  INV_X1 U17975 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14539) );
  NAND2_X1 U17976 ( .A1(n14536), .A2(n14535), .ZN(n14537) );
  NAND2_X1 U17977 ( .A1(n14538), .A2(n14537), .ZN(n15995) );
  OAI222_X1 U17978 ( .A1(n14623), .A2(n14568), .B1(n14539), .B2(n20116), .C1(
        n15995), .C2(n14557), .ZN(P1_U2854) );
  INV_X1 U17979 ( .A(n16005), .ZN(n14540) );
  OAI222_X1 U17980 ( .A1(n14542), .A2(n14732), .B1(n20116), .B2(n14541), .C1(
        n14540), .C2(n14557), .ZN(P1_U2855) );
  NOR2_X1 U17981 ( .A1(n14544), .A2(n14543), .ZN(n14545) );
  OR2_X1 U17982 ( .A1(n14546), .A2(n14545), .ZN(n16020) );
  INV_X1 U17983 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14549) );
  AND2_X1 U17984 ( .A1(n14457), .A2(n14547), .ZN(n14548) );
  OR2_X1 U17985 ( .A1(n14548), .A2(n14444), .ZN(n15929) );
  OAI222_X1 U17986 ( .A1(n16020), .A2(n14557), .B1(n14549), .B2(n20116), .C1(
        n15929), .C2(n14568), .ZN(P1_U2856) );
  OAI22_X1 U17987 ( .A1(n14551), .A2(n14557), .B1(n14550), .B2(n20116), .ZN(
        n14552) );
  AOI21_X1 U17988 ( .B1(n14746), .B2(n20112), .A(n14552), .ZN(n14553) );
  INV_X1 U17989 ( .A(n14553), .ZN(P1_U2857) );
  OAI21_X1 U17990 ( .B1(n14474), .B2(n14554), .A(n14456), .ZN(n15867) );
  INV_X1 U17991 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14558) );
  XNOR2_X1 U17992 ( .A(n14556), .B(n14555), .ZN(n15866) );
  INV_X1 U17993 ( .A(n15866), .ZN(n14877) );
  OAI222_X1 U17994 ( .A1(n15867), .A2(n14568), .B1(n14558), .B2(n20116), .C1(
        n14557), .C2(n14877), .ZN(P1_U2858) );
  NOR2_X1 U17995 ( .A1(n20116), .A2(n14559), .ZN(n14560) );
  AOI21_X1 U17996 ( .B1(n16031), .B2(n20111), .A(n14560), .ZN(n14561) );
  OAI21_X1 U17997 ( .B1(n14641), .B2(n14568), .A(n14561), .ZN(P1_U2859) );
  OAI21_X1 U17998 ( .B1(n14564), .B2(n14563), .A(n14562), .ZN(n15876) );
  XNOR2_X1 U17999 ( .A(n14476), .B(n14565), .ZN(n15875) );
  AOI22_X1 U18000 ( .A1(n15875), .A2(n20111), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14566), .ZN(n14567) );
  OAI21_X1 U18001 ( .B1(n15876), .B2(n14568), .A(n14567), .ZN(P1_U2860) );
  INV_X1 U18002 ( .A(DATAI_14_), .ZN(n14570) );
  MUX2_X1 U18003 ( .A(n14570), .B(n14569), .S(n20256), .Z(n20164) );
  OAI22_X1 U18004 ( .A1(n14630), .A2(n20164), .B1(n14637), .B2(n13632), .ZN(
        n14571) );
  AOI21_X1 U18005 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14625), .A(n14571), .ZN(
        n14573) );
  NAND2_X1 U18006 ( .A1(n14633), .A2(DATAI_30_), .ZN(n14572) );
  OAI211_X1 U18007 ( .C1(n14574), .C2(n14647), .A(n14573), .B(n14572), .ZN(
        P1_U2874) );
  INV_X1 U18008 ( .A(DATAI_12_), .ZN(n14576) );
  INV_X1 U18009 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14575) );
  MUX2_X1 U18010 ( .A(n14576), .B(n14575), .S(n20256), .Z(n20158) );
  OAI22_X1 U18011 ( .A1(n14630), .A2(n20158), .B1(n14637), .B2(n13638), .ZN(
        n14577) );
  AOI21_X1 U18012 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14625), .A(n14577), .ZN(
        n14579) );
  NAND2_X1 U18013 ( .A1(n14633), .A2(DATAI_28_), .ZN(n14578) );
  OAI211_X1 U18014 ( .C1(n14580), .C2(n14647), .A(n14579), .B(n14578), .ZN(
        P1_U2876) );
  INV_X1 U18015 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n15060) );
  NOR2_X1 U18016 ( .A1(n14628), .A2(n15060), .ZN(n14583) );
  INV_X1 U18017 ( .A(DATAI_11_), .ZN(n14581) );
  INV_X1 U18018 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n15055) );
  MUX2_X1 U18019 ( .A(n14581), .B(n15055), .S(n20256), .Z(n20155) );
  OAI22_X1 U18020 ( .A1(n14630), .A2(n20155), .B1(n14637), .B2(n13640), .ZN(
        n14582) );
  NOR2_X1 U18021 ( .A1(n14583), .A2(n14582), .ZN(n14585) );
  NAND2_X1 U18022 ( .A1(n14633), .A2(DATAI_27_), .ZN(n14584) );
  OAI211_X1 U18023 ( .C1(n14675), .C2(n14647), .A(n14585), .B(n14584), .ZN(
        P1_U2877) );
  INV_X1 U18024 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16490) );
  NOR2_X1 U18025 ( .A1(n14628), .A2(n16490), .ZN(n14587) );
  OAI22_X1 U18026 ( .A1(n14630), .A2(n20152), .B1(n14637), .B2(n13634), .ZN(
        n14586) );
  NOR2_X1 U18027 ( .A1(n14587), .A2(n14586), .ZN(n14589) );
  NAND2_X1 U18028 ( .A1(n14633), .A2(DATAI_26_), .ZN(n14588) );
  OAI211_X1 U18029 ( .C1(n14688), .C2(n14647), .A(n14589), .B(n14588), .ZN(
        P1_U2878) );
  INV_X1 U18030 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n15080) );
  NOR2_X1 U18031 ( .A1(n14628), .A2(n15080), .ZN(n14591) );
  OAI22_X1 U18032 ( .A1(n14630), .A2(n20148), .B1(n14637), .B2(n13649), .ZN(
        n14590) );
  NOR2_X1 U18033 ( .A1(n14591), .A2(n14590), .ZN(n14593) );
  NAND2_X1 U18034 ( .A1(n14633), .A2(DATAI_25_), .ZN(n14592) );
  OAI211_X1 U18035 ( .C1(n14594), .C2(n14647), .A(n14593), .B(n14592), .ZN(
        P1_U2879) );
  INV_X1 U18036 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16493) );
  NOR2_X1 U18037 ( .A1(n14628), .A2(n16493), .ZN(n14597) );
  OAI22_X1 U18038 ( .A1(n14630), .A2(n20145), .B1(n14637), .B2(n14595), .ZN(
        n14596) );
  NOR2_X1 U18039 ( .A1(n14597), .A2(n14596), .ZN(n14599) );
  NAND2_X1 U18040 ( .A1(n14633), .A2(DATAI_24_), .ZN(n14598) );
  OAI211_X1 U18041 ( .C1(n14600), .C2(n14647), .A(n14599), .B(n14598), .ZN(
        P1_U2880) );
  OAI22_X1 U18042 ( .A1(n14630), .A2(n20309), .B1(n14637), .B2(n13646), .ZN(
        n14601) );
  AOI21_X1 U18043 ( .B1(n14625), .B2(BUF1_REG_23__SCAN_IN), .A(n14601), .ZN(
        n14603) );
  NAND2_X1 U18044 ( .A1(n14633), .A2(DATAI_23_), .ZN(n14602) );
  OAI211_X1 U18045 ( .C1(n15825), .C2(n14647), .A(n14603), .B(n14602), .ZN(
        P1_U2881) );
  OAI22_X1 U18046 ( .A1(n14630), .A2(n20301), .B1(n14637), .B2(n14604), .ZN(
        n14605) );
  AOI21_X1 U18047 ( .B1(n14625), .B2(BUF1_REG_22__SCAN_IN), .A(n14605), .ZN(
        n14607) );
  NAND2_X1 U18048 ( .A1(n14633), .A2(DATAI_22_), .ZN(n14606) );
  OAI211_X1 U18049 ( .C1(n15894), .C2(n14647), .A(n14607), .B(n14606), .ZN(
        P1_U2882) );
  OAI22_X1 U18050 ( .A1(n14630), .A2(n20297), .B1(n14637), .B2(n13654), .ZN(
        n14608) );
  AOI21_X1 U18051 ( .B1(n14625), .B2(BUF1_REG_21__SCAN_IN), .A(n14608), .ZN(
        n14610) );
  NAND2_X1 U18052 ( .A1(n14633), .A2(DATAI_21_), .ZN(n14609) );
  OAI211_X1 U18053 ( .C1(n14611), .C2(n14647), .A(n14610), .B(n14609), .ZN(
        P1_U2883) );
  OAI22_X1 U18054 ( .A1(n14630), .A2(n20292), .B1(n14637), .B2(n14612), .ZN(
        n14613) );
  AOI21_X1 U18055 ( .B1(n14625), .B2(BUF1_REG_20__SCAN_IN), .A(n14613), .ZN(
        n14615) );
  NAND2_X1 U18056 ( .A1(n14633), .A2(DATAI_20_), .ZN(n14614) );
  OAI211_X1 U18057 ( .C1(n15908), .C2(n14647), .A(n14615), .B(n14614), .ZN(
        P1_U2884) );
  OAI22_X1 U18058 ( .A1(n14630), .A2(n20286), .B1(n14637), .B2(n13644), .ZN(
        n14616) );
  AOI21_X1 U18059 ( .B1(n14625), .B2(BUF1_REG_19__SCAN_IN), .A(n14616), .ZN(
        n14618) );
  NAND2_X1 U18060 ( .A1(n14633), .A2(DATAI_19_), .ZN(n14617) );
  OAI211_X1 U18061 ( .C1(n14722), .C2(n14647), .A(n14618), .B(n14617), .ZN(
        P1_U2885) );
  INV_X1 U18062 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n19355) );
  NOR2_X1 U18063 ( .A1(n14628), .A2(n19355), .ZN(n14620) );
  OAI22_X1 U18064 ( .A1(n14630), .A2(n20282), .B1(n14637), .B2(n13652), .ZN(
        n14619) );
  NOR2_X1 U18065 ( .A1(n14620), .A2(n14619), .ZN(n14622) );
  NAND2_X1 U18066 ( .A1(n14633), .A2(DATAI_18_), .ZN(n14621) );
  OAI211_X1 U18067 ( .C1(n14623), .C2(n14647), .A(n14622), .B(n14621), .ZN(
        P1_U2886) );
  OAI22_X1 U18068 ( .A1(n14630), .A2(n20277), .B1(n14637), .B2(n13636), .ZN(
        n14624) );
  AOI21_X1 U18069 ( .B1(n14625), .B2(BUF1_REG_17__SCAN_IN), .A(n14624), .ZN(
        n14627) );
  NAND2_X1 U18070 ( .A1(n14633), .A2(DATAI_17_), .ZN(n14626) );
  OAI211_X1 U18071 ( .C1(n14732), .C2(n14647), .A(n14627), .B(n14626), .ZN(
        P1_U2887) );
  NOR2_X1 U18072 ( .A1(n14628), .A2(n16503), .ZN(n14632) );
  OAI22_X1 U18073 ( .A1(n14630), .A2(n20267), .B1(n14637), .B2(n14629), .ZN(
        n14631) );
  NOR2_X1 U18074 ( .A1(n14632), .A2(n14631), .ZN(n14635) );
  NAND2_X1 U18075 ( .A1(n14633), .A2(DATAI_16_), .ZN(n14634) );
  OAI211_X1 U18076 ( .C1(n15929), .C2(n14647), .A(n14635), .B(n14634), .ZN(
        P1_U2888) );
  OAI222_X1 U18077 ( .A1(n14638), .A2(n14647), .B1(n14637), .B2(n13625), .C1(
        n14645), .C2(n14636), .ZN(P1_U2889) );
  OAI222_X1 U18078 ( .A1(n15867), .A2(n14647), .B1(n14639), .B2(n14637), .C1(
        n14645), .C2(n20164), .ZN(P1_U2890) );
  OAI222_X1 U18079 ( .A1(n14641), .A2(n14647), .B1(n14640), .B2(n14637), .C1(
        n14645), .C2(n20161), .ZN(P1_U2891) );
  OAI222_X1 U18080 ( .A1(n15876), .A2(n14647), .B1(n14642), .B2(n14637), .C1(
        n14645), .C2(n20158), .ZN(P1_U2892) );
  XOR2_X1 U18081 ( .A(n14644), .B(n14643), .Z(n15947) );
  INV_X1 U18082 ( .A(n15947), .ZN(n14648) );
  INV_X1 U18083 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14646) );
  OAI222_X1 U18084 ( .A1(n14648), .A2(n14647), .B1(n14646), .B2(n14637), .C1(
        n14645), .C2(n20155), .ZN(P1_U2893) );
  INV_X1 U18085 ( .A(n14649), .ZN(n14653) );
  NAND2_X1 U18086 ( .A1(n20209), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14779) );
  NAND2_X1 U18087 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14655) );
  OAI211_X1 U18088 ( .C1(n20193), .C2(n14656), .A(n14779), .B(n14655), .ZN(
        n14657) );
  AOI21_X1 U18089 ( .B1(n14658), .B2(n20189), .A(n14657), .ZN(n14659) );
  OAI21_X1 U18090 ( .B1(n14787), .B2(n20016), .A(n14659), .ZN(P1_U2969) );
  NAND2_X1 U18091 ( .A1(n14684), .A2(n14660), .ZN(n14672) );
  NAND2_X1 U18092 ( .A1(n14862), .A2(n14818), .ZN(n14683) );
  NAND3_X1 U18093 ( .A1(n14709), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14683), .ZN(n14661) );
  NAND2_X1 U18094 ( .A1(n14672), .A2(n14661), .ZN(n14663) );
  INV_X1 U18095 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14807) );
  MUX2_X1 U18096 ( .A(n14807), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n14761), .Z(n14662) );
  NAND2_X1 U18097 ( .A1(n14663), .A2(n14662), .ZN(n14665) );
  INV_X1 U18098 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14664) );
  XNOR2_X1 U18099 ( .A(n14665), .B(n14664), .ZN(n14806) );
  NAND2_X1 U18100 ( .A1(n20209), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14796) );
  NAND2_X1 U18101 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14666) );
  OAI211_X1 U18102 ( .C1(n20193), .C2(n14667), .A(n14796), .B(n14666), .ZN(
        n14668) );
  AOI21_X1 U18103 ( .B1(n14669), .B2(n20189), .A(n14668), .ZN(n14670) );
  OAI21_X1 U18104 ( .B1(n20016), .B2(n14806), .A(n14670), .ZN(P1_U2971) );
  MUX2_X1 U18105 ( .A(n14672), .B(n14671), .S(n14862), .Z(n14673) );
  XNOR2_X1 U18106 ( .A(n14673), .B(n14807), .ZN(n14815) );
  NAND2_X1 U18107 ( .A1(n20209), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14810) );
  OAI21_X1 U18108 ( .B1(n15913), .B2(n14674), .A(n14810), .ZN(n14677) );
  NOR2_X1 U18109 ( .A1(n14675), .A2(n20258), .ZN(n14676) );
  AOI211_X1 U18110 ( .C1(n14678), .C2(n20199), .A(n14677), .B(n14676), .ZN(
        n14679) );
  OAI21_X1 U18111 ( .B1(n14815), .B2(n20016), .A(n14679), .ZN(P1_U2972) );
  NOR2_X1 U18112 ( .A1(n20244), .A2(n14680), .ZN(n14820) );
  NOR2_X1 U18113 ( .A1(n20193), .A2(n14681), .ZN(n14682) );
  AOI211_X1 U18114 ( .C1(n20194), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14820), .B(n14682), .ZN(n14687) );
  OAI211_X1 U18115 ( .C1(n14684), .C2(n14761), .A(n9885), .B(n14683), .ZN(
        n14685) );
  XNOR2_X1 U18116 ( .A(n14685), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14816) );
  NAND2_X1 U18117 ( .A1(n14816), .A2(n20200), .ZN(n14686) );
  OAI211_X1 U18118 ( .C1(n14688), .C2(n20258), .A(n14687), .B(n14686), .ZN(
        P1_U2973) );
  NAND2_X1 U18119 ( .A1(n14761), .A2(n12431), .ZN(n14700) );
  NAND2_X1 U18120 ( .A1(n14709), .A2(n14700), .ZN(n14689) );
  MUX2_X1 U18121 ( .A(n12419), .B(n14689), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n14690) );
  INV_X1 U18122 ( .A(n14690), .ZN(n14692) );
  NAND2_X1 U18123 ( .A1(n14691), .A2(n15943), .ZN(n14701) );
  NAND2_X1 U18124 ( .A1(n14692), .A2(n14701), .ZN(n14693) );
  XNOR2_X1 U18125 ( .A(n14693), .B(n14822), .ZN(n14835) );
  NAND2_X1 U18126 ( .A1(n20199), .A2(n14694), .ZN(n14695) );
  NAND2_X1 U18127 ( .A1(n20209), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14830) );
  OAI211_X1 U18128 ( .C1(n15913), .C2(n14696), .A(n14695), .B(n14830), .ZN(
        n14697) );
  AOI21_X1 U18129 ( .B1(n14698), .B2(n20189), .A(n14697), .ZN(n14699) );
  OAI21_X1 U18130 ( .B1(n20016), .B2(n14835), .A(n14699), .ZN(P1_U2974) );
  NAND3_X1 U18131 ( .A1(n14701), .A2(n9885), .A3(n14700), .ZN(n14703) );
  XNOR2_X1 U18132 ( .A(n14703), .B(n14702), .ZN(n14842) );
  INV_X1 U18133 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14704) );
  NOR2_X1 U18134 ( .A1(n20244), .A2(n14704), .ZN(n14838) );
  AOI21_X1 U18135 ( .B1(n20194), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14838), .ZN(n14705) );
  OAI21_X1 U18136 ( .B1(n20193), .B2(n15821), .A(n14705), .ZN(n14706) );
  AOI21_X1 U18137 ( .B1(n15819), .B2(n20189), .A(n14706), .ZN(n14707) );
  OAI21_X1 U18138 ( .B1(n20016), .B2(n14842), .A(n14707), .ZN(P1_U2975) );
  XNOR2_X1 U18139 ( .A(n14862), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14708) );
  XNOR2_X1 U18140 ( .A(n14709), .B(n14708), .ZN(n15971) );
  INV_X1 U18141 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14710) );
  OAI22_X1 U18142 ( .A1(n15913), .A2(n15829), .B1(n20244), .B2(n14710), .ZN(
        n14712) );
  NOR2_X1 U18143 ( .A1(n15825), .A2(n20258), .ZN(n14711) );
  AOI211_X1 U18144 ( .C1(n20199), .C2(n15822), .A(n14712), .B(n14711), .ZN(
        n14713) );
  OAI21_X1 U18145 ( .B1(n15971), .B2(n20016), .A(n14713), .ZN(P1_U2976) );
  NOR2_X1 U18146 ( .A1(n14761), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14715) );
  MUX2_X1 U18147 ( .A(n14862), .B(n14715), .S(n14714), .Z(n14717) );
  XNOR2_X1 U18148 ( .A(n14717), .B(n14716), .ZN(n15990) );
  NAND2_X1 U18149 ( .A1(n15990), .A2(n20200), .ZN(n14721) );
  OAI22_X1 U18150 ( .A1(n15913), .A2(n11927), .B1(n20244), .B2(n20887), .ZN(
        n14718) );
  AOI21_X1 U18151 ( .B1(n20199), .B2(n14719), .A(n14718), .ZN(n14720) );
  OAI211_X1 U18152 ( .C1(n20258), .C2(n14722), .A(n14721), .B(n14720), .ZN(
        P1_U2980) );
  NOR2_X1 U18153 ( .A1(n14761), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14729) );
  INV_X1 U18154 ( .A(n14723), .ZN(n14752) );
  NOR2_X1 U18155 ( .A1(n14752), .A2(n14724), .ZN(n14861) );
  INV_X1 U18156 ( .A(n14725), .ZN(n14726) );
  AOI21_X1 U18157 ( .B1(n14861), .B2(n14727), .A(n14726), .ZN(n14728) );
  MUX2_X1 U18158 ( .A(n14729), .B(n14761), .S(n14728), .Z(n14730) );
  XNOR2_X1 U18159 ( .A(n14730), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16004) );
  OAI22_X1 U18160 ( .A1(n15913), .A2(n14731), .B1(n20244), .B2(n20883), .ZN(
        n14734) );
  NOR2_X1 U18161 ( .A1(n14732), .A2(n20258), .ZN(n14733) );
  AOI211_X1 U18162 ( .C1(n20199), .C2(n14735), .A(n14734), .B(n14733), .ZN(
        n14736) );
  OAI21_X1 U18163 ( .B1(n20016), .B2(n16004), .A(n14736), .ZN(P1_U2982) );
  INV_X1 U18164 ( .A(n14737), .ZN(n14738) );
  OAI21_X1 U18165 ( .B1(n14723), .B2(n14739), .A(n14738), .ZN(n15923) );
  NAND2_X1 U18166 ( .A1(n14741), .A2(n14740), .ZN(n14742) );
  XNOR2_X1 U18167 ( .A(n15923), .B(n14742), .ZN(n16024) );
  INV_X1 U18168 ( .A(n16024), .ZN(n14748) );
  AOI22_X1 U18169 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14743) );
  OAI21_X1 U18170 ( .B1(n20193), .B2(n14744), .A(n14743), .ZN(n14745) );
  AOI21_X1 U18171 ( .B1(n14746), .B2(n20189), .A(n14745), .ZN(n14747) );
  OAI21_X1 U18172 ( .B1(n14748), .B2(n20016), .A(n14747), .ZN(P1_U2984) );
  NAND2_X1 U18173 ( .A1(n14862), .A2(n14749), .ZN(n14856) );
  INV_X1 U18174 ( .A(n14750), .ZN(n14751) );
  AOI22_X1 U18175 ( .A1(n14752), .A2(n14856), .B1(n15943), .B2(n14751), .ZN(
        n14884) );
  INV_X1 U18176 ( .A(n14857), .ZN(n14753) );
  AOI21_X1 U18177 ( .B1(n15943), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14753), .ZN(n14883) );
  NAND2_X1 U18178 ( .A1(n14884), .A2(n14883), .ZN(n14882) );
  NAND2_X1 U18179 ( .A1(n14882), .A2(n14857), .ZN(n14754) );
  XOR2_X1 U18180 ( .A(n14855), .B(n14754), .Z(n16032) );
  INV_X1 U18181 ( .A(n16032), .ZN(n14760) );
  AOI22_X1 U18182 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14755) );
  OAI21_X1 U18183 ( .B1(n20193), .B2(n14756), .A(n14755), .ZN(n14757) );
  AOI21_X1 U18184 ( .B1(n14758), .B2(n20189), .A(n14757), .ZN(n14759) );
  OAI21_X1 U18185 ( .B1(n14760), .B2(n20016), .A(n14759), .ZN(P1_U2986) );
  AND2_X1 U18186 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14763) );
  XNOR2_X1 U18187 ( .A(n14723), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14762) );
  MUX2_X1 U18188 ( .A(n14763), .B(n14762), .S(n14761), .Z(n14765) );
  NOR3_X1 U18189 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14862), .ZN(n15944) );
  NOR2_X1 U18190 ( .A1(n14765), .A2(n15944), .ZN(n16048) );
  AOI22_X1 U18191 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14766) );
  OAI21_X1 U18192 ( .B1(n20193), .B2(n14767), .A(n14766), .ZN(n14768) );
  AOI21_X1 U18193 ( .B1(n14769), .B2(n20189), .A(n14768), .ZN(n14770) );
  OAI21_X1 U18194 ( .B1(n16048), .B2(n20016), .A(n14770), .ZN(P1_U2989) );
  XNOR2_X1 U18195 ( .A(n14862), .B(n16060), .ZN(n14771) );
  XNOR2_X1 U18196 ( .A(n14772), .B(n14771), .ZN(n16056) );
  NAND2_X1 U18197 ( .A1(n16056), .A2(n20200), .ZN(n14776) );
  OAI22_X1 U18198 ( .A1(n15913), .A2(n14179), .B1(n20244), .B2(n20870), .ZN(
        n14773) );
  AOI21_X1 U18199 ( .B1(n20199), .B2(n14774), .A(n14773), .ZN(n14775) );
  OAI211_X1 U18200 ( .C1(n20258), .C2(n14777), .A(n14776), .B(n14775), .ZN(
        P1_U2990) );
  INV_X1 U18201 ( .A(n14778), .ZN(n14785) );
  INV_X1 U18202 ( .A(n14779), .ZN(n14784) );
  AOI21_X1 U18203 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n14783) );
  AOI211_X1 U18204 ( .C1(n14785), .C2(n20235), .A(n14784), .B(n14783), .ZN(
        n14786) );
  OAI21_X1 U18205 ( .B1(n14787), .B2(n20230), .A(n14786), .ZN(P1_U3001) );
  NAND3_X1 U18206 ( .A1(n14808), .A2(n14798), .A3(n14788), .ZN(n14789) );
  OAI211_X1 U18207 ( .C1(n14791), .C2(n20246), .A(n14790), .B(n14789), .ZN(
        n14792) );
  AOI21_X1 U18208 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14793), .A(
        n14792), .ZN(n14794) );
  OAI21_X1 U18209 ( .B1(n14795), .B2(n20230), .A(n14794), .ZN(P1_U3002) );
  INV_X1 U18210 ( .A(n14796), .ZN(n14801) );
  INV_X1 U18211 ( .A(n14808), .ZN(n14799) );
  NOR3_X1 U18212 ( .A1(n14799), .A2(n14798), .A3(n14797), .ZN(n14800) );
  AOI211_X1 U18213 ( .C1(n14802), .C2(n20235), .A(n14801), .B(n14800), .ZN(
        n14805) );
  INV_X1 U18214 ( .A(n14803), .ZN(n14813) );
  NAND2_X1 U18215 ( .A1(n14813), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14804) );
  OAI211_X1 U18216 ( .C1(n14806), .C2(n20230), .A(n14805), .B(n14804), .ZN(
        P1_U3003) );
  NAND2_X1 U18217 ( .A1(n14808), .A2(n14807), .ZN(n14809) );
  OAI211_X1 U18218 ( .C1(n14811), .C2(n20246), .A(n14810), .B(n14809), .ZN(
        n14812) );
  AOI21_X1 U18219 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14813), .A(
        n14812), .ZN(n14814) );
  OAI21_X1 U18220 ( .B1(n14815), .B2(n20230), .A(n14814), .ZN(P1_U3004) );
  INV_X1 U18221 ( .A(n14816), .ZN(n14827) );
  INV_X1 U18222 ( .A(n14817), .ZN(n14821) );
  NOR3_X1 U18223 ( .A1(n14836), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14818), .ZN(n14819) );
  AOI211_X1 U18224 ( .C1(n14821), .C2(n20235), .A(n14820), .B(n14819), .ZN(
        n14826) );
  AND2_X1 U18225 ( .A1(n14823), .A2(n14822), .ZN(n14824) );
  AND2_X1 U18226 ( .A1(n15970), .A2(n14824), .ZN(n14828) );
  OAI21_X1 U18227 ( .B1(n14833), .B2(n14828), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14825) );
  OAI211_X1 U18228 ( .C1(n14827), .C2(n20230), .A(n14826), .B(n14825), .ZN(
        P1_U3005) );
  INV_X1 U18229 ( .A(n14828), .ZN(n14829) );
  OAI211_X1 U18230 ( .C1(n14831), .C2(n20246), .A(n14830), .B(n14829), .ZN(
        n14832) );
  AOI21_X1 U18231 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14833), .A(
        n14832), .ZN(n14834) );
  OAI21_X1 U18232 ( .B1(n14835), .B2(n20230), .A(n14834), .ZN(P1_U3006) );
  NOR3_X1 U18233 ( .A1(n14836), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n12431), .ZN(n14837) );
  AOI211_X1 U18234 ( .C1(n14839), .C2(n20235), .A(n14838), .B(n14837), .ZN(
        n14841) );
  NAND2_X1 U18235 ( .A1(n15969), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14840) );
  OAI211_X1 U18236 ( .C1(n14842), .C2(n20230), .A(n14841), .B(n14840), .ZN(
        P1_U3007) );
  INV_X1 U18237 ( .A(n14714), .ZN(n14843) );
  NAND3_X1 U18238 ( .A1(n14843), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14761), .ZN(n15794) );
  INV_X1 U18239 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15800) );
  OR2_X1 U18240 ( .A1(n14844), .A2(n14862), .ZN(n15793) );
  AOI22_X1 U18241 ( .A1(n15794), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15800), .B2(n15793), .ZN(n14845) );
  XNOR2_X1 U18242 ( .A(n14845), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15906) );
  OR2_X1 U18243 ( .A1(n15906), .A2(n20230), .ZN(n14854) );
  AOI22_X1 U18244 ( .A1(n14846), .A2(n20235), .B1(n20209), .B2(
        P1_REIP_REG_21__SCAN_IN), .ZN(n14853) );
  NOR2_X1 U18245 ( .A1(n20223), .A2(n16028), .ZN(n14867) );
  INV_X1 U18246 ( .A(n14847), .ZN(n14848) );
  AOI21_X1 U18247 ( .B1(n14902), .B2(n14867), .A(n14848), .ZN(n14872) );
  NOR2_X1 U18248 ( .A1(n14872), .A2(n14849), .ZN(n15796) );
  AOI21_X1 U18249 ( .B1(n14850), .B2(n15798), .A(n15796), .ZN(n15993) );
  NOR2_X1 U18250 ( .A1(n15993), .A2(n15797), .ZN(n15977) );
  NAND2_X1 U18251 ( .A1(n15977), .A2(n15980), .ZN(n14852) );
  NAND2_X1 U18252 ( .A1(n15983), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14851) );
  NAND4_X1 U18253 ( .A1(n14854), .A2(n14853), .A3(n14852), .A4(n14851), .ZN(
        P1_U3010) );
  INV_X1 U18254 ( .A(n14855), .ZN(n14858) );
  NAND3_X1 U18255 ( .A1(n14858), .A2(n14857), .A3(n14856), .ZN(n14860) );
  OAI21_X1 U18256 ( .B1(n14861), .B2(n14860), .A(n14859), .ZN(n14864) );
  XNOR2_X1 U18257 ( .A(n14862), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14863) );
  XNOR2_X1 U18258 ( .A(n14864), .B(n14863), .ZN(n15937) );
  INV_X1 U18259 ( .A(n16046), .ZN(n14866) );
  INV_X1 U18260 ( .A(n20222), .ZN(n16065) );
  INV_X1 U18261 ( .A(n20228), .ZN(n20205) );
  OAI22_X1 U18262 ( .A1(n16065), .A2(n16045), .B1(n20205), .B2(n20229), .ZN(
        n20216) );
  NAND2_X1 U18263 ( .A1(n14865), .A2(n20216), .ZN(n16079) );
  NOR2_X1 U18264 ( .A1(n14866), .A2(n16079), .ZN(n16055) );
  NAND3_X1 U18265 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16055), .ZN(n16043) );
  NOR2_X1 U18266 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16043), .ZN(
        n14880) );
  INV_X1 U18267 ( .A(n14867), .ZN(n14868) );
  NAND2_X1 U18268 ( .A1(n14902), .A2(n14868), .ZN(n14875) );
  INV_X1 U18269 ( .A(n14869), .ZN(n14870) );
  OR2_X1 U18270 ( .A1(n20229), .A2(n14870), .ZN(n14874) );
  AND2_X1 U18271 ( .A1(n15798), .A2(n14871), .ZN(n16029) );
  NOR2_X1 U18272 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14872), .ZN(
        n16034) );
  NOR2_X1 U18273 ( .A1(n16029), .A2(n16034), .ZN(n14873) );
  NAND4_X1 U18274 ( .A1(n14875), .A2(n14874), .A3(n14873), .A4(n20253), .ZN(
        n16033) );
  AOI22_X1 U18275 ( .A1(n16033), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14876) );
  OAI21_X1 U18276 ( .B1(n14877), .B2(n20246), .A(n14876), .ZN(n14878) );
  AOI21_X1 U18277 ( .B1(n14880), .B2(n14879), .A(n14878), .ZN(n14881) );
  OAI21_X1 U18278 ( .B1(n15937), .B2(n20230), .A(n14881), .ZN(P1_U3017) );
  OAI21_X1 U18279 ( .B1(n14884), .B2(n14883), .A(n14882), .ZN(n14885) );
  INV_X1 U18280 ( .A(n14885), .ZN(n15942) );
  NAND2_X1 U18281 ( .A1(n20209), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14892) );
  INV_X1 U18282 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14890) );
  OR2_X1 U18283 ( .A1(n14890), .A2(n14886), .ZN(n14893) );
  OAI21_X1 U18284 ( .B1(n16061), .B2(n14893), .A(n20206), .ZN(n14887) );
  OAI211_X1 U18285 ( .C1(n14889), .C2(n14888), .A(n14887), .B(n16044), .ZN(
        n16039) );
  OAI221_X1 U18286 ( .B1(n16039), .B2(n20222), .C1(n16039), .C2(n14890), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14891) );
  NAND2_X1 U18287 ( .A1(n14892), .A2(n14891), .ZN(n14895) );
  NOR3_X1 U18288 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14893), .A3(
        n16079), .ZN(n14894) );
  AOI211_X1 U18289 ( .C1(n20235), .C2(n15875), .A(n14895), .B(n14894), .ZN(
        n14896) );
  OAI21_X1 U18290 ( .B1(n15942), .B2(n20230), .A(n14896), .ZN(P1_U3019) );
  INV_X1 U18291 ( .A(n14897), .ZN(n14900) );
  INV_X1 U18292 ( .A(n15798), .ZN(n14898) );
  NAND2_X1 U18293 ( .A1(n14898), .A2(n20253), .ZN(n14899) );
  AOI22_X1 U18294 ( .A1(n14900), .A2(n20249), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14899), .ZN(n14905) );
  AOI21_X1 U18295 ( .B1(n20235), .B2(n20098), .A(n14901), .ZN(n14904) );
  OR2_X1 U18296 ( .A1(n20206), .A2(n14902), .ZN(n14903) );
  NAND2_X1 U18297 ( .A1(n14903), .A2(n20223), .ZN(n20252) );
  NAND3_X1 U18298 ( .A1(n14905), .A2(n14904), .A3(n20252), .ZN(P1_U3031) );
  OAI21_X1 U18299 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14911), .A(n20787), 
        .ZN(n14907) );
  OAI21_X1 U18300 ( .B1(n14913), .B2(n14906), .A(n14907), .ZN(n14908) );
  MUX2_X1 U18301 ( .A(n14908), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n20255), .Z(P1_U3477) );
  MUX2_X1 U18302 ( .A(n20732), .B(n20506), .S(n14911), .Z(n14912) );
  NOR3_X1 U18303 ( .A1(n14912), .A2(n20631), .A3(n20418), .ZN(n14916) );
  OAI21_X1 U18304 ( .B1(n20260), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20791), 
        .ZN(n14915) );
  OAI22_X1 U18305 ( .A1(n14916), .A2(n14915), .B1(n14914), .B2(n14913), .ZN(
        n14917) );
  MUX2_X1 U18306 ( .A(n14917), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n20255), .Z(P1_U3475) );
  INV_X1 U18307 ( .A(n14906), .ZN(n20728) );
  INV_X1 U18308 ( .A(n14918), .ZN(n14920) );
  NAND2_X1 U18309 ( .A1(n14920), .A2(n14919), .ZN(n14925) );
  NAND2_X1 U18310 ( .A1(n15750), .A2(n11435), .ZN(n14921) );
  OAI21_X1 U18311 ( .B1(n14922), .B2(n14925), .A(n14921), .ZN(n14923) );
  AOI21_X1 U18312 ( .B1(n20728), .B2(n14924), .A(n14923), .ZN(n15748) );
  INV_X1 U18313 ( .A(n16097), .ZN(n14936) );
  INV_X1 U18314 ( .A(n14925), .ZN(n14929) );
  INV_X1 U18315 ( .A(n14926), .ZN(n14927) );
  AOI22_X1 U18316 ( .A1(n14930), .A2(n14929), .B1(n14928), .B2(n14927), .ZN(
        n14931) );
  OAI21_X1 U18317 ( .B1(n15748), .B2(n14936), .A(n14931), .ZN(n14933) );
  INV_X1 U18318 ( .A(n14932), .ZN(n16101) );
  MUX2_X1 U18319 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14933), .S(
        n16101), .Z(P1_U3473) );
  OAI22_X1 U18320 ( .A1(n14937), .A2(n14936), .B1(n14935), .B2(n14934), .ZN(
        n14938) );
  MUX2_X1 U18321 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14938), .S(
        n16101), .Z(P1_U3469) );
  NOR2_X1 U18322 ( .A1(n9963), .A2(n14939), .ZN(n14941) );
  XNOR2_X1 U18323 ( .A(n14941), .B(n14940), .ZN(n14942) );
  NAND2_X1 U18324 ( .A1(n14942), .A2(n19123), .ZN(n14952) );
  AOI22_X1 U18325 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19130), .B1(n14943), 
        .B2(n19089), .ZN(n14944) );
  INV_X1 U18326 ( .A(n14944), .ZN(n14947) );
  INV_X1 U18327 ( .A(n19146), .ZN(n19115) );
  OAI22_X1 U18328 ( .A1(n19115), .A2(n10281), .B1(n14945), .B2(n19139), .ZN(
        n14946) );
  AOI211_X1 U18329 ( .C1(n19098), .C2(n19198), .A(n14947), .B(n14946), .ZN(
        n14951) );
  NAND2_X1 U18330 ( .A1(n19947), .A2(n19141), .ZN(n14950) );
  NAND2_X1 U18331 ( .A1(n14948), .A2(n19151), .ZN(n14949) );
  NAND4_X1 U18332 ( .A1(n14952), .A2(n14951), .A3(n14950), .A4(n14949), .ZN(
        P2_U2852) );
  OAI22_X1 U18333 ( .A1(n19115), .A2(n10494), .B1(n14953), .B2(n19139), .ZN(
        n14954) );
  AOI21_X1 U18334 ( .B1(n19130), .B2(P2_REIP_REG_1__SCAN_IN), .A(n14954), .ZN(
        n14955) );
  OAI21_X1 U18335 ( .B1(n19149), .B2(n14956), .A(n14955), .ZN(n14957) );
  AOI21_X1 U18336 ( .B1(n19098), .B2(n19965), .A(n14957), .ZN(n14958) );
  OAI21_X1 U18337 ( .B1(n15506), .B2(n19121), .A(n14958), .ZN(n14963) );
  OAI211_X1 U18338 ( .C1(n14961), .C2(n14960), .A(n9704), .B(n14959), .ZN(
        n15507) );
  AOI221_X1 U18339 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n15507), .C1(
        n9704), .C2(n15507), .A(n19847), .ZN(n14962) );
  AOI211_X1 U18340 ( .C1(n19963), .C2(n19141), .A(n14963), .B(n14962), .ZN(
        n14964) );
  INV_X1 U18341 ( .A(n14964), .ZN(P2_U2854) );
  MUX2_X1 U18342 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16116), .S(n15036), .Z(
        P2_U2856) );
  NAND2_X1 U18343 ( .A1(n14966), .A2(n14965), .ZN(n14968) );
  XNOR2_X1 U18344 ( .A(n14968), .B(n14967), .ZN(n15051) );
  AND2_X1 U18345 ( .A1(n14980), .A2(n14969), .ZN(n14971) );
  OR2_X1 U18346 ( .A1(n14971), .A2(n14970), .ZN(n15287) );
  NOR2_X1 U18347 ( .A1(n15287), .A2(n15042), .ZN(n14972) );
  AOI21_X1 U18348 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15042), .A(n14972), .ZN(
        n14973) );
  OAI21_X1 U18349 ( .B1(n15051), .B2(n15044), .A(n14973), .ZN(P2_U2859) );
  AOI21_X1 U18350 ( .B1(n14976), .B2(n14975), .A(n14974), .ZN(n14977) );
  INV_X1 U18351 ( .A(n14977), .ZN(n15064) );
  NAND2_X1 U18352 ( .A1(n14990), .A2(n14978), .ZN(n14979) );
  NAND2_X1 U18353 ( .A1(n14980), .A2(n14979), .ZN(n16146) );
  NOR2_X1 U18354 ( .A1(n16146), .A2(n15042), .ZN(n14981) );
  AOI21_X1 U18355 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15042), .A(n14981), .ZN(
        n14982) );
  OAI21_X1 U18356 ( .B1(n15064), .B2(n15044), .A(n14982), .ZN(P2_U2860) );
  OAI21_X1 U18357 ( .B1(n14986), .B2(n14985), .A(n14984), .ZN(n15072) );
  NAND2_X1 U18358 ( .A1(n14987), .A2(n14988), .ZN(n14989) );
  AND2_X1 U18359 ( .A1(n14990), .A2(n14989), .ZN(n16157) );
  INV_X1 U18360 ( .A(n16157), .ZN(n15320) );
  NOR2_X1 U18361 ( .A1(n15320), .A2(n15042), .ZN(n14991) );
  AOI21_X1 U18362 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15042), .A(n14991), .ZN(
        n14992) );
  OAI21_X1 U18363 ( .B1(n15072), .B2(n15044), .A(n14992), .ZN(P2_U2861) );
  OAI21_X1 U18364 ( .B1(n14993), .B2(n14995), .A(n14994), .ZN(n15085) );
  OR2_X1 U18365 ( .A1(n14309), .A2(n14996), .ZN(n14997) );
  NAND2_X1 U18366 ( .A1(n14987), .A2(n14997), .ZN(n16167) );
  MUX2_X1 U18367 ( .A(n14998), .B(n16167), .S(n15036), .Z(n14999) );
  OAI21_X1 U18368 ( .B1(n15085), .B2(n15044), .A(n14999), .ZN(P2_U2862) );
  AOI21_X1 U18369 ( .B1(n15000), .B2(n15002), .A(n15001), .ZN(n15004) );
  XNOR2_X1 U18370 ( .A(n15004), .B(n15003), .ZN(n16198) );
  NAND2_X1 U18371 ( .A1(n16198), .A2(n15029), .ZN(n15006) );
  NAND2_X1 U18372 ( .A1(n16176), .A2(n15036), .ZN(n15005) );
  OAI211_X1 U18373 ( .C1(n15036), .C2(n9810), .A(n15006), .B(n15005), .ZN(
        P2_U2863) );
  AOI21_X1 U18374 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15010) );
  INV_X1 U18375 ( .A(n15010), .ZN(n15094) );
  OAI21_X1 U18376 ( .B1(n9682), .B2(n15012), .A(n15011), .ZN(n16219) );
  NOR2_X1 U18377 ( .A1(n16219), .A2(n15042), .ZN(n15013) );
  AOI21_X1 U18378 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n15042), .A(n15013), .ZN(
        n15014) );
  OAI21_X1 U18379 ( .B1(n15094), .B2(n15044), .A(n15014), .ZN(P2_U2864) );
  AOI21_X1 U18380 ( .B1(n15018), .B2(n15016), .A(n15017), .ZN(n16204) );
  NAND2_X1 U18381 ( .A1(n16204), .A2(n15029), .ZN(n15021) );
  AOI21_X1 U18382 ( .B1(n10078), .B2(n15019), .A(n9682), .ZN(n15738) );
  NAND2_X1 U18383 ( .A1(n15738), .A2(n15036), .ZN(n15020) );
  OAI211_X1 U18384 ( .C1(n15036), .C2(n10905), .A(n15021), .B(n15020), .ZN(
        P2_U2865) );
  OAI21_X1 U18385 ( .B1(n15022), .B2(n15023), .A(n15016), .ZN(n15104) );
  XOR2_X1 U18386 ( .A(n15024), .B(n15032), .Z(n18945) );
  NOR2_X1 U18387 ( .A1(n15036), .A2(n18942), .ZN(n15025) );
  AOI21_X1 U18388 ( .B1(n18945), .B2(n15036), .A(n15025), .ZN(n15026) );
  OAI21_X1 U18389 ( .B1(n15104), .B2(n15044), .A(n15026), .ZN(P2_U2866) );
  AOI21_X1 U18390 ( .B1(n15028), .B2(n15027), .A(n15022), .ZN(n16208) );
  NAND2_X1 U18391 ( .A1(n16208), .A2(n15029), .ZN(n15034) );
  NOR2_X1 U18392 ( .A1(n15040), .A2(n15030), .ZN(n15031) );
  NOR2_X1 U18393 ( .A1(n15032), .A2(n15031), .ZN(n18954) );
  NAND2_X1 U18394 ( .A1(n18954), .A2(n15036), .ZN(n15033) );
  OAI211_X1 U18395 ( .C1(n15036), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        P2_U2867) );
  OAI21_X1 U18396 ( .B1(n14276), .B2(n15037), .A(n15027), .ZN(n15116) );
  NOR2_X1 U18397 ( .A1(n14272), .A2(n15038), .ZN(n15039) );
  NOR2_X1 U18398 ( .A1(n15040), .A2(n15039), .ZN(n18966) );
  INV_X1 U18399 ( .A(n18966), .ZN(n16231) );
  NOR2_X1 U18400 ( .A1(n16231), .A2(n15042), .ZN(n15041) );
  AOI21_X1 U18401 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15042), .A(n15041), .ZN(
        n15043) );
  OAI21_X1 U18402 ( .B1(n15116), .B2(n15044), .A(n15043), .ZN(P2_U2868) );
  AOI21_X1 U18403 ( .B1(n15046), .B2(n15054), .A(n15045), .ZN(n16135) );
  AOI22_X1 U18404 ( .A1(n19167), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19166), .ZN(n19281) );
  OAI22_X1 U18405 ( .A1(n16196), .A2(n19281), .B1(n19187), .B2(n15047), .ZN(
        n15048) );
  AOI21_X1 U18406 ( .B1(n16135), .B2(n19206), .A(n15048), .ZN(n15050) );
  AOI22_X1 U18407 ( .A1(n19160), .A2(BUF1_REG_28__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15049) );
  OAI211_X1 U18408 ( .C1(n15051), .C2(n19210), .A(n15050), .B(n15049), .ZN(
        P2_U2891) );
  NAND2_X1 U18409 ( .A1(n15066), .A2(n15052), .ZN(n15053) );
  NAND2_X1 U18410 ( .A1(n15054), .A2(n15053), .ZN(n16145) );
  INV_X1 U18411 ( .A(n16145), .ZN(n15306) );
  OR2_X1 U18412 ( .A1(n19166), .A2(n15055), .ZN(n15057) );
  NAND2_X1 U18413 ( .A1(n19166), .A2(BUF2_REG_11__SCAN_IN), .ZN(n15056) );
  AND2_X1 U18414 ( .A1(n15057), .A2(n15056), .ZN(n19279) );
  OAI22_X1 U18415 ( .A1(n16196), .A2(n19279), .B1(n19187), .B2(n15058), .ZN(
        n15062) );
  INV_X1 U18416 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15059) );
  OAI22_X1 U18417 ( .A1(n15112), .A2(n15060), .B1(n15110), .B2(n15059), .ZN(
        n15061) );
  AOI211_X1 U18418 ( .C1(n19206), .C2(n15306), .A(n15062), .B(n15061), .ZN(
        n15063) );
  OAI21_X1 U18419 ( .B1(n15064), .B2(n19210), .A(n15063), .ZN(P2_U2892) );
  AOI21_X1 U18420 ( .B1(n15067), .B2(n15065), .A(n9910), .ZN(n16156) );
  INV_X1 U18421 ( .A(n19178), .ZN(n15068) );
  OAI22_X1 U18422 ( .A1(n16196), .A2(n15068), .B1(n19187), .B2(n13565), .ZN(
        n15069) );
  AOI21_X1 U18423 ( .B1(n19206), .B2(n16156), .A(n15069), .ZN(n15071) );
  AOI22_X1 U18424 ( .A1(n19160), .A2(BUF1_REG_26__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15070) );
  OAI211_X1 U18425 ( .C1(n15072), .C2(n19210), .A(n15071), .B(n15070), .ZN(
        P2_U2893) );
  OR2_X1 U18426 ( .A1(n14312), .A2(n15073), .ZN(n15074) );
  NAND2_X1 U18427 ( .A1(n15065), .A2(n15074), .ZN(n16166) );
  INV_X1 U18428 ( .A(n16166), .ZN(n15083) );
  OR2_X1 U18429 ( .A1(n19166), .A2(n15075), .ZN(n15077) );
  NAND2_X1 U18430 ( .A1(n19166), .A2(BUF2_REG_9__SCAN_IN), .ZN(n15076) );
  AND2_X1 U18431 ( .A1(n15077), .A2(n15076), .ZN(n19277) );
  OAI22_X1 U18432 ( .A1(n16196), .A2(n19277), .B1(n19187), .B2(n15078), .ZN(
        n15082) );
  INV_X1 U18433 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15079) );
  OAI22_X1 U18434 ( .A1(n15112), .A2(n15080), .B1(n15110), .B2(n15079), .ZN(
        n15081) );
  AOI211_X1 U18435 ( .C1(n19206), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15084) );
  OAI21_X1 U18436 ( .B1(n15085), .B2(n19210), .A(n15084), .ZN(P2_U2894) );
  OR2_X1 U18437 ( .A1(n15086), .A2(n9684), .ZN(n15087) );
  NAND2_X1 U18438 ( .A1(n15088), .A2(n15087), .ZN(n15346) );
  INV_X1 U18439 ( .A(n15346), .ZN(n16187) );
  AOI22_X1 U18440 ( .A1(n19167), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19166), .ZN(n19275) );
  OAI22_X1 U18441 ( .A1(n16196), .A2(n19275), .B1(n19187), .B2(n15089), .ZN(
        n15092) );
  AOI22_X1 U18442 ( .A1(n19160), .A2(BUF1_REG_23__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15090) );
  INV_X1 U18443 ( .A(n15090), .ZN(n15091) );
  AOI211_X1 U18444 ( .C1(n19206), .C2(n16187), .A(n15092), .B(n15091), .ZN(
        n15093) );
  OAI21_X1 U18445 ( .B1(n15094), .B2(n19210), .A(n15093), .ZN(P2_U2896) );
  OR2_X1 U18446 ( .A1(n15381), .A2(n15095), .ZN(n15096) );
  NAND2_X1 U18447 ( .A1(n15096), .A2(n15359), .ZN(n18951) );
  INV_X1 U18448 ( .A(n18951), .ZN(n15102) );
  OAI22_X1 U18449 ( .A1(n16196), .A2(n19271), .B1(n19187), .B2(n15097), .ZN(
        n15101) );
  INV_X1 U18450 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15099) );
  INV_X1 U18451 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15098) );
  OAI22_X1 U18452 ( .A1(n15112), .A2(n15099), .B1(n15110), .B2(n15098), .ZN(
        n15100) );
  AOI211_X1 U18453 ( .C1(n19206), .C2(n15102), .A(n15101), .B(n15100), .ZN(
        n15103) );
  OAI21_X1 U18454 ( .B1(n15104), .B2(n19210), .A(n15103), .ZN(P2_U2898) );
  NOR2_X1 U18455 ( .A1(n15106), .A2(n9687), .ZN(n15107) );
  AOI22_X1 U18456 ( .A1(n19167), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19166), .ZN(n19358) );
  OAI22_X1 U18457 ( .A1(n16196), .A2(n19358), .B1(n19187), .B2(n15108), .ZN(
        n15114) );
  INV_X1 U18458 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15111) );
  INV_X1 U18459 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15109) );
  OAI22_X1 U18460 ( .A1(n15112), .A2(n15111), .B1(n15110), .B2(n15109), .ZN(
        n15113) );
  AOI211_X1 U18461 ( .C1(n19206), .C2(n10082), .A(n15114), .B(n15113), .ZN(
        n15115) );
  OAI21_X1 U18462 ( .B1(n15116), .B2(n19210), .A(n15115), .ZN(P2_U2900) );
  NOR2_X1 U18463 ( .A1(n15118), .A2(n15117), .ZN(n15123) );
  INV_X1 U18464 ( .A(n15119), .ZN(n15121) );
  NAND2_X1 U18465 ( .A1(n15121), .A2(n15120), .ZN(n15122) );
  XNOR2_X1 U18466 ( .A(n15123), .B(n15122), .ZN(n15286) );
  XNOR2_X1 U18467 ( .A(n12625), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15283) );
  NOR2_X1 U18468 ( .A1(n19091), .A2(n19925), .ZN(n15277) );
  AOI21_X1 U18469 ( .B1(n19313), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15277), .ZN(n15125) );
  OAI21_X1 U18470 ( .B1(n16118), .B2(n19304), .A(n15125), .ZN(n15126) );
  NAND2_X1 U18471 ( .A1(n10075), .A2(n15127), .ZN(n15128) );
  AOI21_X1 U18472 ( .B1(n15283), .B2(n16265), .A(n15128), .ZN(n15129) );
  OAI21_X1 U18473 ( .B1(n15286), .B2(n19297), .A(n15129), .ZN(P2_U2984) );
  NOR2_X1 U18474 ( .A1(n15131), .A2(n15130), .ZN(n15138) );
  NAND3_X1 U18475 ( .A1(n9930), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n15132), .ZN(
        n15133) );
  AND2_X1 U18476 ( .A1(n15134), .A2(n15133), .ZN(n16144) );
  NAND2_X1 U18477 ( .A1(n16144), .A2(n15135), .ZN(n15137) );
  XNOR2_X1 U18478 ( .A(n15139), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15140) );
  INV_X1 U18479 ( .A(n15141), .ZN(n15161) );
  NAND2_X1 U18480 ( .A1(n15161), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15311) );
  AOI21_X1 U18481 ( .B1(n15142), .B2(n15311), .A(n12624), .ZN(n15296) );
  INV_X1 U18482 ( .A(n15287), .ZN(n16136) );
  NAND2_X1 U18483 ( .A1(n19291), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15291) );
  OAI21_X1 U18484 ( .B1(n19312), .B2(n15143), .A(n15291), .ZN(n15144) );
  AOI21_X1 U18485 ( .B1(n16136), .B2(n19319), .A(n15144), .ZN(n15145) );
  OAI21_X1 U18486 ( .B1(n16139), .B2(n19304), .A(n15145), .ZN(n15146) );
  AOI21_X1 U18487 ( .B1(n15296), .B2(n16265), .A(n15146), .ZN(n15147) );
  OAI21_X1 U18488 ( .B1(n15299), .B2(n19297), .A(n15147), .ZN(P2_U2986) );
  NAND3_X1 U18489 ( .A1(n15301), .A2(n19318), .A3(n15300), .ZN(n15155) );
  NOR2_X1 U18490 ( .A1(n19091), .A2(n19918), .ZN(n15305) );
  AOI21_X1 U18491 ( .B1(n19313), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15305), .ZN(n15149) );
  OAI21_X1 U18492 ( .B1(n16146), .B2(n19305), .A(n15149), .ZN(n15150) );
  AOI21_X1 U18493 ( .B1(n15151), .B2(n19290), .A(n15150), .ZN(n15154) );
  NAND2_X1 U18494 ( .A1(n15141), .A2(n15152), .ZN(n15310) );
  NAND3_X1 U18495 ( .A1(n15311), .A2(n16265), .A3(n15310), .ZN(n15153) );
  NAND3_X1 U18496 ( .A1(n15155), .A2(n15154), .A3(n15153), .ZN(P2_U2987) );
  AOI21_X1 U18497 ( .B1(n15170), .B2(n15168), .A(n15167), .ZN(n15157) );
  XOR2_X1 U18498 ( .A(n15158), .B(n15157), .Z(n15328) );
  INV_X1 U18499 ( .A(n15160), .ZN(n15330) );
  AOI21_X1 U18500 ( .B1(n15323), .B2(n15330), .A(n15161), .ZN(n15315) );
  OR2_X1 U18501 ( .A1(n19328), .A2(n15162), .ZN(n15319) );
  OAI21_X1 U18502 ( .B1(n19312), .B2(n9980), .A(n15319), .ZN(n15163) );
  AOI21_X1 U18503 ( .B1(n16157), .B2(n19319), .A(n15163), .ZN(n15164) );
  OAI21_X1 U18504 ( .B1(n16160), .B2(n19304), .A(n15164), .ZN(n15165) );
  AOI21_X1 U18505 ( .B1(n15315), .B2(n16265), .A(n15165), .ZN(n15166) );
  OAI21_X1 U18506 ( .B1(n19297), .B2(n15328), .A(n15166), .ZN(P2_U2988) );
  NAND2_X1 U18507 ( .A1(n10694), .A2(n15168), .ZN(n15169) );
  XNOR2_X1 U18508 ( .A(n15170), .B(n15169), .ZN(n15340) );
  NAND2_X1 U18509 ( .A1(n15171), .A2(n15322), .ZN(n15329) );
  NAND3_X1 U18510 ( .A1(n15330), .A2(n16265), .A3(n15329), .ZN(n15176) );
  NOR2_X1 U18511 ( .A1(n19091), .A2(n19913), .ZN(n15332) );
  AOI21_X1 U18512 ( .B1(n19313), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15332), .ZN(n15172) );
  OAI21_X1 U18513 ( .B1(n16167), .B2(n19305), .A(n15172), .ZN(n15173) );
  AOI21_X1 U18514 ( .B1(n15174), .B2(n19290), .A(n15173), .ZN(n15175) );
  OAI211_X1 U18515 ( .C1(n15340), .C2(n19297), .A(n15176), .B(n15175), .ZN(
        P2_U2989) );
  NOR2_X1 U18516 ( .A1(n15178), .A2(n9688), .ZN(n15179) );
  XNOR2_X1 U18517 ( .A(n15177), .B(n15179), .ZN(n15367) );
  INV_X1 U18518 ( .A(n15181), .ZN(n15184) );
  INV_X1 U18519 ( .A(n15182), .ZN(n15183) );
  AOI21_X1 U18520 ( .B1(n15357), .B2(n15184), .A(n15183), .ZN(n15365) );
  OAI22_X1 U18521 ( .A1(n10902), .A2(n19328), .B1(n19304), .B2(n15741), .ZN(
        n15187) );
  INV_X1 U18522 ( .A(n15738), .ZN(n15362) );
  INV_X1 U18523 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15185) );
  OAI22_X1 U18524 ( .A1(n15362), .A2(n19305), .B1(n15185), .B2(n19312), .ZN(
        n15186) );
  AOI211_X1 U18525 ( .C1(n15365), .C2(n16265), .A(n15187), .B(n15186), .ZN(
        n15188) );
  OAI21_X1 U18526 ( .B1(n15367), .B2(n19297), .A(n15188), .ZN(P2_U2992) );
  NAND2_X1 U18527 ( .A1(n15190), .A2(n15189), .ZN(n15201) );
  INV_X1 U18528 ( .A(n15452), .ZN(n15192) );
  INV_X1 U18529 ( .A(n16246), .ZN(n15193) );
  INV_X1 U18530 ( .A(n15438), .ZN(n15194) );
  INV_X1 U18531 ( .A(n15195), .ZN(n15196) );
  NAND2_X1 U18532 ( .A1(n15198), .A2(n15197), .ZN(n15223) );
  NAND2_X1 U18533 ( .A1(n19290), .A2(n15202), .ZN(n15203) );
  NAND2_X1 U18534 ( .A1(n19291), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15369) );
  OAI211_X1 U18535 ( .C1(n18941), .C2(n19312), .A(n15203), .B(n15369), .ZN(
        n15204) );
  AOI21_X1 U18536 ( .B1(n18945), .B2(n19319), .A(n15204), .ZN(n15209) );
  OR2_X1 U18537 ( .A1(n15206), .A2(n15207), .ZN(n15216) );
  AOI21_X1 U18538 ( .B1(n21096), .B2(n15216), .A(n15181), .ZN(n15375) );
  NAND2_X1 U18539 ( .A1(n15375), .A2(n16265), .ZN(n15208) );
  OAI211_X1 U18540 ( .C1(n15377), .C2(n19297), .A(n15209), .B(n15208), .ZN(
        P2_U2993) );
  INV_X1 U18541 ( .A(n15210), .ZN(n15214) );
  OAI21_X1 U18542 ( .B1(n15212), .B2(n15214), .A(n15211), .ZN(n15213) );
  OAI21_X1 U18543 ( .B1(n15215), .B2(n15214), .A(n15213), .ZN(n15390) );
  OR2_X1 U18544 ( .A1(n15206), .A2(n20966), .ZN(n15396) );
  INV_X1 U18545 ( .A(n15216), .ZN(n15217) );
  AOI21_X1 U18546 ( .B1(n15378), .B2(n15396), .A(n15217), .ZN(n15388) );
  INV_X1 U18547 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15218) );
  NOR2_X1 U18548 ( .A1(n19091), .A2(n15218), .ZN(n15382) );
  AOI21_X1 U18549 ( .B1(n19313), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15382), .ZN(n15220) );
  NAND2_X1 U18550 ( .A1(n18954), .A2(n19319), .ZN(n15219) );
  OAI211_X1 U18551 ( .C1(n18957), .C2(n19304), .A(n15220), .B(n15219), .ZN(
        n15221) );
  AOI21_X1 U18552 ( .B1(n15388), .B2(n16265), .A(n15221), .ZN(n15222) );
  OAI21_X1 U18553 ( .B1(n15390), .B2(n19297), .A(n15222), .ZN(P2_U2994) );
  XNOR2_X1 U18554 ( .A(n15224), .B(n15223), .ZN(n15436) );
  INV_X1 U18555 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19900) );
  NOR2_X1 U18556 ( .A1(n19900), .A2(n19328), .ZN(n15430) );
  OAI22_X1 U18557 ( .A1(n18985), .A2(n19312), .B1(n19304), .B2(n18992), .ZN(
        n15225) );
  AOI211_X1 U18558 ( .C1(n19319), .C2(n18988), .A(n15430), .B(n15225), .ZN(
        n15230) );
  NAND2_X1 U18559 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15226) );
  INV_X1 U18560 ( .A(n15227), .ZN(n15228) );
  OAI211_X1 U18561 ( .C1(n15426), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15228), .B(n16265), .ZN(n15229) );
  OAI211_X1 U18562 ( .C1(n15436), .C2(n19297), .A(n15230), .B(n15229), .ZN(
        P2_U2997) );
  XOR2_X1 U18563 ( .A(n15232), .B(n15231), .Z(n15733) );
  INV_X1 U18564 ( .A(n15733), .ZN(n15238) );
  INV_X1 U18565 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19898) );
  NOR2_X1 U18566 ( .A1(n19898), .A2(n19328), .ZN(n15234) );
  INV_X1 U18567 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18999) );
  OAI22_X1 U18568 ( .A1(n18999), .A2(n19312), .B1(n19304), .B2(n18998), .ZN(
        n15233) );
  AOI211_X1 U18569 ( .C1(n19319), .C2(n19003), .A(n15234), .B(n15233), .ZN(
        n15237) );
  NOR2_X1 U18570 ( .A1(n16249), .A2(n10874), .ZN(n16240) );
  INV_X1 U18571 ( .A(n15426), .ZN(n15235) );
  OAI211_X1 U18572 ( .C1(n16240), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15235), .B(n16265), .ZN(n15236) );
  OAI211_X1 U18573 ( .C1(n15238), .C2(n19297), .A(n15237), .B(n15236), .ZN(
        P2_U2998) );
  NAND2_X1 U18574 ( .A1(n15240), .A2(n15458), .ZN(n15471) );
  XNOR2_X1 U18575 ( .A(n15471), .B(n16300), .ZN(n16306) );
  XNOR2_X1 U18576 ( .A(n15241), .B(n15242), .ZN(n16303) );
  NAND2_X1 U18577 ( .A1(n16303), .A2(n19318), .ZN(n15248) );
  NOR2_X1 U18578 ( .A1(n15243), .A2(n19305), .ZN(n15246) );
  INV_X1 U18579 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19890) );
  OAI22_X1 U18580 ( .A1(n15244), .A2(n19312), .B1(n19890), .B2(n19328), .ZN(
        n15245) );
  AOI211_X1 U18581 ( .C1(n19290), .C2(n19041), .A(n15246), .B(n15245), .ZN(
        n15247) );
  OAI211_X1 U18582 ( .C1(n19323), .C2(n16306), .A(n15248), .B(n15247), .ZN(
        P2_U3002) );
  XNOR2_X1 U18583 ( .A(n15240), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15500) );
  INV_X1 U18584 ( .A(n15249), .ZN(n16273) );
  NOR2_X1 U18585 ( .A1(n16273), .A2(n15250), .ZN(n15251) );
  XNOR2_X1 U18586 ( .A(n15252), .B(n15251), .ZN(n15498) );
  OAI22_X1 U18587 ( .A1(n9985), .A2(n19312), .B1(n19304), .B2(n19071), .ZN(
        n15255) );
  OAI22_X1 U18588 ( .A1(n19074), .A2(n19305), .B1(n19091), .B2(n15253), .ZN(
        n15254) );
  AOI211_X1 U18589 ( .C1(n15498), .C2(n19318), .A(n15255), .B(n15254), .ZN(
        n15256) );
  OAI21_X1 U18590 ( .B1(n15500), .B2(n19323), .A(n15256), .ZN(P2_U3005) );
  INV_X1 U18591 ( .A(n15257), .ZN(n15258) );
  AOI21_X1 U18592 ( .B1(n14267), .B2(n15259), .A(n15258), .ZN(n15263) );
  NAND2_X1 U18593 ( .A1(n15261), .A2(n15260), .ZN(n15262) );
  XNOR2_X1 U18594 ( .A(n15263), .B(n15262), .ZN(n16333) );
  NAND2_X1 U18595 ( .A1(n15265), .A2(n15264), .ZN(n15266) );
  AND2_X1 U18596 ( .A1(n15267), .A2(n15266), .ZN(n16330) );
  INV_X1 U18597 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19884) );
  OAI22_X1 U18598 ( .A1(n15268), .A2(n19312), .B1(n19884), .B2(n19328), .ZN(
        n15272) );
  INV_X1 U18599 ( .A(n19081), .ZN(n15269) );
  OAI22_X1 U18600 ( .A1(n15270), .A2(n19305), .B1(n19304), .B2(n15269), .ZN(
        n15271) );
  AOI211_X1 U18601 ( .C1(n16330), .C2(n16265), .A(n15272), .B(n15271), .ZN(
        n15273) );
  OAI21_X1 U18602 ( .B1(n16333), .B2(n19297), .A(n15273), .ZN(P2_U3006) );
  AND2_X1 U18603 ( .A1(n15275), .A2(n15274), .ZN(n15276) );
  NOR2_X1 U18604 ( .A1(n15277), .A2(n15276), .ZN(n15280) );
  NAND2_X1 U18605 ( .A1(n15278), .A2(n16350), .ZN(n15279) );
  OAI211_X1 U18606 ( .C1(n15124), .C2(n16341), .A(n15280), .B(n15279), .ZN(
        n15281) );
  AOI21_X1 U18607 ( .B1(n15282), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15281), .ZN(n15285) );
  NAND2_X1 U18608 ( .A1(n15283), .A2(n16329), .ZN(n15284) );
  OAI211_X1 U18609 ( .C1(n15286), .C2(n19331), .A(n15285), .B(n15284), .ZN(
        P2_U3016) );
  NOR2_X1 U18610 ( .A1(n15287), .A2(n16341), .ZN(n15294) );
  INV_X1 U18611 ( .A(n16135), .ZN(n15292) );
  NAND3_X1 U18612 ( .A1(n15289), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15288), .ZN(n15290) );
  OAI211_X1 U18613 ( .C1(n15292), .C2(n19330), .A(n15291), .B(n15290), .ZN(
        n15293) );
  AOI211_X1 U18614 ( .C1(n15295), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15294), .B(n15293), .ZN(n15298) );
  NAND2_X1 U18615 ( .A1(n15296), .A2(n16329), .ZN(n15297) );
  OAI211_X1 U18616 ( .C1(n15299), .C2(n19331), .A(n15298), .B(n15297), .ZN(
        P2_U3018) );
  NAND3_X1 U18617 ( .A1(n15301), .A2(n16344), .A3(n15300), .ZN(n15314) );
  INV_X1 U18618 ( .A(n15302), .ZN(n15309) );
  NOR2_X1 U18619 ( .A1(n15303), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15304) );
  AOI211_X1 U18620 ( .C1(n16350), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15307) );
  OAI21_X1 U18621 ( .B1(n16146), .B2(n16341), .A(n15307), .ZN(n15308) );
  AOI21_X1 U18622 ( .B1(n15309), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15308), .ZN(n15313) );
  NAND3_X1 U18623 ( .A1(n15311), .A2(n16329), .A3(n15310), .ZN(n15312) );
  NAND3_X1 U18624 ( .A1(n15314), .A2(n15313), .A3(n15312), .ZN(P2_U3019) );
  NAND2_X1 U18625 ( .A1(n15315), .A2(n16329), .ZN(n15327) );
  OR3_X1 U18626 ( .A1(n15317), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15316), .ZN(n15318) );
  OAI211_X1 U18627 ( .C1(n15320), .C2(n16341), .A(n15319), .B(n15318), .ZN(
        n15325) );
  NAND3_X1 U18628 ( .A1(n15322), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15321), .ZN(n15334) );
  AOI21_X1 U18629 ( .B1(n15331), .B2(n15334), .A(n15323), .ZN(n15324) );
  AOI211_X1 U18630 ( .C1(n16350), .C2(n16156), .A(n15325), .B(n15324), .ZN(
        n15326) );
  OAI211_X1 U18631 ( .C1(n15328), .C2(n19331), .A(n15327), .B(n15326), .ZN(
        P2_U3020) );
  NAND3_X1 U18632 ( .A1(n15330), .A2(n16329), .A3(n15329), .ZN(n15339) );
  INV_X1 U18633 ( .A(n15331), .ZN(n15337) );
  NOR2_X1 U18634 ( .A1(n19330), .A2(n16166), .ZN(n15336) );
  INV_X1 U18635 ( .A(n15332), .ZN(n15333) );
  OAI211_X1 U18636 ( .C1(n16167), .C2(n16341), .A(n15334), .B(n15333), .ZN(
        n15335) );
  AOI211_X1 U18637 ( .C1(n15337), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15336), .B(n15335), .ZN(n15338) );
  OAI211_X1 U18638 ( .C1(n15340), .C2(n19331), .A(n15339), .B(n15338), .ZN(
        P2_U3021) );
  AOI21_X1 U18639 ( .B1(n15342), .B2(n15182), .A(n14304), .ZN(n16221) );
  INV_X1 U18640 ( .A(n16221), .ZN(n15354) );
  OAI21_X1 U18641 ( .B1(n15368), .B2(n21096), .A(n15473), .ZN(n15358) );
  NAND3_X1 U18642 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15341), .A3(
        n15357), .ZN(n15356) );
  NAND2_X1 U18643 ( .A1(n15358), .A2(n15356), .ZN(n15348) );
  INV_X1 U18644 ( .A(n16219), .ZN(n16188) );
  NAND2_X1 U18645 ( .A1(n16188), .A2(n19338), .ZN(n15345) );
  AOI22_X1 U18646 ( .A1(n19291), .A2(P2_REIP_REG_23__SCAN_IN), .B1(n15343), 
        .B2(n15342), .ZN(n15344) );
  OAI211_X1 U18647 ( .C1(n19330), .C2(n15346), .A(n15345), .B(n15344), .ZN(
        n15347) );
  AOI21_X1 U18648 ( .B1(n15348), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15347), .ZN(n15353) );
  NAND2_X1 U18649 ( .A1(n15351), .A2(n15350), .ZN(n16217) );
  NAND3_X1 U18650 ( .A1(n15349), .A2(n16217), .A3(n16344), .ZN(n15352) );
  OAI211_X1 U18651 ( .C1(n15354), .C2(n19343), .A(n15353), .B(n15352), .ZN(
        P2_U3023) );
  NAND2_X1 U18652 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19291), .ZN(n15355) );
  OAI211_X1 U18653 ( .C1(n15358), .C2(n15357), .A(n15356), .B(n15355), .ZN(
        n15364) );
  AOI21_X1 U18654 ( .B1(n15360), .B2(n15359), .A(n9684), .ZN(n16203) );
  INV_X1 U18655 ( .A(n16203), .ZN(n15361) );
  OAI22_X1 U18656 ( .A1(n15362), .A2(n16341), .B1(n19330), .B2(n15361), .ZN(
        n15363) );
  AOI211_X1 U18657 ( .C1(n15365), .C2(n16329), .A(n15364), .B(n15363), .ZN(
        n15366) );
  OAI21_X1 U18658 ( .B1(n15367), .B2(n19331), .A(n15366), .ZN(P2_U3024) );
  NAND2_X1 U18659 ( .A1(n15368), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15372) );
  OAI21_X1 U18660 ( .B1(n19330), .B2(n18951), .A(n15369), .ZN(n15370) );
  AOI21_X1 U18661 ( .B1(n18945), .B2(n19338), .A(n15370), .ZN(n15371) );
  OAI211_X1 U18662 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15373), .A(
        n15372), .B(n15371), .ZN(n15374) );
  AOI21_X1 U18663 ( .B1(n15375), .B2(n16329), .A(n15374), .ZN(n15376) );
  OAI21_X1 U18664 ( .B1(n15377), .B2(n19331), .A(n15376), .ZN(P2_U3025) );
  INV_X1 U18665 ( .A(n15473), .ZN(n15425) );
  NOR3_X1 U18666 ( .A1(n15397), .A2(n15425), .A3(n15378), .ZN(n15387) );
  XNOR2_X1 U18667 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15385) );
  NOR2_X1 U18668 ( .A1(n15105), .A2(n15379), .ZN(n15380) );
  NOR2_X1 U18669 ( .A1(n15381), .A2(n15380), .ZN(n18953) );
  AOI21_X1 U18670 ( .B1(n16350), .B2(n18953), .A(n15382), .ZN(n15384) );
  NAND2_X1 U18671 ( .A1(n18954), .A2(n19338), .ZN(n15383) );
  OAI211_X1 U18672 ( .C1(n15400), .C2(n15385), .A(n15384), .B(n15383), .ZN(
        n15386) );
  AOI211_X1 U18673 ( .C1(n15388), .C2(n16329), .A(n15387), .B(n15386), .ZN(
        n15389) );
  OAI21_X1 U18674 ( .B1(n15390), .B2(n19331), .A(n15389), .ZN(P2_U3026) );
  NAND2_X1 U18675 ( .A1(n15407), .A2(n15405), .ZN(n15410) );
  NAND2_X1 U18676 ( .A1(n15410), .A2(n15406), .ZN(n15394) );
  NAND2_X1 U18677 ( .A1(n15392), .A2(n15391), .ZN(n15393) );
  XNOR2_X1 U18678 ( .A(n15394), .B(n15393), .ZN(n16228) );
  INV_X1 U18679 ( .A(n16228), .ZN(n15404) );
  NAND2_X1 U18680 ( .A1(n15206), .A2(n20966), .ZN(n15395) );
  AND2_X1 U18681 ( .A1(n15396), .A2(n15395), .ZN(n16227) );
  NOR3_X1 U18682 ( .A1(n15397), .A2(n15425), .A3(n20966), .ZN(n15402) );
  INV_X1 U18683 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19903) );
  OAI22_X1 U18684 ( .A1(n16231), .A2(n16341), .B1(n19903), .B2(n19091), .ZN(
        n15398) );
  AOI21_X1 U18685 ( .B1(n16350), .B2(n10082), .A(n15398), .ZN(n15399) );
  OAI21_X1 U18686 ( .B1(n15400), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15399), .ZN(n15401) );
  AOI211_X1 U18687 ( .C1(n16227), .C2(n16329), .A(n15402), .B(n15401), .ZN(
        n15403) );
  OAI21_X1 U18688 ( .B1(n15404), .B2(n19331), .A(n15403), .ZN(P2_U3027) );
  INV_X1 U18689 ( .A(n15406), .ZN(n15409) );
  AND2_X1 U18690 ( .A1(n15406), .A2(n15405), .ZN(n15408) );
  OAI22_X1 U18691 ( .A1(n15410), .A2(n15409), .B1(n15408), .B2(n15407), .ZN(
        n16233) );
  OR2_X1 U18692 ( .A1(n15227), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15411) );
  NAND2_X1 U18693 ( .A1(n15206), .A2(n15411), .ZN(n16232) );
  AOI21_X1 U18694 ( .B1(n15413), .B2(n15412), .A(n9687), .ZN(n18976) );
  AOI22_X1 U18695 ( .A1(n16350), .A2(n18976), .B1(n18977), .B2(n19338), .ZN(
        n15421) );
  NAND2_X1 U18696 ( .A1(n15473), .A2(n15414), .ZN(n15416) );
  NAND2_X1 U18697 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n19291), .ZN(n15415) );
  OAI221_X1 U18698 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15418), 
        .C1(n15417), .C2(n15416), .A(n15415), .ZN(n15419) );
  INV_X1 U18699 ( .A(n15419), .ZN(n15420) );
  OAI211_X1 U18700 ( .C1(n16232), .C2(n19343), .A(n15421), .B(n15420), .ZN(
        n15422) );
  INV_X1 U18701 ( .A(n15422), .ZN(n15423) );
  OAI21_X1 U18702 ( .B1(n16233), .B2(n19331), .A(n15423), .ZN(P2_U3028) );
  INV_X1 U18703 ( .A(n18989), .ZN(n15431) );
  NOR2_X1 U18704 ( .A1(n15425), .A2(n15424), .ZN(n15443) );
  AOI21_X1 U18705 ( .B1(n19343), .B2(n15427), .A(n15426), .ZN(n15428) );
  INV_X1 U18706 ( .A(n15442), .ZN(n15432) );
  OAI21_X1 U18707 ( .B1(n16249), .B2(n19343), .A(n15432), .ZN(n15732) );
  NAND3_X1 U18708 ( .A1(n15732), .A2(n15433), .A3(n10882), .ZN(n15434) );
  OAI211_X1 U18709 ( .C1(n15436), .C2(n19331), .A(n15435), .B(n15434), .ZN(
        P2_U3029) );
  NAND2_X1 U18710 ( .A1(n15438), .A2(n15437), .ZN(n15440) );
  XOR2_X1 U18711 ( .A(n15440), .B(n15439), .Z(n16242) );
  NAND2_X1 U18712 ( .A1(n16249), .A2(n10874), .ZN(n16238) );
  NAND2_X1 U18713 ( .A1(n16238), .A2(n16329), .ZN(n15449) );
  INV_X1 U18714 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19896) );
  NOR2_X1 U18715 ( .A1(n19896), .A2(n19328), .ZN(n15441) );
  AOI221_X1 U18716 ( .B1(n15443), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), 
        .C1(n15442), .C2(n10874), .A(n15441), .ZN(n15448) );
  OAI21_X1 U18717 ( .B1(n15444), .B2(n15445), .A(n15729), .ZN(n19168) );
  OAI22_X1 U18718 ( .A1(n19168), .A2(n19330), .B1(n16341), .B2(n19013), .ZN(
        n15446) );
  INV_X1 U18719 ( .A(n15446), .ZN(n15447) );
  OAI211_X1 U18720 ( .C1(n16240), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        n15450) );
  AOI21_X1 U18721 ( .B1(n16242), .B2(n16344), .A(n15450), .ZN(n15451) );
  INV_X1 U18722 ( .A(n15451), .ZN(P2_U3031) );
  INV_X1 U18723 ( .A(n16259), .ZN(n15466) );
  OAI21_X1 U18724 ( .B1(n15471), .B2(n16300), .A(n10648), .ZN(n15454) );
  AND2_X1 U18725 ( .A1(n9644), .A2(n15454), .ZN(n16258) );
  OAI21_X1 U18726 ( .B1(n15455), .B2(n15457), .A(n15456), .ZN(n19173) );
  INV_X1 U18727 ( .A(n15458), .ZN(n15459) );
  OAI21_X1 U18728 ( .B1(n15459), .B2(n15492), .A(n15473), .ZN(n16301) );
  INV_X1 U18729 ( .A(n16287), .ZN(n16307) );
  NAND3_X1 U18730 ( .A1(n15458), .A2(n16307), .A3(n16300), .ZN(n16299) );
  NAND2_X1 U18731 ( .A1(n16301), .A2(n16299), .ZN(n16291) );
  NOR3_X1 U18732 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15459), .A3(
        n16287), .ZN(n16292) );
  INV_X1 U18733 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19892) );
  NOR2_X1 U18734 ( .A1(n19892), .A2(n19328), .ZN(n15460) );
  AOI21_X1 U18735 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16292), .A(
        n15460), .ZN(n15461) );
  OAI21_X1 U18736 ( .B1(n16341), .B2(n19033), .A(n15461), .ZN(n15462) );
  AOI21_X1 U18737 ( .B1(n16291), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15462), .ZN(n15463) );
  OAI21_X1 U18738 ( .B1(n19173), .B2(n19330), .A(n15463), .ZN(n15464) );
  AOI21_X1 U18739 ( .B1(n16258), .B2(n16329), .A(n15464), .ZN(n15465) );
  OAI21_X1 U18740 ( .B1(n15466), .B2(n19331), .A(n15465), .ZN(P2_U3033) );
  XOR2_X1 U18741 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15468), .Z(
        n15469) );
  XNOR2_X1 U18742 ( .A(n15467), .B(n15469), .ZN(n16264) );
  INV_X1 U18743 ( .A(n16264), .ZN(n15487) );
  AND2_X1 U18744 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15470) );
  NAND2_X1 U18745 ( .A1(n15240), .A2(n15470), .ZN(n16271) );
  NAND2_X1 U18746 ( .A1(n16271), .A2(n10612), .ZN(n15472) );
  AND2_X1 U18747 ( .A1(n15472), .A2(n15471), .ZN(n16266) );
  OAI21_X1 U18748 ( .B1(n15493), .B2(n15492), .A(n15473), .ZN(n16309) );
  OAI21_X1 U18749 ( .B1(n15474), .B2(n15476), .A(n15475), .ZN(n19176) );
  INV_X1 U18750 ( .A(n19176), .ZN(n15483) );
  INV_X1 U18751 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19889) );
  NOR2_X1 U18752 ( .A1(n19889), .A2(n19328), .ZN(n15480) );
  AOI211_X1 U18753 ( .C1(n16269), .C2(n10612), .A(n15493), .B(n16287), .ZN(
        n15477) );
  AND2_X1 U18754 ( .A1(n15478), .A2(n15477), .ZN(n15479) );
  NOR2_X1 U18755 ( .A1(n15480), .A2(n15479), .ZN(n15481) );
  OAI21_X1 U18756 ( .B1(n19054), .B2(n16341), .A(n15481), .ZN(n15482) );
  AOI21_X1 U18757 ( .B1(n15483), .B2(n16350), .A(n15482), .ZN(n15484) );
  OAI21_X1 U18758 ( .B1(n16309), .B2(n10612), .A(n15484), .ZN(n15485) );
  AOI21_X1 U18759 ( .B1(n16266), .B2(n16329), .A(n15485), .ZN(n15486) );
  OAI21_X1 U18760 ( .B1(n15487), .B2(n19331), .A(n15486), .ZN(P2_U3035) );
  OAI21_X1 U18761 ( .B1(n15488), .B2(n15490), .A(n15489), .ZN(n19181) );
  NOR2_X1 U18762 ( .A1(n15253), .A2(n19328), .ZN(n15491) );
  AOI221_X1 U18763 ( .B1(n16307), .B2(n15493), .C1(n15492), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15491), .ZN(n15496) );
  NAND2_X1 U18764 ( .A1(n15494), .A2(n19338), .ZN(n15495) );
  OAI211_X1 U18765 ( .C1(n19181), .C2(n19330), .A(n15496), .B(n15495), .ZN(
        n15497) );
  AOI21_X1 U18766 ( .B1(n15498), .B2(n16344), .A(n15497), .ZN(n15499) );
  OAI21_X1 U18767 ( .B1(n15500), .B2(n19343), .A(n15499), .ZN(P2_U3037) );
  NOR3_X1 U18768 ( .A1(n15501), .A2(n10329), .A3(n10330), .ZN(n15502) );
  AOI21_X1 U18769 ( .B1(n15504), .B2(n15503), .A(n15502), .ZN(n15505) );
  OAI21_X1 U18770 ( .B1(n15506), .B2(n15524), .A(n15505), .ZN(n16368) );
  OAI21_X1 U18771 ( .B1(n9704), .B2(n15508), .A(n15507), .ZN(n15527) );
  INV_X1 U18772 ( .A(n15527), .ZN(n15510) );
  NOR2_X1 U18773 ( .A1(n15509), .A2(n15803), .ZN(n15526) );
  AOI222_X1 U18774 ( .A1(n16368), .A2(n19940), .B1(n15525), .B2(n19963), .C1(
        n15510), .C2(n15526), .ZN(n15512) );
  NAND2_X1 U18775 ( .A1(n15696), .A2(n15516), .ZN(n15511) );
  OAI21_X1 U18776 ( .B1(n15512), .B2(n15696), .A(n15511), .ZN(P2_U3600) );
  NAND2_X1 U18777 ( .A1(n15514), .A2(n15513), .ZN(n15521) );
  AOI21_X1 U18778 ( .B1(n15516), .B2(n16364), .A(n15515), .ZN(n15517) );
  OAI22_X1 U18779 ( .A1(n15519), .A2(n15521), .B1(n15518), .B2(n15517), .ZN(
        n15520) );
  AOI21_X1 U18780 ( .B1(n15522), .B2(n15521), .A(n15520), .ZN(n15523) );
  OAI21_X1 U18781 ( .B1(n10289), .B2(n15524), .A(n15523), .ZN(n16373) );
  AOI222_X1 U18782 ( .A1(n16373), .A2(n19940), .B1(n15527), .B2(n15526), .C1(
        n15525), .C2(n19955), .ZN(n15529) );
  NAND2_X1 U18783 ( .A1(n15696), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15528) );
  OAI21_X1 U18784 ( .B1(n15529), .B2(n15696), .A(n15528), .ZN(P2_U3599) );
  INV_X1 U18785 ( .A(n19400), .ZN(n15530) );
  INV_X1 U18786 ( .A(n19938), .ZN(n19989) );
  NOR3_X1 U18787 ( .A1(n19837), .A2(n19387), .A3(n19989), .ZN(n15531) );
  AND2_X1 U18788 ( .A1(n19938), .A2(n18922), .ZN(n19941) );
  NOR2_X1 U18789 ( .A1(n15531), .A2(n19941), .ZN(n15534) );
  NOR2_X1 U18790 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19431) );
  INV_X1 U18791 ( .A(n19431), .ZN(n16375) );
  NOR2_X1 U18792 ( .A1(n19684), .A2(n16375), .ZN(n19373) );
  NOR2_X1 U18793 ( .A1(n19833), .A2(n19373), .ZN(n15537) );
  INV_X1 U18794 ( .A(n10544), .ZN(n15532) );
  OAI21_X1 U18795 ( .B1(n15532), .B2(n19373), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15533) );
  INV_X1 U18796 ( .A(n19374), .ZN(n15549) );
  INV_X1 U18797 ( .A(n19821), .ZN(n15542) );
  INV_X1 U18798 ( .A(n15534), .ZN(n15538) );
  AOI21_X1 U18799 ( .B1(n10544), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n15535) );
  OAI21_X1 U18800 ( .B1(n15535), .B2(n19373), .A(n19788), .ZN(n15536) );
  INV_X1 U18801 ( .A(n19378), .ZN(n15546) );
  INV_X1 U18802 ( .A(n19763), .ZN(n19825) );
  INV_X1 U18803 ( .A(n19837), .ZN(n19800) );
  AOI22_X1 U18804 ( .A1(n19822), .A2(n19387), .B1(n19820), .B2(n19373), .ZN(
        n15539) );
  OAI21_X1 U18805 ( .B1(n19825), .B2(n19800), .A(n15539), .ZN(n15540) );
  AOI21_X1 U18806 ( .B1(n15546), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15540), .ZN(n15541) );
  OAI21_X1 U18807 ( .B1(n15549), .B2(n15542), .A(n15541), .ZN(P2_U3053) );
  OAI22_X1 U18808 ( .A1(n19166), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19167), .ZN(n19273) );
  NOR2_X2 U18809 ( .A1(n19273), .A2(n19601), .ZN(n19827) );
  INV_X1 U18810 ( .A(n19827), .ZN(n15548) );
  AOI22_X1 U18811 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19361), .ZN(n19529) );
  NOR2_X2 U18812 ( .A1(n15543), .A2(n19363), .ZN(n19826) );
  AOI22_X1 U18813 ( .A1(n19828), .A2(n19387), .B1(n19373), .B2(n19826), .ZN(
        n15544) );
  OAI21_X1 U18814 ( .B1(n19831), .B2(n19800), .A(n15544), .ZN(n15545) );
  AOI21_X1 U18815 ( .B1(n15546), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15545), .ZN(n15547) );
  OAI21_X1 U18816 ( .B1(n15549), .B2(n15548), .A(n15547), .ZN(P2_U3054) );
  NAND2_X1 U18817 ( .A1(n10498), .A2(n19431), .ZN(n15557) );
  NOR2_X1 U18818 ( .A1(n19950), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19967) );
  OR3_X1 U18819 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19600), .A3(n19542), 
        .ZN(n15550) );
  OAI21_X1 U18820 ( .B1(n15557), .B2(n19967), .A(n15550), .ZN(n15554) );
  NOR2_X1 U18821 ( .A1(n19973), .A2(n15557), .ZN(n19394) );
  INV_X1 U18822 ( .A(n19394), .ZN(n15561) );
  AND2_X1 U18823 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15561), .ZN(n15551) );
  NAND2_X1 U18824 ( .A1(n15552), .A2(n15551), .ZN(n15555) );
  AND2_X1 U18825 ( .A1(n15555), .A2(n19788), .ZN(n15553) );
  NAND2_X1 U18826 ( .A1(n15554), .A2(n15553), .ZN(n19396) );
  INV_X1 U18827 ( .A(n19396), .ZN(n19382) );
  INV_X1 U18828 ( .A(n15555), .ZN(n15556) );
  AOI211_X2 U18829 ( .C1(n15557), .C2(n19777), .A(n19721), .B(n15556), .ZN(
        n19395) );
  NOR2_X2 U18830 ( .A1(n19275), .A2(n19601), .ZN(n19834) );
  NAND2_X1 U18831 ( .A1(n15558), .A2(n19352), .ZN(n19372) );
  INV_X1 U18832 ( .A(n19600), .ZN(n15559) );
  NAND2_X1 U18833 ( .A1(n15559), .A2(n19548), .ZN(n19423) );
  INV_X1 U18834 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n21103) );
  INV_X1 U18835 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18292) );
  OAI22_X2 U18836 ( .A1(n21103), .A2(n19368), .B1(n18292), .B2(n19366), .ZN(
        n19836) );
  AOI22_X1 U18837 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19361), .ZN(n19842) );
  AOI22_X1 U18838 ( .A1(n19426), .A2(n19836), .B1(n19387), .B2(n19770), .ZN(
        n15560) );
  OAI21_X1 U18839 ( .B1(n19372), .B2(n15561), .A(n15560), .ZN(n15562) );
  AOI21_X1 U18840 ( .B1(n19395), .B2(n19834), .A(n15562), .ZN(n15563) );
  OAI21_X1 U18841 ( .B1(n19382), .B2(n15564), .A(n15563), .ZN(P2_U3063) );
  AOI21_X1 U18842 ( .B1(n19520), .B2(n19563), .A(n18922), .ZN(n15565) );
  NAND2_X1 U18843 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19536), .ZN(
        n19544) );
  NOR2_X1 U18844 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19544), .ZN(
        n19530) );
  AOI221_X1 U18845 ( .B1(n19510), .B2(n19950), .C1(n15565), .C2(n19950), .A(
        n19530), .ZN(n15568) );
  INV_X1 U18846 ( .A(n15566), .ZN(n15569) );
  NOR3_X1 U18847 ( .A1(n15569), .A2(n19530), .A3(n19777), .ZN(n15567) );
  INV_X1 U18848 ( .A(n19533), .ZN(n15576) );
  INV_X1 U18849 ( .A(n19536), .ZN(n19461) );
  OAI21_X1 U18850 ( .B1(n15569), .B2(n19530), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15570) );
  OAI21_X1 U18851 ( .B1(n19461), .B2(n19632), .A(n15570), .ZN(n19531) );
  INV_X1 U18852 ( .A(n19530), .ZN(n15572) );
  INV_X1 U18853 ( .A(n19563), .ZN(n19565) );
  AOI22_X1 U18854 ( .A1(n19565), .A2(n19790), .B1(n19532), .B2(n19695), .ZN(
        n15571) );
  OAI21_X1 U18855 ( .B1(n15582), .B2(n15572), .A(n15571), .ZN(n15573) );
  AOI21_X1 U18856 ( .B1(n19531), .B2(n19782), .A(n15573), .ZN(n15574) );
  OAI21_X1 U18857 ( .B1(n15576), .B2(n15575), .A(n15574), .ZN(P2_U3096) );
  NOR3_X1 U18858 ( .A1(n19797), .A2(n19771), .A3(n19989), .ZN(n15578) );
  NOR2_X1 U18859 ( .A1(n15578), .A2(n19941), .ZN(n15587) );
  INV_X1 U18860 ( .A(n15587), .ZN(n15580) );
  NAND2_X1 U18861 ( .A1(n19463), .A2(n19719), .ZN(n15586) );
  INV_X1 U18862 ( .A(n10431), .ZN(n15584) );
  NAND2_X1 U18863 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19719), .ZN(
        n19786) );
  NOR2_X1 U18864 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19786), .ZN(
        n19769) );
  AOI211_X1 U18865 ( .C1(n15584), .C2(n19950), .A(n19938), .B(n19769), .ZN(
        n15579) );
  INV_X1 U18866 ( .A(n19769), .ZN(n15581) );
  OAI22_X1 U18867 ( .A1(n19841), .A2(n19698), .B1(n15582), .B2(n15581), .ZN(
        n15583) );
  AOI21_X1 U18868 ( .B1(n19771), .B2(n19695), .A(n15583), .ZN(n15589) );
  OAI21_X1 U18869 ( .B1(n15584), .B2(n19769), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15585) );
  NAND2_X1 U18870 ( .A1(n19772), .A2(n19782), .ZN(n15588) );
  OAI211_X1 U18871 ( .C1(n19775), .C2(n15590), .A(n15589), .B(n15588), .ZN(
        P2_U3160) );
  INV_X1 U18872 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16645) );
  NOR3_X1 U18873 ( .A1(n15592), .A2(n17340), .A3(n15591), .ZN(n15594) );
  INV_X1 U18874 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17269) );
  NAND3_X1 U18875 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17268) );
  NOR4_X1 U18876 ( .A1(n16864), .A2(n17269), .A3(n15596), .A4(n17268), .ZN(
        n15597) );
  NAND3_X1 U18877 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n15597), .ZN(n15690) );
  NAND2_X1 U18878 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .ZN(n15689) );
  NAND4_X1 U18879 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n17132)
         );
  NOR3_X1 U18880 ( .A1(n15690), .A2(n15689), .A3(n17132), .ZN(n15598) );
  NAND4_X1 U18881 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n15598), .ZN(n17112) );
  NOR2_X1 U18882 ( .A1(n17114), .A2(n17112), .ZN(n17087) );
  NAND2_X1 U18883 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17087), .ZN(n17086) );
  NAND2_X1 U18884 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17083), .ZN(n17082) );
  NOR2_X1 U18885 ( .A1(n17340), .A2(n17082), .ZN(n17070) );
  NAND2_X1 U18886 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17070), .ZN(n17056) );
  NAND2_X1 U18887 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17029), .ZN(n17022) );
  NAND2_X1 U18888 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17028), .ZN(n17012) );
  NAND2_X1 U18889 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17017), .ZN(n17002) );
  NAND2_X1 U18890 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17007), .ZN(n17001) );
  INV_X1 U18891 ( .A(n17001), .ZN(n15677) );
  INV_X2 U18892 ( .A(n17296), .ZN(n17290) );
  AOI21_X1 U18893 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17290), .A(n17007), .ZN(
        n15676) );
  AOI22_X1 U18894 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15599) );
  OAI21_X1 U18895 ( .B1(n13126), .B2(n17060), .A(n15599), .ZN(n15610) );
  AOI22_X1 U18896 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15607) );
  AOI22_X1 U18897 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15600) );
  OAI21_X1 U18898 ( .B1(n17229), .B2(n15601), .A(n15600), .ZN(n15605) );
  AOI22_X1 U18899 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15603) );
  AOI22_X1 U18900 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15602) );
  OAI211_X1 U18901 ( .C1(n9629), .C2(n17172), .A(n15603), .B(n15602), .ZN(
        n15604) );
  AOI211_X1 U18902 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n15605), .B(n15604), .ZN(n15606) );
  OAI211_X1 U18903 ( .C1(n13156), .C2(n15608), .A(n15607), .B(n15606), .ZN(
        n15609) );
  AOI211_X1 U18904 ( .C1(n9639), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n15610), .B(n15609), .ZN(n17004) );
  AOI22_X1 U18905 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15611) );
  OAI21_X1 U18906 ( .B1(n17058), .B2(n17289), .A(n15611), .ZN(n15620) );
  INV_X1 U18907 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U18908 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18909 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15612) );
  OAI21_X1 U18910 ( .B1(n17250), .B2(n20947), .A(n15612), .ZN(n15616) );
  AOI22_X1 U18911 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U18912 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15613) );
  OAI211_X1 U18913 ( .C1(n17229), .C2(n17218), .A(n15614), .B(n15613), .ZN(
        n15615) );
  AOI211_X1 U18914 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n15616), .B(n15615), .ZN(n15617) );
  OAI211_X1 U18915 ( .C1(n13131), .C2(n17207), .A(n15618), .B(n15617), .ZN(
        n15619) );
  AOI211_X1 U18916 ( .C1(n9632), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n15620), .B(n15619), .ZN(n17014) );
  INV_X1 U18917 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15622) );
  AOI22_X1 U18918 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15621) );
  OAI21_X1 U18919 ( .B1(n17208), .B2(n15622), .A(n15621), .ZN(n15631) );
  INV_X1 U18920 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U18921 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15629) );
  OAI22_X1 U18922 ( .A1(n13126), .A2(n17122), .B1(n13194), .B2(n17126), .ZN(
        n15627) );
  AOI22_X1 U18923 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15625) );
  AOI22_X1 U18924 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U18925 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15623) );
  NAND3_X1 U18926 ( .A1(n15625), .A2(n15624), .A3(n15623), .ZN(n15626) );
  AOI211_X1 U18927 ( .C1(n17255), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n15627), .B(n15626), .ZN(n15628) );
  OAI211_X1 U18928 ( .C1(n17264), .C2(n17249), .A(n15629), .B(n15628), .ZN(
        n15630) );
  AOI211_X1 U18929 ( .C1(n9639), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n15631), .B(n15630), .ZN(n17024) );
  AOI22_X1 U18930 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n13141), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17254), .ZN(n15632) );
  OAI21_X1 U18931 ( .B1(n21077), .B2(n17208), .A(n15632), .ZN(n15643) );
  INV_X1 U18932 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15641) );
  AOI22_X1 U18933 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15639) );
  AOI22_X1 U18934 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17236), .B1(
        n13171), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15633) );
  OAI21_X1 U18935 ( .B1(n17264), .B2(n17270), .A(n15633), .ZN(n15637) );
  INV_X1 U18936 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U18937 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13196), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U18938 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17230), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15634) );
  OAI211_X1 U18939 ( .C1(n17139), .C2(n9629), .A(n15635), .B(n15634), .ZN(
        n15636) );
  AOI211_X1 U18940 ( .C1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .C2(n13138), .A(
        n15637), .B(n15636), .ZN(n15638) );
  OAI211_X1 U18941 ( .C1(n15641), .C2(n15640), .A(n15639), .B(n15638), .ZN(
        n15642) );
  AOI211_X1 U18942 ( .C1(n17255), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n15643), .B(n15642), .ZN(n17025) );
  NOR2_X1 U18943 ( .A1(n17024), .A2(n17025), .ZN(n17023) );
  AOI22_X1 U18944 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15653) );
  AOI22_X1 U18945 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U18946 ( .A1(n17236), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15651) );
  OAI22_X1 U18947 ( .A1(n13194), .A2(n17102), .B1(n17199), .B2(n17101), .ZN(
        n15649) );
  AOI22_X1 U18948 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15647) );
  AOI22_X1 U18949 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U18950 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13171), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15645) );
  NAND2_X1 U18951 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n15644) );
  NAND4_X1 U18952 ( .A1(n15647), .A2(n15646), .A3(n15645), .A4(n15644), .ZN(
        n15648) );
  AOI211_X1 U18953 ( .C1(n17255), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n15649), .B(n15648), .ZN(n15650) );
  NAND4_X1 U18954 ( .A1(n15653), .A2(n15652), .A3(n15651), .A4(n15650), .ZN(
        n17019) );
  NAND2_X1 U18955 ( .A1(n17023), .A2(n17019), .ZN(n17018) );
  NOR2_X1 U18956 ( .A1(n17014), .A2(n17018), .ZN(n17013) );
  AOI22_X1 U18957 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U18958 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15654) );
  OAI21_X1 U18959 ( .B1(n13126), .B2(n17198), .A(n15654), .ZN(n15662) );
  AOI22_X1 U18960 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15660) );
  INV_X1 U18961 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U18962 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18963 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15655) );
  OAI211_X1 U18964 ( .C1(n17250), .C2(n15657), .A(n15656), .B(n15655), .ZN(
        n15658) );
  AOI21_X1 U18965 ( .B1(n17244), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n15658), .ZN(n15659) );
  OAI211_X1 U18966 ( .C1(n17229), .C2(n21072), .A(n15660), .B(n15659), .ZN(
        n15661) );
  AOI211_X1 U18967 ( .C1(n17255), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n15662), .B(n15661), .ZN(n15663) );
  OAI211_X1 U18968 ( .C1(n17058), .C2(n17283), .A(n15664), .B(n15663), .ZN(
        n17009) );
  NAND2_X1 U18969 ( .A1(n17013), .A2(n17009), .ZN(n17008) );
  NOR2_X1 U18970 ( .A1(n17004), .A2(n17008), .ZN(n17003) );
  AOI22_X1 U18971 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15674) );
  INV_X1 U18972 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U18973 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U18974 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15665) );
  OAI211_X1 U18975 ( .C1(n9629), .C2(n17044), .A(n15666), .B(n15665), .ZN(
        n15672) );
  AOI22_X1 U18976 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15670) );
  AOI22_X1 U18977 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15669) );
  AOI22_X1 U18978 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9632), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15668) );
  NAND2_X1 U18979 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n15667) );
  NAND4_X1 U18980 ( .A1(n15670), .A2(n15669), .A3(n15668), .A4(n15667), .ZN(
        n15671) );
  AOI211_X1 U18981 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15672), .B(n15671), .ZN(n15673) );
  OAI211_X1 U18982 ( .C1(n17229), .C2(n21120), .A(n15674), .B(n15673), .ZN(
        n15675) );
  NAND2_X1 U18983 ( .A1(n17003), .A2(n15675), .ZN(n16997) );
  OAI21_X1 U18984 ( .B1(n17003), .B2(n15675), .A(n16997), .ZN(n17314) );
  OAI22_X1 U18985 ( .A1(n15677), .A2(n15676), .B1(n17314), .B2(n17290), .ZN(
        P3_U2675) );
  INV_X1 U18986 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U18987 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15678) );
  OAI21_X1 U18988 ( .B1(n13156), .B2(n15679), .A(n15678), .ZN(n15688) );
  AOI22_X1 U18989 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18990 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17245), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15680) );
  OAI21_X1 U18991 ( .B1(n9629), .B2(n17277), .A(n15680), .ZN(n15684) );
  INV_X1 U18992 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n21058) );
  AOI22_X1 U18993 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15682) );
  AOI22_X1 U18994 ( .A1(n17253), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15681) );
  OAI211_X1 U18995 ( .C1(n17229), .C2(n21058), .A(n15682), .B(n15681), .ZN(
        n15683) );
  AOI211_X1 U18996 ( .C1(n17236), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15684), .B(n15683), .ZN(n15685) );
  OAI211_X1 U18997 ( .C1(n13131), .C2(n17044), .A(n15686), .B(n15685), .ZN(
        n15687) );
  AOI211_X1 U18998 ( .C1(n9639), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n15688), .B(n15687), .ZN(n17391) );
  INV_X1 U18999 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17184) );
  INV_X1 U19000 ( .A(n15689), .ZN(n17185) );
  NAND3_X1 U19001 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17272), .ZN(n17242) );
  NAND2_X1 U19002 ( .A1(n17185), .A2(n17202), .ZN(n17203) );
  NOR2_X1 U19003 ( .A1(n17184), .A2(n17203), .ZN(n17151) );
  AND2_X1 U19004 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17151), .ZN(n17169) );
  NOR2_X1 U19005 ( .A1(n17296), .A2(n17169), .ZN(n17168) );
  OAI21_X1 U19006 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17151), .A(n17168), .ZN(
        n15691) );
  OAI21_X1 U19007 ( .B1(n17391), .B2(n17290), .A(n15691), .ZN(P3_U2690) );
  NAND2_X1 U19008 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18407) );
  AOI221_X1 U19009 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18407), .C1(n15693), 
        .C2(n18407), .A(n15692), .ZN(n18258) );
  NOR2_X1 U19010 ( .A1(n15694), .A2(n18714), .ZN(n15695) );
  OAI21_X1 U19011 ( .B1(n15695), .B2(n18604), .A(n18259), .ZN(n18256) );
  AOI22_X1 U19012 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18258), .B1(
        n18256), .B2(n18255), .ZN(P3_U2865) );
  INV_X1 U19013 ( .A(n15696), .ZN(n15701) );
  NOR4_X1 U19014 ( .A1(n10767), .A2(n16380), .A3(n19997), .A4(n15697), .ZN(
        n15698) );
  NAND2_X1 U19015 ( .A1(n15701), .A2(n15698), .ZN(n15699) );
  OAI21_X1 U19016 ( .B1(n15701), .B2(n15700), .A(n15699), .ZN(P2_U3595) );
  INV_X1 U19017 ( .A(n15702), .ZN(n18220) );
  INV_X1 U19018 ( .A(n18696), .ZN(n15707) );
  OAI21_X1 U19019 ( .B1(n18273), .B2(n18268), .A(n18891), .ZN(n15703) );
  OAI21_X1 U19020 ( .B1(n15704), .B2(n15703), .A(n18904), .ZN(n16575) );
  OR3_X1 U19021 ( .A1(n15709), .A2(n16576), .A3(n16575), .ZN(n15705) );
  OAI211_X1 U19022 ( .C1(n15708), .C2(n15707), .A(n15706), .B(n15705), .ZN(
        n15710) );
  NOR3_X1 U19023 ( .A1(n18160), .A2(n18155), .A3(n18154), .ZN(n18043) );
  AOI21_X1 U19024 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18216) );
  NAND3_X1 U19025 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18042) );
  NOR2_X1 U19026 ( .A1(n18216), .A2(n18042), .ZN(n18153) );
  NAND2_X1 U19027 ( .A1(n18043), .A2(n18153), .ZN(n18138) );
  NAND2_X1 U19028 ( .A1(n18039), .A2(n17992), .ZN(n16459) );
  NOR2_X1 U19029 ( .A1(n18138), .A2(n16459), .ZN(n18034) );
  NAND2_X1 U19030 ( .A1(n17958), .A2(n18034), .ZN(n17980) );
  NOR2_X1 U19031 ( .A1(n16460), .A2(n17980), .ZN(n15715) );
  INV_X1 U19032 ( .A(n18712), .ZN(n18243) );
  OAI21_X1 U19033 ( .B1(n17934), .B2(n18876), .A(n18243), .ZN(n18217) );
  NOR2_X1 U19034 ( .A1(n18227), .A2(n18861), .ZN(n18194) );
  INV_X1 U19035 ( .A(n18194), .ZN(n18040) );
  NOR2_X1 U19036 ( .A1(n18040), .A2(n18042), .ZN(n18150) );
  NAND2_X1 U19037 ( .A1(n18150), .A2(n18043), .ZN(n18137) );
  OR2_X1 U19038 ( .A1(n18045), .A2(n18137), .ZN(n18036) );
  NOR2_X1 U19039 ( .A1(n15711), .A2(n18036), .ZN(n15717) );
  AOI22_X1 U19040 ( .A1(n18691), .A2(n15715), .B1(n18217), .B2(n15717), .ZN(
        n15712) );
  NOR2_X1 U19041 ( .A1(n15712), .A2(n18235), .ZN(n16450) );
  NAND2_X1 U19042 ( .A1(n17416), .A2(n18171), .ZN(n18064) );
  NOR2_X1 U19043 ( .A1(n18235), .A2(n18064), .ZN(n18163) );
  INV_X1 U19044 ( .A(n18163), .ZN(n15718) );
  NOR2_X1 U19045 ( .A1(n17942), .A2(n15718), .ZN(n15713) );
  AOI211_X1 U19046 ( .C1(n18246), .C2(n17940), .A(n16450), .B(n15713), .ZN(
        n15789) );
  INV_X1 U19047 ( .A(n16436), .ZN(n16423) );
  NAND2_X1 U19048 ( .A1(n16423), .A2(n16425), .ZN(n15727) );
  INV_X1 U19049 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17566) );
  NOR2_X1 U19050 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16469) );
  AOI21_X1 U19051 ( .B1(n18156), .B2(n17566), .A(n16469), .ZN(n15720) );
  NAND2_X1 U19052 ( .A1(n15782), .A2(n17940), .ZN(n16417) );
  NOR2_X2 U19053 ( .A1(n9633), .A2(n18242), .ZN(n18237) );
  NOR2_X1 U19054 ( .A1(n17934), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18212) );
  AOI21_X1 U19055 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15717), .A(
        n17934), .ZN(n15714) );
  NOR3_X1 U19056 ( .A1(n18237), .A2(n18212), .A3(n15714), .ZN(n15716) );
  OR2_X1 U19057 ( .A1(n18731), .A2(n15715), .ZN(n17938) );
  OAI211_X1 U19058 ( .C1(n18243), .C2(n15717), .A(n15716), .B(n17938), .ZN(
        n16468) );
  NAND2_X1 U19059 ( .A1(n18229), .A2(n16468), .ZN(n16446) );
  OAI21_X1 U19060 ( .B1(n16437), .B2(n15718), .A(n16446), .ZN(n15719) );
  AOI21_X1 U19061 ( .B1(n18246), .B2(n16417), .A(n15719), .ZN(n15786) );
  OAI21_X1 U19062 ( .B1(n9633), .B2(n15720), .A(n15786), .ZN(n15725) );
  INV_X1 U19063 ( .A(n18171), .ZN(n18697) );
  NOR3_X4 U19064 ( .A1(n17416), .A2(n18697), .A3(n18235), .ZN(n18145) );
  NOR2_X1 U19065 ( .A1(n15722), .A2(n15721), .ZN(n15723) );
  XOR2_X1 U19066 ( .A(n15723), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16441) );
  INV_X1 U19067 ( .A(n16441), .ZN(n15724) );
  AOI22_X1 U19068 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15725), .B1(
        n18145), .B2(n15724), .ZN(n15726) );
  NAND2_X1 U19069 ( .A1(n9633), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16430) );
  OAI211_X1 U19070 ( .C1(n15789), .C2(n15727), .A(n15726), .B(n16430), .ZN(
        P3_U2833) );
  AOI21_X1 U19071 ( .B1(n15729), .B2(n15728), .A(n14195), .ZN(n19161) );
  AOI22_X1 U19072 ( .A1(n19161), .A2(n16350), .B1(n19338), .B2(n19003), .ZN(
        n15736) );
  INV_X1 U19073 ( .A(n15730), .ZN(n15734) );
  NOR2_X1 U19074 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n10874), .ZN(
        n15731) );
  AOI222_X1 U19075 ( .A1(n15734), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), 
        .B1(n16344), .B2(n15733), .C1(n15732), .C2(n15731), .ZN(n15735) );
  OAI211_X1 U19076 ( .C1(n19898), .C2(n19091), .A(n15736), .B(n15735), .ZN(
        P2_U3030) );
  AOI22_X1 U19077 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19130), .B1(n15737), 
        .B2(n19089), .ZN(n15745) );
  AOI22_X1 U19078 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19127), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19146), .ZN(n15744) );
  AOI22_X1 U19079 ( .A1(n15738), .A2(n19151), .B1(n16203), .B2(n19098), .ZN(
        n15743) );
  OAI211_X1 U19080 ( .C1(n15741), .C2(n15740), .A(n19123), .B(n15739), .ZN(
        n15742) );
  NAND4_X1 U19081 ( .A1(n15745), .A2(n15744), .A3(n15743), .A4(n15742), .ZN(
        P2_U2833) );
  INV_X1 U19082 ( .A(n15746), .ZN(n15756) );
  OR2_X1 U19083 ( .A1(n15748), .A2(n15747), .ZN(n15752) );
  AOI21_X1 U19084 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15750), .A(
        n15749), .ZN(n15751) );
  OAI211_X1 U19085 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15752), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15751), .ZN(n15754) );
  NAND2_X1 U19086 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15752), .ZN(
        n15753) );
  NAND2_X1 U19087 ( .A1(n15754), .A2(n15753), .ZN(n15755) );
  AOI222_X1 U19088 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15756), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15755), .C1(n15756), 
        .C2(n15755), .ZN(n15757) );
  AOI222_X1 U19089 ( .A1(n15758), .A2(n15757), .B1(n15758), .B2(n20590), .C1(
        n15757), .C2(n20590), .ZN(n15764) );
  OR2_X1 U19090 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15760) );
  AOI21_X1 U19091 ( .B1(n15761), .B2(n15760), .A(n15759), .ZN(n15762) );
  OAI211_X1 U19092 ( .C1(n15764), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15763), .B(n15762), .ZN(n15765) );
  NOR3_X1 U19093 ( .A1(n15767), .A2(n15766), .A3(n15765), .ZN(n15781) );
  AOI21_X1 U19094 ( .B1(n15768), .B2(n20671), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n16109) );
  NAND2_X1 U19095 ( .A1(n15768), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16102) );
  INV_X1 U19096 ( .A(n15769), .ZN(n15772) );
  AND2_X1 U19097 ( .A1(n15770), .A2(n20418), .ZN(n20934) );
  INV_X1 U19098 ( .A(n16102), .ZN(n20937) );
  INV_X1 U19099 ( .A(n20938), .ZN(n15771) );
  AND2_X1 U19100 ( .A1(n15779), .A2(n15771), .ZN(n20840) );
  AOI211_X1 U19101 ( .C1(n15772), .C2(n20934), .A(n20937), .B(n20840), .ZN(
        n16105) );
  OAI221_X1 U19102 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15781), 
        .A(n16105), .ZN(n15776) );
  NAND2_X1 U19103 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15776), .ZN(n16110) );
  AOI211_X1 U19104 ( .C1(n16109), .C2(n16102), .A(n15773), .B(n16110), .ZN(
        n15780) );
  NAND2_X1 U19105 ( .A1(n15775), .A2(n15774), .ZN(n15777) );
  AOI21_X1 U19106 ( .B1(n15777), .B2(n15776), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n15778) );
  AOI221_X1 U19107 ( .B1(n15781), .B2(n15780), .C1(n15779), .C2(n15780), .A(
        n15778), .ZN(P1_U3161) );
  NAND2_X1 U19108 ( .A1(n15782), .A2(n16444), .ZN(n16422) );
  NAND2_X1 U19109 ( .A1(n15784), .A2(n15783), .ZN(n15785) );
  XNOR2_X1 U19110 ( .A(n15785), .B(n16444), .ZN(n16418) );
  NAND2_X1 U19111 ( .A1(n18156), .A2(n18242), .ZN(n18230) );
  INV_X1 U19112 ( .A(n18230), .ZN(n18196) );
  NAND2_X1 U19113 ( .A1(n18196), .A2(n16445), .ZN(n16447) );
  AOI21_X1 U19114 ( .B1(n15786), .B2(n16447), .A(n16444), .ZN(n15787) );
  AOI21_X1 U19115 ( .B1(n18145), .B2(n16418), .A(n15787), .ZN(n15788) );
  NAND2_X1 U19116 ( .A1(n9633), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16413) );
  OAI211_X1 U19117 ( .C1(n15789), .C2(n16422), .A(n15788), .B(n16413), .ZN(
        P3_U2832) );
  INV_X1 U19118 ( .A(HOLD), .ZN(n19861) );
  NAND2_X1 U19119 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20841) );
  OAI21_X1 U19120 ( .B1(n19861), .B2(n20008), .A(n20841), .ZN(n15790) );
  OAI21_X1 U19121 ( .B1(n19861), .B2(n20857), .A(n15790), .ZN(n15792) );
  NAND2_X1 U19122 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20850), .ZN(n20848) );
  NAND3_X1 U19123 ( .A1(n15792), .A2(n15791), .A3(n20848), .ZN(P1_U3195) );
  INV_X1 U19124 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16566) );
  NOR2_X1 U19125 ( .A1(n20123), .A2(n16566), .ZN(P1_U2905) );
  NAND2_X1 U19126 ( .A1(n15794), .A2(n15793), .ZN(n15795) );
  XNOR2_X1 U19127 ( .A(n15795), .B(n15800), .ZN(n15910) );
  AOI221_X1 U19128 ( .B1(n15798), .B2(n15797), .C1(n15796), .C2(n15797), .A(
        n15988), .ZN(n15799) );
  AOI221_X1 U19129 ( .B1(n15993), .B2(n15800), .C1(n14716), .C2(n15800), .A(
        n15799), .ZN(n15801) );
  AOI21_X1 U19130 ( .B1(n15910), .B2(n20249), .A(n15801), .ZN(n15802) );
  NAND2_X1 U19131 ( .A1(n20209), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15911) );
  OAI211_X1 U19132 ( .C1(n20246), .C2(n15848), .A(n15802), .B(n15911), .ZN(
        P1_U3011) );
  NOR2_X1 U19133 ( .A1(n19864), .A2(n13085), .ZN(n19844) );
  AOI21_X1 U19134 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n13085), .A(n19844), 
        .ZN(n15804) );
  AOI221_X1 U19135 ( .B1(n15804), .B2(n19777), .C1(n15803), .C2(n19777), .A(
        n16411), .ZN(P2_U3178) );
  AOI221_X1 U19136 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16411), .C1(n19977), .C2(
        n16411), .A(n19788), .ZN(n19974) );
  INV_X1 U19137 ( .A(n19974), .ZN(n19971) );
  NOR2_X1 U19138 ( .A1(n16376), .A2(n19971), .ZN(P2_U3047) );
  NAND2_X1 U19139 ( .A1(n18296), .A2(n15811), .ZN(n17414) );
  INV_X1 U19140 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17510) );
  INV_X1 U19141 ( .A(n18708), .ZN(n15809) );
  AOI22_X1 U19142 ( .A1(n17442), .A2(BUF2_REG_0__SCAN_IN), .B1(n17423), .B2(
        n17926), .ZN(n15810) );
  OAI221_X1 U19143 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17414), .C1(n17510), 
        .C2(n15811), .A(n15810), .ZN(P3_U2735) );
  INV_X1 U19144 ( .A(n15823), .ZN(n15814) );
  NOR2_X1 U19145 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n20071), .ZN(n15812) );
  AOI22_X1 U19146 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15814), .B1(n15813), 
        .B2(n15812), .ZN(n15816) );
  AOI22_X1 U19147 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20103), .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n15815) );
  OAI211_X1 U19148 ( .C1(n15817), .C2(n20088), .A(n15816), .B(n15815), .ZN(
        n15818) );
  AOI21_X1 U19149 ( .B1(n15819), .B2(n20052), .A(n15818), .ZN(n15820) );
  OAI21_X1 U19150 ( .B1(n15821), .B2(n20101), .A(n15820), .ZN(P1_U2816) );
  AOI22_X1 U19151 ( .A1(n15877), .A2(n15822), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n20103), .ZN(n15828) );
  INV_X1 U19152 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20892) );
  NOR2_X1 U19153 ( .A1(n20892), .A2(n20890), .ZN(n15832) );
  AOI21_X1 U19154 ( .B1(n15832), .B2(n15830), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15824) );
  OAI22_X1 U19155 ( .A1(n15825), .A2(n15859), .B1(n15824), .B2(n15823), .ZN(
        n15826) );
  AOI21_X1 U19156 ( .B1(n20099), .B2(n15972), .A(n15826), .ZN(n15827) );
  OAI211_X1 U19157 ( .C1(n15829), .C2(n20102), .A(n15828), .B(n15827), .ZN(
        P1_U2817) );
  INV_X1 U19158 ( .A(n15830), .ZN(n15831) );
  AOI211_X1 U19159 ( .C1(n20892), .C2(n20890), .A(n15832), .B(n15831), .ZN(
        n15835) );
  OAI22_X1 U19160 ( .A1(n15840), .A2(n20892), .B1(n15833), .B2(n20034), .ZN(
        n15834) );
  AOI211_X1 U19161 ( .C1(n20095), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15835), .B(n15834), .ZN(n15838) );
  OAI22_X1 U19162 ( .A1(n15894), .A2(n15859), .B1(n20088), .B2(n15987), .ZN(
        n15836) );
  INV_X1 U19163 ( .A(n15836), .ZN(n15837) );
  OAI211_X1 U19164 ( .C1(n15901), .C2(n20101), .A(n15838), .B(n15837), .ZN(
        P1_U2818) );
  AOI21_X1 U19165 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15839), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n15841) );
  NOR2_X1 U19166 ( .A1(n15841), .A2(n15840), .ZN(n15845) );
  INV_X1 U19167 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15914) );
  INV_X1 U19168 ( .A(n15907), .ZN(n15842) );
  AOI22_X1 U19169 ( .A1(n15877), .A2(n15842), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n20103), .ZN(n15843) );
  OAI21_X1 U19170 ( .B1(n20102), .B2(n15914), .A(n15843), .ZN(n15844) );
  AOI211_X1 U19171 ( .C1(n15846), .C2(n20052), .A(n15845), .B(n15844), .ZN(
        n15847) );
  OAI21_X1 U19172 ( .B1(n20088), .B2(n15848), .A(n15847), .ZN(P1_U2820) );
  AOI21_X1 U19173 ( .B1(n20095), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20209), .ZN(n15850) );
  NAND2_X1 U19174 ( .A1(n20103), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n15849) );
  OAI211_X1 U19175 ( .C1(n20101), .C2(n15921), .A(n15850), .B(n15849), .ZN(
        n15852) );
  AOI211_X1 U19176 ( .C1(n15853), .C2(P1_REIP_REG_18__SCAN_IN), .A(n15852), 
        .B(n15851), .ZN(n15854) );
  INV_X1 U19177 ( .A(n15854), .ZN(n15855) );
  AOI21_X1 U19178 ( .B1(n15918), .B2(n20052), .A(n15855), .ZN(n15856) );
  OAI21_X1 U19179 ( .B1(n20088), .B2(n15995), .A(n15856), .ZN(P1_U2822) );
  AOI21_X1 U19180 ( .B1(n20095), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20209), .ZN(n15858) );
  NAND2_X1 U19181 ( .A1(n20103), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15857) );
  OAI211_X1 U19182 ( .C1(n20101), .C2(n15928), .A(n15858), .B(n15857), .ZN(
        n15861) );
  NOR2_X1 U19183 ( .A1(n15929), .A2(n15859), .ZN(n15860) );
  AOI211_X1 U19184 ( .C1(n15869), .C2(P1_REIP_REG_16__SCAN_IN), .A(n15861), 
        .B(n15860), .ZN(n15865) );
  OAI211_X1 U19185 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n15863), .B(n15862), .ZN(n15864) );
  OAI211_X1 U19186 ( .C1(n16020), .C2(n20088), .A(n15865), .B(n15864), .ZN(
        P1_U2824) );
  AOI22_X1 U19187 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20103), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n15874) );
  AOI21_X1 U19188 ( .B1(n15866), .B2(n20099), .A(n20209), .ZN(n15873) );
  INV_X1 U19189 ( .A(n15867), .ZN(n15934) );
  AOI22_X1 U19190 ( .A1(n15934), .A2(n20052), .B1(n15877), .B2(n15933), .ZN(
        n15872) );
  INV_X1 U19191 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20877) );
  NOR2_X1 U19192 ( .A1(n20877), .A2(n15868), .ZN(n15870) );
  OAI221_X1 U19193 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n15870), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(n15888), .A(n15869), .ZN(n15871) );
  NAND4_X1 U19194 ( .A1(n15874), .A2(n15873), .A3(n15872), .A4(n15871), .ZN(
        P1_U2826) );
  AOI22_X1 U19195 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20103), .B2(P1_EBX_REG_12__SCAN_IN), .ZN(n15882) );
  AOI21_X1 U19196 ( .B1(n15875), .B2(n20099), .A(n20209), .ZN(n15881) );
  INV_X1 U19197 ( .A(n15876), .ZN(n15938) );
  AOI22_X1 U19198 ( .A1(n15939), .A2(n15877), .B1(n20052), .B2(n15938), .ZN(
        n15880) );
  OAI221_X1 U19199 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n15888), .A(n15878), .ZN(n15879) );
  NAND4_X1 U19200 ( .A1(n15882), .A2(n15881), .A3(n15880), .A4(n15879), .ZN(
        P1_U2828) );
  OAI21_X1 U19201 ( .B1(n15884), .B2(n15883), .A(n14476), .ZN(n15891) );
  AOI22_X1 U19202 ( .A1(n20103), .A2(P1_EBX_REG_11__SCAN_IN), .B1(n15885), 
        .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15886) );
  OAI21_X1 U19203 ( .B1(n15891), .B2(n20088), .A(n15886), .ZN(n15887) );
  AOI211_X1 U19204 ( .C1(n20095), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20209), .B(n15887), .ZN(n15890) );
  INV_X1 U19205 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U19206 ( .A1(n15947), .A2(n20052), .B1(n15888), .B2(n20873), .ZN(
        n15889) );
  OAI211_X1 U19207 ( .C1(n15950), .C2(n20101), .A(n15890), .B(n15889), .ZN(
        P1_U2829) );
  INV_X1 U19208 ( .A(n15891), .ZN(n16038) );
  AOI22_X1 U19209 ( .A1(n15947), .A2(n20112), .B1(n20111), .B2(n16038), .ZN(
        n15892) );
  OAI21_X1 U19210 ( .B1(n20116), .B2(n15893), .A(n15892), .ZN(P1_U2861) );
  AOI22_X1 U19211 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15900) );
  INV_X1 U19212 ( .A(n15894), .ZN(n15898) );
  NAND2_X1 U19213 ( .A1(n15896), .A2(n15895), .ZN(n15897) );
  XNOR2_X1 U19214 ( .A(n15897), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15984) );
  AOI22_X1 U19215 ( .A1(n15898), .A2(n20189), .B1(n15984), .B2(n20200), .ZN(
        n15899) );
  OAI211_X1 U19216 ( .C1(n20193), .C2(n15901), .A(n15900), .B(n15899), .ZN(
        P1_U2977) );
  AOI22_X1 U19217 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15905) );
  AOI22_X1 U19218 ( .A1(n15903), .A2(n20189), .B1(n20199), .B2(n15902), .ZN(
        n15904) );
  OAI211_X1 U19219 ( .C1(n15906), .C2(n20016), .A(n15905), .B(n15904), .ZN(
        P1_U2978) );
  OAI22_X1 U19220 ( .A1(n15908), .A2(n20258), .B1(n15907), .B2(n20193), .ZN(
        n15909) );
  AOI21_X1 U19221 ( .B1(n20200), .B2(n15910), .A(n15909), .ZN(n15912) );
  OAI211_X1 U19222 ( .C1(n15914), .C2(n15913), .A(n15912), .B(n15911), .ZN(
        P1_U2979) );
  AOI22_X1 U19223 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15920) );
  OR2_X1 U19224 ( .A1(n15916), .A2(n15915), .ZN(n15917) );
  AND2_X1 U19225 ( .A1(n14714), .A2(n15917), .ZN(n15997) );
  AOI22_X1 U19226 ( .A1(n15918), .A2(n20189), .B1(n20200), .B2(n15997), .ZN(
        n15919) );
  OAI211_X1 U19227 ( .C1(n20193), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        P1_U2981) );
  NOR2_X1 U19228 ( .A1(n15923), .A2(n15922), .ZN(n15925) );
  NOR2_X1 U19229 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16012) );
  NOR2_X1 U19230 ( .A1(n15925), .A2(n16012), .ZN(n15927) );
  OAI22_X1 U19231 ( .A1(n15927), .A2(n15926), .B1(n15925), .B2(n15924), .ZN(
        n16016) );
  AOI22_X1 U19232 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15932) );
  OAI22_X1 U19233 ( .A1(n15929), .A2(n20258), .B1(n15928), .B2(n20193), .ZN(
        n15930) );
  INV_X1 U19234 ( .A(n15930), .ZN(n15931) );
  OAI211_X1 U19235 ( .C1(n20016), .C2(n16016), .A(n15932), .B(n15931), .ZN(
        P1_U2983) );
  AOI22_X1 U19236 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15936) );
  AOI22_X1 U19237 ( .A1(n15934), .A2(n20189), .B1(n20199), .B2(n15933), .ZN(
        n15935) );
  OAI211_X1 U19238 ( .C1(n15937), .C2(n20016), .A(n15936), .B(n15935), .ZN(
        P1_U2985) );
  AOI22_X1 U19239 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15941) );
  AOI22_X1 U19240 ( .A1(n20199), .A2(n15939), .B1(n20189), .B2(n15938), .ZN(
        n15940) );
  OAI211_X1 U19241 ( .C1(n15942), .C2(n20016), .A(n15941), .B(n15940), .ZN(
        P1_U2987) );
  AOI22_X1 U19242 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15949) );
  INV_X1 U19243 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16053) );
  NOR3_X1 U19244 ( .A1(n14723), .A2(n15943), .A3(n16053), .ZN(n15945) );
  NOR2_X1 U19245 ( .A1(n15945), .A2(n15944), .ZN(n15946) );
  XNOR2_X1 U19246 ( .A(n15946), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16040) );
  AOI22_X1 U19247 ( .A1(n20200), .A2(n16040), .B1(n20189), .B2(n15947), .ZN(
        n15948) );
  OAI211_X1 U19248 ( .C1(n20193), .C2(n15950), .A(n15949), .B(n15948), .ZN(
        P1_U2988) );
  AOI22_X1 U19249 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15956) );
  NAND2_X1 U19250 ( .A1(n15952), .A2(n15951), .ZN(n15953) );
  XNOR2_X1 U19251 ( .A(n15954), .B(n15953), .ZN(n16074) );
  AOI22_X1 U19252 ( .A1(n16074), .A2(n20200), .B1(n20189), .B2(n20041), .ZN(
        n15955) );
  OAI211_X1 U19253 ( .C1(n20193), .C2(n20044), .A(n15956), .B(n15955), .ZN(
        P1_U2992) );
  AOI22_X1 U19254 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15961) );
  XNOR2_X1 U19255 ( .A(n15957), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15958) );
  XNOR2_X1 U19256 ( .A(n15959), .B(n15958), .ZN(n16083) );
  AOI22_X1 U19257 ( .A1(n16083), .A2(n20200), .B1(n20189), .B2(n20051), .ZN(
        n15960) );
  OAI211_X1 U19258 ( .C1(n20193), .C2(n20054), .A(n15961), .B(n15960), .ZN(
        P1_U2993) );
  AOI22_X1 U19259 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15968) );
  OAI21_X1 U19260 ( .B1(n15964), .B2(n15963), .A(n15962), .ZN(n15965) );
  INV_X1 U19261 ( .A(n15965), .ZN(n16090) );
  INV_X1 U19262 ( .A(n15966), .ZN(n20113) );
  AOI22_X1 U19263 ( .A1(n16090), .A2(n20200), .B1(n20189), .B2(n20113), .ZN(
        n15967) );
  OAI211_X1 U19264 ( .C1(n20193), .C2(n20063), .A(n15968), .B(n15967), .ZN(
        P1_U2994) );
  INV_X1 U19265 ( .A(n15969), .ZN(n15976) );
  AOI22_X1 U19266 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n20209), .B1(n15970), 
        .B2(n12431), .ZN(n15975) );
  INV_X1 U19267 ( .A(n15971), .ZN(n15973) );
  AOI22_X1 U19268 ( .A1(n15973), .A2(n20249), .B1(n20235), .B2(n15972), .ZN(
        n15974) );
  OAI211_X1 U19269 ( .C1(n15976), .C2(n12431), .A(n15975), .B(n15974), .ZN(
        P1_U3008) );
  INV_X1 U19270 ( .A(n15977), .ZN(n15978) );
  AOI21_X1 U19271 ( .B1(n15980), .B2(n15979), .A(n15978), .ZN(n15982) );
  AOI22_X1 U19272 ( .A1(n20209), .A2(P1_REIP_REG_22__SCAN_IN), .B1(n15982), 
        .B2(n15981), .ZN(n15986) );
  AOI22_X1 U19273 ( .A1(n15984), .A2(n20249), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15983), .ZN(n15985) );
  OAI211_X1 U19274 ( .C1(n20246), .C2(n15987), .A(n15986), .B(n15985), .ZN(
        P1_U3009) );
  AOI22_X1 U19275 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15988), .B1(
        n20209), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15992) );
  AOI22_X1 U19276 ( .A1(n15990), .A2(n20249), .B1(n20235), .B2(n15989), .ZN(
        n15991) );
  OAI211_X1 U19277 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15993), .A(
        n15992), .B(n15991), .ZN(P1_U3012) );
  NAND2_X1 U19278 ( .A1(n15994), .A2(n16002), .ZN(n16000) );
  AOI21_X1 U19279 ( .B1(n16013), .B2(n16001), .A(n16033), .ZN(n16010) );
  OAI22_X1 U19280 ( .A1(n15995), .A2(n20246), .B1(n16010), .B2(n15994), .ZN(
        n15996) );
  AOI21_X1 U19281 ( .B1(n15997), .B2(n20249), .A(n15996), .ZN(n15999) );
  NAND2_X1 U19282 ( .A1(n20209), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15998) );
  OAI211_X1 U19283 ( .C1(n16001), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        P1_U3013) );
  NAND2_X1 U19284 ( .A1(n16002), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16027) );
  INV_X1 U19285 ( .A(n16027), .ZN(n16003) );
  AOI21_X1 U19286 ( .B1(n16011), .B2(n16003), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16009) );
  INV_X1 U19287 ( .A(n16004), .ZN(n16006) );
  AOI22_X1 U19288 ( .A1(n16006), .A2(n20249), .B1(n20235), .B2(n16005), .ZN(
        n16008) );
  NAND2_X1 U19289 ( .A1(n20209), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16007) );
  OAI211_X1 U19290 ( .C1(n16010), .C2(n16009), .A(n16008), .B(n16007), .ZN(
        P1_U3014) );
  NOR3_X1 U19291 ( .A1(n16012), .A2(n16011), .A3(n16027), .ZN(n16018) );
  AOI21_X1 U19292 ( .B1(n16014), .B2(n16013), .A(n16033), .ZN(n16021) );
  OAI22_X1 U19293 ( .A1(n16016), .A2(n20230), .B1(n16021), .B2(n16015), .ZN(
        n16017) );
  AOI211_X1 U19294 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(n20209), .A(n16018), 
        .B(n16017), .ZN(n16019) );
  OAI21_X1 U19295 ( .B1(n20246), .B2(n16020), .A(n16019), .ZN(P1_U3015) );
  INV_X1 U19296 ( .A(n16021), .ZN(n16022) );
  AOI22_X1 U19297 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16022), .B1(
        n20209), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16026) );
  AOI22_X1 U19298 ( .A1(n16024), .A2(n20249), .B1(n20235), .B2(n16023), .ZN(
        n16025) );
  OAI211_X1 U19299 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16027), .A(
        n16026), .B(n16025), .ZN(P1_U3016) );
  INV_X1 U19300 ( .A(n16028), .ZN(n16030) );
  AOI22_X1 U19301 ( .A1(n20209), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n16030), 
        .B2(n16029), .ZN(n16037) );
  AOI22_X1 U19302 ( .A1(n16032), .A2(n20249), .B1(n20235), .B2(n16031), .ZN(
        n16036) );
  OAI21_X1 U19303 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16034), .A(
        n16033), .ZN(n16035) );
  NAND3_X1 U19304 ( .A1(n16037), .A2(n16036), .A3(n16035), .ZN(P1_U3018) );
  AOI22_X1 U19305 ( .A1(n20209), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20235), 
        .B2(n16038), .ZN(n16042) );
  AOI22_X1 U19306 ( .A1(n16040), .A2(n20249), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16039), .ZN(n16041) );
  OAI211_X1 U19307 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16043), .A(
        n16042), .B(n16041), .ZN(P1_U3020) );
  INV_X1 U19308 ( .A(n16044), .ZN(n20224) );
  AOI21_X1 U19309 ( .B1(n20226), .B2(n16045), .A(n20224), .ZN(n16062) );
  NAND2_X1 U19310 ( .A1(n16046), .A2(n16062), .ZN(n16047) );
  OAI21_X1 U19311 ( .B1(n16061), .B2(n16047), .A(n16066), .ZN(n16059) );
  INV_X1 U19312 ( .A(n16048), .ZN(n16050) );
  AOI222_X1 U19313 ( .A1(n16050), .A2(n20249), .B1(n20235), .B2(n16049), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(n20209), .ZN(n16052) );
  OAI221_X1 U19314 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16053), .C2(n16060), .A(
        n16055), .ZN(n16051) );
  OAI211_X1 U19315 ( .C1(n16053), .C2(n16059), .A(n16052), .B(n16051), .ZN(
        P1_U3021) );
  AOI22_X1 U19316 ( .A1(n20209), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20235), 
        .B2(n16054), .ZN(n16058) );
  AOI22_X1 U19317 ( .A1(n16056), .A2(n20249), .B1(n16055), .B2(n16060), .ZN(
        n16057) );
  OAI211_X1 U19318 ( .C1(n16060), .C2(n16059), .A(n16058), .B(n16057), .ZN(
        P1_U3022) );
  NOR2_X1 U19319 ( .A1(n20210), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16089) );
  INV_X1 U19320 ( .A(n16089), .ZN(n16064) );
  AND2_X1 U19321 ( .A1(n16061), .A2(n20206), .ZN(n16063) );
  INV_X1 U19322 ( .A(n16062), .ZN(n20204) );
  AOI211_X1 U19323 ( .C1(n20226), .C2(n20210), .A(n16063), .B(n20204), .ZN(
        n16094) );
  OAI211_X1 U19324 ( .C1(n16065), .C2(n16064), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16094), .ZN(n16081) );
  NAND2_X1 U19325 ( .A1(n16066), .A2(n16081), .ZN(n16077) );
  OAI222_X1 U19326 ( .A1(n16068), .A2(n20246), .B1(n20244), .B2(n14095), .C1(
        n20230), .C2(n16067), .ZN(n16069) );
  INV_X1 U19327 ( .A(n16069), .ZN(n16071) );
  NOR2_X1 U19328 ( .A1(n16080), .A2(n16079), .ZN(n16073) );
  OAI221_X1 U19329 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16072), .C2(n16078), .A(
        n16073), .ZN(n16070) );
  OAI211_X1 U19330 ( .C1(n16077), .C2(n16072), .A(n16071), .B(n16070), .ZN(
        P1_U3023) );
  AOI22_X1 U19331 ( .A1(n20209), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20235), 
        .B2(n20037), .ZN(n16076) );
  AOI22_X1 U19332 ( .A1(n16074), .A2(n20249), .B1(n16073), .B2(n16078), .ZN(
        n16075) );
  OAI211_X1 U19333 ( .C1(n16078), .C2(n16077), .A(n16076), .B(n16075), .ZN(
        P1_U3024) );
  NAND2_X1 U19334 ( .A1(n16080), .A2(n16079), .ZN(n16082) );
  AOI22_X1 U19335 ( .A1(n16083), .A2(n20249), .B1(n16082), .B2(n16081), .ZN(
        n16085) );
  NAND2_X1 U19336 ( .A1(n20209), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n16084) );
  OAI211_X1 U19337 ( .C1(n20246), .C2(n20047), .A(n16085), .B(n16084), .ZN(
        P1_U3025) );
  AND2_X1 U19338 ( .A1(n16087), .A2(n16086), .ZN(n16088) );
  NOR2_X1 U19339 ( .A1(n14070), .A2(n16088), .ZN(n20110) );
  AOI22_X1 U19340 ( .A1(n20209), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20235), 
        .B2(n20110), .ZN(n16092) );
  AOI22_X1 U19341 ( .A1(n16090), .A2(n20249), .B1(n16089), .B2(n20216), .ZN(
        n16091) );
  OAI211_X1 U19342 ( .C1(n16094), .C2(n16093), .A(n16092), .B(n16091), .ZN(
        P1_U3026) );
  INV_X1 U19343 ( .A(n16095), .ZN(n16098) );
  NAND3_X1 U19344 ( .A1(n16098), .A2(n16097), .A3(n16096), .ZN(n16099) );
  OAI21_X1 U19345 ( .B1(n16101), .B2(n16100), .A(n16099), .ZN(P1_U3468) );
  NOR3_X1 U19346 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n9758), .A3(n16102), 
        .ZN(n16103) );
  NOR2_X1 U19347 ( .A1(n16104), .A2(n16103), .ZN(n20839) );
  AOI21_X1 U19348 ( .B1(n20839), .B2(n16106), .A(n16105), .ZN(n16107) );
  AOI221_X1 U19349 ( .B1(n16109), .B2(n16108), .C1(n16110), .C2(n16108), .A(
        n16107), .ZN(P1_U3162) );
  INV_X1 U19350 ( .A(n16110), .ZN(n16112) );
  OAI21_X1 U19351 ( .B1(n16112), .B2(n20671), .A(n16111), .ZN(P1_U3466) );
  AOI22_X1 U19352 ( .A1(n16113), .A2(n19089), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n19130), .ZN(n16122) );
  AOI22_X1 U19353 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19127), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n16114), .ZN(n16121) );
  INV_X1 U19354 ( .A(n16115), .ZN(n19154) );
  AOI22_X1 U19355 ( .A1(n19098), .A2(n19154), .B1(n19151), .B2(n16116), .ZN(
        n16120) );
  NAND4_X1 U19356 ( .A1(n19123), .A2(n16118), .A3(n9704), .A4(n16117), .ZN(
        n16119) );
  NAND4_X1 U19357 ( .A1(n16122), .A2(n16121), .A3(n16120), .A4(n16119), .ZN(
        P2_U2824) );
  AOI22_X1 U19358 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19130), .B1(n16123), 
        .B2(n19089), .ZN(n16133) );
  AOI22_X1 U19359 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19127), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19146), .ZN(n16132) );
  OAI22_X1 U19360 ( .A1(n16125), .A2(n19121), .B1(n16124), .B2(n19144), .ZN(
        n16126) );
  INV_X1 U19361 ( .A(n16126), .ZN(n16131) );
  OAI211_X1 U19362 ( .C1(n16129), .C2(n16128), .A(n19123), .B(n16127), .ZN(
        n16130) );
  NAND4_X1 U19363 ( .A1(n16133), .A2(n16132), .A3(n16131), .A4(n16130), .ZN(
        P2_U2826) );
  AOI22_X1 U19364 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19130), .B1(n16134), 
        .B2(n19089), .ZN(n16143) );
  AOI22_X1 U19365 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19146), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19127), .ZN(n16142) );
  AOI22_X1 U19366 ( .A1(n16136), .A2(n19151), .B1(n16135), .B2(n19098), .ZN(
        n16141) );
  OAI211_X1 U19367 ( .C1(n16139), .C2(n16138), .A(n19123), .B(n16137), .ZN(
        n16140) );
  NAND4_X1 U19368 ( .A1(n16143), .A2(n16142), .A3(n16141), .A4(n16140), .ZN(
        P2_U2827) );
  AOI22_X1 U19369 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19146), .B1(n16144), 
        .B2(n19089), .ZN(n16154) );
  AOI22_X1 U19370 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19127), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19130), .ZN(n16153) );
  OAI22_X1 U19371 ( .A1(n16146), .A2(n19121), .B1(n16145), .B2(n19144), .ZN(
        n16147) );
  INV_X1 U19372 ( .A(n16147), .ZN(n16152) );
  OAI211_X1 U19373 ( .C1(n16150), .C2(n16149), .A(n19123), .B(n16148), .ZN(
        n16151) );
  NAND4_X1 U19374 ( .A1(n16154), .A2(n16153), .A3(n16152), .A4(n16151), .ZN(
        P2_U2828) );
  AOI22_X1 U19375 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19130), .B1(n16155), 
        .B2(n19089), .ZN(n16164) );
  AOI22_X1 U19376 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19146), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19127), .ZN(n16163) );
  AOI22_X1 U19377 ( .A1(n16157), .A2(n19151), .B1(n16156), .B2(n19098), .ZN(
        n16162) );
  OAI211_X1 U19378 ( .C1(n16160), .C2(n16159), .A(n19123), .B(n16158), .ZN(
        n16161) );
  NAND4_X1 U19379 ( .A1(n16164), .A2(n16163), .A3(n16162), .A4(n16161), .ZN(
        P2_U2829) );
  AOI22_X1 U19380 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19130), .B1(n16165), 
        .B2(n19089), .ZN(n16175) );
  AOI22_X1 U19381 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19146), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19127), .ZN(n16174) );
  OAI22_X1 U19382 ( .A1(n16167), .A2(n19121), .B1(n16166), .B2(n19144), .ZN(
        n16168) );
  INV_X1 U19383 ( .A(n16168), .ZN(n16173) );
  OAI211_X1 U19384 ( .C1(n16171), .C2(n16170), .A(n19123), .B(n16169), .ZN(
        n16172) );
  NAND4_X1 U19385 ( .A1(n16175), .A2(n16174), .A3(n16173), .A4(n16172), .ZN(
        P2_U2830) );
  INV_X1 U19386 ( .A(n16177), .ZN(n16178) );
  OAI22_X1 U19387 ( .A1(n16178), .A2(n19149), .B1(n19911), .B2(n19142), .ZN(
        n16180) );
  OAI22_X1 U19388 ( .A1(n19115), .A2(n9810), .B1(n9979), .B2(n19139), .ZN(
        n16179) );
  AOI211_X1 U19389 ( .C1(n16197), .C2(n19098), .A(n16180), .B(n16179), .ZN(
        n16185) );
  OAI211_X1 U19390 ( .C1(n16183), .C2(n16182), .A(n19123), .B(n16181), .ZN(
        n16184) );
  OAI211_X1 U19391 ( .C1(n19121), .C2(n14316), .A(n16185), .B(n16184), .ZN(
        P2_U2831) );
  AOI22_X1 U19392 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19130), .B1(n16186), 
        .B2(n19089), .ZN(n16195) );
  AOI22_X1 U19393 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19127), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19146), .ZN(n16194) );
  AOI22_X1 U19394 ( .A1(n16188), .A2(n19151), .B1(n16187), .B2(n19098), .ZN(
        n16193) );
  OAI211_X1 U19395 ( .C1(n16191), .C2(n16190), .A(n19123), .B(n16189), .ZN(
        n16192) );
  NAND4_X1 U19396 ( .A1(n16195), .A2(n16194), .A3(n16193), .A4(n16192), .ZN(
        P2_U2832) );
  INV_X1 U19397 ( .A(n16196), .ZN(n19158) );
  AOI22_X1 U19398 ( .A1(n19158), .A2(n19183), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19205), .ZN(n16201) );
  AOI22_X1 U19399 ( .A1(n19160), .A2(BUF1_REG_24__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16200) );
  AOI22_X1 U19400 ( .A1(n16198), .A2(n19191), .B1(n19206), .B2(n16197), .ZN(
        n16199) );
  NAND3_X1 U19401 ( .A1(n16201), .A2(n16200), .A3(n16199), .ZN(P2_U2895) );
  INV_X1 U19402 ( .A(n19273), .ZN(n16202) );
  AOI22_X1 U19403 ( .A1(n19158), .A2(n16202), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19205), .ZN(n16207) );
  AOI22_X1 U19404 ( .A1(n19160), .A2(BUF1_REG_22__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16206) );
  AOI22_X1 U19405 ( .A1(n16204), .A2(n19191), .B1(n19206), .B2(n16203), .ZN(
        n16205) );
  NAND3_X1 U19406 ( .A1(n16207), .A2(n16206), .A3(n16205), .ZN(P2_U2897) );
  AOI22_X1 U19407 ( .A1(n19158), .A2(n19255), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19205), .ZN(n16211) );
  AOI22_X1 U19408 ( .A1(n19160), .A2(BUF1_REG_20__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16210) );
  AOI22_X1 U19409 ( .A1(n16208), .A2(n19191), .B1(n19206), .B2(n18953), .ZN(
        n16209) );
  NAND3_X1 U19410 ( .A1(n16211), .A2(n16210), .A3(n16209), .ZN(P2_U2899) );
  AOI22_X1 U19411 ( .A1(n19158), .A2(n19252), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19205), .ZN(n16215) );
  AOI22_X1 U19412 ( .A1(n19160), .A2(BUF1_REG_18__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16214) );
  AOI22_X1 U19413 ( .A1(n16212), .A2(n19191), .B1(n19206), .B2(n18976), .ZN(
        n16213) );
  NAND3_X1 U19414 ( .A1(n16215), .A2(n16214), .A3(n16213), .ZN(P2_U2901) );
  AOI22_X1 U19415 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19291), .B1(n19290), 
        .B2(n16216), .ZN(n16223) );
  NAND3_X1 U19416 ( .A1(n15349), .A2(n16217), .A3(n19318), .ZN(n16218) );
  OAI21_X1 U19417 ( .B1(n19305), .B2(n16219), .A(n16218), .ZN(n16220) );
  AOI21_X1 U19418 ( .B1(n16221), .B2(n16265), .A(n16220), .ZN(n16222) );
  OAI211_X1 U19419 ( .C1(n16224), .C2(n19312), .A(n16223), .B(n16222), .ZN(
        P2_U2991) );
  OAI22_X1 U19420 ( .A1(n18963), .A2(n19312), .B1(n19903), .B2(n19328), .ZN(
        n16225) );
  AOI21_X1 U19421 ( .B1(n19290), .B2(n16226), .A(n16225), .ZN(n16230) );
  AOI22_X1 U19422 ( .A1(n16228), .A2(n19318), .B1(n16265), .B2(n16227), .ZN(
        n16229) );
  OAI211_X1 U19423 ( .C1(n19305), .C2(n16231), .A(n16230), .B(n16229), .ZN(
        P2_U2995) );
  AOI22_X1 U19424 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19313), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19291), .ZN(n16236) );
  OAI22_X1 U19425 ( .A1(n16233), .A2(n19297), .B1(n19323), .B2(n16232), .ZN(
        n16234) );
  AOI21_X1 U19426 ( .B1(n19319), .B2(n18977), .A(n16234), .ZN(n16235) );
  OAI211_X1 U19427 ( .C1(n19304), .C2(n18980), .A(n16236), .B(n16235), .ZN(
        P2_U2996) );
  AOI22_X1 U19428 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19291), .B1(n19290), 
        .B2(n16237), .ZN(n16244) );
  NAND2_X1 U19429 ( .A1(n16238), .A2(n16265), .ZN(n16239) );
  OAI22_X1 U19430 ( .A1(n16240), .A2(n16239), .B1(n19305), .B2(n19013), .ZN(
        n16241) );
  AOI21_X1 U19431 ( .B1(n16242), .B2(n19318), .A(n16241), .ZN(n16243) );
  OAI211_X1 U19432 ( .C1(n19008), .C2(n19312), .A(n16244), .B(n16243), .ZN(
        P2_U2999) );
  AOI22_X1 U19433 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19291), .B1(n19290), 
        .B2(n19020), .ZN(n16255) );
  NAND2_X1 U19434 ( .A1(n16246), .A2(n16245), .ZN(n16247) );
  XNOR2_X1 U19435 ( .A(n16248), .B(n16247), .ZN(n16290) );
  INV_X1 U19436 ( .A(n16249), .ZN(n16250) );
  AOI21_X1 U19437 ( .B1(n16251), .B2(n9644), .A(n16250), .ZN(n16289) );
  AOI22_X1 U19438 ( .A1(n16290), .A2(n19318), .B1(n16265), .B2(n16289), .ZN(
        n16252) );
  INV_X1 U19439 ( .A(n16252), .ZN(n16253) );
  AOI21_X1 U19440 ( .B1(n19319), .B2(n19024), .A(n16253), .ZN(n16254) );
  OAI211_X1 U19441 ( .C1(n16256), .C2(n19312), .A(n16255), .B(n16254), .ZN(
        P2_U3000) );
  INV_X1 U19442 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19038) );
  OAI22_X1 U19443 ( .A1(n19038), .A2(n19312), .B1(n19304), .B2(n19032), .ZN(
        n16257) );
  AOI21_X1 U19444 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n19291), .A(n16257), 
        .ZN(n16261) );
  AOI22_X1 U19445 ( .A1(n16259), .A2(n19318), .B1(n16265), .B2(n16258), .ZN(
        n16260) );
  OAI211_X1 U19446 ( .C1(n19305), .C2(n19033), .A(n16261), .B(n16260), .ZN(
        P2_U3001) );
  INV_X1 U19447 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16262) );
  OAI22_X1 U19448 ( .A1(n16262), .A2(n19312), .B1(n19304), .B2(n19051), .ZN(
        n16263) );
  AOI21_X1 U19449 ( .B1(P2_REIP_REG_11__SCAN_IN), .B2(n19291), .A(n16263), 
        .ZN(n16268) );
  AOI22_X1 U19450 ( .A1(n16266), .A2(n16265), .B1(n19318), .B2(n16264), .ZN(
        n16267) );
  OAI211_X1 U19451 ( .C1(n19305), .C2(n19054), .A(n16268), .B(n16267), .ZN(
        P2_U3003) );
  AOI22_X1 U19452 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19291), .B1(n19290), 
        .B2(n19064), .ZN(n16283) );
  NAND2_X1 U19453 ( .A1(n15240), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16270) );
  NAND2_X1 U19454 ( .A1(n16270), .A2(n16269), .ZN(n16272) );
  INV_X1 U19455 ( .A(n16316), .ZN(n16279) );
  NOR2_X1 U19456 ( .A1(n16274), .A2(n16273), .ZN(n16278) );
  NAND2_X1 U19457 ( .A1(n16276), .A2(n16275), .ZN(n16277) );
  XNOR2_X1 U19458 ( .A(n16278), .B(n16277), .ZN(n16318) );
  OAI22_X1 U19459 ( .A1(n16279), .A2(n19323), .B1(n16318), .B2(n19297), .ZN(
        n16280) );
  AOI21_X1 U19460 ( .B1(n19319), .B2(n16281), .A(n16280), .ZN(n16282) );
  OAI211_X1 U19461 ( .C1(n16284), .C2(n19312), .A(n16283), .B(n16282), .ZN(
        P2_U3004) );
  AOI21_X1 U19462 ( .B1(n15456), .B2(n16285), .A(n15444), .ZN(n19169) );
  NOR3_X1 U19463 ( .A1(n16287), .A2(n16286), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16288) );
  AOI21_X1 U19464 ( .B1(n19169), .B2(n16350), .A(n16288), .ZN(n16296) );
  AOI222_X1 U19465 ( .A1(n16290), .A2(n16344), .B1(n19338), .B2(n19024), .C1(
        n16329), .C2(n16289), .ZN(n16295) );
  NAND2_X1 U19466 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19291), .ZN(n16294) );
  OAI21_X1 U19467 ( .B1(n16292), .B2(n16291), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16293) );
  NAND4_X1 U19468 ( .A1(n16296), .A2(n16295), .A3(n16294), .A4(n16293), .ZN(
        P2_U3032) );
  AOI21_X1 U19469 ( .B1(n15475), .B2(n16297), .A(n15455), .ZN(n19174) );
  NAND2_X1 U19470 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19291), .ZN(n16298) );
  OAI211_X1 U19471 ( .C1(n16301), .C2(n16300), .A(n16299), .B(n16298), .ZN(
        n16302) );
  AOI21_X1 U19472 ( .B1(n16350), .B2(n19174), .A(n16302), .ZN(n16305) );
  AOI22_X1 U19473 ( .A1(n16303), .A2(n16344), .B1(n19338), .B2(n19045), .ZN(
        n16304) );
  OAI211_X1 U19474 ( .C1(n19343), .C2(n16306), .A(n16305), .B(n16304), .ZN(
        P2_U3034) );
  NAND2_X1 U19475 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16307), .ZN(
        n16310) );
  NAND2_X1 U19476 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19291), .ZN(n16308) );
  OAI221_X1 U19477 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16310), 
        .C1(n16269), .C2(n16309), .A(n16308), .ZN(n16314) );
  AOI21_X1 U19478 ( .B1(n15489), .B2(n16311), .A(n15474), .ZN(n19177) );
  NAND2_X1 U19479 ( .A1(n19177), .A2(n16350), .ZN(n16312) );
  OAI21_X1 U19480 ( .B1(n16341), .B2(n19068), .A(n16312), .ZN(n16313) );
  OR2_X1 U19481 ( .A1(n16314), .A2(n16313), .ZN(n16315) );
  AOI21_X1 U19482 ( .B1(n16316), .B2(n16329), .A(n16315), .ZN(n16317) );
  OAI21_X1 U19483 ( .B1(n16318), .B2(n19331), .A(n16317), .ZN(P2_U3036) );
  AOI21_X1 U19484 ( .B1(n16320), .B2(n16319), .A(n15488), .ZN(n19182) );
  NOR2_X1 U19485 ( .A1(n19091), .A2(n19884), .ZN(n16328) );
  OAI21_X1 U19486 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16334), .ZN(n16325) );
  INV_X1 U19487 ( .A(n16321), .ZN(n16322) );
  NOR2_X1 U19488 ( .A1(n16323), .A2(n16322), .ZN(n16336) );
  OAI22_X1 U19489 ( .A1(n16326), .A2(n16325), .B1(n16336), .B2(n16324), .ZN(
        n16327) );
  AOI211_X1 U19490 ( .C1(n16350), .C2(n19182), .A(n16328), .B(n16327), .ZN(
        n16332) );
  AOI22_X1 U19491 ( .A1(n16330), .A2(n16329), .B1(n19338), .B2(n19085), .ZN(
        n16331) );
  OAI211_X1 U19492 ( .C1(n16333), .C2(n19331), .A(n16332), .B(n16331), .ZN(
        P2_U3038) );
  INV_X1 U19493 ( .A(n16334), .ZN(n16338) );
  NAND2_X1 U19494 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19291), .ZN(n16335) );
  OAI221_X1 U19495 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16338), .C1(
        n16337), .C2(n16336), .A(n16335), .ZN(n16343) );
  XOR2_X1 U19496 ( .A(n16339), .B(n16340), .Z(n19097) );
  INV_X1 U19497 ( .A(n19097), .ZN(n19186) );
  OAI22_X1 U19498 ( .A1(n19186), .A2(n19330), .B1(n16341), .B2(n19102), .ZN(
        n16342) );
  AOI211_X1 U19499 ( .C1(n16345), .C2(n16344), .A(n16343), .B(n16342), .ZN(
        n16346) );
  OAI21_X1 U19500 ( .B1(n19343), .B2(n16347), .A(n16346), .ZN(P2_U3039) );
  AOI22_X1 U19501 ( .A1(n16350), .A2(n16349), .B1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16348), .ZN(n16358) );
  NOR2_X1 U19502 ( .A1(n19091), .A2(n10242), .ZN(n19316) );
  NAND2_X1 U19503 ( .A1(n19148), .A2(n16351), .ZN(n16352) );
  NAND2_X1 U19504 ( .A1(n16353), .A2(n16352), .ZN(n19315) );
  OAI21_X1 U19505 ( .B1(n16355), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16354), .ZN(n19324) );
  OAI22_X1 U19506 ( .A1(n19331), .A2(n19315), .B1(n19343), .B2(n19324), .ZN(
        n16356) );
  AOI211_X1 U19507 ( .C1(n19338), .C2(n19320), .A(n19316), .B(n16356), .ZN(
        n16357) );
  OAI211_X1 U19508 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16359), .A(
        n16358), .B(n16357), .ZN(P2_U3046) );
  OAI21_X1 U19509 ( .B1(n16392), .B2(n16360), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16361) );
  OAI21_X1 U19510 ( .B1(n16362), .B2(n16392), .A(n16361), .ZN(n16363) );
  INV_X1 U19511 ( .A(n16363), .ZN(n16396) );
  NAND2_X1 U19512 ( .A1(n16392), .A2(n16364), .ZN(n16365) );
  OAI21_X1 U19513 ( .B1(n16373), .B2(n16392), .A(n16365), .ZN(n16395) );
  INV_X1 U19514 ( .A(n16366), .ZN(n16371) );
  OAI21_X1 U19515 ( .B1(n16368), .B2(n19973), .A(n16367), .ZN(n16370) );
  NOR2_X1 U19516 ( .A1(n16368), .A2(n10498), .ZN(n16369) );
  AOI211_X1 U19517 ( .C1(n16371), .C2(n16370), .A(n16392), .B(n16369), .ZN(
        n16372) );
  OAI21_X1 U19518 ( .B1(n19957), .B2(n16373), .A(n16372), .ZN(n16374) );
  AOI21_X1 U19519 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16396), .A(
        n16374), .ZN(n16378) );
  OAI22_X1 U19520 ( .A1(n16396), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n16375), .B2(n16395), .ZN(n16377) );
  OAI21_X1 U19521 ( .B1(n16378), .B2(n16377), .A(n16376), .ZN(n16394) );
  OAI21_X1 U19522 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16379), .ZN(n16382) );
  OR3_X1 U19523 ( .A1(n10767), .A2(n16380), .A3(n19997), .ZN(n16381) );
  OAI211_X1 U19524 ( .C1(n16384), .C2(n16383), .A(n16382), .B(n16381), .ZN(
        n16391) );
  INV_X1 U19525 ( .A(n16385), .ZN(n16390) );
  AOI22_X1 U19526 ( .A1(n16389), .A2(n16387), .B1(n11189), .B2(n16386), .ZN(
        n16388) );
  OAI21_X1 U19527 ( .B1(n16390), .B2(n16389), .A(n16388), .ZN(n19981) );
  AOI211_X1 U19528 ( .C1(n16392), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16391), .B(n19981), .ZN(n16393) );
  OAI211_X1 U19529 ( .C1(n16396), .C2(n16395), .A(n16394), .B(n16393), .ZN(
        n16407) );
  OAI21_X1 U19530 ( .B1(n16407), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16400) );
  AOI211_X1 U19531 ( .C1(n16398), .C2(n16397), .A(n19987), .B(n19777), .ZN(
        n16399) );
  AND2_X1 U19532 ( .A1(n16400), .A2(n16399), .ZN(n19849) );
  INV_X1 U19533 ( .A(n16401), .ZN(n16403) );
  NOR2_X1 U19534 ( .A1(n16403), .A2(n16402), .ZN(n19968) );
  AOI211_X1 U19535 ( .C1(n19864), .C2(n19777), .A(n19849), .B(n19968), .ZN(
        n16410) );
  AOI21_X1 U19536 ( .B1(n13085), .B2(n16404), .A(n19992), .ZN(n16405) );
  AOI21_X1 U19537 ( .B1(n19849), .B2(n19864), .A(n16405), .ZN(n16406) );
  AOI21_X1 U19538 ( .B1(n19843), .B2(n16407), .A(n16406), .ZN(n16409) );
  OAI211_X1 U19539 ( .C1(n16410), .C2(n13085), .A(n16409), .B(n16408), .ZN(
        P2_U3176) );
  AOI221_X1 U19540 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13085), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19849), .A(n16411), .ZN(n16412) );
  INV_X1 U19541 ( .A(n16412), .ZN(P2_U3593) );
  INV_X1 U19542 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17625) );
  INV_X1 U19543 ( .A(n17623), .ZN(n17624) );
  INV_X1 U19544 ( .A(n18117), .ZN(n17778) );
  AOI22_X2 U19545 ( .A1(n17842), .A2(n17777), .B1(n17916), .B2(n17778), .ZN(
        n17832) );
  NOR2_X2 U19546 ( .A1(n17832), .A2(n18045), .ZN(n17723) );
  INV_X1 U19547 ( .A(n17723), .ZN(n17738) );
  NAND2_X1 U19548 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17592), .ZN(
        n17564) );
  XOR2_X1 U19549 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16426), .Z(
        n16609) );
  INV_X1 U19550 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16610) );
  OAI221_X1 U19551 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16415), .C1(
        n16610), .C2(n16414), .A(n16413), .ZN(n16416) );
  AOI21_X1 U19552 ( .B1(n17789), .B2(n16609), .A(n16416), .ZN(n16421) );
  INV_X1 U19553 ( .A(n17842), .ZN(n17761) );
  NAND2_X1 U19554 ( .A1(n17916), .A2(n16417), .ZN(n16424) );
  OAI21_X1 U19555 ( .B1(n16437), .B2(n17761), .A(n16424), .ZN(n16419) );
  AOI22_X1 U19556 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16419), .B1(
        n17829), .B2(n16418), .ZN(n16420) );
  OAI211_X1 U19557 ( .C1(n17564), .C2(n16422), .A(n16421), .B(n16420), .ZN(
        P3_U2800) );
  NAND2_X1 U19558 ( .A1(n16423), .A2(n17940), .ZN(n16470) );
  AOI21_X1 U19559 ( .B1(n16425), .B2(n16470), .A(n16424), .ZN(n16434) );
  INV_X1 U19560 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16620) );
  INV_X1 U19561 ( .A(n16595), .ZN(n16427) );
  AOI21_X1 U19562 ( .B1(n16620), .B2(n16427), .A(n16426), .ZN(n16619) );
  OAI21_X1 U19563 ( .B1(n16428), .B2(n17789), .A(n16619), .ZN(n16429) );
  OAI211_X1 U19564 ( .C1(n16432), .C2(n16431), .A(n16430), .B(n16429), .ZN(
        n16433) );
  AOI211_X1 U19565 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16435), .A(
        n16434), .B(n16433), .ZN(n16440) );
  NOR2_X1 U19566 ( .A1(n17942), .A2(n16436), .ZN(n16472) );
  NOR2_X1 U19567 ( .A1(n16437), .A2(n17761), .ZN(n16438) );
  OAI21_X1 U19568 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16472), .A(
        n16438), .ZN(n16439) );
  OAI211_X1 U19569 ( .C1(n16441), .C2(n17845), .A(n16440), .B(n16439), .ZN(
        P3_U2801) );
  INV_X1 U19570 ( .A(n18246), .ZN(n18240) );
  OAI21_X1 U19571 ( .B1(n16442), .B2(n18230), .A(n18240), .ZN(n16443) );
  INV_X1 U19572 ( .A(n16443), .ZN(n16456) );
  NOR3_X1 U19573 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16445), .A3(
        n16444), .ZN(n16451) );
  INV_X1 U19574 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18860) );
  AOI21_X1 U19575 ( .B1(n16447), .B2(n16446), .A(n18860), .ZN(n16448) );
  AOI211_X1 U19576 ( .C1(n16451), .C2(n16450), .A(n16449), .B(n16448), .ZN(
        n16455) );
  AOI22_X1 U19577 ( .A1(n16453), .A2(n18163), .B1(n16452), .B2(n18145), .ZN(
        n16454) );
  OAI211_X1 U19578 ( .C1(n16457), .C2(n16456), .A(n16455), .B(n16454), .ZN(
        P3_U2831) );
  NAND2_X1 U19579 ( .A1(n9633), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17577) );
  NOR2_X1 U19580 ( .A1(n17834), .A2(n16458), .ZN(n16461) );
  AOI22_X1 U19581 ( .A1(n15702), .A2(n17778), .B1(n17777), .B2(n18116), .ZN(
        n18044) );
  NOR2_X1 U19582 ( .A1(n18137), .A2(n16459), .ZN(n17935) );
  AOI22_X1 U19583 ( .A1(n18691), .A2(n18034), .B1(n18217), .B2(n17935), .ZN(
        n17960) );
  OAI21_X1 U19584 ( .B1(n18044), .B2(n16459), .A(n17960), .ZN(n18001) );
  NAND2_X1 U19585 ( .A1(n17958), .A2(n18001), .ZN(n17987) );
  NOR2_X1 U19586 ( .A1(n16460), .A2(n17987), .ZN(n17945) );
  NOR2_X1 U19587 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17944), .ZN(
        n17573) );
  OAI211_X1 U19588 ( .C1(n16461), .C2(n17945), .A(n18242), .B(n17573), .ZN(
        n16477) );
  OAI21_X1 U19589 ( .B1(n17745), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16462), .ZN(n17569) );
  NAND3_X1 U19590 ( .A1(n18145), .A2(n16463), .A3(n17569), .ZN(n16476) );
  INV_X1 U19591 ( .A(n17581), .ZN(n16467) );
  NOR2_X1 U19592 ( .A1(n17570), .A2(n17569), .ZN(n17568) );
  NAND2_X1 U19593 ( .A1(n18171), .A2(n16464), .ZN(n16465) );
  AOI211_X1 U19594 ( .C1(n16467), .C2(n16466), .A(n17568), .B(n16465), .ZN(
        n16474) );
  AOI211_X1 U19595 ( .C1(n15702), .C2(n16470), .A(n16469), .B(n16468), .ZN(
        n16471) );
  OAI21_X1 U19596 ( .B1(n16472), .B2(n18064), .A(n16471), .ZN(n16473) );
  OAI211_X1 U19597 ( .C1(n16474), .C2(n16473), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18229), .ZN(n16475) );
  NAND4_X1 U19598 ( .A1(n17577), .A2(n16477), .A3(n16476), .A4(n16475), .ZN(
        P3_U2834) );
  NOR3_X1 U19599 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16479) );
  NOR4_X1 U19600 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16478) );
  NAND4_X1 U19601 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16479), .A3(n16478), .A4(
        U215), .ZN(U213) );
  INV_X1 U19602 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19215) );
  INV_X2 U19603 ( .A(U214), .ZN(n16525) );
  NOR2_X1 U19604 ( .A1(n16525), .A2(n16480), .ZN(n16523) );
  OAI222_X1 U19605 ( .A1(U212), .A2(n19215), .B1(n16528), .B2(n16481), .C1(
        U214), .C2(n16566), .ZN(U216) );
  INV_X1 U19606 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16483) );
  INV_X1 U19607 ( .A(U212), .ZN(n16526) );
  AOI22_X1 U19608 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16525), .ZN(n16482) );
  OAI21_X1 U19609 ( .B1(n16483), .B2(n16528), .A(n16482), .ZN(U217) );
  AOI22_X1 U19610 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16525), .ZN(n16484) );
  OAI21_X1 U19611 ( .B1(n16485), .B2(n16528), .A(n16484), .ZN(U218) );
  INV_X1 U19612 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16487) );
  AOI22_X1 U19613 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16525), .ZN(n16486) );
  OAI21_X1 U19614 ( .B1(n16487), .B2(n16528), .A(n16486), .ZN(U219) );
  AOI22_X1 U19615 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16525), .ZN(n16488) );
  OAI21_X1 U19616 ( .B1(n15060), .B2(n16528), .A(n16488), .ZN(U220) );
  AOI22_X1 U19617 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16525), .ZN(n16489) );
  OAI21_X1 U19618 ( .B1(n16490), .B2(n16528), .A(n16489), .ZN(U221) );
  AOI222_X1 U19619 ( .A1(n16525), .A2(P1_DATAO_REG_25__SCAN_IN), .B1(n16523), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n16526), .C2(P2_DATAO_REG_25__SCAN_IN), 
        .ZN(n16491) );
  INV_X1 U19620 ( .A(n16491), .ZN(U222) );
  AOI22_X1 U19621 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16525), .ZN(n16492) );
  OAI21_X1 U19622 ( .B1(n16493), .B2(n16528), .A(n16492), .ZN(U223) );
  AOI22_X1 U19623 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16525), .ZN(n16494) );
  OAI21_X1 U19624 ( .B1(n21103), .B2(n16528), .A(n16494), .ZN(U224) );
  INV_X1 U19625 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16496) );
  AOI22_X1 U19626 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16525), .ZN(n16495) );
  OAI21_X1 U19627 ( .B1(n16496), .B2(n16528), .A(n16495), .ZN(U225) );
  AOI22_X1 U19628 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16525), .ZN(n16497) );
  OAI21_X1 U19629 ( .B1(n15099), .B2(n16528), .A(n16497), .ZN(U226) );
  INV_X1 U19630 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19369) );
  AOI22_X1 U19631 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16525), .ZN(n16498) );
  OAI21_X1 U19632 ( .B1(n19369), .B2(n16528), .A(n16498), .ZN(U227) );
  AOI22_X1 U19633 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16525), .ZN(n16499) );
  OAI21_X1 U19634 ( .B1(n15111), .B2(n16528), .A(n16499), .ZN(U228) );
  AOI22_X1 U19635 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16525), .ZN(n16500) );
  OAI21_X1 U19636 ( .B1(n19355), .B2(n16528), .A(n16500), .ZN(U229) );
  AOI22_X1 U19637 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16525), .ZN(n16501) );
  OAI21_X1 U19638 ( .B1(n14200), .B2(n16528), .A(n16501), .ZN(U230) );
  AOI22_X1 U19639 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16525), .ZN(n16502) );
  OAI21_X1 U19640 ( .B1(n16503), .B2(n16528), .A(n16502), .ZN(U231) );
  AOI22_X1 U19641 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16525), .ZN(n16504) );
  OAI21_X1 U19642 ( .B1(n13622), .B2(n16528), .A(n16504), .ZN(U232) );
  AOI22_X1 U19643 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16525), .ZN(n16505) );
  OAI21_X1 U19644 ( .B1(n14569), .B2(n16528), .A(n16505), .ZN(U233) );
  AOI22_X1 U19645 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16525), .ZN(n16506) );
  OAI21_X1 U19646 ( .B1(n14349), .B2(n16528), .A(n16506), .ZN(U234) );
  INV_X1 U19647 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n21055) );
  AOI22_X1 U19648 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16523), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16526), .ZN(n16507) );
  OAI21_X1 U19649 ( .B1(n21055), .B2(U214), .A(n16507), .ZN(U235) );
  INV_X1 U19650 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16542) );
  AOI22_X1 U19651 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16523), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16525), .ZN(n16508) );
  OAI21_X1 U19652 ( .B1(n16542), .B2(U212), .A(n16508), .ZN(U236) );
  AOI22_X1 U19653 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16525), .ZN(n16509) );
  OAI21_X1 U19654 ( .B1(n16510), .B2(n16528), .A(n16509), .ZN(U237) );
  INV_X1 U19655 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16540) );
  AOI22_X1 U19656 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16523), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16525), .ZN(n16511) );
  OAI21_X1 U19657 ( .B1(n16540), .B2(U212), .A(n16511), .ZN(U238) );
  AOI22_X1 U19658 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16525), .ZN(n16512) );
  OAI21_X1 U19659 ( .B1(n16513), .B2(n16528), .A(n16512), .ZN(U239) );
  INV_X1 U19660 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16537) );
  AOI22_X1 U19661 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16523), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16525), .ZN(n16514) );
  OAI21_X1 U19662 ( .B1(n16537), .B2(U212), .A(n16514), .ZN(U240) );
  INV_X1 U19663 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16516) );
  AOI22_X1 U19664 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16525), .ZN(n16515) );
  OAI21_X1 U19665 ( .B1(n16516), .B2(n16528), .A(n16515), .ZN(U241) );
  INV_X1 U19666 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16535) );
  AOI22_X1 U19667 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16523), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16525), .ZN(n16517) );
  OAI21_X1 U19668 ( .B1(n16535), .B2(U212), .A(n16517), .ZN(U242) );
  AOI22_X1 U19669 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16525), .ZN(n16518) );
  OAI21_X1 U19670 ( .B1(n16519), .B2(n16528), .A(n16518), .ZN(U243) );
  INV_X1 U19671 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16533) );
  AOI22_X1 U19672 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16523), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16525), .ZN(n16520) );
  OAI21_X1 U19673 ( .B1(n16533), .B2(U212), .A(n16520), .ZN(U244) );
  AOI22_X1 U19674 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16525), .ZN(n16521) );
  OAI21_X1 U19675 ( .B1(n16522), .B2(n16528), .A(n16521), .ZN(U245) );
  INV_X1 U19676 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16531) );
  AOI22_X1 U19677 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16523), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16525), .ZN(n16524) );
  OAI21_X1 U19678 ( .B1(n16531), .B2(U212), .A(n16524), .ZN(U246) );
  AOI22_X1 U19679 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16526), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16525), .ZN(n16527) );
  OAI21_X1 U19680 ( .B1(n16529), .B2(n16528), .A(n16527), .ZN(U247) );
  INV_X1 U19681 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16530) );
  AOI22_X1 U19682 ( .A1(n16563), .A2(n16530), .B1(n18263), .B2(U215), .ZN(U251) );
  INV_X1 U19683 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n21108) );
  AOI22_X1 U19684 ( .A1(n16563), .A2(n16531), .B1(n21108), .B2(U215), .ZN(U252) );
  INV_X1 U19685 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16532) );
  AOI22_X1 U19686 ( .A1(n16563), .A2(n16532), .B1(n18271), .B2(U215), .ZN(U253) );
  INV_X1 U19687 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U19688 ( .A1(n16563), .A2(n16533), .B1(n18276), .B2(U215), .ZN(U254) );
  INV_X1 U19689 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16534) );
  AOI22_X1 U19690 ( .A1(n16563), .A2(n16534), .B1(n18280), .B2(U215), .ZN(U255) );
  INV_X1 U19691 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18284) );
  AOI22_X1 U19692 ( .A1(n16563), .A2(n16535), .B1(n18284), .B2(U215), .ZN(U256) );
  INV_X1 U19693 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16536) );
  INV_X1 U19694 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18288) );
  AOI22_X1 U19695 ( .A1(n16557), .A2(n16536), .B1(n18288), .B2(U215), .ZN(U257) );
  INV_X1 U19696 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18293) );
  AOI22_X1 U19697 ( .A1(n16557), .A2(n16537), .B1(n18293), .B2(U215), .ZN(U258) );
  INV_X1 U19698 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16538) );
  AOI22_X1 U19699 ( .A1(n16563), .A2(n16538), .B1(n17541), .B2(U215), .ZN(U259) );
  INV_X1 U19700 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n16539) );
  AOI22_X1 U19701 ( .A1(n16563), .A2(n16540), .B1(n16539), .B2(U215), .ZN(U260) );
  INV_X1 U19702 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16541) );
  INV_X1 U19703 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17546) );
  AOI22_X1 U19704 ( .A1(n16557), .A2(n16541), .B1(n17546), .B2(U215), .ZN(U261) );
  INV_X1 U19705 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17548) );
  AOI22_X1 U19706 ( .A1(n16563), .A2(n16542), .B1(n17548), .B2(U215), .ZN(U262) );
  INV_X1 U19707 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16543) );
  INV_X1 U19708 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U19709 ( .A1(n16557), .A2(n16543), .B1(n17550), .B2(U215), .ZN(U263) );
  INV_X1 U19710 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16544) );
  INV_X1 U19711 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U19712 ( .A1(n16563), .A2(n16544), .B1(n17554), .B2(U215), .ZN(U264) );
  OAI22_X1 U19713 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16563), .ZN(n16545) );
  INV_X1 U19714 ( .A(n16545), .ZN(U265) );
  OAI22_X1 U19715 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16557), .ZN(n16546) );
  INV_X1 U19716 ( .A(n16546), .ZN(U266) );
  INV_X1 U19717 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n16547) );
  AOI22_X1 U19718 ( .A1(n16557), .A2(n16547), .B1(n18265), .B2(U215), .ZN(U267) );
  OAI22_X1 U19719 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16563), .ZN(n16548) );
  INV_X1 U19720 ( .A(n16548), .ZN(U268) );
  INV_X1 U19721 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16549) );
  INV_X1 U19722 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19354) );
  AOI22_X1 U19723 ( .A1(n16563), .A2(n16549), .B1(n19354), .B2(U215), .ZN(U269) );
  INV_X1 U19724 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n16550) );
  AOI22_X1 U19725 ( .A1(n16557), .A2(n16550), .B1(n15109), .B2(U215), .ZN(U270) );
  INV_X1 U19726 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16551) );
  INV_X1 U19727 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19367) );
  AOI22_X1 U19728 ( .A1(n16557), .A2(n16551), .B1(n19367), .B2(U215), .ZN(U271) );
  OAI22_X1 U19729 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16563), .ZN(n16552) );
  INV_X1 U19730 ( .A(n16552), .ZN(U272) );
  OAI22_X1 U19731 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16563), .ZN(n16553) );
  INV_X1 U19732 ( .A(n16553), .ZN(U273) );
  INV_X1 U19733 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16554) );
  AOI22_X1 U19734 ( .A1(n16563), .A2(n16554), .B1(n18292), .B2(U215), .ZN(U274) );
  OAI22_X1 U19735 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16557), .ZN(n16555) );
  INV_X1 U19736 ( .A(n16555), .ZN(U275) );
  AOI22_X1 U19737 ( .A1(n16563), .A2(n16556), .B1(n15079), .B2(U215), .ZN(U276) );
  OAI22_X1 U19738 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16557), .ZN(n16558) );
  INV_X1 U19739 ( .A(n16558), .ZN(U277) );
  OAI22_X1 U19740 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16563), .ZN(n16559) );
  INV_X1 U19741 ( .A(n16559), .ZN(U278) );
  OAI22_X1 U19742 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16563), .ZN(n16560) );
  INV_X1 U19743 ( .A(n16560), .ZN(U279) );
  INV_X1 U19744 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16561) );
  AOI22_X1 U19745 ( .A1(n16563), .A2(n16561), .B1(n17310), .B2(U215), .ZN(U280) );
  OAI22_X1 U19746 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16563), .ZN(n16562) );
  INV_X1 U19747 ( .A(n16562), .ZN(U281) );
  OAI22_X1 U19748 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16563), .ZN(n16564) );
  INV_X1 U19749 ( .A(n16564), .ZN(U282) );
  INV_X1 U19750 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16565) );
  AOI222_X1 U19751 ( .A1(n19215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16566), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16565), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16567) );
  INV_X2 U19752 ( .A(n16569), .ZN(n16568) );
  INV_X1 U19753 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18795) );
  INV_X1 U19754 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U19755 ( .A1(n16568), .A2(n18795), .B1(n19888), .B2(n16569), .ZN(
        U347) );
  INV_X1 U19756 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18793) );
  INV_X1 U19757 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19886) );
  AOI22_X1 U19758 ( .A1(n16568), .A2(n18793), .B1(n19886), .B2(n16569), .ZN(
        U348) );
  INV_X1 U19759 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18791) );
  INV_X1 U19760 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U19761 ( .A1(n16568), .A2(n18791), .B1(n19885), .B2(n16569), .ZN(
        U349) );
  INV_X1 U19762 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18789) );
  INV_X1 U19763 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U19764 ( .A1(n16568), .A2(n18789), .B1(n19883), .B2(n16569), .ZN(
        U350) );
  INV_X1 U19765 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18787) );
  INV_X1 U19766 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19767 ( .A1(n16568), .A2(n18787), .B1(n19881), .B2(n16569), .ZN(
        U351) );
  INV_X1 U19768 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18785) );
  INV_X1 U19769 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19770 ( .A1(n16568), .A2(n18785), .B1(n19879), .B2(n16569), .ZN(
        U352) );
  INV_X1 U19771 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18783) );
  INV_X1 U19772 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U19773 ( .A1(n16568), .A2(n18783), .B1(n19878), .B2(n16569), .ZN(
        U353) );
  INV_X1 U19774 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18781) );
  AOI22_X1 U19775 ( .A1(n16568), .A2(n18781), .B1(n19876), .B2(n16569), .ZN(
        U354) );
  INV_X1 U19776 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18834) );
  INV_X1 U19777 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19926) );
  AOI22_X1 U19778 ( .A1(n16568), .A2(n18834), .B1(n19926), .B2(n16569), .ZN(
        U355) );
  INV_X1 U19779 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18832) );
  INV_X1 U19780 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19922) );
  AOI22_X1 U19781 ( .A1(n16568), .A2(n18832), .B1(n19922), .B2(n16569), .ZN(
        U356) );
  INV_X1 U19782 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18829) );
  INV_X1 U19783 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19920) );
  AOI22_X1 U19784 ( .A1(n16568), .A2(n18829), .B1(n19920), .B2(n16569), .ZN(
        U357) );
  INV_X1 U19785 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18828) );
  INV_X1 U19786 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19917) );
  AOI22_X1 U19787 ( .A1(n16568), .A2(n18828), .B1(n19917), .B2(n16569), .ZN(
        U358) );
  INV_X1 U19788 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18825) );
  INV_X1 U19789 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U19790 ( .A1(n16568), .A2(n18825), .B1(n19915), .B2(n16569), .ZN(
        U359) );
  INV_X1 U19791 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18823) );
  INV_X1 U19792 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U19793 ( .A1(n16568), .A2(n18823), .B1(n19914), .B2(n16569), .ZN(
        U360) );
  INV_X1 U19794 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18821) );
  INV_X1 U19795 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19912) );
  AOI22_X1 U19796 ( .A1(n16568), .A2(n18821), .B1(n19912), .B2(n16569), .ZN(
        U361) );
  INV_X1 U19797 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18819) );
  INV_X1 U19798 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19910) );
  AOI22_X1 U19799 ( .A1(n16568), .A2(n18819), .B1(n19910), .B2(n16569), .ZN(
        U362) );
  INV_X1 U19800 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18817) );
  INV_X1 U19801 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19908) );
  AOI22_X1 U19802 ( .A1(n16568), .A2(n18817), .B1(n19908), .B2(n16569), .ZN(
        U363) );
  INV_X1 U19803 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18815) );
  INV_X1 U19804 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U19805 ( .A1(n16568), .A2(n18815), .B1(n19907), .B2(n16569), .ZN(
        U364) );
  INV_X1 U19806 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18779) );
  INV_X1 U19807 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U19808 ( .A1(n16568), .A2(n18779), .B1(n19875), .B2(n16569), .ZN(
        U365) );
  INV_X1 U19809 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18813) );
  INV_X1 U19810 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19811 ( .A1(n16568), .A2(n18813), .B1(n19905), .B2(n16569), .ZN(
        U366) );
  INV_X1 U19812 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18812) );
  INV_X1 U19813 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U19814 ( .A1(n16568), .A2(n18812), .B1(n19904), .B2(n16569), .ZN(
        U367) );
  INV_X1 U19815 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18810) );
  INV_X1 U19816 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U19817 ( .A1(n16568), .A2(n18810), .B1(n19902), .B2(n16569), .ZN(
        U368) );
  INV_X1 U19818 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18807) );
  INV_X1 U19819 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U19820 ( .A1(n16568), .A2(n18807), .B1(n19901), .B2(n16569), .ZN(
        U369) );
  INV_X1 U19821 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18806) );
  INV_X1 U19822 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U19823 ( .A1(n16568), .A2(n18806), .B1(n19899), .B2(n16569), .ZN(
        U370) );
  INV_X1 U19824 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n21118) );
  INV_X1 U19825 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19826 ( .A1(n16568), .A2(n21118), .B1(n19897), .B2(n16569), .ZN(
        U371) );
  INV_X1 U19827 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18802) );
  INV_X1 U19828 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19895) );
  AOI22_X1 U19829 ( .A1(n16568), .A2(n18802), .B1(n19895), .B2(n16569), .ZN(
        U372) );
  INV_X1 U19830 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18801) );
  INV_X1 U19831 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U19832 ( .A1(n16568), .A2(n18801), .B1(n19893), .B2(n16569), .ZN(
        U373) );
  INV_X1 U19833 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18799) );
  INV_X1 U19834 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19835 ( .A1(n16568), .A2(n18799), .B1(n19891), .B2(n16569), .ZN(
        U374) );
  INV_X1 U19836 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18797) );
  INV_X1 U19837 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20959) );
  AOI22_X1 U19838 ( .A1(n16568), .A2(n18797), .B1(n20959), .B2(n16569), .ZN(
        U375) );
  INV_X1 U19839 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18777) );
  INV_X1 U19840 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19873) );
  AOI22_X1 U19841 ( .A1(n16568), .A2(n18777), .B1(n19873), .B2(n16569), .ZN(
        U376) );
  INV_X1 U19842 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16570) );
  NOR2_X1 U19843 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18768), .ZN(n18767) );
  NOR2_X1 U19844 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18764) );
  AOI21_X1 U19845 ( .B1(n18767), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18764), 
        .ZN(n18760) );
  INV_X1 U19846 ( .A(n18760), .ZN(n18847) );
  INV_X1 U19847 ( .A(n18847), .ZN(n18761) );
  OAI21_X1 U19848 ( .B1(n18768), .B2(n16570), .A(n18761), .ZN(P3_U2633) );
  NAND2_X1 U19849 ( .A1(n18910), .A2(n18850), .ZN(n16573) );
  AND2_X1 U19850 ( .A1(n17512), .A2(n16578), .ZN(n16571) );
  OAI21_X1 U19851 ( .B1(n16571), .B2(n17511), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16572) );
  OAI21_X1 U19852 ( .B1(n16573), .B2(n18754), .A(n16572), .ZN(P3_U2634) );
  INV_X1 U19853 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18776) );
  AOI21_X1 U19854 ( .B1(n18768), .B2(n18776), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16574) );
  AOI22_X1 U19855 ( .A1(n18843), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16574), 
        .B2(n18908), .ZN(P3_U2635) );
  NOR2_X1 U19856 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18762) );
  OAI21_X1 U19857 ( .B1(n18762), .B2(BS16), .A(n18847), .ZN(n18845) );
  OAI21_X1 U19858 ( .B1(n18847), .B2(n18893), .A(n18845), .ZN(P3_U2636) );
  INV_X1 U19859 ( .A(n16575), .ZN(n16577) );
  AOI211_X1 U19860 ( .C1(n17512), .C2(n16578), .A(n16577), .B(n16576), .ZN(
        n18737) );
  NOR2_X1 U19861 ( .A1(n18737), .A2(n18750), .ZN(n18889) );
  OAI21_X1 U19862 ( .B1(n18889), .B2(n18253), .A(n16579), .ZN(P3_U2637) );
  NOR4_X1 U19863 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16583) );
  NOR4_X1 U19864 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16582) );
  NOR4_X1 U19865 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16581) );
  NOR4_X1 U19866 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16580) );
  NAND4_X1 U19867 ( .A1(n16583), .A2(n16582), .A3(n16581), .A4(n16580), .ZN(
        n16589) );
  NOR4_X1 U19868 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16587) );
  AOI211_X1 U19869 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_12__SCAN_IN), .B(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16586) );
  NOR4_X1 U19870 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16585) );
  NOR4_X1 U19871 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16584) );
  NAND4_X1 U19872 ( .A1(n16587), .A2(n16586), .A3(n16585), .A4(n16584), .ZN(
        n16588) );
  NOR2_X1 U19873 ( .A1(n16589), .A2(n16588), .ZN(n18887) );
  INV_X1 U19874 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18841) );
  NOR3_X1 U19875 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16591) );
  OAI21_X1 U19876 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16591), .A(n18887), .ZN(
        n16590) );
  OAI21_X1 U19877 ( .B1(n18887), .B2(n18841), .A(n16590), .ZN(P3_U2638) );
  INV_X1 U19878 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18881) );
  INV_X1 U19879 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18846) );
  AOI21_X1 U19880 ( .B1(n18881), .B2(n18846), .A(n16591), .ZN(n16592) );
  INV_X1 U19881 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18838) );
  INV_X1 U19882 ( .A(n18887), .ZN(n18883) );
  AOI22_X1 U19883 ( .A1(n18887), .A2(n16592), .B1(n18838), .B2(n18883), .ZN(
        P3_U2639) );
  INV_X1 U19884 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18835) );
  NAND4_X1 U19885 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16637), .ZN(n16600) );
  NOR3_X1 U19886 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18835), .A3(n16600), 
        .ZN(n16594) );
  AOI21_X1 U19887 ( .B1(n16956), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16594), .ZN(
        n16605) );
  NAND2_X1 U19888 ( .A1(n16646), .A2(n16645), .ZN(n16644) );
  NOR2_X1 U19889 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16644), .ZN(n16628) );
  INV_X1 U19890 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16964) );
  NAND2_X1 U19891 ( .A1(n16628), .A2(n16964), .ZN(n16607) );
  NOR2_X1 U19892 ( .A1(n16954), .A2(n16607), .ZN(n16614) );
  INV_X1 U19893 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16969) );
  INV_X1 U19894 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16636) );
  NAND2_X1 U19895 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16598), .ZN(
        n16597) );
  AOI21_X1 U19896 ( .B1(n16636), .B2(n16597), .A(n16595), .ZN(n17563) );
  OAI21_X1 U19897 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16598), .A(
        n16597), .ZN(n17583) );
  INV_X1 U19898 ( .A(n17583), .ZN(n16640) );
  NOR2_X1 U19899 ( .A1(n16638), .A2(n16884), .ZN(n16630) );
  NAND2_X1 U19900 ( .A1(n13498), .A2(n16935), .ZN(n16945) );
  NOR3_X1 U19901 ( .A1(n16609), .A2(n16608), .A3(n16945), .ZN(n16603) );
  NAND3_X1 U19902 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16599) );
  AOI21_X1 U19903 ( .B1(n16599), .B2(n16957), .A(n16643), .ZN(n16621) );
  NOR2_X1 U19904 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16600), .ZN(n16612) );
  INV_X1 U19905 ( .A(n16612), .ZN(n16601) );
  AOI21_X1 U19906 ( .B1(n16621), .B2(n16601), .A(n18833), .ZN(n16602) );
  AOI211_X1 U19907 ( .C1(n16614), .C2(n16969), .A(n16603), .B(n16602), .ZN(
        n16604) );
  OAI211_X1 U19908 ( .C1(n16606), .C2(n16944), .A(n16605), .B(n16604), .ZN(
        P3_U2640) );
  NAND2_X1 U19909 ( .A1(n16955), .A2(n16607), .ZN(n16626) );
  XOR2_X1 U19910 ( .A(n16609), .B(n16608), .Z(n16613) );
  OAI22_X1 U19911 ( .A1(n16621), .A2(n18835), .B1(n16610), .B2(n16944), .ZN(
        n16611) );
  OAI21_X1 U19912 ( .B1(n16956), .B2(n16614), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16615) );
  NOR2_X1 U19913 ( .A1(n16628), .A2(n16964), .ZN(n16627) );
  AOI211_X1 U19914 ( .C1(n16619), .C2(n16618), .A(n16617), .B(n18757), .ZN(
        n16623) );
  INV_X1 U19915 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18831) );
  OAI22_X1 U19916 ( .A1(n16621), .A2(n18831), .B1(n16620), .B2(n16944), .ZN(
        n16622) );
  AOI211_X1 U19917 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16956), .A(n16623), .B(
        n16622), .ZN(n16625) );
  NAND4_X1 U19918 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16637), .A4(n18831), .ZN(n16624) );
  OAI211_X1 U19919 ( .C1(n16627), .C2(n16626), .A(n16625), .B(n16624), .ZN(
        P3_U2642) );
  AOI22_X1 U19920 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16643), .B1(n16956), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16635) );
  INV_X1 U19921 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18827) );
  INV_X1 U19922 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21059) );
  AOI22_X1 U19923 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .B1(n18827), .B2(n21059), .ZN(n16633) );
  AOI211_X1 U19924 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16644), .A(n16628), .B(
        n16954), .ZN(n16632) );
  AOI211_X1 U19925 ( .C1(n17563), .C2(n16630), .A(n16629), .B(n18757), .ZN(
        n16631) );
  AOI211_X1 U19926 ( .C1(n16637), .C2(n16633), .A(n16632), .B(n16631), .ZN(
        n16634) );
  OAI211_X1 U19927 ( .C1(n16636), .C2(n16944), .A(n16635), .B(n16634), .ZN(
        P3_U2643) );
  INV_X1 U19928 ( .A(n16637), .ZN(n16649) );
  AOI211_X1 U19929 ( .C1(n16640), .C2(n16639), .A(n16638), .B(n18757), .ZN(
        n16642) );
  INV_X1 U19930 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17586) );
  OAI22_X1 U19931 ( .A1(n17586), .A2(n16944), .B1(n16947), .B2(n16645), .ZN(
        n16641) );
  AOI211_X1 U19932 ( .C1(n16643), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16642), 
        .B(n16641), .ZN(n16648) );
  OAI211_X1 U19933 ( .C1(n16646), .C2(n16645), .A(n16955), .B(n16644), .ZN(
        n16647) );
  OAI211_X1 U19934 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16649), .A(n16648), 
        .B(n16647), .ZN(P3_U2644) );
  OR2_X1 U19935 ( .A1(n16954), .A2(n16650), .ZN(n16663) );
  AOI21_X1 U19936 ( .B1(n16955), .B2(n16650), .A(n16956), .ZN(n16660) );
  AOI211_X1 U19937 ( .C1(n17603), .C2(n16652), .A(n16651), .B(n18757), .ZN(
        n16657) );
  NAND3_X1 U19938 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16957), .A3(n16653), 
        .ZN(n16654) );
  OAI21_X1 U19939 ( .B1(n16944), .B2(n16655), .A(n16654), .ZN(n16656) );
  AOI211_X1 U19940 ( .C1(n16658), .C2(n18822), .A(n16657), .B(n16656), .ZN(
        n16659) );
  OAI221_X1 U19941 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16663), .C1(n21056), 
        .C2(n16660), .A(n16659), .ZN(P3_U2646) );
  AOI22_X1 U19942 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16923), .B1(
        n16956), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16669) );
  NOR2_X1 U19943 ( .A1(n16662), .A2(n16661), .ZN(n16677) );
  AOI21_X1 U19944 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16678), .A(n16663), .ZN(
        n16667) );
  AOI211_X1 U19945 ( .C1(n17617), .C2(n16665), .A(n16664), .B(n18757), .ZN(
        n16666) );
  AOI211_X1 U19946 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16677), .A(n16667), 
        .B(n16666), .ZN(n16668) );
  OAI211_X1 U19947 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16670), .A(n16669), 
        .B(n16668), .ZN(P3_U2647) );
  INV_X1 U19948 ( .A(n16671), .ZN(n16701) );
  NAND2_X1 U19949 ( .A1(n16925), .A2(n16701), .ZN(n16699) );
  OAI21_X1 U19950 ( .B1(n16682), .B2(n16699), .A(n18818), .ZN(n16676) );
  AOI211_X1 U19951 ( .C1(n17632), .C2(n16673), .A(n16672), .B(n18757), .ZN(
        n16675) );
  OAI22_X1 U19952 ( .A1(n9843), .A2(n16944), .B1(n16947), .B2(n16679), .ZN(
        n16674) );
  AOI211_X1 U19953 ( .C1(n16677), .C2(n16676), .A(n16675), .B(n16674), .ZN(
        n16681) );
  OAI211_X1 U19954 ( .C1(n16683), .C2(n16679), .A(n16955), .B(n16678), .ZN(
        n16680) );
  NAND2_X1 U19955 ( .A1(n16681), .A2(n16680), .ZN(P3_U2648) );
  OAI21_X1 U19956 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(P3_REIP_REG_22__SCAN_IN), 
        .A(n16682), .ZN(n16690) );
  AOI22_X1 U19957 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16923), .B1(
        n16956), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16689) );
  OAI21_X1 U19958 ( .B1(n16701), .B2(n16948), .A(n16958), .ZN(n16700) );
  AOI211_X1 U19959 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16695), .A(n16683), .B(
        n16954), .ZN(n16687) );
  AOI211_X1 U19960 ( .C1(n17653), .C2(n16685), .A(n16684), .B(n18757), .ZN(
        n16686) );
  AOI211_X1 U19961 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16700), .A(n16687), 
        .B(n16686), .ZN(n16688) );
  OAI211_X1 U19962 ( .C1(n16699), .C2(n16690), .A(n16689), .B(n16688), .ZN(
        P3_U2649) );
  AOI211_X1 U19963 ( .C1(n17671), .C2(n16692), .A(n16691), .B(n18757), .ZN(
        n16694) );
  OAI22_X1 U19964 ( .A1(n17668), .A2(n16944), .B1(n16947), .B2(n16696), .ZN(
        n16693) );
  AOI211_X1 U19965 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16700), .A(n16694), 
        .B(n16693), .ZN(n16698) );
  OAI211_X1 U19966 ( .C1(n16704), .C2(n16696), .A(n16955), .B(n16695), .ZN(
        n16697) );
  OAI211_X1 U19967 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16699), .A(n16698), 
        .B(n16697), .ZN(P3_U2650) );
  INV_X1 U19968 ( .A(n16700), .ZN(n16711) );
  INV_X1 U19969 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18814) );
  AOI22_X1 U19970 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16923), .B1(
        n16956), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16710) );
  NOR2_X1 U19971 ( .A1(n16701), .A2(n16948), .ZN(n16708) );
  AOI211_X1 U19972 ( .C1(n17681), .C2(n16703), .A(n16702), .B(n18757), .ZN(
        n16706) );
  AOI211_X1 U19973 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16720), .A(n16704), .B(
        n16954), .ZN(n16705) );
  AOI211_X1 U19974 ( .C1(n16708), .C2(n16707), .A(n16706), .B(n16705), .ZN(
        n16709) );
  OAI211_X1 U19975 ( .C1(n16711), .C2(n18814), .A(n16710), .B(n16709), .ZN(
        P3_U2651) );
  INV_X1 U19976 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18811) );
  INV_X1 U19977 ( .A(n16958), .ZN(n16943) );
  AOI21_X1 U19978 ( .B1(n16925), .B2(n16736), .A(n16943), .ZN(n16740) );
  INV_X1 U19979 ( .A(n16725), .ZN(n16712) );
  OAI21_X1 U19980 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16712), .A(
        n17645), .ZN(n17697) );
  INV_X1 U19981 ( .A(n16715), .ZN(n16714) );
  INV_X1 U19982 ( .A(n17697), .ZN(n16713) );
  OAI221_X1 U19983 ( .B1(n16715), .B2(n17697), .C1(n16714), .C2(n16713), .A(
        n16935), .ZN(n16717) );
  AOI22_X1 U19984 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16923), .B1(
        n16956), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16716) );
  OAI211_X1 U19985 ( .C1(n18811), .C2(n16740), .A(n16717), .B(n16716), .ZN(
        n16718) );
  INV_X1 U19986 ( .A(n16718), .ZN(n16724) );
  NOR2_X1 U19987 ( .A1(n16948), .A2(n16736), .ZN(n16729) );
  OAI211_X1 U19988 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16729), .B(n16719), .ZN(n16723) );
  OAI211_X1 U19989 ( .C1(n16728), .C2(n16721), .A(n16955), .B(n16720), .ZN(
        n16722) );
  NAND4_X1 U19990 ( .A1(n16724), .A2(n18229), .A3(n16723), .A4(n16722), .ZN(
        P3_U2652) );
  OAI21_X1 U19991 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17693), .A(
        n16725), .ZN(n17704) );
  INV_X1 U19992 ( .A(n17693), .ZN(n16726) );
  OAI21_X1 U19993 ( .B1(n16726), .B2(n16750), .A(n13498), .ZN(n16727) );
  XNOR2_X1 U19994 ( .A(n17704), .B(n16727), .ZN(n16734) );
  AOI211_X1 U19995 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16743), .A(n16728), .B(
        n16954), .ZN(n16732) );
  INV_X1 U19996 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18809) );
  AOI22_X1 U19997 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16923), .B1(
        n16729), .B2(n18809), .ZN(n16730) );
  OAI211_X1 U19998 ( .C1(n16740), .C2(n18809), .A(n16730), .B(n18229), .ZN(
        n16731) );
  AOI211_X1 U19999 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16956), .A(n16732), .B(
        n16731), .ZN(n16733) );
  OAI21_X1 U20000 ( .B1(n16734), .B2(n18757), .A(n16733), .ZN(P3_U2653) );
  AOI21_X1 U20001 ( .B1(n9840), .B2(n16746), .A(n17693), .ZN(n17720) );
  OAI21_X1 U20002 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16746), .A(
        n13498), .ZN(n16735) );
  XNOR2_X1 U20003 ( .A(n17720), .B(n16735), .ZN(n16742) );
  INV_X1 U20004 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18808) );
  AND2_X1 U20005 ( .A1(n16736), .A2(n16925), .ZN(n16737) );
  AOI22_X1 U20006 ( .A1(n16956), .A2(P3_EBX_REG_17__SCAN_IN), .B1(n16738), 
        .B2(n16737), .ZN(n16739) );
  OAI211_X1 U20007 ( .C1(n16740), .C2(n18808), .A(n16739), .B(n18229), .ZN(
        n16741) );
  AOI21_X1 U20008 ( .B1(n16935), .B2(n16742), .A(n16741), .ZN(n16745) );
  OAI211_X1 U20009 ( .C1(n16749), .C2(n17114), .A(n16955), .B(n16743), .ZN(
        n16744) );
  OAI211_X1 U20010 ( .C1(n16944), .C2(n9840), .A(n16745), .B(n16744), .ZN(
        P3_U2654) );
  INV_X1 U20011 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18805) );
  AOI21_X1 U20012 ( .B1(n16925), .B2(n16775), .A(n16943), .ZN(n16784) );
  OAI21_X1 U20013 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16747), .A(
        n16746), .ZN(n17734) );
  AOI211_X1 U20014 ( .C1(n13498), .C2(n16750), .A(n18757), .B(n17734), .ZN(
        n16748) );
  AOI211_X1 U20015 ( .C1(n16956), .C2(P3_EBX_REG_16__SCAN_IN), .A(n9633), .B(
        n16748), .ZN(n16758) );
  INV_X1 U20016 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18804) );
  NAND3_X1 U20017 ( .A1(n16925), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16776), 
        .ZN(n16769) );
  AOI21_X1 U20018 ( .B1(n18805), .B2(n18804), .A(n16769), .ZN(n16756) );
  AOI211_X1 U20019 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16763), .A(n16749), .B(
        n16954), .ZN(n16754) );
  INV_X1 U20020 ( .A(n17734), .ZN(n16752) );
  NAND3_X1 U20021 ( .A1(n16935), .A2(n13498), .A3(n16750), .ZN(n16760) );
  INV_X1 U20022 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16751) );
  OAI22_X1 U20023 ( .A1(n16752), .A2(n16760), .B1(n16751), .B2(n16944), .ZN(
        n16753) );
  AOI211_X1 U20024 ( .C1(n16756), .C2(n16755), .A(n16754), .B(n16753), .ZN(
        n16757) );
  OAI211_X1 U20025 ( .C1(n18805), .C2(n16784), .A(n16758), .B(n16757), .ZN(
        P3_U2655) );
  OAI21_X1 U20026 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17729), .A(
        n16759), .ZN(n17739) );
  INV_X1 U20027 ( .A(n17739), .ZN(n16762) );
  INV_X1 U20028 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17742) );
  AOI21_X1 U20029 ( .B1(n13498), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18757), .ZN(n16951) );
  OAI21_X1 U20030 ( .B1(n17742), .B2(n16884), .A(n16951), .ZN(n16761) );
  AOI22_X1 U20031 ( .A1(n16762), .A2(n16761), .B1(n16760), .B2(n17739), .ZN(
        n16767) );
  OAI211_X1 U20032 ( .C1(n16770), .C2(n16765), .A(n16955), .B(n16763), .ZN(
        n16764) );
  OAI211_X1 U20033 ( .C1(n16947), .C2(n16765), .A(n18229), .B(n16764), .ZN(
        n16766) );
  AOI211_X1 U20034 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16923), .A(
        n16767), .B(n16766), .ZN(n16768) );
  OAI221_X1 U20035 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16769), .C1(n18804), 
        .C2(n16784), .A(n16768), .ZN(P3_U2656) );
  INV_X1 U20036 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18803) );
  AOI211_X1 U20037 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16792), .A(n16770), .B(
        n16954), .ZN(n16771) );
  AOI21_X1 U20038 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16956), .A(n16771), .ZN(
        n16783) );
  INV_X1 U20039 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16777) );
  INV_X1 U20040 ( .A(n16772), .ZN(n17836) );
  NAND2_X1 U20041 ( .A1(n17836), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16859) );
  NOR2_X1 U20042 ( .A1(n16773), .A2(n16859), .ZN(n17768) );
  NAND2_X1 U20043 ( .A1(n17771), .A2(n17768), .ZN(n16787) );
  AOI21_X1 U20044 ( .B1(n16777), .B2(n16787), .A(n17729), .ZN(n17756) );
  NOR2_X1 U20045 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17923), .ZN(
        n16936) );
  NAND3_X1 U20046 ( .A1(n17800), .A2(n17771), .A3(n16936), .ZN(n16788) );
  NAND2_X1 U20047 ( .A1(n13498), .A2(n16788), .ZN(n16774) );
  XNOR2_X1 U20048 ( .A(n17756), .B(n16774), .ZN(n16781) );
  INV_X1 U20049 ( .A(n16775), .ZN(n16779) );
  NAND2_X1 U20050 ( .A1(n16925), .A2(n16776), .ZN(n16778) );
  OAI22_X1 U20051 ( .A1(n16779), .A2(n16778), .B1(n16777), .B2(n16944), .ZN(
        n16780) );
  AOI211_X1 U20052 ( .C1(n16935), .C2(n16781), .A(n9633), .B(n16780), .ZN(
        n16782) );
  OAI211_X1 U20053 ( .C1(n18803), .C2(n16784), .A(n16783), .B(n16782), .ZN(
        P3_U2657) );
  NOR3_X1 U20054 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16948), .A3(n16785), 
        .ZN(n16786) );
  AOI211_X1 U20055 ( .C1(n16956), .C2(P3_EBX_REG_13__SCAN_IN), .A(n9633), .B(
        n16786), .ZN(n16796) );
  OAI21_X1 U20056 ( .B1(n16800), .B2(n16948), .A(n16958), .ZN(n16817) );
  NOR2_X1 U20057 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16948), .ZN(n16799) );
  INV_X1 U20058 ( .A(n17768), .ZN(n16802) );
  NOR2_X1 U20059 ( .A1(n17773), .A2(n16802), .ZN(n16801) );
  OAI21_X1 U20060 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16801), .A(
        n16787), .ZN(n17783) );
  NAND2_X1 U20061 ( .A1(n17783), .A2(n16788), .ZN(n16789) );
  OAI22_X1 U20062 ( .A1(n17772), .A2(n16944), .B1(n16945), .B2(n16789), .ZN(
        n16790) );
  AOI221_X1 U20063 ( .B1(n16817), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16799), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16790), .ZN(n16795) );
  INV_X1 U20064 ( .A(n17783), .ZN(n16791) );
  OAI211_X1 U20065 ( .C1(n16801), .C2(n16884), .A(n16791), .B(n16951), .ZN(
        n16794) );
  OAI211_X1 U20066 ( .C1(n16797), .C2(n17150), .A(n16955), .B(n16792), .ZN(
        n16793) );
  NAND4_X1 U20067 ( .A1(n16796), .A2(n16795), .A3(n16794), .A4(n16793), .ZN(
        P3_U2658) );
  AOI211_X1 U20068 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16811), .A(n16797), .B(
        n16954), .ZN(n16798) );
  AOI21_X1 U20069 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16956), .A(n16798), .ZN(
        n16807) );
  AOI22_X1 U20070 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16923), .B1(
        n16800), .B2(n16799), .ZN(n16806) );
  AOI21_X1 U20071 ( .B1(n17773), .B2(n16802), .A(n16801), .ZN(n17788) );
  AOI21_X1 U20072 ( .B1(n17800), .B2(n16936), .A(n16884), .ZN(n16803) );
  XOR2_X1 U20073 ( .A(n17788), .B(n16803), .Z(n16804) );
  AOI22_X1 U20074 ( .A1(n16935), .A2(n16804), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16817), .ZN(n16805) );
  NAND4_X1 U20075 ( .A1(n16807), .A2(n16806), .A3(n16805), .A4(n18229), .ZN(
        P3_U2659) );
  OAI21_X1 U20076 ( .B1(n16948), .B2(n16808), .A(n18796), .ZN(n16816) );
  INV_X1 U20077 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16814) );
  NAND2_X1 U20078 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16826) );
  NOR2_X1 U20079 ( .A1(n16826), .A2(n16859), .ZN(n16833) );
  NAND2_X1 U20080 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16833), .ZN(
        n16825) );
  AOI21_X1 U20081 ( .B1(n16814), .B2(n16825), .A(n17768), .ZN(n17803) );
  OAI21_X1 U20082 ( .B1(n16825), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n13498), .ZN(n16809) );
  INV_X1 U20083 ( .A(n16809), .ZN(n16827) );
  INV_X1 U20084 ( .A(n17803), .ZN(n16810) );
  OAI221_X1 U20085 ( .B1(n17803), .B2(n16827), .C1(n16810), .C2(n16809), .A(
        n16935), .ZN(n16813) );
  OAI211_X1 U20086 ( .C1(n16820), .C2(n16819), .A(n16955), .B(n16811), .ZN(
        n16812) );
  OAI211_X1 U20087 ( .C1(n16944), .C2(n16814), .A(n16813), .B(n16812), .ZN(
        n16815) );
  AOI21_X1 U20088 ( .B1(n16817), .B2(n16816), .A(n16815), .ZN(n16818) );
  OAI211_X1 U20089 ( .C1(n16947), .C2(n16819), .A(n16818), .B(n18229), .ZN(
        P3_U2660) );
  AOI221_X1 U20090 ( .B1(n18792), .B2(n16925), .C1(n16832), .C2(n16925), .A(
        n16943), .ZN(n16831) );
  INV_X1 U20091 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18794) );
  AOI211_X1 U20092 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16843), .A(n16820), .B(
        n16954), .ZN(n16824) );
  INV_X1 U20093 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17222) );
  NAND3_X1 U20094 ( .A1(n16925), .A2(n16821), .A3(n18794), .ZN(n16822) );
  OAI211_X1 U20095 ( .C1(n16947), .C2(n17222), .A(n18229), .B(n16822), .ZN(
        n16823) );
  AOI211_X1 U20096 ( .C1(n16923), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16824), .B(n16823), .ZN(n16830) );
  OAI21_X1 U20097 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16833), .A(
        n16825), .ZN(n17819) );
  INV_X1 U20098 ( .A(n17819), .ZN(n16828) );
  OR2_X1 U20099 ( .A1(n16859), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16852) );
  OAI21_X1 U20100 ( .B1(n16826), .B2(n16852), .A(n13498), .ZN(n16838) );
  OAI221_X1 U20101 ( .B1(n16828), .B2(n16827), .C1(n17819), .C2(n16838), .A(
        n16935), .ZN(n16829) );
  OAI211_X1 U20102 ( .C1(n16831), .C2(n18794), .A(n16830), .B(n16829), .ZN(
        P3_U2661) );
  INV_X1 U20103 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17824) );
  INV_X1 U20104 ( .A(n16832), .ZN(n16839) );
  OAI21_X1 U20105 ( .B1(n16839), .B2(n16948), .A(n16958), .ZN(n16854) );
  NAND2_X1 U20106 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17835) );
  NAND2_X1 U20107 ( .A1(n9725), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16860) );
  NOR2_X1 U20108 ( .A1(n17835), .A2(n16860), .ZN(n16851) );
  INV_X1 U20109 ( .A(n16833), .ZN(n16834) );
  OAI21_X1 U20110 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16851), .A(
        n16834), .ZN(n17826) );
  INV_X1 U20111 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20983) );
  INV_X1 U20112 ( .A(n17826), .ZN(n16835) );
  OAI21_X1 U20113 ( .B1(n20983), .B2(n16852), .A(n16835), .ZN(n16836) );
  OAI21_X1 U20114 ( .B1(n16884), .B2(n16836), .A(n16935), .ZN(n16837) );
  AOI21_X1 U20115 ( .B1(n17826), .B2(n16838), .A(n16837), .ZN(n16842) );
  NAND3_X1 U20116 ( .A1(n16925), .A2(n16839), .A3(n18792), .ZN(n16840) );
  OAI211_X1 U20117 ( .C1(n16947), .C2(n16844), .A(n18229), .B(n16840), .ZN(
        n16841) );
  AOI211_X1 U20118 ( .C1(n16854), .C2(P3_REIP_REG_9__SCAN_IN), .A(n16842), .B(
        n16841), .ZN(n16846) );
  OAI211_X1 U20119 ( .C1(n16847), .C2(n16844), .A(n16955), .B(n16843), .ZN(
        n16845) );
  OAI211_X1 U20120 ( .C1(n16944), .C2(n17824), .A(n16846), .B(n16845), .ZN(
        P3_U2662) );
  AOI211_X1 U20121 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16862), .A(n16847), .B(
        n16954), .ZN(n16848) );
  AOI21_X1 U20122 ( .B1(n16923), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16848), .ZN(n16858) );
  NOR2_X1 U20123 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16948), .ZN(n16849) );
  AOI22_X1 U20124 ( .A1(n16956), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n16850), .B2(
        n16849), .ZN(n16857) );
  AOI21_X1 U20125 ( .B1(n20983), .B2(n16859), .A(n16851), .ZN(n17839) );
  NAND2_X1 U20126 ( .A1(n13498), .A2(n16852), .ZN(n16853) );
  XNOR2_X1 U20127 ( .A(n17839), .B(n16853), .ZN(n16855) );
  AOI22_X1 U20128 ( .A1(n16935), .A2(n16855), .B1(P3_REIP_REG_8__SCAN_IN), 
        .B2(n16854), .ZN(n16856) );
  NAND4_X1 U20129 ( .A1(n16858), .A2(n16857), .A3(n16856), .A4(n18229), .ZN(
        P3_U2663) );
  INV_X1 U20130 ( .A(n16860), .ZN(n16874) );
  OAI21_X1 U20131 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16874), .A(
        n16859), .ZN(n17856) );
  OAI21_X1 U20132 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16860), .A(
        n13498), .ZN(n16876) );
  XNOR2_X1 U20133 ( .A(n17856), .B(n16876), .ZN(n16870) );
  NOR3_X1 U20134 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16948), .A3(n16861), .ZN(
        n16866) );
  OAI211_X1 U20135 ( .C1(n16871), .C2(n16864), .A(n16955), .B(n16862), .ZN(
        n16863) );
  OAI211_X1 U20136 ( .C1(n16947), .C2(n16864), .A(n18229), .B(n16863), .ZN(
        n16865) );
  AOI211_X1 U20137 ( .C1(n16923), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16866), .B(n16865), .ZN(n16869) );
  INV_X1 U20138 ( .A(n16867), .ZN(n16888) );
  NOR3_X1 U20139 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16948), .A3(n16888), .ZN(
        n16873) );
  OAI21_X1 U20140 ( .B1(n16867), .B2(n16948), .A(n16958), .ZN(n16892) );
  OAI21_X1 U20141 ( .B1(n16873), .B2(n16892), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n16868) );
  OAI211_X1 U20142 ( .C1(n16870), .C2(n18757), .A(n16869), .B(n16868), .ZN(
        P3_U2664) );
  AOI211_X1 U20143 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16886), .A(n16871), .B(
        n16954), .ZN(n16872) );
  AOI211_X1 U20144 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16956), .A(n16873), .B(
        n16872), .ZN(n16882) );
  NOR2_X1 U20145 ( .A1(n17857), .A2(n17923), .ZN(n16883) );
  INV_X1 U20146 ( .A(n16883), .ZN(n16875) );
  AOI21_X1 U20147 ( .B1(n16877), .B2(n16875), .A(n16874), .ZN(n17863) );
  NOR3_X1 U20148 ( .A1(n17863), .A2(n18757), .A3(n16876), .ZN(n16879) );
  NOR2_X1 U20149 ( .A1(n16877), .A2(n16944), .ZN(n16878) );
  AOI211_X1 U20150 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n16892), .A(n16879), .B(
        n16878), .ZN(n16881) );
  OAI211_X1 U20151 ( .C1(n16883), .C2(n16884), .A(n17863), .B(n16951), .ZN(
        n16880) );
  NAND4_X1 U20152 ( .A1(n16882), .A2(n16881), .A3(n18229), .A4(n16880), .ZN(
        P3_U2665) );
  NAND2_X1 U20153 ( .A1(n9823), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16896) );
  AOI21_X1 U20154 ( .B1(n9826), .B2(n16896), .A(n16883), .ZN(n17875) );
  AOI21_X1 U20155 ( .B1(n9823), .B2(n16936), .A(n16884), .ZN(n16899) );
  XNOR2_X1 U20156 ( .A(n17875), .B(n16899), .ZN(n16895) );
  INV_X1 U20157 ( .A(n16900), .ZN(n16885) );
  AOI21_X1 U20158 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16885), .A(n16954), .ZN(
        n16887) );
  AOI22_X1 U20159 ( .A1(n16956), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n16887), .B2(
        n16886), .ZN(n16894) );
  NAND2_X1 U20160 ( .A1(n16925), .A2(n16888), .ZN(n16889) );
  OAI22_X1 U20161 ( .A1(n9826), .A2(n16944), .B1(n16890), .B2(n16889), .ZN(
        n16891) );
  AOI211_X1 U20162 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n16892), .A(n9633), .B(
        n16891), .ZN(n16893) );
  OAI211_X1 U20163 ( .C1(n18757), .C2(n16895), .A(n16894), .B(n16893), .ZN(
        P3_U2666) );
  NOR2_X1 U20164 ( .A1(n17885), .A2(n17923), .ZN(n16909) );
  OAI21_X1 U20165 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16909), .A(
        n16896), .ZN(n17888) );
  INV_X1 U20166 ( .A(n16936), .ZN(n16897) );
  OR2_X1 U20167 ( .A1(n17885), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17892) );
  OAI22_X1 U20168 ( .A1(n13498), .A2(n17888), .B1(n16897), .B2(n17892), .ZN(
        n16898) );
  AOI21_X1 U20169 ( .B1(n16899), .B2(n17888), .A(n16898), .ZN(n16908) );
  AOI22_X1 U20170 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16923), .B1(
        n16956), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16907) );
  OAI21_X1 U20171 ( .B1(n16901), .B2(n16948), .A(n16958), .ZN(n16917) );
  AOI211_X1 U20172 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16918), .A(n16900), .B(
        n16954), .ZN(n16905) );
  NAND2_X1 U20173 ( .A1(n16925), .A2(n16901), .ZN(n16903) );
  NOR2_X1 U20174 ( .A1(n18262), .A2(n18900), .ZN(n18915) );
  OAI21_X1 U20175 ( .B1(n17236), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18915), .ZN(n16902) );
  OAI211_X1 U20176 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16903), .A(n18229), .B(
        n16902), .ZN(n16904) );
  AOI211_X1 U20177 ( .C1(n16917), .C2(P3_REIP_REG_4__SCAN_IN), .A(n16905), .B(
        n16904), .ZN(n16906) );
  OAI211_X1 U20178 ( .C1(n16908), .C2(n18757), .A(n16907), .B(n16906), .ZN(
        P3_U2667) );
  INV_X1 U20179 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16922) );
  OAI21_X1 U20180 ( .B1(n16948), .B2(n16926), .A(n18780), .ZN(n16916) );
  NAND2_X1 U20181 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16924) );
  AOI21_X1 U20182 ( .B1(n16922), .B2(n16924), .A(n16909), .ZN(n17899) );
  OAI21_X1 U20183 ( .B1(n16924), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n13498), .ZN(n16910) );
  INV_X1 U20184 ( .A(n16910), .ZN(n16934) );
  OAI21_X1 U20185 ( .B1(n17899), .B2(n16934), .A(n16935), .ZN(n16911) );
  AOI21_X1 U20186 ( .B1(n17899), .B2(n16934), .A(n16911), .ZN(n16915) );
  INV_X1 U20187 ( .A(n18722), .ZN(n18704) );
  NOR2_X1 U20188 ( .A1(n18879), .A2(n18704), .ZN(n18703) );
  OAI21_X1 U20189 ( .B1(n18856), .B2(n18703), .A(n16912), .ZN(n18854) );
  AOI22_X1 U20190 ( .A1(n18854), .A2(n18915), .B1(n16956), .B2(
        P3_EBX_REG_3__SCAN_IN), .ZN(n16913) );
  INV_X1 U20191 ( .A(n16913), .ZN(n16914) );
  AOI211_X1 U20192 ( .C1(n16917), .C2(n16916), .A(n16915), .B(n16914), .ZN(
        n16921) );
  OAI211_X1 U20193 ( .C1(n16928), .C2(n16919), .A(n16955), .B(n16918), .ZN(
        n16920) );
  OAI211_X1 U20194 ( .C1(n16944), .C2(n16922), .A(n16921), .B(n16920), .ZN(
        P3_U2668) );
  AOI22_X1 U20195 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16923), .B1(
        n16956), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20196 ( .A1(n18722), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n18865), .B2(n18701), .ZN(n18862) );
  AOI22_X1 U20197 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16943), .B1(n18862), 
        .B2(n18915), .ZN(n16939) );
  NOR2_X1 U20198 ( .A1(n13498), .A2(n18757), .ZN(n16933) );
  OAI21_X1 U20199 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16924), .ZN(n17909) );
  INV_X1 U20200 ( .A(n17909), .ZN(n16932) );
  OAI211_X1 U20201 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16926), .B(n16925), .ZN(n16927) );
  INV_X1 U20202 ( .A(n16927), .ZN(n16931) );
  INV_X1 U20203 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n21061) );
  INV_X1 U20204 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17292) );
  NAND2_X1 U20205 ( .A1(n21061), .A2(n17292), .ZN(n16929) );
  AOI211_X1 U20206 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16929), .A(n16928), .B(
        n16954), .ZN(n16930) );
  AOI211_X1 U20207 ( .C1(n16933), .C2(n16932), .A(n16931), .B(n16930), .ZN(
        n16938) );
  OAI211_X1 U20208 ( .C1(n16936), .C2(n17909), .A(n16935), .B(n16934), .ZN(
        n16937) );
  NAND4_X1 U20209 ( .A1(n16940), .A2(n16939), .A3(n16938), .A4(n16937), .ZN(
        P3_U2669) );
  NOR2_X1 U20210 ( .A1(n21061), .A2(n17292), .ZN(n17286) );
  INV_X1 U20211 ( .A(n17286), .ZN(n16941) );
  OAI21_X1 U20212 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n16941), .ZN(n17293) );
  INV_X1 U20213 ( .A(n18701), .ZN(n18719) );
  NOR2_X1 U20214 ( .A1(n16942), .A2(n18719), .ZN(n18870) );
  AOI22_X1 U20215 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16943), .B1(n18870), 
        .B2(n18915), .ZN(n16953) );
  OAI21_X1 U20216 ( .B1(n16946), .B2(n16945), .A(n16944), .ZN(n16950) );
  OAI22_X1 U20217 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16948), .B1(n16947), 
        .B2(n17292), .ZN(n16949) );
  AOI221_X1 U20218 ( .B1(n16951), .B2(n17923), .C1(n16950), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16949), .ZN(n16952) );
  OAI211_X1 U20219 ( .C1(n16954), .C2(n17293), .A(n16953), .B(n16952), .ZN(
        P3_U2670) );
  NOR2_X1 U20220 ( .A1(n16956), .A2(n16955), .ZN(n16961) );
  AOI22_X1 U20221 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16957), .B1(n18915), 
        .B2(n18879), .ZN(n16960) );
  NAND3_X1 U20222 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18851), .A3(
        n16958), .ZN(n16959) );
  OAI211_X1 U20223 ( .C1(n16961), .C2(n21061), .A(n16960), .B(n16959), .ZN(
        P3_U2671) );
  INV_X1 U20224 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16962) );
  NOR2_X1 U20225 ( .A1(n16962), .A2(n17082), .ZN(n17043) );
  INV_X1 U20226 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21125) );
  NAND4_X1 U20227 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16963)
         );
  NOR4_X1 U20228 ( .A1(n16964), .A2(n21056), .A3(n21125), .A4(n16963), .ZN(
        n16965) );
  NAND4_X1 U20229 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17043), .A4(n16965), .ZN(n16968) );
  NOR2_X1 U20230 ( .A1(n16969), .A2(n16968), .ZN(n16995) );
  NAND2_X1 U20231 ( .A1(n17290), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16967) );
  NAND2_X1 U20232 ( .A1(n16995), .A2(n18296), .ZN(n16966) );
  OAI22_X1 U20233 ( .A1(n16995), .A2(n16967), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16966), .ZN(P3_U2672) );
  NAND2_X1 U20234 ( .A1(n16969), .A2(n16968), .ZN(n16970) );
  NAND2_X1 U20235 ( .A1(n16970), .A2(n17290), .ZN(n16994) );
  AOI22_X1 U20236 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16971) );
  OAI21_X1 U20237 ( .B1(n17058), .B2(n17274), .A(n16971), .ZN(n16981) );
  AOI22_X1 U20238 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16978) );
  INV_X1 U20239 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17159) );
  OAI22_X1 U20240 ( .A1(n17229), .A2(n21086), .B1(n17250), .B2(n17159), .ZN(
        n16976) );
  AOI22_X1 U20241 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20242 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20243 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16972) );
  NAND3_X1 U20244 ( .A1(n16974), .A2(n16973), .A3(n16972), .ZN(n16975) );
  AOI211_X1 U20245 ( .C1(n16984), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n16976), .B(n16975), .ZN(n16977) );
  OAI211_X1 U20246 ( .C1(n13194), .C2(n16979), .A(n16978), .B(n16977), .ZN(
        n16980) );
  AOI211_X1 U20247 ( .C1(n9632), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n16981), .B(n16980), .ZN(n16998) );
  NOR2_X1 U20248 ( .A1(n16998), .A2(n16997), .ZN(n16996) );
  AOI22_X1 U20249 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n13155), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16992) );
  INV_X1 U20250 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17138) );
  AOI22_X1 U20251 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20252 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17246), .ZN(n16982) );
  OAI211_X1 U20253 ( .C1(n17250), .C2(n17138), .A(n16983), .B(n16982), .ZN(
        n16990) );
  AOI22_X1 U20254 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20255 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17230), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17253), .ZN(n16987) );
  AOI22_X1 U20256 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n13171), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n16984), .ZN(n16986) );
  NAND2_X1 U20257 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17245), .ZN(
        n16985) );
  NAND4_X1 U20258 ( .A1(n16988), .A2(n16987), .A3(n16986), .A4(n16985), .ZN(
        n16989) );
  AOI211_X1 U20259 ( .C1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n17244), .A(
        n16990), .B(n16989), .ZN(n16991) );
  OAI211_X1 U20260 ( .C1(n17137), .C2(n17219), .A(n16992), .B(n16991), .ZN(
        n16993) );
  XNOR2_X1 U20261 ( .A(n16996), .B(n16993), .ZN(n17304) );
  OAI22_X1 U20262 ( .A1(n16995), .A2(n16994), .B1(n17304), .B2(n17290), .ZN(
        P3_U2673) );
  AOI21_X1 U20263 ( .B1(n16998), .B2(n16997), .A(n16996), .ZN(n17305) );
  INV_X1 U20264 ( .A(n17305), .ZN(n17000) );
  NAND3_X1 U20265 ( .A1(n17001), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17290), 
        .ZN(n16999) );
  OAI221_X1 U20266 ( .B1(n17001), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17290), 
        .C2(n17000), .A(n16999), .ZN(P3_U2674) );
  INV_X1 U20267 ( .A(n17002), .ZN(n17011) );
  AOI21_X1 U20268 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17290), .A(n17011), .ZN(
        n17006) );
  AOI21_X1 U20269 ( .B1(n17004), .B2(n17008), .A(n17003), .ZN(n17318) );
  INV_X1 U20270 ( .A(n17318), .ZN(n17005) );
  OAI22_X1 U20271 ( .A1(n17007), .A2(n17006), .B1(n17005), .B2(n17290), .ZN(
        P3_U2676) );
  AOI21_X1 U20272 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17290), .A(n17017), .ZN(
        n17010) );
  OAI21_X1 U20273 ( .B1(n17013), .B2(n17009), .A(n17008), .ZN(n17324) );
  OAI22_X1 U20274 ( .A1(n17011), .A2(n17010), .B1(n17324), .B2(n17290), .ZN(
        P3_U2677) );
  INV_X1 U20275 ( .A(n17012), .ZN(n17021) );
  AOI21_X1 U20276 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17290), .A(n17021), .ZN(
        n17016) );
  AOI21_X1 U20277 ( .B1(n17014), .B2(n17018), .A(n17013), .ZN(n17325) );
  INV_X1 U20278 ( .A(n17325), .ZN(n17015) );
  OAI22_X1 U20279 ( .A1(n17017), .A2(n17016), .B1(n17290), .B2(n17015), .ZN(
        P3_U2678) );
  AOI21_X1 U20280 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17290), .A(n17028), .ZN(
        n17020) );
  OAI21_X1 U20281 ( .B1(n17023), .B2(n17019), .A(n17018), .ZN(n17334) );
  OAI22_X1 U20282 ( .A1(n17021), .A2(n17020), .B1(n17290), .B2(n17334), .ZN(
        P3_U2679) );
  INV_X1 U20283 ( .A(n17022), .ZN(n17042) );
  AOI21_X1 U20284 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17290), .A(n17042), .ZN(
        n17027) );
  AOI21_X1 U20285 ( .B1(n17025), .B2(n17024), .A(n17023), .ZN(n17335) );
  INV_X1 U20286 ( .A(n17335), .ZN(n17026) );
  OAI22_X1 U20287 ( .A1(n17028), .A2(n17027), .B1(n17290), .B2(n17026), .ZN(
        P3_U2680) );
  AOI21_X1 U20288 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17290), .A(n17029), .ZN(
        n17041) );
  AOI22_X1 U20289 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20290 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20291 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17037) );
  OAI22_X1 U20292 ( .A1(n17264), .A2(n17274), .B1(n17199), .B2(n21086), .ZN(
        n17035) );
  AOI22_X1 U20293 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9632), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20294 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20295 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17031) );
  NAND2_X1 U20296 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n17030) );
  NAND4_X1 U20297 ( .A1(n17033), .A2(n17032), .A3(n17031), .A4(n17030), .ZN(
        n17034) );
  AOI211_X1 U20298 ( .C1(n17253), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17035), .B(n17034), .ZN(n17036) );
  NAND4_X1 U20299 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17341) );
  INV_X1 U20300 ( .A(n17341), .ZN(n17040) );
  OAI22_X1 U20301 ( .A1(n17042), .A2(n17041), .B1(n17040), .B2(n17290), .ZN(
        P3_U2681) );
  NOR2_X1 U20302 ( .A1(n17296), .A2(n17043), .ZN(n17069) );
  AOI22_X1 U20303 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20304 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20305 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17052) );
  OAI22_X1 U20306 ( .A1(n17264), .A2(n17277), .B1(n17250), .B2(n17044), .ZN(
        n17050) );
  AOI22_X1 U20307 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20308 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U20309 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17046) );
  NAND2_X1 U20310 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n17045) );
  NAND4_X1 U20311 ( .A1(n17048), .A2(n17047), .A3(n17046), .A4(n17045), .ZN(
        n17049) );
  AOI211_X1 U20312 ( .C1(n13171), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17050), .B(n17049), .ZN(n17051) );
  NAND4_X1 U20313 ( .A1(n17054), .A2(n17053), .A3(n17052), .A4(n17051), .ZN(
        n17347) );
  AOI22_X1 U20314 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17069), .B1(n17296), 
        .B2(n17347), .ZN(n17055) );
  OAI21_X1 U20315 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17056), .A(n17055), .ZN(
        P3_U2682) );
  AOI22_X1 U20316 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17057) );
  OAI21_X1 U20317 ( .B1(n17058), .B2(n17181), .A(n17057), .ZN(n17068) );
  AOI22_X1 U20318 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20319 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17059) );
  OAI21_X1 U20320 ( .B1(n17229), .B2(n17060), .A(n17059), .ZN(n17064) );
  AOI22_X1 U20321 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20322 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17061) );
  OAI211_X1 U20323 ( .C1(n17250), .C2(n17172), .A(n17062), .B(n17061), .ZN(
        n17063) );
  AOI211_X1 U20324 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17064), .B(n17063), .ZN(n17065) );
  OAI211_X1 U20325 ( .C1(n13126), .C2(n17174), .A(n17066), .B(n17065), .ZN(
        n17067) );
  AOI211_X1 U20326 ( .C1(n9639), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n17068), .B(n17067), .ZN(n17352) );
  OAI21_X1 U20327 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17070), .A(n17069), .ZN(
        n17071) );
  OAI21_X1 U20328 ( .B1(n17352), .B2(n17290), .A(n17071), .ZN(P3_U2683) );
  AOI22_X1 U20329 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20330 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20331 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17072) );
  OAI211_X1 U20332 ( .C1(n17229), .C2(n17198), .A(n17073), .B(n17072), .ZN(
        n17079) );
  AOI22_X1 U20333 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20334 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U20335 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17075) );
  NAND2_X1 U20336 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n17074) );
  NAND4_X1 U20337 ( .A1(n17077), .A2(n17076), .A3(n17075), .A4(n17074), .ZN(
        n17078) );
  AOI211_X1 U20338 ( .C1(n17244), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17079), .B(n17078), .ZN(n17080) );
  OAI211_X1 U20339 ( .C1(n17264), .C2(n17283), .A(n17081), .B(n17080), .ZN(
        n17356) );
  INV_X1 U20340 ( .A(n17356), .ZN(n17085) );
  OAI21_X1 U20341 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17083), .A(n17082), .ZN(
        n17084) );
  AOI22_X1 U20342 ( .A1(n17296), .A2(n17085), .B1(n17084), .B2(n17290), .ZN(
        P3_U2684) );
  NAND2_X1 U20343 ( .A1(n18296), .A2(n17298), .ZN(n17294) );
  OAI21_X1 U20344 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17087), .A(n17086), .ZN(
        n17099) );
  AOI22_X1 U20345 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20346 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U20347 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17088) );
  OAI211_X1 U20348 ( .C1(n13098), .C2(n17207), .A(n17089), .B(n17088), .ZN(
        n17095) );
  AOI22_X1 U20349 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20350 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20351 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17091) );
  NAND2_X1 U20352 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n17090) );
  NAND4_X1 U20353 ( .A1(n17093), .A2(n17092), .A3(n17091), .A4(n17090), .ZN(
        n17094) );
  AOI211_X1 U20354 ( .C1(n17236), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17095), .B(n17094), .ZN(n17096) );
  OAI211_X1 U20355 ( .C1(n17264), .C2(n17289), .A(n17097), .B(n17096), .ZN(
        n17363) );
  AOI22_X1 U20356 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17113), .B1(n17296), 
        .B2(n17363), .ZN(n17098) );
  OAI21_X1 U20357 ( .B1(n17294), .B2(n17099), .A(n17098), .ZN(P3_U2685) );
  AOI22_X1 U20358 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20359 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17100) );
  OAI21_X1 U20360 ( .B1(n17219), .B2(n17101), .A(n17100), .ZN(n17109) );
  OAI22_X1 U20361 ( .A1(n17226), .A2(n17102), .B1(n13194), .B2(n17225), .ZN(
        n17103) );
  AOI21_X1 U20362 ( .B1(n17255), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17103), .ZN(n17107) );
  AOI22_X1 U20363 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20364 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20365 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17104) );
  NAND4_X1 U20366 ( .A1(n17107), .A2(n17106), .A3(n17105), .A4(n17104), .ZN(
        n17108) );
  AOI211_X1 U20367 ( .C1(n9632), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17109), .B(n17108), .ZN(n17110) );
  OAI211_X1 U20368 ( .C1(n17264), .C2(n17291), .A(n17111), .B(n17110), .ZN(
        n17367) );
  INV_X1 U20369 ( .A(n17367), .ZN(n17118) );
  INV_X1 U20370 ( .A(n17112), .ZN(n17115) );
  NOR2_X1 U20371 ( .A1(n17115), .A2(n17340), .ZN(n17133) );
  OAI21_X1 U20372 ( .B1(n17133), .B2(n17113), .A(P3_EBX_REG_17__SCAN_IN), .ZN(
        n17117) );
  INV_X1 U20373 ( .A(n17294), .ZN(n17295) );
  NAND3_X1 U20374 ( .A1(n17115), .A2(n17295), .A3(n17114), .ZN(n17116) );
  OAI211_X1 U20375 ( .C1(n17118), .C2(n17290), .A(n17117), .B(n17116), .ZN(
        P3_U2686) );
  INV_X1 U20376 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17136) );
  OAI21_X1 U20377 ( .B1(n17132), .B2(n17203), .A(n17290), .ZN(n17153) );
  AOI22_X1 U20378 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20379 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17130) );
  OAI22_X1 U20380 ( .A1(n17264), .A2(n17119), .B1(n9629), .B2(n17249), .ZN(
        n17128) );
  AOI22_X1 U20381 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20382 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20383 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17120) );
  OAI211_X1 U20384 ( .C1(n17229), .C2(n17122), .A(n17121), .B(n17120), .ZN(
        n17123) );
  AOI21_X1 U20385 ( .B1(n17236), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17123), .ZN(n17124) );
  OAI211_X1 U20386 ( .C1(n17226), .C2(n17126), .A(n17125), .B(n17124), .ZN(
        n17127) );
  AOI211_X1 U20387 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17128), .B(n17127), .ZN(n17129) );
  NAND3_X1 U20388 ( .A1(n17131), .A2(n17130), .A3(n17129), .ZN(n17373) );
  NOR2_X1 U20389 ( .A1(n17132), .A2(n17203), .ZN(n17134) );
  AOI22_X1 U20390 ( .A1(n17296), .A2(n17373), .B1(n17134), .B2(n17133), .ZN(
        n17135) );
  OAI21_X1 U20391 ( .B1(n17136), .B2(n17153), .A(n17135), .ZN(P3_U2687) );
  OAI22_X1 U20392 ( .A1(n17264), .A2(n17137), .B1(n21077), .B2(n13156), .ZN(
        n17149) );
  AOI22_X1 U20393 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20394 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17254), .ZN(n17146) );
  OAI22_X1 U20395 ( .A1(n17139), .A2(n17250), .B1(n13098), .B2(n17138), .ZN(
        n17144) );
  AOI22_X1 U20396 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17253), .ZN(n17142) );
  AOI22_X1 U20397 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n13141), .B1(
        n9632), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20398 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17244), .ZN(n17140) );
  NAND3_X1 U20399 ( .A1(n17142), .A2(n17141), .A3(n17140), .ZN(n17143) );
  AOI211_X1 U20400 ( .C1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .C2(n13155), .A(
        n17144), .B(n17143), .ZN(n17145) );
  NAND3_X1 U20401 ( .A1(n17147), .A2(n17146), .A3(n17145), .ZN(n17148) );
  AOI211_X1 U20402 ( .C1(n17255), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17149), .B(n17148), .ZN(n17383) );
  INV_X1 U20403 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17167) );
  NOR2_X1 U20404 ( .A1(n17167), .A2(n17150), .ZN(n17152) );
  AOI21_X1 U20405 ( .B1(n17152), .B2(n17151), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n17154) );
  OAI22_X1 U20406 ( .A1(n17383), .A2(n17290), .B1(n17154), .B2(n17153), .ZN(
        P3_U2688) );
  OAI22_X1 U20407 ( .A1(n17264), .A2(n17155), .B1(n17219), .B2(n21086), .ZN(
        n17166) );
  AOI22_X1 U20408 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20409 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20410 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17156) );
  OAI21_X1 U20411 ( .B1(n9629), .B2(n17274), .A(n17156), .ZN(n17161) );
  AOI22_X1 U20412 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20413 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17157) );
  OAI211_X1 U20414 ( .C1(n13098), .C2(n17159), .A(n17158), .B(n17157), .ZN(
        n17160) );
  AOI211_X1 U20415 ( .C1(n17236), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17161), .B(n17160), .ZN(n17162) );
  NAND3_X1 U20416 ( .A1(n17164), .A2(n17163), .A3(n17162), .ZN(n17165) );
  AOI211_X1 U20417 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n17166), .B(n17165), .ZN(n17388) );
  OAI222_X1 U20418 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18296), .B1(
        P3_EBX_REG_14__SCAN_IN), .B2(n17169), .C1(n17168), .C2(n17167), .ZN(
        n17170) );
  OAI21_X1 U20419 ( .B1(n17388), .B2(n17290), .A(n17170), .ZN(P3_U2689) );
  AOI22_X1 U20420 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20421 ( .B1(n13131), .B2(n17172), .A(n17171), .ZN(n17183) );
  AOI22_X1 U20422 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20423 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U20424 ( .B1(n17229), .B2(n17174), .A(n17173), .ZN(n17178) );
  AOI22_X1 U20425 ( .A1(n17230), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20426 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17175) );
  OAI211_X1 U20427 ( .C1(n9629), .C2(n17280), .A(n17176), .B(n17175), .ZN(
        n17177) );
  AOI211_X1 U20428 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17178), .B(n17177), .ZN(n17179) );
  OAI211_X1 U20429 ( .C1(n17264), .C2(n17181), .A(n17180), .B(n17179), .ZN(
        n17182) );
  AOI211_X1 U20430 ( .C1(n13196), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17183), .B(n17182), .ZN(n17395) );
  NAND3_X1 U20431 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17290), .A3(n17203), 
        .ZN(n17187) );
  NAND4_X1 U20432 ( .A1(n18296), .A2(n17185), .A3(n17202), .A4(n17184), .ZN(
        n17186) );
  OAI211_X1 U20433 ( .C1(n17395), .C2(n17290), .A(n17187), .B(n17186), .ZN(
        P3_U2691) );
  INV_X1 U20434 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20435 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17188) );
  OAI21_X1 U20436 ( .B1(n13156), .B2(n17189), .A(n17188), .ZN(n17201) );
  AOI22_X1 U20437 ( .A1(n16984), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17197) );
  INV_X1 U20438 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U20439 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17190) );
  OAI21_X1 U20440 ( .B1(n17250), .B2(n17191), .A(n17190), .ZN(n17195) );
  AOI22_X1 U20441 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20442 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17192) );
  OAI211_X1 U20443 ( .C1(n9629), .C2(n17283), .A(n17193), .B(n17192), .ZN(
        n17194) );
  AOI211_X1 U20444 ( .C1(n17245), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17195), .B(n17194), .ZN(n17196) );
  OAI211_X1 U20445 ( .C1(n17199), .C2(n17198), .A(n17197), .B(n17196), .ZN(
        n17200) );
  AOI211_X1 U20446 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n17201), .B(n17200), .ZN(n17398) );
  AOI21_X1 U20447 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17202), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n17205) );
  NAND2_X1 U20448 ( .A1(n17290), .A2(n17203), .ZN(n17204) );
  OAI22_X1 U20449 ( .A1(n17398), .A2(n17290), .B1(n17205), .B2(n17204), .ZN(
        P3_U2692) );
  AOI22_X1 U20450 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17206) );
  OAI21_X1 U20451 ( .B1(n17208), .B2(n17207), .A(n17206), .ZN(n17221) );
  AOI22_X1 U20452 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17217) );
  INV_X1 U20453 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20454 ( .A1(n13171), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17236), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17209) );
  OAI21_X1 U20455 ( .B1(n17264), .B2(n17210), .A(n17209), .ZN(n17214) );
  AOI22_X1 U20456 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9632), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20457 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17254), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17211) );
  OAI211_X1 U20458 ( .C1(n9629), .C2(n17289), .A(n17212), .B(n17211), .ZN(
        n17213) );
  AOI211_X1 U20459 ( .C1(n17215), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17214), .B(n17213), .ZN(n17216) );
  OAI211_X1 U20460 ( .C1(n17219), .C2(n17218), .A(n17217), .B(n17216), .ZN(
        n17220) );
  AOI211_X1 U20461 ( .C1(n9639), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n17221), .B(n17220), .ZN(n17401) );
  AOI22_X1 U20462 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17242), .B1(n17202), 
        .B2(n17222), .ZN(n17223) );
  AOI22_X1 U20463 ( .A1(n17296), .A2(n17401), .B1(n17223), .B2(n17290), .ZN(
        P3_U2693) );
  AOI22_X1 U20464 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17224) );
  OAI21_X1 U20465 ( .B1(n17226), .B2(n17225), .A(n17224), .ZN(n17241) );
  AOI22_X1 U20466 ( .A1(n17246), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17238) );
  INV_X1 U20467 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20468 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13155), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17227) );
  OAI21_X1 U20469 ( .B1(n17229), .B2(n17228), .A(n17227), .ZN(n17235) );
  AOI22_X1 U20470 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17230), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U20471 ( .A1(n17255), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17231) );
  OAI211_X1 U20472 ( .C1(n9629), .C2(n17291), .A(n17232), .B(n17231), .ZN(
        n17234) );
  AOI211_X1 U20473 ( .C1(n17236), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n17235), .B(n17234), .ZN(n17237) );
  OAI211_X1 U20474 ( .C1(n17264), .C2(n17239), .A(n17238), .B(n17237), .ZN(
        n17240) );
  AOI211_X1 U20475 ( .C1(n9632), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n17241), .B(n17240), .ZN(n17408) );
  AND2_X1 U20476 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17272), .ZN(n17266) );
  OAI21_X1 U20477 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17266), .A(n17242), .ZN(
        n17243) );
  AOI22_X1 U20478 ( .A1(n17296), .A2(n17408), .B1(n17243), .B2(n17290), .ZN(
        P3_U2694) );
  AOI22_X1 U20479 ( .A1(n17245), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17244), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U20480 ( .A1(n13196), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17246), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20481 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13141), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17247) );
  OAI211_X1 U20482 ( .C1(n17250), .C2(n17249), .A(n17248), .B(n17247), .ZN(
        n17261) );
  AOI22_X1 U20483 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17251), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20484 ( .A1(n17254), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17253), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20485 ( .A1(n9632), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17255), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17257) );
  NAND2_X1 U20486 ( .A1(n13155), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n17256) );
  NAND4_X1 U20487 ( .A1(n17259), .A2(n17258), .A3(n17257), .A4(n17256), .ZN(
        n17260) );
  AOI211_X1 U20488 ( .C1(n13171), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17261), .B(n17260), .ZN(n17262) );
  OAI211_X1 U20489 ( .C1(n17264), .C2(n21110), .A(n17263), .B(n17262), .ZN(
        n17410) );
  INV_X1 U20490 ( .A(n17410), .ZN(n17267) );
  OAI21_X1 U20491 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17272), .A(n17290), .ZN(
        n17265) );
  OAI22_X1 U20492 ( .A1(n17267), .A2(n17290), .B1(n17266), .B2(n17265), .ZN(
        P3_U2695) );
  NOR2_X1 U20493 ( .A1(n17268), .A2(n17294), .ZN(n17287) );
  NAND2_X1 U20494 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17282), .ZN(n17273) );
  NOR2_X1 U20495 ( .A1(n17269), .A2(n17273), .ZN(n17276) );
  AOI21_X1 U20496 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17290), .A(n17276), .ZN(
        n17271) );
  OAI22_X1 U20497 ( .A1(n17272), .A2(n17271), .B1(n17270), .B2(n17290), .ZN(
        P3_U2696) );
  INV_X1 U20498 ( .A(n17273), .ZN(n17279) );
  AOI21_X1 U20499 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17290), .A(n17279), .ZN(
        n17275) );
  OAI22_X1 U20500 ( .A1(n17276), .A2(n17275), .B1(n17274), .B2(n17290), .ZN(
        P3_U2697) );
  AOI21_X1 U20501 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17290), .A(n17282), .ZN(
        n17278) );
  OAI22_X1 U20502 ( .A1(n17279), .A2(n17278), .B1(n17277), .B2(n17290), .ZN(
        P3_U2698) );
  AOI21_X1 U20503 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17290), .A(n17285), .ZN(
        n17281) );
  OAI22_X1 U20504 ( .A1(n17282), .A2(n17281), .B1(n17280), .B2(n17290), .ZN(
        P3_U2699) );
  AOI21_X1 U20505 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17290), .A(n17287), .ZN(
        n17284) );
  OAI22_X1 U20506 ( .A1(n17285), .A2(n17284), .B1(n17283), .B2(n17290), .ZN(
        P3_U2700) );
  AOI221_X1 U20507 ( .B1(n17286), .B2(n17298), .C1(n17340), .C2(n17298), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17288) );
  AOI211_X1 U20508 ( .C1(n17296), .C2(n17289), .A(n17288), .B(n17287), .ZN(
        P3_U2701) );
  OAI222_X1 U20509 ( .A1(n17294), .A2(n17293), .B1(n17292), .B2(n17298), .C1(
        n17291), .C2(n17290), .ZN(P3_U2702) );
  AOI22_X1 U20510 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17296), .B1(
        n17295), .B2(n21061), .ZN(n17297) );
  OAI21_X1 U20511 ( .B1(n17298), .B2(n21061), .A(n17297), .ZN(P3_U2703) );
  INV_X1 U20512 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17454) );
  INV_X1 U20513 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17458) );
  INV_X1 U20514 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17462) );
  INV_X1 U20515 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17468) );
  INV_X1 U20516 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17477) );
  INV_X1 U20517 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17560) );
  INV_X1 U20518 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17544) );
  NAND2_X1 U20519 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17443) );
  NAND2_X1 U20520 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17415) );
  NAND4_X1 U20521 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17299) );
  NOR3_X1 U20522 ( .A1(n17443), .A2(n17415), .A3(n17299), .ZN(n17409) );
  NAND2_X1 U20523 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17409), .ZN(n17405) );
  NOR2_X1 U20524 ( .A1(n17544), .A2(n17405), .ZN(n17389) );
  INV_X1 U20525 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17486) );
  INV_X1 U20526 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17488) );
  INV_X1 U20527 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17490) );
  NOR3_X1 U20528 ( .A1(n17486), .A2(n17488), .A3(n17490), .ZN(n17390) );
  NAND3_X1 U20529 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17389), .A3(n17390), 
        .ZN(n17384) );
  NAND4_X1 U20530 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n17346)
         );
  NAND2_X1 U20531 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17337), .ZN(n17336) );
  NAND2_X1 U20532 ( .A1(n17306), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20533 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17374), .ZN(n17303) );
  OAI211_X1 U20534 ( .C1(n17306), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17437), .B(
        n17301), .ZN(n17302) );
  OAI211_X1 U20535 ( .C1(n17304), .C2(n17447), .A(n17303), .B(n17302), .ZN(
        P3_U2705) );
  INV_X1 U20536 ( .A(n17374), .ZN(n17362) );
  AOI22_X1 U20537 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17357), .B1(n17423), .B2(
        n17305), .ZN(n17309) );
  AOI211_X1 U20538 ( .C1(n17454), .C2(n17311), .A(n17306), .B(n17425), .ZN(
        n17307) );
  INV_X1 U20539 ( .A(n17307), .ZN(n17308) );
  OAI211_X1 U20540 ( .C1(n17362), .C2(n17310), .A(n17309), .B(n17308), .ZN(
        P3_U2706) );
  AOI22_X1 U20541 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17374), .ZN(n17313) );
  OAI211_X1 U20542 ( .C1(n17315), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17437), .B(
        n17311), .ZN(n17312) );
  OAI211_X1 U20543 ( .C1(n17314), .C2(n17447), .A(n17313), .B(n17312), .ZN(
        P3_U2707) );
  INV_X1 U20544 ( .A(n17315), .ZN(n17317) );
  OAI21_X1 U20545 ( .B1(n17425), .B2(n17458), .A(n17321), .ZN(n17316) );
  AOI22_X1 U20546 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17374), .B1(n17317), .B2(
        n17316), .ZN(n17320) );
  AOI22_X1 U20547 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17357), .B1(n17423), .B2(
        n17318), .ZN(n17319) );
  NAND2_X1 U20548 ( .A1(n17320), .A2(n17319), .ZN(P3_U2708) );
  AOI22_X1 U20549 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17374), .ZN(n17323) );
  OAI211_X1 U20550 ( .C1(n17326), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17437), .B(
        n17321), .ZN(n17322) );
  OAI211_X1 U20551 ( .C1(n17324), .C2(n17447), .A(n17323), .B(n17322), .ZN(
        P3_U2709) );
  AOI22_X1 U20552 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17357), .B1(n17423), .B2(
        n17325), .ZN(n17329) );
  AOI211_X1 U20553 ( .C1(n17462), .C2(n17330), .A(n17326), .B(n17425), .ZN(
        n17327) );
  INV_X1 U20554 ( .A(n17327), .ZN(n17328) );
  OAI211_X1 U20555 ( .C1(n17362), .C2(n15079), .A(n17329), .B(n17328), .ZN(
        P3_U2710) );
  AOI22_X1 U20556 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17374), .ZN(n17333) );
  OAI211_X1 U20557 ( .C1(n17331), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17437), .B(
        n17330), .ZN(n17332) );
  OAI211_X1 U20558 ( .C1(n17334), .C2(n17447), .A(n17333), .B(n17332), .ZN(
        P3_U2711) );
  AOI22_X1 U20559 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17357), .B1(n17423), .B2(
        n17335), .ZN(n17339) );
  OAI211_X1 U20560 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17337), .A(n17437), .B(
        n17336), .ZN(n17338) );
  OAI211_X1 U20561 ( .C1(n17362), .C2(n18292), .A(n17339), .B(n17338), .ZN(
        P3_U2712) );
  NAND2_X1 U20562 ( .A1(n17368), .A2(n17468), .ZN(n17345) );
  AOI22_X1 U20563 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17374), .B1(n17423), .B2(
        n17341), .ZN(n17344) );
  INV_X1 U20564 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17473) );
  NAND2_X1 U20565 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17368), .ZN(n17364) );
  NAND2_X1 U20566 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17358), .ZN(n17351) );
  NAND2_X1 U20567 ( .A1(n17437), .A2(n17351), .ZN(n17348) );
  OAI21_X1 U20568 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17414), .A(n17348), .ZN(
        n17342) );
  AOI22_X1 U20569 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17357), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17342), .ZN(n17343) );
  OAI211_X1 U20570 ( .C1(n17346), .C2(n17345), .A(n17344), .B(n17343), .ZN(
        P3_U2713) );
  AOI22_X1 U20571 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17374), .B1(n17423), .B2(
        n17347), .ZN(n17350) );
  INV_X1 U20572 ( .A(n17348), .ZN(n17354) );
  AOI22_X1 U20573 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17357), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17354), .ZN(n17349) );
  OAI211_X1 U20574 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17351), .A(n17350), .B(
        n17349), .ZN(P3_U2714) );
  INV_X1 U20575 ( .A(n17357), .ZN(n17378) );
  INV_X1 U20576 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17471) );
  OAI22_X1 U20577 ( .A1(n17352), .A2(n17447), .B1(n19367), .B2(n17362), .ZN(
        n17353) );
  AOI221_X1 U20578 ( .B1(n17354), .B2(P3_EAX_REG_20__SCAN_IN), .C1(n17358), 
        .C2(n17471), .A(n17353), .ZN(n17355) );
  OAI21_X1 U20579 ( .B1(n18280), .B2(n17378), .A(n17355), .ZN(P3_U2715) );
  AOI22_X1 U20580 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17357), .B1(n17423), .B2(
        n17356), .ZN(n17361) );
  AOI211_X1 U20581 ( .C1(n17473), .C2(n17364), .A(n17358), .B(n17425), .ZN(
        n17359) );
  INV_X1 U20582 ( .A(n17359), .ZN(n17360) );
  OAI211_X1 U20583 ( .C1(n17362), .C2(n15109), .A(n17361), .B(n17360), .ZN(
        P3_U2716) );
  AOI22_X1 U20584 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17374), .B1(n17423), .B2(
        n17363), .ZN(n17366) );
  OAI211_X1 U20585 ( .C1(n17368), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17437), .B(
        n17364), .ZN(n17365) );
  OAI211_X1 U20586 ( .C1(n17378), .C2(n18271), .A(n17366), .B(n17365), .ZN(
        P3_U2717) );
  AOI22_X1 U20587 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n17374), .B1(n17423), .B2(
        n17367), .ZN(n17372) );
  INV_X1 U20588 ( .A(n17375), .ZN(n17370) );
  INV_X1 U20589 ( .A(n17368), .ZN(n17369) );
  OAI211_X1 U20590 ( .C1(n17370), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17437), .B(
        n17369), .ZN(n17371) );
  OAI211_X1 U20591 ( .C1(n17378), .C2(n21108), .A(n17372), .B(n17371), .ZN(
        P3_U2718) );
  AOI22_X1 U20592 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17374), .B1(n17423), .B2(
        n17373), .ZN(n17377) );
  OAI211_X1 U20593 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17379), .A(n17437), .B(
        n17375), .ZN(n17376) );
  OAI211_X1 U20594 ( .C1(n17378), .C2(n18263), .A(n17377), .B(n17376), .ZN(
        P3_U2719) );
  AOI211_X1 U20595 ( .C1(n17560), .C2(n17380), .A(n17425), .B(n17379), .ZN(
        n17381) );
  AOI21_X1 U20596 ( .B1(n17442), .B2(BUF2_REG_15__SCAN_IN), .A(n17381), .ZN(
        n17382) );
  OAI21_X1 U20597 ( .B1(n17383), .B2(n17447), .A(n17382), .ZN(P3_U2720) );
  NOR2_X1 U20598 ( .A1(n17384), .A2(n17414), .ZN(n17393) );
  INV_X1 U20599 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U20600 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17442), .B1(n17393), .B2(
        n17556), .ZN(n17387) );
  OR3_X1 U20601 ( .A1(n17556), .A2(n17425), .A3(n17385), .ZN(n17386) );
  OAI211_X1 U20602 ( .C1(n17388), .C2(n17447), .A(n17387), .B(n17386), .ZN(
        P3_U2721) );
  INV_X1 U20603 ( .A(n17414), .ZN(n17444) );
  NAND2_X1 U20604 ( .A1(n17389), .A2(n17444), .ZN(n17394) );
  INV_X1 U20605 ( .A(n17394), .ZN(n17404) );
  AND2_X1 U20606 ( .A1(n17390), .A2(n17404), .ZN(n17397) );
  AOI21_X1 U20607 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17437), .A(n17397), .ZN(
        n17392) );
  OAI222_X1 U20608 ( .A1(n17440), .A2(n17554), .B1(n17393), .B2(n17392), .C1(
        n17447), .C2(n17391), .ZN(P3_U2722) );
  NOR2_X1 U20609 ( .A1(n17490), .A2(n17394), .ZN(n17403) );
  AND2_X1 U20610 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17403), .ZN(n17400) );
  AOI21_X1 U20611 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17437), .A(n17400), .ZN(
        n17396) );
  OAI222_X1 U20612 ( .A1(n17440), .A2(n17550), .B1(n17397), .B2(n17396), .C1(
        n17447), .C2(n17395), .ZN(P3_U2723) );
  AOI21_X1 U20613 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17437), .A(n17403), .ZN(
        n17399) );
  OAI222_X1 U20614 ( .A1(n17440), .A2(n17548), .B1(n17400), .B2(n17399), .C1(
        n17447), .C2(n17398), .ZN(P3_U2724) );
  AOI21_X1 U20615 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17437), .A(n17404), .ZN(
        n17402) );
  OAI222_X1 U20616 ( .A1(n17440), .A2(n17546), .B1(n17403), .B2(n17402), .C1(
        n17447), .C2(n17401), .ZN(P3_U2725) );
  AOI221_X1 U20617 ( .B1(n17441), .B2(n17544), .C1(n17405), .C2(n17544), .A(
        n17404), .ZN(n17406) );
  AOI22_X1 U20618 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17442), .B1(n17406), .B2(
        n17437), .ZN(n17407) );
  OAI21_X1 U20619 ( .B1(n17408), .B2(n17447), .A(n17407), .ZN(P3_U2726) );
  NAND2_X1 U20620 ( .A1(n17409), .A2(n17444), .ZN(n17413) );
  NAND2_X1 U20621 ( .A1(n17413), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20622 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17442), .B1(n17423), .B2(
        n17410), .ZN(n17411) );
  OAI221_X1 U20623 ( .B1(n17413), .B2(P3_EAX_REG_8__SCAN_IN), .C1(n17412), 
        .C2(n17425), .A(n17411), .ZN(P3_U2727) );
  INV_X1 U20624 ( .A(n17413), .ZN(n17418) );
  INV_X1 U20625 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17502) );
  NOR2_X1 U20626 ( .A1(n17443), .A2(n17414), .ZN(n17436) );
  NAND2_X1 U20627 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17436), .ZN(n17431) );
  NAND2_X1 U20628 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17435), .ZN(n17427) );
  NOR2_X1 U20629 ( .A1(n17415), .A2(n17427), .ZN(n17421) );
  AOI21_X1 U20630 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17437), .A(n17421), .ZN(
        n17417) );
  OAI222_X1 U20631 ( .A1(n17440), .A2(n18293), .B1(n17418), .B2(n17417), .C1(
        n17447), .C2(n17416), .ZN(P3_U2728) );
  INV_X1 U20632 ( .A(n17427), .ZN(n17430) );
  AOI22_X1 U20633 ( .A1(n17430), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17437), .ZN(n17420) );
  OAI222_X1 U20634 ( .A1(n17440), .A2(n18288), .B1(n17421), .B2(n17420), .C1(
        n17447), .C2(n17419), .ZN(P3_U2729) );
  NAND2_X1 U20635 ( .A1(n17427), .A2(P3_EAX_REG_5__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20636 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17442), .B1(n17423), .B2(
        n17422), .ZN(n17424) );
  OAI221_X1 U20637 ( .B1(n17427), .B2(P3_EAX_REG_5__SCAN_IN), .C1(n17426), 
        .C2(n17425), .A(n17424), .ZN(P3_U2730) );
  AOI21_X1 U20638 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17437), .A(n17435), .ZN(
        n17429) );
  OAI222_X1 U20639 ( .A1(n17440), .A2(n18280), .B1(n17430), .B2(n17429), .C1(
        n17447), .C2(n17428), .ZN(P3_U2731) );
  INV_X1 U20640 ( .A(n17431), .ZN(n17439) );
  AOI21_X1 U20641 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17437), .A(n17439), .ZN(
        n17434) );
  INV_X1 U20642 ( .A(n17432), .ZN(n17433) );
  OAI222_X1 U20643 ( .A1(n18276), .A2(n17440), .B1(n17435), .B2(n17434), .C1(
        n17447), .C2(n17433), .ZN(P3_U2732) );
  AOI21_X1 U20644 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17437), .A(n17436), .ZN(
        n17438) );
  OAI222_X1 U20645 ( .A1(n18271), .A2(n17440), .B1(n17439), .B2(n17438), .C1(
        n17447), .C2(n10083), .ZN(P3_U2733) );
  AOI22_X1 U20646 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17442), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17441), .ZN(n17446) );
  OAI211_X1 U20647 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17444), .B(n17443), .ZN(n17445) );
  OAI211_X1 U20648 ( .C1(n17448), .C2(n17447), .A(n17446), .B(n17445), .ZN(
        P3_U2734) );
  NOR2_X2 U20649 ( .A1(n18859), .A2(n17928), .ZN(n18905) );
  NOR2_X4 U20650 ( .A1(n18905), .A2(n17451), .ZN(n17492) );
  AND2_X1 U20651 ( .A1(n17492), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20652 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17530) );
  AOI22_X1 U20653 ( .A1(n18905), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20654 ( .B1(n17530), .B2(n17479), .A(n17452), .ZN(P3_U2737) );
  AOI22_X1 U20655 ( .A1(n18905), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17453) );
  OAI21_X1 U20656 ( .B1(n17454), .B2(n17479), .A(n17453), .ZN(P3_U2738) );
  INV_X1 U20657 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20658 ( .A1(n18905), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17455) );
  OAI21_X1 U20659 ( .B1(n17456), .B2(n17479), .A(n17455), .ZN(P3_U2739) );
  AOI22_X1 U20660 ( .A1(n18905), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U20661 ( .B1(n17458), .B2(n17479), .A(n17457), .ZN(P3_U2740) );
  INV_X1 U20662 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20663 ( .A1(n18905), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20664 ( .B1(n17460), .B2(n17479), .A(n17459), .ZN(P3_U2741) );
  AOI22_X1 U20665 ( .A1(P3_UWORD_REG_9__SCAN_IN), .A2(n18905), .B1(n17492), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17461) );
  OAI21_X1 U20666 ( .B1(n17462), .B2(n17479), .A(n17461), .ZN(P3_U2742) );
  INV_X1 U20667 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U20668 ( .A1(n18905), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U20669 ( .B1(n17464), .B2(n17479), .A(n17463), .ZN(P3_U2743) );
  INV_X1 U20670 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U20671 ( .A1(n18905), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20672 ( .B1(n17466), .B2(n17479), .A(n17465), .ZN(P3_U2744) );
  AOI22_X1 U20673 ( .A1(n17507), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20674 ( .B1(n17468), .B2(n17479), .A(n17467), .ZN(P3_U2745) );
  INV_X1 U20675 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U20676 ( .A1(n17507), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20677 ( .B1(n17519), .B2(n17479), .A(n17469), .ZN(P3_U2746) );
  AOI22_X1 U20678 ( .A1(n17507), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17470) );
  OAI21_X1 U20679 ( .B1(n17471), .B2(n17479), .A(n17470), .ZN(P3_U2747) );
  AOI22_X1 U20680 ( .A1(n17507), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17472) );
  OAI21_X1 U20681 ( .B1(n17473), .B2(n17479), .A(n17472), .ZN(P3_U2748) );
  INV_X1 U20682 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17475) );
  AOI22_X1 U20683 ( .A1(n17507), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17474) );
  OAI21_X1 U20684 ( .B1(n17475), .B2(n17479), .A(n17474), .ZN(P3_U2749) );
  AOI22_X1 U20685 ( .A1(n17507), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17476) );
  OAI21_X1 U20686 ( .B1(n17477), .B2(n17479), .A(n17476), .ZN(P3_U2750) );
  INV_X1 U20687 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17480) );
  AOI22_X1 U20688 ( .A1(n17507), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17478) );
  OAI21_X1 U20689 ( .B1(n17480), .B2(n17479), .A(n17478), .ZN(P3_U2751) );
  AOI22_X1 U20690 ( .A1(n17507), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17481) );
  OAI21_X1 U20691 ( .B1(n17560), .B2(n17509), .A(n17481), .ZN(P3_U2752) );
  AOI22_X1 U20692 ( .A1(n17507), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17482) );
  OAI21_X1 U20693 ( .B1(n17556), .B2(n17509), .A(n17482), .ZN(P3_U2753) );
  INV_X1 U20694 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20695 ( .A1(n17507), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20696 ( .B1(n17484), .B2(n17509), .A(n17483), .ZN(P3_U2754) );
  AOI22_X1 U20697 ( .A1(n17507), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17485) );
  OAI21_X1 U20698 ( .B1(n17486), .B2(n17509), .A(n17485), .ZN(P3_U2755) );
  AOI22_X1 U20699 ( .A1(n17507), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17487) );
  OAI21_X1 U20700 ( .B1(n17488), .B2(n17509), .A(n17487), .ZN(P3_U2756) );
  AOI22_X1 U20701 ( .A1(n17507), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17489) );
  OAI21_X1 U20702 ( .B1(n17490), .B2(n17509), .A(n17489), .ZN(P3_U2757) );
  AOI22_X1 U20703 ( .A1(n17507), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17491) );
  OAI21_X1 U20704 ( .B1(n17544), .B2(n17509), .A(n17491), .ZN(P3_U2758) );
  INV_X1 U20705 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21090) );
  AOI22_X1 U20706 ( .A1(n17507), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17493) );
  OAI21_X1 U20707 ( .B1(n21090), .B2(n17509), .A(n17493), .ZN(P3_U2759) );
  INV_X1 U20708 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U20709 ( .A1(n17507), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17494) );
  OAI21_X1 U20710 ( .B1(n17495), .B2(n17509), .A(n17494), .ZN(P3_U2760) );
  INV_X1 U20711 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U20712 ( .A1(n17507), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17496) );
  OAI21_X1 U20713 ( .B1(n17497), .B2(n17509), .A(n17496), .ZN(P3_U2761) );
  INV_X1 U20714 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U20715 ( .A1(n17507), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17498) );
  OAI21_X1 U20716 ( .B1(n17537), .B2(n17509), .A(n17498), .ZN(P3_U2762) );
  INV_X1 U20717 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U20718 ( .A1(n17507), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17499) );
  OAI21_X1 U20719 ( .B1(n17500), .B2(n17509), .A(n17499), .ZN(P3_U2763) );
  AOI22_X1 U20720 ( .A1(n17507), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17501) );
  OAI21_X1 U20721 ( .B1(n17502), .B2(n17509), .A(n17501), .ZN(P3_U2764) );
  INV_X1 U20722 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17504) );
  AOI22_X1 U20723 ( .A1(n17507), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17503) );
  OAI21_X1 U20724 ( .B1(n17504), .B2(n17509), .A(n17503), .ZN(P3_U2765) );
  INV_X1 U20725 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17506) );
  AOI22_X1 U20726 ( .A1(n17507), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17505) );
  OAI21_X1 U20727 ( .B1(n17506), .B2(n17509), .A(n17505), .ZN(P3_U2766) );
  AOI22_X1 U20728 ( .A1(n17507), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17492), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U20729 ( .B1(n17510), .B2(n17509), .A(n17508), .ZN(P3_U2767) );
  OR3_X1 U20730 ( .A1(n18268), .A2(n17512), .A3(n17511), .ZN(n17559) );
  INV_X2 U20731 ( .A(n17559), .ZN(n17551) );
  AOI22_X1 U20732 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17542), .ZN(n17513) );
  OAI21_X1 U20733 ( .B1(n18263), .B2(n17553), .A(n17513), .ZN(P3_U2768) );
  AOI22_X1 U20734 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17542), .ZN(n17514) );
  OAI21_X1 U20735 ( .B1(n21108), .B2(n17553), .A(n17514), .ZN(P3_U2769) );
  AOI22_X1 U20736 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17542), .ZN(n17515) );
  OAI21_X1 U20737 ( .B1(n18271), .B2(n17553), .A(n17515), .ZN(P3_U2770) );
  AOI22_X1 U20738 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17542), .ZN(n17516) );
  OAI21_X1 U20739 ( .B1(n18276), .B2(n17553), .A(n17516), .ZN(P3_U2771) );
  AOI22_X1 U20740 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17542), .ZN(n17517) );
  OAI21_X1 U20741 ( .B1(n18280), .B2(n17553), .A(n17517), .ZN(P3_U2772) );
  AOI22_X1 U20742 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17557), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17542), .ZN(n17518) );
  OAI21_X1 U20743 ( .B1(n17519), .B2(n17559), .A(n17518), .ZN(P3_U2773) );
  AOI22_X1 U20744 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17542), .ZN(n17520) );
  OAI21_X1 U20745 ( .B1(n18288), .B2(n17553), .A(n17520), .ZN(P3_U2774) );
  AOI22_X1 U20746 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17542), .ZN(n17521) );
  OAI21_X1 U20747 ( .B1(n18293), .B2(n17553), .A(n17521), .ZN(P3_U2775) );
  AOI22_X1 U20748 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17542), .ZN(n17522) );
  OAI21_X1 U20749 ( .B1(n17541), .B2(n17553), .A(n17522), .ZN(P3_U2776) );
  INV_X1 U20750 ( .A(P3_UWORD_REG_9__SCAN_IN), .ZN(n21123) );
  AOI22_X1 U20751 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17557), .B1(
        P3_EAX_REG_25__SCAN_IN), .B2(n17551), .ZN(n17523) );
  OAI21_X1 U20752 ( .B1(n17524), .B2(n21123), .A(n17523), .ZN(P3_U2777) );
  AOI22_X1 U20753 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17542), .ZN(n17525) );
  OAI21_X1 U20754 ( .B1(n17546), .B2(n17553), .A(n17525), .ZN(P3_U2778) );
  AOI22_X1 U20755 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17542), .ZN(n17526) );
  OAI21_X1 U20756 ( .B1(n17548), .B2(n17553), .A(n17526), .ZN(P3_U2779) );
  AOI22_X1 U20757 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17542), .ZN(n17527) );
  OAI21_X1 U20758 ( .B1(n17550), .B2(n17553), .A(n17527), .ZN(P3_U2780) );
  AOI22_X1 U20759 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17551), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17542), .ZN(n17528) );
  OAI21_X1 U20760 ( .B1(n17554), .B2(n17553), .A(n17528), .ZN(P3_U2781) );
  AOI22_X1 U20761 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17557), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17542), .ZN(n17529) );
  OAI21_X1 U20762 ( .B1(n17530), .B2(n17559), .A(n17529), .ZN(P3_U2782) );
  AOI22_X1 U20763 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17542), .ZN(n17531) );
  OAI21_X1 U20764 ( .B1(n18263), .B2(n17553), .A(n17531), .ZN(P3_U2783) );
  AOI22_X1 U20765 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17542), .ZN(n17532) );
  OAI21_X1 U20766 ( .B1(n21108), .B2(n17553), .A(n17532), .ZN(P3_U2784) );
  AOI22_X1 U20767 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17542), .ZN(n17533) );
  OAI21_X1 U20768 ( .B1(n18271), .B2(n17553), .A(n17533), .ZN(P3_U2785) );
  AOI22_X1 U20769 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17542), .ZN(n17534) );
  OAI21_X1 U20770 ( .B1(n18276), .B2(n17553), .A(n17534), .ZN(P3_U2786) );
  AOI22_X1 U20771 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17542), .ZN(n17535) );
  OAI21_X1 U20772 ( .B1(n18280), .B2(n17553), .A(n17535), .ZN(P3_U2787) );
  AOI22_X1 U20773 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17557), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17542), .ZN(n17536) );
  OAI21_X1 U20774 ( .B1(n17537), .B2(n17559), .A(n17536), .ZN(P3_U2788) );
  AOI22_X1 U20775 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17542), .ZN(n17538) );
  OAI21_X1 U20776 ( .B1(n18288), .B2(n17553), .A(n17538), .ZN(P3_U2789) );
  AOI22_X1 U20777 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17542), .ZN(n17539) );
  OAI21_X1 U20778 ( .B1(n18293), .B2(n17553), .A(n17539), .ZN(P3_U2790) );
  AOI22_X1 U20779 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17542), .ZN(n17540) );
  OAI21_X1 U20780 ( .B1(n17541), .B2(n17553), .A(n17540), .ZN(P3_U2791) );
  AOI22_X1 U20781 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17557), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17542), .ZN(n17543) );
  OAI21_X1 U20782 ( .B1(n17544), .B2(n17559), .A(n17543), .ZN(P3_U2792) );
  AOI22_X1 U20783 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17542), .ZN(n17545) );
  OAI21_X1 U20784 ( .B1(n17546), .B2(n17553), .A(n17545), .ZN(P3_U2793) );
  AOI22_X1 U20785 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17542), .ZN(n17547) );
  OAI21_X1 U20786 ( .B1(n17548), .B2(n17553), .A(n17547), .ZN(P3_U2794) );
  AOI22_X1 U20787 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17542), .ZN(n17549) );
  OAI21_X1 U20788 ( .B1(n17550), .B2(n17553), .A(n17549), .ZN(P3_U2795) );
  AOI22_X1 U20789 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17551), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17542), .ZN(n17552) );
  OAI21_X1 U20790 ( .B1(n17554), .B2(n17553), .A(n17552), .ZN(P3_U2796) );
  AOI22_X1 U20791 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17557), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17542), .ZN(n17555) );
  OAI21_X1 U20792 ( .B1(n17556), .B2(n17559), .A(n17555), .ZN(P3_U2797) );
  AOI22_X1 U20793 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17557), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17542), .ZN(n17558) );
  OAI21_X1 U20794 ( .B1(n17560), .B2(n17559), .A(n17558), .ZN(P3_U2798) );
  OAI21_X1 U20795 ( .B1(n17561), .B2(n17928), .A(n17927), .ZN(n17562) );
  AOI21_X1 U20796 ( .B1(n17886), .B2(n17574), .A(n17562), .ZN(n17601) );
  OAI21_X1 U20797 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17715), .A(
        n17601), .ZN(n17585) );
  AOI22_X1 U20798 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17585), .B1(
        n17789), .B2(n17563), .ZN(n17579) );
  INV_X1 U20799 ( .A(n17564), .ZN(n17588) );
  NOR2_X1 U20800 ( .A1(n17842), .A2(n17916), .ZN(n17687) );
  OAI22_X1 U20801 ( .A1(n17565), .A2(n17761), .B1(n17940), .B2(n17932), .ZN(
        n17597) );
  NOR2_X1 U20802 ( .A1(n17944), .A2(n17597), .ZN(n17567) );
  NOR3_X1 U20803 ( .A1(n17687), .A2(n17567), .A3(n17566), .ZN(n17572) );
  AOI211_X1 U20804 ( .C1(n17570), .C2(n17569), .A(n17568), .B(n17845), .ZN(
        n17571) );
  AOI211_X1 U20805 ( .C1(n17573), .C2(n17588), .A(n17572), .B(n17571), .ZN(
        n17578) );
  NOR2_X1 U20806 ( .A1(n17769), .A2(n17574), .ZN(n17587) );
  OAI211_X1 U20807 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17587), .B(n17575), .ZN(n17576) );
  NAND4_X1 U20808 ( .A1(n17579), .A2(n17578), .A3(n17577), .A4(n17576), .ZN(
        P3_U2802) );
  NAND2_X1 U20809 ( .A1(n17581), .A2(n17580), .ZN(n17582) );
  XNOR2_X1 U20810 ( .A(n17745), .B(n17582), .ZN(n17948) );
  OAI22_X1 U20811 ( .A1(n18229), .A2(n18827), .B1(n17784), .B2(n17583), .ZN(
        n17584) );
  AOI221_X1 U20812 ( .B1(n17587), .B2(n17586), .C1(n17585), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17584), .ZN(n17590) );
  AOI22_X1 U20813 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17597), .B1(
        n17588), .B2(n17944), .ZN(n17589) );
  OAI211_X1 U20814 ( .C1(n17948), .C2(n17845), .A(n17590), .B(n17589), .ZN(
        P3_U2803) );
  AOI21_X1 U20815 ( .B1(n18636), .B2(n9726), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17600) );
  NOR2_X1 U20816 ( .A1(n18229), .A2(n18824), .ZN(n17954) );
  AOI221_X1 U20817 ( .B1(n17789), .B2(n17591), .C1(n17680), .C2(n17591), .A(
        n17954), .ZN(n17599) );
  INV_X1 U20818 ( .A(n17592), .ZN(n17595) );
  AOI21_X1 U20819 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17594), .A(
        n17593), .ZN(n17956) );
  OAI22_X1 U20820 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17595), .B1(
        n17956), .B2(n17845), .ZN(n17596) );
  AOI21_X1 U20821 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17597), .A(
        n17596), .ZN(n17598) );
  OAI211_X1 U20822 ( .C1(n17601), .C2(n17600), .A(n17599), .B(n17598), .ZN(
        P3_U2804) );
  AND2_X1 U20823 ( .A1(n17610), .A2(n18636), .ZN(n17637) );
  AOI211_X1 U20824 ( .C1(n17646), .C2(n17602), .A(n17884), .B(n17637), .ZN(
        n17635) );
  OAI21_X1 U20825 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17715), .A(
        n17635), .ZN(n17620) );
  AOI22_X1 U20826 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17620), .B1(
        n17789), .B2(n17603), .ZN(n17614) );
  NAND3_X1 U20827 ( .A1(n18065), .A2(n17623), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17604) );
  XNOR2_X1 U20828 ( .A(n17604), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17971) );
  NOR2_X1 U20829 ( .A1(n18075), .A2(n17624), .ZN(n17979) );
  NAND2_X1 U20830 ( .A1(n17979), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17605) );
  XNOR2_X1 U20831 ( .A(n17605), .B(n17949), .ZN(n17969) );
  OAI21_X1 U20832 ( .B1(n17834), .B2(n17607), .A(n17606), .ZN(n17608) );
  XNOR2_X1 U20833 ( .A(n17608), .B(n17949), .ZN(n17973) );
  OAI22_X1 U20834 ( .A1(n17932), .A2(n17969), .B1(n17845), .B2(n17973), .ZN(
        n17609) );
  AOI21_X1 U20835 ( .B1(n17842), .B2(n17971), .A(n17609), .ZN(n17613) );
  NAND2_X1 U20836 ( .A1(n9633), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17967) );
  NOR2_X1 U20837 ( .A1(n17769), .A2(n17610), .ZN(n17622) );
  OAI211_X1 U20838 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17622), .B(n17611), .ZN(n17612) );
  NAND4_X1 U20839 ( .A1(n17614), .A2(n17613), .A3(n17967), .A4(n17612), .ZN(
        P3_U2805) );
  AOI21_X1 U20840 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17616), .A(
        n17615), .ZN(n17985) );
  AOI22_X1 U20841 ( .A1(n9633), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17789), 
        .B2(n17617), .ZN(n17618) );
  INV_X1 U20842 ( .A(n17618), .ZN(n17619) );
  AOI221_X1 U20843 ( .B1(n17622), .B2(n17621), .C1(n17620), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17619), .ZN(n17628) );
  NAND2_X1 U20844 ( .A1(n18065), .A2(n17623), .ZN(n17976) );
  NAND2_X1 U20845 ( .A1(n17842), .A2(n17976), .ZN(n17640) );
  OAI21_X1 U20846 ( .B1(n17979), .B2(n17932), .A(n17640), .ZN(n17641) );
  NOR2_X1 U20847 ( .A1(n17624), .A2(n17738), .ZN(n17626) );
  AOI22_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17641), .B1(
        n17626), .B2(n17625), .ZN(n17627) );
  OAI211_X1 U20849 ( .C1(n17985), .C2(n17845), .A(n17628), .B(n17627), .ZN(
        P3_U2806) );
  AOI22_X1 U20850 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17834), .B1(
        n17629), .B2(n17655), .ZN(n17630) );
  NAND2_X1 U20851 ( .A1(n17676), .A2(n17630), .ZN(n17631) );
  XNOR2_X1 U20852 ( .A(n17631), .B(n17986), .ZN(n17991) );
  NAND2_X1 U20853 ( .A1(n9633), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17634) );
  OAI21_X1 U20854 ( .B1(n17789), .B2(n17680), .A(n17632), .ZN(n17633) );
  OAI211_X1 U20855 ( .C1(n17635), .C2(n9843), .A(n17634), .B(n17633), .ZN(
        n17636) );
  AOI21_X1 U20856 ( .B1(n17638), .B2(n17637), .A(n17636), .ZN(n17644) );
  OR2_X1 U20857 ( .A1(n17932), .A2(n17979), .ZN(n17639) );
  OAI22_X1 U20858 ( .A1(n17995), .A2(n17640), .B1(n18075), .B2(n17639), .ZN(
        n17642) );
  AOI22_X1 U20859 ( .A1(n17993), .A2(n17642), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17641), .ZN(n17643) );
  OAI211_X1 U20860 ( .C1(n17845), .C2(n17991), .A(n17644), .B(n17643), .ZN(
        P3_U2807) );
  AOI22_X1 U20861 ( .A1(n17646), .A2(n17645), .B1(n17886), .B2(n17648), .ZN(
        n17647) );
  NAND2_X1 U20862 ( .A1(n17647), .A2(n17927), .ZN(n17686) );
  AOI21_X1 U20863 ( .B1(n17680), .B2(n9836), .A(n17686), .ZN(n17667) );
  OR2_X1 U20864 ( .A1(n17648), .A2(n17769), .ZN(n17669) );
  OAI21_X1 U20865 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17649), .ZN(n17650) );
  OAI22_X1 U20866 ( .A1(n17667), .A2(n17651), .B1(n17669), .B2(n17650), .ZN(
        n17652) );
  AOI21_X1 U20867 ( .B1(n17789), .B2(n17653), .A(n17652), .ZN(n17661) );
  INV_X1 U20868 ( .A(n18002), .ZN(n17656) );
  NOR2_X1 U20869 ( .A1(n17712), .A2(n17656), .ZN(n17994) );
  AOI22_X1 U20870 ( .A1(n17842), .A2(n17995), .B1(n17916), .B2(n18075), .ZN(
        n17737) );
  OAI21_X1 U20871 ( .B1(n17687), .B2(n17994), .A(n17737), .ZN(n17673) );
  INV_X1 U20872 ( .A(n17676), .ZN(n17654) );
  AOI221_X1 U20873 ( .B1(n17656), .B2(n17655), .C1(n17662), .C2(n17655), .A(
        n17654), .ZN(n17657) );
  XOR2_X1 U20874 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17657), .Z(
        n18003) );
  AOI22_X1 U20875 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17673), .B1(
        n17829), .B2(n18003), .ZN(n17660) );
  NAND2_X1 U20876 ( .A1(n9633), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18004) );
  INV_X1 U20877 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17658) );
  NAND3_X1 U20878 ( .A1(n17723), .A2(n17994), .A3(n17658), .ZN(n17659) );
  NAND4_X1 U20879 ( .A1(n17661), .A2(n17660), .A3(n18004), .A4(n17659), .ZN(
        P3_U2808) );
  INV_X1 U20880 ( .A(n17672), .ZN(n18015) );
  NOR3_X1 U20881 ( .A1(n17834), .A2(n21089), .A3(n17662), .ZN(n17690) );
  INV_X1 U20882 ( .A(n17710), .ZN(n17691) );
  AOI22_X1 U20883 ( .A1(n18015), .A2(n17690), .B1(n17691), .B2(n17663), .ZN(
        n17665) );
  XNOR2_X1 U20884 ( .A(n17665), .B(n17664), .ZN(n18020) );
  NAND2_X1 U20885 ( .A1(n9633), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17666) );
  OAI221_X1 U20886 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17669), .C1(
        n17668), .C2(n17667), .A(n17666), .ZN(n17670) );
  AOI21_X1 U20887 ( .B1(n17789), .B2(n17671), .A(n17670), .ZN(n17675) );
  NOR2_X1 U20888 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17672), .ZN(
        n18009) );
  NOR2_X1 U20889 ( .A1(n17712), .A2(n21089), .ZN(n18011) );
  AND2_X1 U20890 ( .A1(n17723), .A2(n18011), .ZN(n17699) );
  AOI22_X1 U20891 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17673), .B1(
        n18009), .B2(n17699), .ZN(n17674) );
  OAI211_X1 U20892 ( .C1(n18020), .C2(n17845), .A(n17675), .B(n17674), .ZN(
        P3_U2809) );
  OAI221_X1 U20893 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17709), 
        .C1(n18028), .C2(n17690), .A(n17676), .ZN(n17677) );
  XOR2_X1 U20894 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17677), .Z(
        n18027) );
  AOI21_X1 U20895 ( .B1(n17678), .B2(n18636), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17679) );
  INV_X1 U20896 ( .A(n17679), .ZN(n17685) );
  NOR2_X1 U20897 ( .A1(n18229), .A2(n18814), .ZN(n17684) );
  INV_X1 U20898 ( .A(n17681), .ZN(n17682) );
  AOI21_X1 U20899 ( .B1(n17784), .B2(n17715), .A(n17682), .ZN(n17683) );
  AOI211_X1 U20900 ( .C1(n17686), .C2(n17685), .A(n17684), .B(n17683), .ZN(
        n17689) );
  NAND2_X1 U20901 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18011), .ZN(
        n17996) );
  INV_X1 U20902 ( .A(n17996), .ZN(n18022) );
  OAI21_X1 U20903 ( .B1(n17687), .B2(n18022), .A(n17737), .ZN(n17700) );
  NOR2_X1 U20904 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18028), .ZN(
        n18021) );
  AOI22_X1 U20905 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17700), .B1(
        n18021), .B2(n17699), .ZN(n17688) );
  OAI211_X1 U20906 ( .C1(n17845), .C2(n18027), .A(n17689), .B(n17688), .ZN(
        P3_U2810) );
  AOI21_X1 U20907 ( .B1(n17691), .B2(n17709), .A(n17690), .ZN(n17692) );
  XNOR2_X1 U20908 ( .A(n17692), .B(n18028), .ZN(n18033) );
  AOI21_X1 U20909 ( .B1(n17886), .B2(n17694), .A(n17884), .ZN(n17717) );
  OAI21_X1 U20910 ( .B1(n17693), .B2(n17928), .A(n17717), .ZN(n17706) );
  NAND2_X1 U20911 ( .A1(n9633), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18031) );
  NOR2_X1 U20912 ( .A1(n17769), .A2(n17694), .ZN(n17708) );
  OAI211_X1 U20913 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17708), .B(n17695), .ZN(n17696) );
  OAI211_X1 U20914 ( .C1(n17784), .C2(n17697), .A(n18031), .B(n17696), .ZN(
        n17698) );
  AOI21_X1 U20915 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17706), .A(
        n17698), .ZN(n17702) );
  AOI22_X1 U20916 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17700), .B1(
        n17699), .B2(n18028), .ZN(n17701) );
  OAI211_X1 U20917 ( .C1(n18033), .C2(n17845), .A(n17702), .B(n17701), .ZN(
        P3_U2811) );
  INV_X1 U20918 ( .A(n17737), .ZN(n17703) );
  AOI21_X1 U20919 ( .B1(n17723), .B2(n17712), .A(n17703), .ZN(n17726) );
  INV_X1 U20920 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17707) );
  OAI22_X1 U20921 ( .A1(n18229), .A2(n18809), .B1(n17784), .B2(n17704), .ZN(
        n17705) );
  AOI221_X1 U20922 ( .B1(n17708), .B2(n17707), .C1(n17706), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17705), .ZN(n17714) );
  AOI21_X1 U20923 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17745), .A(
        n17709), .ZN(n17711) );
  XNOR2_X1 U20924 ( .A(n17711), .B(n17710), .ZN(n18047) );
  NOR2_X1 U20925 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17712), .ZN(
        n18046) );
  AOI22_X1 U20926 ( .A1(n17829), .A2(n18047), .B1(n17723), .B2(n18046), .ZN(
        n17713) );
  OAI211_X1 U20927 ( .C1(n17726), .C2(n21089), .A(n17714), .B(n17713), .ZN(
        P3_U2812) );
  AOI21_X1 U20928 ( .B1(n17716), .B2(n18636), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17718) );
  OAI22_X1 U20929 ( .A1(n17718), .A2(n17717), .B1(n18229), .B2(n18808), .ZN(
        n17719) );
  AOI21_X1 U20930 ( .B1(n17720), .B2(n17919), .A(n17719), .ZN(n17725) );
  OAI21_X1 U20931 ( .B1(n17722), .B2(n21117), .A(n17721), .ZN(n18052) );
  NOR2_X1 U20932 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18059), .ZN(
        n18051) );
  AOI22_X1 U20933 ( .A1(n17829), .A2(n18052), .B1(n17723), .B2(n18051), .ZN(
        n17724) );
  OAI211_X1 U20934 ( .C1(n17726), .C2(n21117), .A(n17725), .B(n17724), .ZN(
        P3_U2813) );
  NAND2_X1 U20935 ( .A1(n17745), .A2(n13354), .ZN(n17820) );
  OAI22_X1 U20936 ( .A1(n17745), .A2(n17727), .B1(n17820), .B2(n18045), .ZN(
        n17728) );
  XNOR2_X1 U20937 ( .A(n18059), .B(n17728), .ZN(n18061) );
  AOI21_X1 U20938 ( .B1(n17886), .B2(n17730), .A(n17884), .ZN(n17766) );
  OAI21_X1 U20939 ( .B1(n17729), .B2(n17928), .A(n17766), .ZN(n17741) );
  AOI22_X1 U20940 ( .A1(n9633), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17741), .ZN(n17733) );
  NOR2_X1 U20941 ( .A1(n17769), .A2(n17730), .ZN(n17743) );
  OAI211_X1 U20942 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17743), .B(n17731), .ZN(n17732) );
  OAI211_X1 U20943 ( .C1(n17734), .C2(n17784), .A(n17733), .B(n17732), .ZN(
        n17735) );
  AOI21_X1 U20944 ( .B1(n17829), .B2(n18061), .A(n17735), .ZN(n17736) );
  OAI221_X1 U20945 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17738), 
        .C1(n18059), .C2(n17737), .A(n17736), .ZN(P3_U2814) );
  NOR2_X1 U20946 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18076), .ZN(
        n17754) );
  NAND2_X1 U20947 ( .A1(n17916), .A2(n18075), .ZN(n17753) );
  OAI22_X1 U20948 ( .A1(n18229), .A2(n18804), .B1(n17784), .B2(n17739), .ZN(
        n17740) );
  AOI221_X1 U20949 ( .B1(n17743), .B2(n17742), .C1(n17741), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17740), .ZN(n17752) );
  NOR2_X1 U20950 ( .A1(n17745), .A2(n17744), .ZN(n17811) );
  AOI22_X1 U20951 ( .A1(n13354), .A2(n17747), .B1(n17785), .B2(n17779), .ZN(
        n17748) );
  AOI221_X1 U20952 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17796), 
        .C1(n17834), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17748), .ZN(
        n17749) );
  XNOR2_X1 U20953 ( .A(n17749), .B(n18072), .ZN(n18074) );
  NOR2_X1 U20954 ( .A1(n18065), .A2(n17761), .ZN(n17750) );
  NAND2_X1 U20955 ( .A1(n17759), .A2(n18072), .ZN(n18070) );
  AOI22_X1 U20956 ( .A1(n17829), .A2(n18074), .B1(n17750), .B2(n18070), .ZN(
        n17751) );
  OAI211_X1 U20957 ( .C1(n17754), .C2(n17753), .A(n17752), .B(n17751), .ZN(
        P3_U2815) );
  INV_X1 U20958 ( .A(n17800), .ZN(n17770) );
  NOR2_X1 U20959 ( .A1(n18363), .A2(n17770), .ZN(n17755) );
  AOI21_X1 U20960 ( .B1(n17771), .B2(n17755), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U20961 ( .A1(n9633), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17756), 
        .B2(n17919), .ZN(n17764) );
  AOI221_X1 U20962 ( .B1(n18117), .B2(n18086), .C1(n18067), .C2(n18086), .A(
        n18076), .ZN(n18090) );
  INV_X1 U20963 ( .A(n18067), .ZN(n18080) );
  INV_X1 U20964 ( .A(n17820), .ZN(n17812) );
  AOI22_X1 U20965 ( .A1(n18080), .A2(n17812), .B1(n17757), .B2(n17785), .ZN(
        n17758) );
  XNOR2_X1 U20966 ( .A(n17758), .B(n18086), .ZN(n18094) );
  OAI21_X1 U20967 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17760), .A(
        n17759), .ZN(n18089) );
  OAI22_X1 U20968 ( .A1(n18094), .A2(n17845), .B1(n17761), .B2(n18089), .ZN(
        n17762) );
  AOI21_X1 U20969 ( .B1(n17916), .B2(n18090), .A(n17762), .ZN(n17763) );
  OAI211_X1 U20970 ( .C1(n17766), .C2(n17765), .A(n17764), .B(n17763), .ZN(
        P3_U2816) );
  AOI21_X1 U20971 ( .B1(n17886), .B2(n17770), .A(n17884), .ZN(n17767) );
  OAI21_X1 U20972 ( .B1(n17768), .B2(n17928), .A(n17767), .ZN(n17790) );
  NOR2_X1 U20973 ( .A1(n18229), .A2(n18800), .ZN(n17775) );
  OR2_X1 U20974 ( .A1(n17770), .A2(n17769), .ZN(n17792) );
  AOI211_X1 U20975 ( .C1(n17773), .C2(n17772), .A(n17771), .B(n17792), .ZN(
        n17774) );
  AOI211_X1 U20976 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17790), .A(
        n17775), .B(n17774), .ZN(n17782) );
  NOR2_X1 U20977 ( .A1(n18096), .A2(n17820), .ZN(n17786) );
  AOI22_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17786), .B1(
        n17785), .B2(n17796), .ZN(n17776) );
  XNOR2_X1 U20979 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17776), .ZN(
        n18095) );
  NAND2_X1 U20980 ( .A1(n18106), .A2(n17779), .ZN(n18104) );
  NAND2_X1 U20981 ( .A1(n17777), .A2(n18106), .ZN(n18097) );
  NAND2_X1 U20982 ( .A1(n18106), .A2(n17778), .ZN(n18098) );
  AOI22_X1 U20983 ( .A1(n17842), .A2(n18097), .B1(n17916), .B2(n18098), .ZN(
        n17797) );
  OAI22_X1 U20984 ( .A1(n17832), .A2(n18104), .B1(n17797), .B2(n17779), .ZN(
        n17780) );
  AOI21_X1 U20985 ( .B1(n17829), .B2(n18095), .A(n17780), .ZN(n17781) );
  OAI211_X1 U20986 ( .C1(n17784), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        P3_U2817) );
  NOR2_X1 U20987 ( .A1(n17786), .A2(n17785), .ZN(n17787) );
  XNOR2_X1 U20988 ( .A(n17787), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18109) );
  NOR3_X1 U20989 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17832), .A3(
        n18096), .ZN(n17794) );
  AOI22_X1 U20990 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17790), .B1(
        n17789), .B2(n17788), .ZN(n17791) );
  NAND2_X1 U20991 ( .A1(n9633), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18110) );
  OAI211_X1 U20992 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17792), .A(
        n17791), .B(n18110), .ZN(n17793) );
  AOI211_X1 U20993 ( .C1(n17829), .C2(n18109), .A(n17794), .B(n17793), .ZN(
        n17795) );
  OAI21_X1 U20994 ( .B1(n17797), .B2(n17796), .A(n17795), .ZN(P3_U2818) );
  INV_X1 U20995 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17798) );
  NAND2_X1 U20996 ( .A1(n18123), .A2(n17798), .ZN(n18128) );
  NAND4_X1 U20997 ( .A1(n18636), .A2(n9725), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17825) );
  NOR2_X1 U20998 ( .A1(n17824), .A2(n17825), .ZN(n17823) );
  NAND2_X1 U20999 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17823), .ZN(
        n17810) );
  NAND2_X1 U21000 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17868), .ZN(
        n17799) );
  AOI22_X1 U21001 ( .A1(n18636), .A2(n17800), .B1(n17810), .B2(n17799), .ZN(
        n17802) );
  NOR2_X1 U21002 ( .A1(n18229), .A2(n18796), .ZN(n17801) );
  AOI211_X1 U21003 ( .C1(n17803), .C2(n17919), .A(n17802), .B(n17801), .ZN(
        n17807) );
  AOI22_X1 U21004 ( .A1(n17842), .A2(n18115), .B1(n17916), .B2(n18117), .ZN(
        n17831) );
  OAI21_X1 U21005 ( .B1(n18123), .B2(n17832), .A(n17831), .ZN(n17805) );
  INV_X1 U21006 ( .A(n17811), .ZN(n17821) );
  OAI33_X1 U21007 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n17821), .B1(n18148), .B2(
        n17820), .B3(n17814), .ZN(n17804) );
  XOR2_X1 U21008 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17804), .Z(
        n18114) );
  AOI22_X1 U21009 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17805), .B1(
        n17829), .B2(n18114), .ZN(n17806) );
  OAI211_X1 U21010 ( .C1(n17832), .C2(n18128), .A(n17807), .B(n17806), .ZN(
        P3_U2819) );
  AOI21_X1 U21011 ( .B1(n17868), .B2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17823), .ZN(n17808) );
  INV_X1 U21012 ( .A(n17808), .ZN(n17809) );
  AOI22_X1 U21013 ( .A1(n9633), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17810), 
        .B2(n17809), .ZN(n17818) );
  AOI22_X1 U21014 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17812), .B1(
        n17811), .B2(n18148), .ZN(n17813) );
  XNOR2_X1 U21015 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17813), .ZN(
        n18134) );
  AOI22_X1 U21016 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17814), .B1(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18148), .ZN(n17815) );
  OAI22_X1 U21017 ( .A1(n17832), .A2(n17815), .B1(n17831), .B2(n17814), .ZN(
        n17816) );
  AOI21_X1 U21018 ( .B1(n17829), .B2(n18134), .A(n17816), .ZN(n17817) );
  OAI211_X1 U21019 ( .C1(n17910), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        P3_U2820) );
  NAND2_X1 U21020 ( .A1(n17821), .A2(n17820), .ZN(n17822) );
  XNOR2_X1 U21021 ( .A(n17822), .B(n18148), .ZN(n18144) );
  AOI211_X1 U21022 ( .C1(n17825), .C2(n17824), .A(n17924), .B(n17823), .ZN(
        n17828) );
  OAI22_X1 U21023 ( .A1(n17910), .A2(n17826), .B1(n18229), .B2(n18792), .ZN(
        n17827) );
  AOI211_X1 U21024 ( .C1(n17829), .C2(n18144), .A(n17828), .B(n17827), .ZN(
        n17830) );
  OAI221_X1 U21025 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17832), .C1(
        n18148), .C2(n17831), .A(n17830), .ZN(P3_U2821) );
  OAI21_X1 U21026 ( .B1(n18164), .B2(n17834), .A(n17833), .ZN(n18167) );
  INV_X1 U21027 ( .A(n9725), .ZN(n17847) );
  AOI21_X1 U21028 ( .B1(n17886), .B2(n17847), .A(n17884), .ZN(n17846) );
  OAI211_X1 U21029 ( .C1(n17836), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n18636), .B(n17835), .ZN(n17837) );
  NAND2_X1 U21030 ( .A1(n9633), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18157) );
  OAI211_X1 U21031 ( .C1(n20983), .C2(n17846), .A(n17837), .B(n18157), .ZN(
        n17838) );
  AOI21_X1 U21032 ( .B1(n17839), .B2(n17919), .A(n17838), .ZN(n17844) );
  AOI21_X1 U21033 ( .B1(n17841), .B2(n18160), .A(n17840), .ZN(n18162) );
  AOI22_X1 U21034 ( .A1(n17842), .A2(n18164), .B1(n17916), .B2(n18162), .ZN(
        n17843) );
  OAI211_X1 U21035 ( .C1(n17845), .C2(n18167), .A(n17844), .B(n17843), .ZN(
        P3_U2822) );
  INV_X1 U21036 ( .A(n17846), .ZN(n17848) );
  NOR2_X1 U21037 ( .A1(n18363), .A2(n17847), .ZN(n17867) );
  NOR2_X1 U21038 ( .A1(n18229), .A2(n18788), .ZN(n18170) );
  AOI221_X1 U21039 ( .B1(n17848), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17867), .C2(n9822), .A(n18170), .ZN(n17855) );
  AOI21_X1 U21040 ( .B1(n18154), .B2(n17850), .A(n17849), .ZN(n18172) );
  NAND2_X1 U21041 ( .A1(n17852), .A2(n17851), .ZN(n17853) );
  XNOR2_X1 U21042 ( .A(n17853), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18173) );
  AOI22_X1 U21043 ( .A1(n17920), .A2(n18172), .B1(n17916), .B2(n18173), .ZN(
        n17854) );
  OAI211_X1 U21044 ( .C1(n17910), .C2(n17856), .A(n17855), .B(n17854), .ZN(
        P3_U2823) );
  NOR2_X1 U21045 ( .A1(n18363), .A2(n17857), .ZN(n17879) );
  AOI21_X1 U21046 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17868), .A(
        n17879), .ZN(n17866) );
  AOI21_X1 U21047 ( .B1(n17860), .B2(n17859), .A(n17858), .ZN(n18180) );
  AOI22_X1 U21048 ( .A1(n17920), .A2(n18180), .B1(n9633), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17865) );
  AOI21_X1 U21049 ( .B1(n18155), .B2(n17862), .A(n17861), .ZN(n18181) );
  AOI22_X1 U21050 ( .A1(n17916), .A2(n18181), .B1(n17863), .B2(n17919), .ZN(
        n17864) );
  OAI211_X1 U21051 ( .C1(n17867), .C2(n17866), .A(n17865), .B(n17864), .ZN(
        P3_U2824) );
  OAI221_X1 U21052 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n9823), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17927), .A(n17868), .ZN(n17878) );
  AOI21_X1 U21053 ( .B1(n17870), .B2(n17869), .A(n9723), .ZN(n17871) );
  XNOR2_X1 U21054 ( .A(n17871), .B(n9867), .ZN(n18186) );
  AOI22_X1 U21055 ( .A1(n17920), .A2(n18186), .B1(n9633), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17877) );
  AOI21_X1 U21056 ( .B1(n17874), .B2(n17873), .A(n17872), .ZN(n18187) );
  AOI22_X1 U21057 ( .A1(n17916), .A2(n18187), .B1(n17875), .B2(n17919), .ZN(
        n17876) );
  OAI211_X1 U21058 ( .C1(n17879), .C2(n17878), .A(n17877), .B(n17876), .ZN(
        P3_U2825) );
  AOI21_X1 U21059 ( .B1(n18202), .B2(n17881), .A(n17880), .ZN(n18199) );
  AOI22_X1 U21060 ( .A1(n17916), .A2(n18199), .B1(n9633), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n17891) );
  AOI21_X1 U21061 ( .B1(n17886), .B2(n17885), .A(n17884), .ZN(n17903) );
  OAI22_X1 U21062 ( .A1(n17910), .A2(n17888), .B1(n17903), .B2(n17887), .ZN(
        n17889) );
  AOI21_X1 U21063 ( .B1(n17920), .B2(n18197), .A(n17889), .ZN(n17890) );
  OAI211_X1 U21064 ( .C1(n18363), .C2(n17892), .A(n17891), .B(n17890), .ZN(
        P3_U2826) );
  AOI21_X1 U21065 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17927), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17902) );
  AOI21_X1 U21066 ( .B1(n17895), .B2(n17894), .A(n17893), .ZN(n18205) );
  AOI22_X1 U21067 ( .A1(n17916), .A2(n18205), .B1(n9633), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17901) );
  AOI21_X1 U21068 ( .B1(n17898), .B2(n17897), .A(n17896), .ZN(n18204) );
  AOI22_X1 U21069 ( .A1(n17920), .A2(n18204), .B1(n17899), .B2(n17919), .ZN(
        n17900) );
  OAI211_X1 U21070 ( .C1(n17903), .C2(n17902), .A(n17901), .B(n17900), .ZN(
        P3_U2827) );
  INV_X1 U21071 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17913) );
  AOI21_X1 U21072 ( .B1(n17906), .B2(n17905), .A(n17904), .ZN(n18222) );
  INV_X1 U21073 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18778) );
  NOR2_X1 U21074 ( .A1(n18229), .A2(n18778), .ZN(n18224) );
  XNOR2_X1 U21075 ( .A(n17908), .B(n17907), .ZN(n18221) );
  OAI22_X1 U21076 ( .A1(n17910), .A2(n17909), .B1(n17932), .B2(n18221), .ZN(
        n17911) );
  AOI211_X1 U21077 ( .C1(n17920), .C2(n18222), .A(n18224), .B(n17911), .ZN(
        n17912) );
  OAI221_X1 U21078 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18363), .C1(
        n17913), .C2(n17927), .A(n17912), .ZN(P3_U2828) );
  NOR2_X1 U21079 ( .A1(n17926), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17914) );
  XOR2_X1 U21080 ( .A(n17914), .B(n17918), .Z(n18241) );
  INV_X1 U21081 ( .A(n18241), .ZN(n17915) );
  AOI22_X1 U21082 ( .A1(n17916), .A2(n17915), .B1(n9633), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17922) );
  AOI21_X1 U21083 ( .B1(n17925), .B2(n17918), .A(n17917), .ZN(n18234) );
  AOI22_X1 U21084 ( .A1(n17920), .A2(n18234), .B1(n17923), .B2(n17919), .ZN(
        n17921) );
  OAI211_X1 U21085 ( .C1(n17924), .C2(n17923), .A(n17922), .B(n17921), .ZN(
        P3_U2829) );
  OAI21_X1 U21086 ( .B1(n17926), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17925), .ZN(n18249) );
  INV_X1 U21087 ( .A(n18249), .ZN(n17933) );
  NAND3_X1 U21088 ( .A1(n18859), .A2(n17928), .A3(n17927), .ZN(n17929) );
  AOI22_X1 U21089 ( .A1(n9633), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17929), .ZN(n17930) );
  OAI221_X1 U21090 ( .B1(n17933), .B2(n17932), .C1(n18249), .C2(n17931), .A(
        n17930), .ZN(P3_U2830) );
  AOI22_X1 U21091 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18237), .B1(
        n9633), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17947) );
  INV_X1 U21092 ( .A(n17962), .ZN(n17957) );
  NOR2_X1 U21093 ( .A1(n18712), .A2(n18723), .ZN(n18195) );
  AOI21_X1 U21094 ( .B1(n17935), .B2(n17958), .A(n18195), .ZN(n17936) );
  NOR2_X1 U21095 ( .A1(n18212), .A2(n17936), .ZN(n17978) );
  OAI21_X1 U21096 ( .B1(n17957), .B2(n18195), .A(n17978), .ZN(n17961) );
  AOI22_X1 U21097 ( .A1(n18712), .A2(n17949), .B1(n18723), .B2(n17937), .ZN(
        n17939) );
  OAI211_X1 U21098 ( .C1(n17940), .C2(n18220), .A(n17939), .B(n17938), .ZN(
        n17941) );
  AOI211_X1 U21099 ( .C1(n18116), .C2(n17942), .A(n17961), .B(n17941), .ZN(
        n17952) );
  OAI21_X1 U21100 ( .B1(n18243), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17952), .ZN(n17943) );
  OAI221_X1 U21101 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17945), 
        .C1(n17944), .C2(n17943), .A(n18242), .ZN(n17946) );
  OAI211_X1 U21102 ( .C1(n17948), .C2(n18168), .A(n17947), .B(n17946), .ZN(
        P3_U2835) );
  NAND2_X1 U21103 ( .A1(n18242), .A2(n18001), .ZN(n18008) );
  NOR4_X1 U21104 ( .A1(n17974), .A2(n17962), .A3(n17949), .A4(n18008), .ZN(
        n17950) );
  AOI21_X1 U21105 ( .B1(n18242), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17950), .ZN(n17951) );
  AOI21_X1 U21106 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17952), .A(
        n17951), .ZN(n17953) );
  AOI211_X1 U21107 ( .C1(n18237), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17954), .B(n17953), .ZN(n17955) );
  OAI21_X1 U21108 ( .B1(n17956), .B2(n18168), .A(n17955), .ZN(P3_U2836) );
  NAND2_X1 U21109 ( .A1(n17958), .A2(n17957), .ZN(n17959) );
  NOR2_X1 U21110 ( .A1(n17960), .A2(n17959), .ZN(n17965) );
  AOI221_X1 U21111 ( .B1(n17962), .B2(n18691), .C1(n17980), .C2(n18691), .A(
        n17961), .ZN(n17963) );
  INV_X1 U21112 ( .A(n17963), .ZN(n17964) );
  MUX2_X1 U21113 ( .A(n17965), .B(n17964), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n17966) );
  AOI22_X1 U21114 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18237), .B1(
        n18242), .B2(n17966), .ZN(n17968) );
  OAI211_X1 U21115 ( .C1(n17969), .C2(n18240), .A(n17968), .B(n17967), .ZN(
        n17970) );
  AOI21_X1 U21116 ( .B1(n18163), .B2(n17971), .A(n17970), .ZN(n17972) );
  OAI21_X1 U21117 ( .B1(n18168), .B2(n17973), .A(n17972), .ZN(P3_U2837) );
  NOR4_X1 U21118 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17986), .A3(
        n17974), .A4(n18008), .ZN(n17975) );
  AOI21_X1 U21119 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n9633), .A(n17975), .ZN(
        n17984) );
  AOI21_X1 U21120 ( .B1(n18116), .B2(n17976), .A(n18237), .ZN(n17977) );
  OAI211_X1 U21121 ( .C1(n17979), .C2(n18220), .A(n17978), .B(n17977), .ZN(
        n17982) );
  AOI211_X1 U21122 ( .C1(n18691), .C2(n17980), .A(n17986), .B(n17982), .ZN(
        n17981) );
  NOR2_X1 U21123 ( .A1(n9633), .A2(n17981), .ZN(n17989) );
  OAI211_X1 U21124 ( .C1(n18156), .C2(n17982), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17989), .ZN(n17983) );
  OAI211_X1 U21125 ( .C1(n17985), .C2(n18168), .A(n17984), .B(n17983), .ZN(
        P3_U2838) );
  OAI21_X1 U21126 ( .B1(n18237), .B2(n17987), .A(n17986), .ZN(n17988) );
  AOI22_X1 U21127 ( .A1(n9633), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17989), 
        .B2(n17988), .ZN(n17990) );
  OAI21_X1 U21128 ( .B1(n18168), .B2(n17991), .A(n17990), .ZN(P3_U2839) );
  NOR2_X1 U21129 ( .A1(n18876), .A2(n18137), .ZN(n18141) );
  NAND2_X1 U21130 ( .A1(n17992), .A2(n18141), .ZN(n18055) );
  INV_X1 U21131 ( .A(n18055), .ZN(n18010) );
  AOI22_X1 U21132 ( .A1(n17934), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n17993), .B2(n18010), .ZN(n18000) );
  NOR2_X1 U21133 ( .A1(n15702), .A2(n18116), .ZN(n18122) );
  OAI22_X1 U21134 ( .A1(n18129), .A2(n18015), .B1(n18122), .B2(n17994), .ZN(
        n18017) );
  AOI22_X1 U21135 ( .A1(n15702), .A2(n18075), .B1(n18116), .B2(n17995), .ZN(
        n18012) );
  OAI21_X1 U21136 ( .B1(n18036), .B2(n17996), .A(n18712), .ZN(n17997) );
  OAI221_X1 U21137 ( .B1(n18731), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n18731), .C2(n18034), .A(n17997), .ZN(n18013) );
  INV_X1 U21138 ( .A(n18013), .ZN(n17998) );
  OAI211_X1 U21139 ( .C1(n18129), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n18012), .B(n17998), .ZN(n17999) );
  NOR3_X1 U21140 ( .A1(n18000), .A2(n18017), .A3(n17999), .ZN(n18007) );
  OAI221_X1 U21141 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18002), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18001), .A(n18242), .ZN(
        n18006) );
  AOI22_X1 U21142 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18237), .B1(
        n18145), .B2(n18003), .ZN(n18005) );
  OAI211_X1 U21143 ( .C1(n18007), .C2(n18006), .A(n18005), .B(n18004), .ZN(
        P3_U2840) );
  NOR2_X1 U21144 ( .A1(n21089), .A2(n18008), .ZN(n18029) );
  AOI22_X1 U21145 ( .A1(n9633), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18029), 
        .B2(n18009), .ZN(n18019) );
  AOI21_X1 U21146 ( .B1(n18011), .B2(n18010), .A(n17934), .ZN(n18014) );
  NAND2_X1 U21147 ( .A1(n18242), .A2(n18012), .ZN(n18058) );
  NOR3_X1 U21148 ( .A1(n18014), .A2(n18058), .A3(n18013), .ZN(n18023) );
  OAI21_X1 U21149 ( .B1(n17934), .B2(n18015), .A(n18023), .ZN(n18016) );
  OAI211_X1 U21150 ( .C1(n18017), .C2(n18016), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18229), .ZN(n18018) );
  OAI211_X1 U21151 ( .C1(n18020), .C2(n18168), .A(n18019), .B(n18018), .ZN(
        P3_U2841) );
  AOI22_X1 U21152 ( .A1(n9633), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18029), 
        .B2(n18021), .ZN(n18026) );
  AOI221_X1 U21153 ( .B1(n18122), .B2(n18023), .C1(n18022), .C2(n18023), .A(
        n9633), .ZN(n18030) );
  NOR2_X1 U21154 ( .A1(n18691), .A2(n18723), .ZN(n18236) );
  NOR3_X1 U21155 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18236), .A3(
        n18910), .ZN(n18024) );
  OAI21_X1 U21156 ( .B1(n18030), .B2(n18024), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18025) );
  OAI211_X1 U21157 ( .C1(n18027), .C2(n18168), .A(n18026), .B(n18025), .ZN(
        P3_U2842) );
  AOI22_X1 U21158 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18030), .B1(
        n18029), .B2(n18028), .ZN(n18032) );
  OAI211_X1 U21159 ( .C1(n18033), .C2(n18168), .A(n18032), .B(n18031), .ZN(
        P3_U2843) );
  INV_X1 U21160 ( .A(n18034), .ZN(n18035) );
  AOI211_X1 U21161 ( .C1(n18691), .C2(n18035), .A(n18212), .B(n18058), .ZN(
        n18038) );
  INV_X1 U21162 ( .A(n18195), .ZN(n18211) );
  OAI21_X1 U21163 ( .B1(n18059), .B2(n18036), .A(n18211), .ZN(n18037) );
  OAI211_X1 U21164 ( .C1(n18039), .C2(n18122), .A(n18038), .B(n18037), .ZN(
        n18050) );
  OAI221_X1 U21165 ( .B1(n18050), .B2(n21117), .C1(n18050), .C2(n18211), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18049) );
  INV_X1 U21166 ( .A(n18217), .ZN(n18041) );
  OAI22_X1 U21167 ( .A1(n18731), .A2(n18216), .B1(n18041), .B2(n18040), .ZN(
        n18207) );
  INV_X1 U21168 ( .A(n18207), .ZN(n18188) );
  NOR2_X1 U21169 ( .A1(n18188), .A2(n18042), .ZN(n18169) );
  NAND2_X1 U21170 ( .A1(n18043), .A2(n18169), .ZN(n18066) );
  NAND2_X1 U21171 ( .A1(n18044), .A2(n18066), .ZN(n18105) );
  NAND2_X1 U21172 ( .A1(n18242), .A2(n18105), .ZN(n18149) );
  NOR2_X1 U21173 ( .A1(n18045), .A2(n18149), .ZN(n18060) );
  AOI22_X1 U21174 ( .A1(n18145), .A2(n18047), .B1(n18060), .B2(n18046), .ZN(
        n18048) );
  OAI221_X1 U21175 ( .B1(n9633), .B2(n18049), .C1(n18229), .C2(n18809), .A(
        n18048), .ZN(P3_U2844) );
  NAND2_X1 U21176 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18050), .ZN(
        n18054) );
  AOI22_X1 U21177 ( .A1(n18145), .A2(n18052), .B1(n18060), .B2(n18051), .ZN(
        n18053) );
  OAI221_X1 U21178 ( .B1(n9633), .B2(n18054), .C1(n18229), .C2(n18808), .A(
        n18053), .ZN(P3_U2845) );
  AOI22_X1 U21179 ( .A1(n18691), .A2(n18138), .B1(n18712), .B2(n18137), .ZN(
        n18121) );
  OAI21_X1 U21180 ( .B1(n18072), .B2(n18723), .A(n18055), .ZN(n18056) );
  OAI211_X1 U21181 ( .C1(n18129), .C2(n18057), .A(n18121), .B(n18056), .ZN(
        n18069) );
  OAI221_X1 U21182 ( .B1(n18058), .B2(n18156), .C1(n18058), .C2(n18069), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18063) );
  AOI22_X1 U21183 ( .A1(n18145), .A2(n18061), .B1(n18060), .B2(n18059), .ZN(
        n18062) );
  OAI221_X1 U21184 ( .B1(n9633), .B2(n18063), .C1(n18229), .C2(n18805), .A(
        n18062), .ZN(P3_U2846) );
  NOR2_X1 U21185 ( .A1(n18065), .A2(n18064), .ZN(n18071) );
  OR2_X1 U21186 ( .A1(n18067), .A2(n18066), .ZN(n18085) );
  OAI21_X1 U21187 ( .B1(n18086), .B2(n18085), .A(n18072), .ZN(n18068) );
  AOI22_X1 U21188 ( .A1(n18071), .A2(n18070), .B1(n18069), .B2(n18068), .ZN(
        n18079) );
  INV_X1 U21189 ( .A(n18237), .ZN(n18228) );
  OAI22_X1 U21190 ( .A1(n18072), .A2(n18228), .B1(n18229), .B2(n18804), .ZN(
        n18073) );
  AOI21_X1 U21191 ( .B1(n18145), .B2(n18074), .A(n18073), .ZN(n18078) );
  OAI211_X1 U21192 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18076), .A(
        n18246), .B(n18075), .ZN(n18077) );
  OAI211_X1 U21193 ( .C1(n18079), .C2(n18235), .A(n18078), .B(n18077), .ZN(
        P3_U2847) );
  NOR2_X1 U21194 ( .A1(n18229), .A2(n18803), .ZN(n18088) );
  OAI22_X1 U21195 ( .A1(n18243), .A2(n18080), .B1(n18106), .B2(n18731), .ZN(
        n18083) );
  INV_X1 U21196 ( .A(n18106), .ZN(n18081) );
  INV_X1 U21197 ( .A(n18141), .ZN(n18119) );
  OAI21_X1 U21198 ( .B1(n18081), .B2(n18119), .A(n18723), .ZN(n18100) );
  OAI211_X1 U21199 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18236), .A(
        n18121), .B(n18100), .ZN(n18082) );
  NOR3_X1 U21200 ( .A1(n18086), .A2(n18083), .A3(n18082), .ZN(n18084) );
  AOI211_X1 U21201 ( .C1(n18086), .C2(n18085), .A(n18084), .B(n18235), .ZN(
        n18087) );
  AOI211_X1 U21202 ( .C1(n18237), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18088), .B(n18087), .ZN(n18093) );
  INV_X1 U21203 ( .A(n18089), .ZN(n18091) );
  AOI22_X1 U21204 ( .A1(n18163), .A2(n18091), .B1(n18246), .B2(n18090), .ZN(
        n18092) );
  OAI211_X1 U21205 ( .C1(n18094), .C2(n18168), .A(n18093), .B(n18092), .ZN(
        P3_U2848) );
  AOI22_X1 U21206 ( .A1(n9633), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18145), 
        .B2(n18095), .ZN(n18103) );
  INV_X1 U21207 ( .A(n18096), .ZN(n18124) );
  AOI22_X1 U21208 ( .A1(n15702), .A2(n18098), .B1(n18116), .B2(n18097), .ZN(
        n18099) );
  OAI211_X1 U21209 ( .C1(n18129), .C2(n18124), .A(n18121), .B(n18099), .ZN(
        n18107) );
  OAI211_X1 U21210 ( .C1(n18129), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18242), .B(n18100), .ZN(n18101) );
  OAI211_X1 U21211 ( .C1(n18107), .C2(n18101), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18229), .ZN(n18102) );
  OAI211_X1 U21212 ( .C1(n18104), .C2(n18149), .A(n18103), .B(n18102), .ZN(
        P3_U2849) );
  AOI21_X1 U21213 ( .B1(n18124), .B2(n18105), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18113) );
  AOI22_X1 U21214 ( .A1(n17934), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18106), .B2(n18141), .ZN(n18108) );
  OAI21_X1 U21215 ( .B1(n18108), .B2(n18107), .A(n18242), .ZN(n18112) );
  AOI22_X1 U21216 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18237), .B1(
        n18145), .B2(n18109), .ZN(n18111) );
  OAI211_X1 U21217 ( .C1(n18113), .C2(n18112), .A(n18111), .B(n18110), .ZN(
        P3_U2850) );
  AOI22_X1 U21218 ( .A1(n9633), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18145), 
        .B2(n18114), .ZN(n18127) );
  AOI22_X1 U21219 ( .A1(n15702), .A2(n18117), .B1(n18116), .B2(n18115), .ZN(
        n18118) );
  NAND2_X1 U21220 ( .A1(n18242), .A2(n18118), .ZN(n18143) );
  AOI221_X1 U21221 ( .B1(n18148), .B2(n18723), .C1(n18119), .C2(n18723), .A(
        n18143), .ZN(n18120) );
  OAI211_X1 U21222 ( .C1(n18123), .C2(n18122), .A(n18121), .B(n18120), .ZN(
        n18131) );
  OAI22_X1 U21223 ( .A1(n18129), .A2(n18124), .B1(n17934), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18125) );
  OAI211_X1 U21224 ( .C1(n18131), .C2(n18125), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18229), .ZN(n18126) );
  OAI211_X1 U21225 ( .C1(n18149), .C2(n18128), .A(n18127), .B(n18126), .ZN(
        P3_U2851) );
  INV_X1 U21226 ( .A(n18129), .ZN(n18130) );
  OAI221_X1 U21227 ( .B1(n18131), .B2(n18130), .C1(n18131), .C2(n18148), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18136) );
  INV_X1 U21228 ( .A(n18149), .ZN(n18133) );
  NOR2_X1 U21229 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18148), .ZN(
        n18132) );
  AOI22_X1 U21230 ( .A1(n18145), .A2(n18134), .B1(n18133), .B2(n18132), .ZN(
        n18135) );
  OAI221_X1 U21231 ( .B1(n9633), .B2(n18136), .C1(n18229), .C2(n18794), .A(
        n18135), .ZN(P3_U2852) );
  NAND2_X1 U21232 ( .A1(n18712), .A2(n18137), .ZN(n18140) );
  NAND2_X1 U21233 ( .A1(n18691), .A2(n18138), .ZN(n18139) );
  OAI211_X1 U21234 ( .C1(n18141), .C2(n17934), .A(n18140), .B(n18139), .ZN(
        n18142) );
  OAI21_X1 U21235 ( .B1(n18143), .B2(n18142), .A(n18229), .ZN(n18147) );
  AOI22_X1 U21236 ( .A1(n9633), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18145), .B2(
        n18144), .ZN(n18146) );
  OAI221_X1 U21237 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18149), .C1(
        n18148), .C2(n18147), .A(n18146), .ZN(P3_U2853) );
  NAND2_X1 U21238 ( .A1(n18242), .A2(n18169), .ZN(n18184) );
  NOR3_X1 U21239 ( .A1(n18155), .A2(n18154), .A3(n18184), .ZN(n18161) );
  INV_X1 U21240 ( .A(n18150), .ZN(n18151) );
  AOI21_X1 U21241 ( .B1(n18211), .B2(n18151), .A(n18212), .ZN(n18152) );
  OAI21_X1 U21242 ( .B1(n18153), .B2(n18731), .A(n18152), .ZN(n18178) );
  AOI211_X1 U21243 ( .C1(n18156), .C2(n18155), .A(n18154), .B(n18178), .ZN(
        n18177) );
  OAI21_X1 U21244 ( .B1(n18177), .B2(n18230), .A(n18228), .ZN(n18159) );
  INV_X1 U21245 ( .A(n18157), .ZN(n18158) );
  AOI221_X1 U21246 ( .B1(n18161), .B2(n18160), .C1(n18159), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18158), .ZN(n18166) );
  AOI22_X1 U21247 ( .A1(n18164), .A2(n18163), .B1(n18246), .B2(n18162), .ZN(
        n18165) );
  OAI211_X1 U21248 ( .C1(n18168), .C2(n18167), .A(n18166), .B(n18165), .ZN(
        P3_U2854) );
  OAI221_X1 U21249 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18169), .A(n18242), .ZN(
        n18176) );
  AOI21_X1 U21250 ( .B1(n18237), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18170), .ZN(n18175) );
  NAND2_X1 U21251 ( .A1(n18171), .A2(n18242), .ZN(n18250) );
  AOI22_X1 U21252 ( .A1(n18246), .A2(n18173), .B1(n18233), .B2(n18172), .ZN(
        n18174) );
  OAI211_X1 U21253 ( .C1(n18177), .C2(n18176), .A(n18175), .B(n18174), .ZN(
        P3_U2855) );
  INV_X1 U21254 ( .A(n18178), .ZN(n18179) );
  OAI21_X1 U21255 ( .B1(n18179), .B2(n18235), .A(n18228), .ZN(n18185) );
  AOI22_X1 U21256 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18185), .B1(
        n9633), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18183) );
  AOI22_X1 U21257 ( .A1(n18246), .A2(n18181), .B1(n18233), .B2(n18180), .ZN(
        n18182) );
  OAI211_X1 U21258 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18184), .A(
        n18183), .B(n18182), .ZN(P3_U2856) );
  AOI22_X1 U21259 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18185), .B1(
        n9633), .B2(P3_REIP_REG_5__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U21260 ( .A1(n18246), .A2(n18187), .B1(n18233), .B2(n18186), .ZN(
        n18190) );
  NOR3_X1 U21261 ( .A1(n18188), .A2(n18235), .A3(n18192), .ZN(n18198) );
  NAND3_X1 U21262 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18198), .A3(
        n9867), .ZN(n18189) );
  NAND3_X1 U21263 ( .A1(n18191), .A2(n18190), .A3(n18189), .ZN(P3_U2857) );
  AOI211_X1 U21264 ( .C1(n18691), .C2(n18216), .A(n18212), .B(n18192), .ZN(
        n18193) );
  OAI21_X1 U21265 ( .B1(n18195), .B2(n18194), .A(n18193), .ZN(n18206) );
  AOI21_X1 U21266 ( .B1(n18196), .B2(n18206), .A(n18237), .ZN(n18203) );
  AOI22_X1 U21267 ( .A1(n9633), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18233), .B2(
        n18197), .ZN(n18201) );
  AOI22_X1 U21268 ( .A1(n18199), .A2(n18246), .B1(n18198), .B2(n18202), .ZN(
        n18200) );
  OAI211_X1 U21269 ( .C1(n18203), .C2(n18202), .A(n18201), .B(n18200), .ZN(
        P3_U2858) );
  AOI22_X1 U21270 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18237), .B1(
        n9633), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U21271 ( .A1(n18246), .A2(n18205), .B1(n18233), .B2(n18204), .ZN(
        n18209) );
  OAI211_X1 U21272 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18207), .A(
        n18242), .B(n18206), .ZN(n18208) );
  NAND3_X1 U21273 ( .A1(n18210), .A2(n18209), .A3(n18208), .ZN(P3_U2859) );
  NAND2_X1 U21274 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18214) );
  OAI21_X1 U21275 ( .B1(n18212), .B2(n18861), .A(n18211), .ZN(n18213) );
  OAI21_X1 U21276 ( .B1(n18214), .B2(n18731), .A(n18213), .ZN(n18215) );
  AOI22_X1 U21277 ( .A1(n18691), .A2(n18216), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18215), .ZN(n18219) );
  NAND3_X1 U21278 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18217), .A3(
        n18227), .ZN(n18218) );
  OAI211_X1 U21279 ( .C1(n18221), .C2(n18220), .A(n18219), .B(n18218), .ZN(
        n18223) );
  AOI22_X1 U21280 ( .A1(n18242), .A2(n18223), .B1(n18233), .B2(n18222), .ZN(
        n18226) );
  INV_X1 U21281 ( .A(n18224), .ZN(n18225) );
  OAI211_X1 U21282 ( .C1(n18228), .C2(n18227), .A(n18226), .B(n18225), .ZN(
        P3_U2860) );
  NOR2_X1 U21283 ( .A1(n18229), .A2(n18881), .ZN(n18232) );
  AOI211_X1 U21284 ( .C1(n18243), .C2(n18876), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18230), .ZN(n18231) );
  AOI211_X1 U21285 ( .C1(n18234), .C2(n18233), .A(n18232), .B(n18231), .ZN(
        n18239) );
  NOR3_X1 U21286 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18236), .A3(
        n18235), .ZN(n18245) );
  OAI21_X1 U21287 ( .B1(n18237), .B2(n18245), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18238) );
  OAI211_X1 U21288 ( .C1(n18241), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        P3_U2861) );
  AOI211_X1 U21289 ( .C1(n18243), .C2(n18242), .A(n9633), .B(n18876), .ZN(
        n18244) );
  AOI211_X1 U21290 ( .C1(n18246), .C2(n18249), .A(n18245), .B(n18244), .ZN(
        n18248) );
  NAND2_X1 U21291 ( .A1(n9633), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18247) );
  OAI211_X1 U21292 ( .C1(n18250), .C2(n18249), .A(n18248), .B(n18247), .ZN(
        P3_U2862) );
  AOI21_X1 U21293 ( .B1(n18253), .B2(n18252), .A(n18251), .ZN(n18747) );
  INV_X1 U21294 ( .A(n18430), .ZN(n18300) );
  OAI21_X1 U21295 ( .B1(n18747), .B2(n18300), .A(n18259), .ZN(n18254) );
  OAI221_X1 U21296 ( .B1(n18713), .B2(n18901), .C1(n18713), .C2(n18259), .A(
        n18254), .ZN(P3_U2863) );
  INV_X1 U21297 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18734) );
  NOR2_X1 U21298 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18734), .ZN(
        n18476) );
  NOR2_X1 U21299 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18255), .ZN(
        n18432) );
  NOR2_X1 U21300 ( .A1(n18476), .A2(n18432), .ZN(n18257) );
  OAI22_X1 U21301 ( .A1(n18258), .A2(n18734), .B1(n18257), .B2(n18256), .ZN(
        P3_U2866) );
  NOR2_X1 U21302 ( .A1(n21095), .A2(n18259), .ZN(P3_U2867) );
  NOR2_X1 U21303 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18717) );
  NOR2_X1 U21304 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18340) );
  NAND2_X1 U21305 ( .A1(n18717), .A2(n18340), .ZN(n18361) );
  NOR2_X1 U21306 ( .A1(n18261), .A2(n18260), .ZN(n18272) );
  NAND2_X1 U21307 ( .A1(n18272), .A2(n18262), .ZN(n18640) );
  NAND2_X1 U21308 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18571) );
  INV_X1 U21309 ( .A(n18571), .ZN(n18573) );
  NOR2_X1 U21310 ( .A1(n18713), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18475) );
  NAND2_X1 U21311 ( .A1(n18573), .A2(n18475), .ZN(n18667) );
  INV_X1 U21312 ( .A(n18667), .ZN(n18683) );
  AND2_X1 U21313 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18636), .ZN(n18632) );
  NOR2_X2 U21314 ( .A1(n18362), .A2(n18263), .ZN(n18631) );
  NOR2_X1 U21315 ( .A1(n18734), .A2(n18407), .ZN(n18634) );
  INV_X1 U21316 ( .A(n18634), .ZN(n18630) );
  NOR2_X2 U21317 ( .A1(n18713), .A2(n18630), .ZN(n18685) );
  INV_X1 U21318 ( .A(n18361), .ZN(n18351) );
  NOR2_X1 U21319 ( .A1(n18685), .A2(n18351), .ZN(n18320) );
  NOR2_X1 U21320 ( .A1(n18752), .A2(n18320), .ZN(n18294) );
  AOI22_X1 U21321 ( .A1(n18683), .A2(n18632), .B1(n18631), .B2(n18294), .ZN(
        n18267) );
  NAND2_X1 U21322 ( .A1(n18634), .A2(n18713), .ZN(n18610) );
  NAND2_X1 U21323 ( .A1(n18667), .A2(n18610), .ZN(n18605) );
  AOI21_X1 U21324 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18362), .ZN(n18602) );
  INV_X1 U21325 ( .A(n18320), .ZN(n18264) );
  AOI22_X1 U21326 ( .A1(n18636), .A2(n18605), .B1(n18602), .B2(n18264), .ZN(
        n18297) );
  INV_X1 U21327 ( .A(n18610), .ZN(n18625) );
  NOR2_X2 U21328 ( .A1(n18363), .A2(n18265), .ZN(n18637) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18297), .B1(
        n18625), .B2(n18637), .ZN(n18266) );
  OAI211_X1 U21330 ( .C1(n18361), .C2(n18640), .A(n18267), .B(n18266), .ZN(
        P3_U2868) );
  NAND2_X1 U21331 ( .A1(n18272), .A2(n18268), .ZN(n18646) );
  AND2_X1 U21332 ( .A1(n18636), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18642) );
  NOR2_X2 U21333 ( .A1(n18362), .A2(n21108), .ZN(n18641) );
  AOI22_X1 U21334 ( .A1(n18625), .A2(n18642), .B1(n18294), .B2(n18641), .ZN(
        n18270) );
  NOR2_X2 U21335 ( .A1(n15079), .A2(n18363), .ZN(n18643) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18297), .B1(
        n18683), .B2(n18643), .ZN(n18269) );
  OAI211_X1 U21337 ( .C1(n18361), .C2(n18646), .A(n18270), .B(n18269), .ZN(
        P3_U2869) );
  NAND2_X1 U21338 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18636), .ZN(n18653) );
  NOR2_X2 U21339 ( .A1(n18363), .A2(n19354), .ZN(n18649) );
  NOR2_X2 U21340 ( .A1(n18362), .A2(n18271), .ZN(n18648) );
  AOI22_X1 U21341 ( .A1(n18625), .A2(n18649), .B1(n18294), .B2(n18648), .ZN(
        n18275) );
  NOR2_X1 U21342 ( .A1(n18273), .A2(n18295), .ZN(n18650) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18297), .B1(
        n18351), .B2(n18650), .ZN(n18274) );
  OAI211_X1 U21344 ( .C1(n18667), .C2(n18653), .A(n18275), .B(n18274), .ZN(
        P3_U2870) );
  NAND2_X1 U21345 ( .A1(n18636), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18659) );
  NAND2_X1 U21346 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18636), .ZN(n18584) );
  INV_X1 U21347 ( .A(n18584), .ZN(n18655) );
  NOR2_X2 U21348 ( .A1(n18362), .A2(n18276), .ZN(n18654) );
  AOI22_X1 U21349 ( .A1(n18683), .A2(n18655), .B1(n18294), .B2(n18654), .ZN(
        n18279) );
  NOR2_X2 U21350 ( .A1(n18277), .A2(n18295), .ZN(n18656) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18297), .B1(
        n18351), .B2(n18656), .ZN(n18278) );
  OAI211_X1 U21352 ( .C1(n18610), .C2(n18659), .A(n18279), .B(n18278), .ZN(
        P3_U2871) );
  NAND2_X1 U21353 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18636), .ZN(n18666) );
  NAND2_X1 U21354 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18636), .ZN(n18588) );
  INV_X1 U21355 ( .A(n18588), .ZN(n18662) );
  NOR2_X2 U21356 ( .A1(n18280), .A2(n18362), .ZN(n18660) );
  AOI22_X1 U21357 ( .A1(n18683), .A2(n18662), .B1(n18294), .B2(n18660), .ZN(
        n18283) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18297), .B1(
        n18351), .B2(n9625), .ZN(n18282) );
  OAI211_X1 U21359 ( .C1(n18610), .C2(n18666), .A(n18283), .B(n18282), .ZN(
        P3_U2872) );
  NAND2_X1 U21360 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18636), .ZN(n18673) );
  NAND2_X1 U21361 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18636), .ZN(n18593) );
  INV_X1 U21362 ( .A(n18593), .ZN(n18669) );
  NOR2_X2 U21363 ( .A1(n18284), .A2(n18362), .ZN(n18668) );
  AOI22_X1 U21364 ( .A1(n18625), .A2(n18669), .B1(n18294), .B2(n18668), .ZN(
        n18287) );
  NOR2_X2 U21365 ( .A1(n18285), .A2(n18295), .ZN(n18670) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18297), .B1(
        n18351), .B2(n18670), .ZN(n18286) );
  OAI211_X1 U21367 ( .C1(n18667), .C2(n18673), .A(n18287), .B(n18286), .ZN(
        P3_U2873) );
  NAND2_X1 U21368 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18636), .ZN(n18679) );
  NAND2_X1 U21369 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18636), .ZN(n18623) );
  INV_X1 U21370 ( .A(n18623), .ZN(n18675) );
  NOR2_X2 U21371 ( .A1(n18288), .A2(n18362), .ZN(n18674) );
  AOI22_X1 U21372 ( .A1(n18625), .A2(n18675), .B1(n18294), .B2(n18674), .ZN(
        n18291) );
  NOR2_X2 U21373 ( .A1(n18289), .A2(n18295), .ZN(n18676) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18297), .B1(
        n18351), .B2(n18676), .ZN(n18290) );
  OAI211_X1 U21375 ( .C1(n18667), .C2(n18679), .A(n18291), .B(n18290), .ZN(
        P3_U2874) );
  NAND2_X1 U21376 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18636), .ZN(n18690) );
  NOR2_X2 U21377 ( .A1(n18292), .A2(n18363), .ZN(n18682) );
  NOR2_X2 U21378 ( .A1(n18293), .A2(n18362), .ZN(n18681) );
  AOI22_X1 U21379 ( .A1(n18625), .A2(n18682), .B1(n18294), .B2(n18681), .ZN(
        n18299) );
  NOR2_X2 U21380 ( .A1(n18296), .A2(n18295), .ZN(n18684) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18297), .B1(
        n18351), .B2(n18684), .ZN(n18298) );
  OAI211_X1 U21382 ( .C1(n18667), .C2(n18690), .A(n18299), .B(n18298), .ZN(
        P3_U2875) );
  NAND2_X1 U21383 ( .A1(n18475), .A2(n18340), .ZN(n18354) );
  INV_X1 U21384 ( .A(n18340), .ZN(n18319) );
  NAND2_X1 U21385 ( .A1(n18714), .A2(n18600), .ZN(n18570) );
  NOR2_X1 U21386 ( .A1(n18319), .A2(n18570), .ZN(n18315) );
  AOI22_X1 U21387 ( .A1(n18685), .A2(n18637), .B1(n18631), .B2(n18315), .ZN(
        n18302) );
  NOR2_X1 U21388 ( .A1(n18362), .A2(n18300), .ZN(n18633) );
  AND2_X1 U21389 ( .A1(n18714), .A2(n18633), .ZN(n18572) );
  AOI22_X1 U21390 ( .A1(n18636), .A2(n18634), .B1(n18340), .B2(n18572), .ZN(
        n18316) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18316), .B1(
        n18625), .B2(n18632), .ZN(n18301) );
  OAI211_X1 U21392 ( .C1(n18640), .C2(n18354), .A(n18302), .B(n18301), .ZN(
        P3_U2876) );
  AOI22_X1 U21393 ( .A1(n18685), .A2(n18642), .B1(n18641), .B2(n18315), .ZN(
        n18304) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18316), .B1(
        n18625), .B2(n18643), .ZN(n18303) );
  OAI211_X1 U21395 ( .C1(n18646), .C2(n18354), .A(n18304), .B(n18303), .ZN(
        P3_U2877) );
  INV_X1 U21396 ( .A(n18650), .ZN(n18555) );
  INV_X1 U21397 ( .A(n18653), .ZN(n18552) );
  AOI22_X1 U21398 ( .A1(n18625), .A2(n18552), .B1(n18648), .B2(n18315), .ZN(
        n18306) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18316), .B1(
        n18685), .B2(n18649), .ZN(n18305) );
  OAI211_X1 U21400 ( .C1(n18555), .C2(n18354), .A(n18306), .B(n18305), .ZN(
        P3_U2878) );
  INV_X1 U21401 ( .A(n18685), .ZN(n18647) );
  AOI22_X1 U21402 ( .A1(n18625), .A2(n18655), .B1(n18654), .B2(n18315), .ZN(
        n18308) );
  INV_X1 U21403 ( .A(n18354), .ZN(n18381) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18316), .B1(
        n18656), .B2(n18381), .ZN(n18307) );
  OAI211_X1 U21405 ( .C1(n18647), .C2(n18659), .A(n18308), .B(n18307), .ZN(
        P3_U2879) );
  AOI22_X1 U21406 ( .A1(n18625), .A2(n18662), .B1(n18660), .B2(n18315), .ZN(
        n18310) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18316), .B1(
        n9625), .B2(n18381), .ZN(n18309) );
  OAI211_X1 U21408 ( .C1(n18647), .C2(n18666), .A(n18310), .B(n18309), .ZN(
        P3_U2880) );
  INV_X1 U21409 ( .A(n18673), .ZN(n18590) );
  AOI22_X1 U21410 ( .A1(n18625), .A2(n18590), .B1(n18668), .B2(n18315), .ZN(
        n18312) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18316), .B1(
        n18670), .B2(n18381), .ZN(n18311) );
  OAI211_X1 U21412 ( .C1(n18647), .C2(n18593), .A(n18312), .B(n18311), .ZN(
        P3_U2881) );
  INV_X1 U21413 ( .A(n18679), .ZN(n18620) );
  AOI22_X1 U21414 ( .A1(n18625), .A2(n18620), .B1(n18674), .B2(n18315), .ZN(
        n18314) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18316), .B1(
        n18676), .B2(n18381), .ZN(n18313) );
  OAI211_X1 U21416 ( .C1(n18647), .C2(n18623), .A(n18314), .B(n18313), .ZN(
        P3_U2882) );
  AOI22_X1 U21417 ( .A1(n18685), .A2(n18682), .B1(n18681), .B2(n18315), .ZN(
        n18318) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18316), .B1(
        n18684), .B2(n18381), .ZN(n18317) );
  OAI211_X1 U21419 ( .C1(n18610), .C2(n18690), .A(n18318), .B(n18317), .ZN(
        P3_U2883) );
  NOR2_X1 U21420 ( .A1(n18714), .A2(n18319), .ZN(n18386) );
  NAND2_X1 U21421 ( .A1(n18386), .A2(n18713), .ZN(n18406) );
  NOR2_X1 U21422 ( .A1(n18381), .A2(n18399), .ZN(n18364) );
  NOR2_X1 U21423 ( .A1(n18752), .A2(n18364), .ZN(n18336) );
  AOI22_X1 U21424 ( .A1(n18351), .A2(n18637), .B1(n18631), .B2(n18336), .ZN(
        n18323) );
  INV_X1 U21425 ( .A(n18604), .ZN(n18544) );
  OAI21_X1 U21426 ( .B1(n18320), .B2(n18544), .A(n18364), .ZN(n18321) );
  OAI211_X1 U21427 ( .C1(n18399), .C2(n18850), .A(n18547), .B(n18321), .ZN(
        n18337) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18337), .B1(
        n18685), .B2(n18632), .ZN(n18322) );
  OAI211_X1 U21429 ( .C1(n18640), .C2(n18406), .A(n18323), .B(n18322), .ZN(
        P3_U2884) );
  AOI22_X1 U21430 ( .A1(n18351), .A2(n18642), .B1(n18641), .B2(n18336), .ZN(
        n18325) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18337), .B1(
        n18685), .B2(n18643), .ZN(n18324) );
  OAI211_X1 U21432 ( .C1(n18646), .C2(n18406), .A(n18325), .B(n18324), .ZN(
        P3_U2885) );
  AOI22_X1 U21433 ( .A1(n18351), .A2(n18649), .B1(n18648), .B2(n18336), .ZN(
        n18327) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18337), .B1(
        n18650), .B2(n18399), .ZN(n18326) );
  OAI211_X1 U21435 ( .C1(n18647), .C2(n18653), .A(n18327), .B(n18326), .ZN(
        P3_U2886) );
  AOI22_X1 U21436 ( .A1(n18685), .A2(n18655), .B1(n18654), .B2(n18336), .ZN(
        n18329) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18337), .B1(
        n18656), .B2(n18399), .ZN(n18328) );
  OAI211_X1 U21438 ( .C1(n18361), .C2(n18659), .A(n18329), .B(n18328), .ZN(
        P3_U2887) );
  INV_X1 U21439 ( .A(n18666), .ZN(n18585) );
  AOI22_X1 U21440 ( .A1(n18351), .A2(n18585), .B1(n18660), .B2(n18336), .ZN(
        n18331) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18337), .B1(
        n9625), .B2(n18399), .ZN(n18330) );
  OAI211_X1 U21442 ( .C1(n18647), .C2(n18588), .A(n18331), .B(n18330), .ZN(
        P3_U2888) );
  AOI22_X1 U21443 ( .A1(n18685), .A2(n18590), .B1(n18668), .B2(n18336), .ZN(
        n18333) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18337), .B1(
        n18670), .B2(n18399), .ZN(n18332) );
  OAI211_X1 U21445 ( .C1(n18361), .C2(n18593), .A(n18333), .B(n18332), .ZN(
        P3_U2889) );
  AOI22_X1 U21446 ( .A1(n18685), .A2(n18620), .B1(n18674), .B2(n18336), .ZN(
        n18335) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18337), .B1(
        n18676), .B2(n18399), .ZN(n18334) );
  OAI211_X1 U21448 ( .C1(n18361), .C2(n18623), .A(n18335), .B(n18334), .ZN(
        P3_U2890) );
  AOI22_X1 U21449 ( .A1(n18351), .A2(n18682), .B1(n18681), .B2(n18336), .ZN(
        n18339) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18337), .B1(
        n18684), .B2(n18399), .ZN(n18338) );
  OAI211_X1 U21451 ( .C1(n18647), .C2(n18690), .A(n18339), .B(n18338), .ZN(
        P3_U2891) );
  NAND2_X1 U21452 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18386), .ZN(
        n18429) );
  AND2_X1 U21453 ( .A1(n18600), .A2(n18386), .ZN(n18357) );
  AOI22_X1 U21454 ( .A1(n18637), .A2(n18381), .B1(n18631), .B2(n18357), .ZN(
        n18342) );
  AOI21_X1 U21455 ( .B1(n18714), .B2(n18544), .A(n18362), .ZN(n18431) );
  OAI211_X1 U21456 ( .C1(n18422), .C2(n18850), .A(n18340), .B(n18431), .ZN(
        n18358) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18358), .B1(
        n18351), .B2(n18632), .ZN(n18341) );
  OAI211_X1 U21458 ( .C1(n18640), .C2(n18429), .A(n18342), .B(n18341), .ZN(
        P3_U2892) );
  AOI22_X1 U21459 ( .A1(n18642), .A2(n18381), .B1(n18641), .B2(n18357), .ZN(
        n18344) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18358), .B1(
        n18351), .B2(n18643), .ZN(n18343) );
  OAI211_X1 U21461 ( .C1(n18646), .C2(n18429), .A(n18344), .B(n18343), .ZN(
        P3_U2893) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18358), .B1(
        n18648), .B2(n18357), .ZN(n18346) );
  AOI22_X1 U21463 ( .A1(n18650), .A2(n18422), .B1(n18649), .B2(n18381), .ZN(
        n18345) );
  OAI211_X1 U21464 ( .C1(n18361), .C2(n18653), .A(n18346), .B(n18345), .ZN(
        P3_U2894) );
  INV_X1 U21465 ( .A(n18659), .ZN(n18581) );
  AOI22_X1 U21466 ( .A1(n18581), .A2(n18381), .B1(n18654), .B2(n18357), .ZN(
        n18348) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18358), .B1(
        n18656), .B2(n18422), .ZN(n18347) );
  OAI211_X1 U21468 ( .C1(n18361), .C2(n18584), .A(n18348), .B(n18347), .ZN(
        P3_U2895) );
  AOI22_X1 U21469 ( .A1(n18585), .A2(n18381), .B1(n18660), .B2(n18357), .ZN(
        n18350) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18358), .B1(
        n9625), .B2(n18422), .ZN(n18349) );
  OAI211_X1 U21471 ( .C1(n18361), .C2(n18588), .A(n18350), .B(n18349), .ZN(
        P3_U2896) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18358), .B1(
        n18668), .B2(n18357), .ZN(n18353) );
  AOI22_X1 U21473 ( .A1(n18351), .A2(n18590), .B1(n18670), .B2(n18422), .ZN(
        n18352) );
  OAI211_X1 U21474 ( .C1(n18593), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        P3_U2897) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18358), .B1(
        n18674), .B2(n18357), .ZN(n18356) );
  AOI22_X1 U21476 ( .A1(n18676), .A2(n18422), .B1(n18675), .B2(n18381), .ZN(
        n18355) );
  OAI211_X1 U21477 ( .C1(n18361), .C2(n18679), .A(n18356), .B(n18355), .ZN(
        P3_U2898) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18358), .B1(
        n18681), .B2(n18357), .ZN(n18360) );
  AOI22_X1 U21479 ( .A1(n18684), .A2(n18422), .B1(n18682), .B2(n18381), .ZN(
        n18359) );
  OAI211_X1 U21480 ( .C1(n18361), .C2(n18690), .A(n18360), .B(n18359), .ZN(
        P3_U2899) );
  NAND2_X1 U21481 ( .A1(n18717), .A2(n18432), .ZN(n18447) );
  INV_X1 U21482 ( .A(n18447), .ZN(n18449) );
  NOR2_X1 U21483 ( .A1(n18422), .A2(n18449), .ZN(n18408) );
  NOR2_X1 U21484 ( .A1(n18752), .A2(n18408), .ZN(n18380) );
  AOI22_X1 U21485 ( .A1(n18632), .A2(n18381), .B1(n18631), .B2(n18380), .ZN(
        n18367) );
  OAI22_X1 U21486 ( .A1(n18364), .A2(n18363), .B1(n18408), .B2(n18362), .ZN(
        n18365) );
  OAI21_X1 U21487 ( .B1(n18449), .B2(n18850), .A(n18365), .ZN(n18382) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18382), .B1(
        n18637), .B2(n18399), .ZN(n18366) );
  OAI211_X1 U21489 ( .C1(n18640), .C2(n18447), .A(n18367), .B(n18366), .ZN(
        P3_U2900) );
  AOI22_X1 U21490 ( .A1(n18643), .A2(n18381), .B1(n18641), .B2(n18380), .ZN(
        n18369) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18382), .B1(
        n18642), .B2(n18399), .ZN(n18368) );
  OAI211_X1 U21492 ( .C1(n18646), .C2(n18447), .A(n18369), .B(n18368), .ZN(
        P3_U2901) );
  AOI22_X1 U21493 ( .A1(n18552), .A2(n18381), .B1(n18648), .B2(n18380), .ZN(
        n18371) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18382), .B1(
        n18649), .B2(n18399), .ZN(n18370) );
  OAI211_X1 U21495 ( .C1(n18555), .C2(n18447), .A(n18371), .B(n18370), .ZN(
        P3_U2902) );
  AOI22_X1 U21496 ( .A1(n18655), .A2(n18381), .B1(n18654), .B2(n18380), .ZN(
        n18373) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18382), .B1(
        n18656), .B2(n18449), .ZN(n18372) );
  OAI211_X1 U21498 ( .C1(n18659), .C2(n18406), .A(n18373), .B(n18372), .ZN(
        P3_U2903) );
  AOI22_X1 U21499 ( .A1(n18662), .A2(n18381), .B1(n18660), .B2(n18380), .ZN(
        n18375) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18382), .B1(
        n9625), .B2(n18449), .ZN(n18374) );
  OAI211_X1 U21501 ( .C1(n18666), .C2(n18406), .A(n18375), .B(n18374), .ZN(
        P3_U2904) );
  AOI22_X1 U21502 ( .A1(n18590), .A2(n18381), .B1(n18668), .B2(n18380), .ZN(
        n18377) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18382), .B1(
        n18670), .B2(n18449), .ZN(n18376) );
  OAI211_X1 U21504 ( .C1(n18593), .C2(n18406), .A(n18377), .B(n18376), .ZN(
        P3_U2905) );
  AOI22_X1 U21505 ( .A1(n18620), .A2(n18381), .B1(n18674), .B2(n18380), .ZN(
        n18379) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18382), .B1(
        n18676), .B2(n18449), .ZN(n18378) );
  OAI211_X1 U21507 ( .C1(n18623), .C2(n18406), .A(n18379), .B(n18378), .ZN(
        P3_U2906) );
  INV_X1 U21508 ( .A(n18682), .ZN(n18543) );
  INV_X1 U21509 ( .A(n18690), .ZN(n18539) );
  AOI22_X1 U21510 ( .A1(n18539), .A2(n18381), .B1(n18681), .B2(n18380), .ZN(
        n18384) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18382), .B1(
        n18684), .B2(n18449), .ZN(n18383) );
  OAI211_X1 U21512 ( .C1(n18543), .C2(n18406), .A(n18384), .B(n18383), .ZN(
        P3_U2907) );
  NAND2_X1 U21513 ( .A1(n18432), .A2(n18475), .ZN(n18474) );
  INV_X1 U21514 ( .A(n18432), .ZN(n18385) );
  NOR2_X1 U21515 ( .A1(n18385), .A2(n18570), .ZN(n18402) );
  AOI22_X1 U21516 ( .A1(n18632), .A2(n18399), .B1(n18631), .B2(n18402), .ZN(
        n18388) );
  AOI22_X1 U21517 ( .A1(n18636), .A2(n18386), .B1(n18432), .B2(n18572), .ZN(
        n18403) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18403), .B1(
        n18637), .B2(n18422), .ZN(n18387) );
  OAI211_X1 U21519 ( .C1(n18640), .C2(n18474), .A(n18388), .B(n18387), .ZN(
        P3_U2908) );
  AOI22_X1 U21520 ( .A1(n18642), .A2(n18422), .B1(n18641), .B2(n18402), .ZN(
        n18390) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18403), .B1(
        n18643), .B2(n18399), .ZN(n18389) );
  OAI211_X1 U21522 ( .C1(n18646), .C2(n18474), .A(n18390), .B(n18389), .ZN(
        P3_U2909) );
  AOI22_X1 U21523 ( .A1(n18648), .A2(n18402), .B1(n18649), .B2(n18422), .ZN(
        n18392) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18403), .B1(
        n18552), .B2(n18399), .ZN(n18391) );
  OAI211_X1 U21525 ( .C1(n18555), .C2(n18474), .A(n18392), .B(n18391), .ZN(
        P3_U2910) );
  AOI22_X1 U21526 ( .A1(n18655), .A2(n18399), .B1(n18654), .B2(n18402), .ZN(
        n18394) );
  INV_X1 U21527 ( .A(n18474), .ZN(n18465) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18403), .B1(
        n18656), .B2(n18465), .ZN(n18393) );
  OAI211_X1 U21529 ( .C1(n18659), .C2(n18429), .A(n18394), .B(n18393), .ZN(
        P3_U2911) );
  AOI22_X1 U21530 ( .A1(n18585), .A2(n18422), .B1(n18660), .B2(n18402), .ZN(
        n18396) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18403), .B1(
        n9625), .B2(n18465), .ZN(n18395) );
  OAI211_X1 U21532 ( .C1(n18588), .C2(n18406), .A(n18396), .B(n18395), .ZN(
        P3_U2912) );
  AOI22_X1 U21533 ( .A1(n18590), .A2(n18399), .B1(n18668), .B2(n18402), .ZN(
        n18398) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18403), .B1(
        n18670), .B2(n18465), .ZN(n18397) );
  OAI211_X1 U21535 ( .C1(n18593), .C2(n18429), .A(n18398), .B(n18397), .ZN(
        P3_U2913) );
  AOI22_X1 U21536 ( .A1(n18620), .A2(n18399), .B1(n18674), .B2(n18402), .ZN(
        n18401) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18403), .B1(
        n18676), .B2(n18465), .ZN(n18400) );
  OAI211_X1 U21538 ( .C1(n18623), .C2(n18429), .A(n18401), .B(n18400), .ZN(
        P3_U2914) );
  AOI22_X1 U21539 ( .A1(n18682), .A2(n18422), .B1(n18681), .B2(n18402), .ZN(
        n18405) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18403), .B1(
        n18684), .B2(n18465), .ZN(n18404) );
  OAI211_X1 U21541 ( .C1(n18690), .C2(n18406), .A(n18405), .B(n18404), .ZN(
        P3_U2915) );
  NOR2_X1 U21542 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18407), .ZN(
        n18477) );
  NAND2_X1 U21543 ( .A1(n18477), .A2(n18713), .ZN(n18497) );
  NAND2_X1 U21544 ( .A1(n18474), .A2(n18497), .ZN(n18453) );
  AND2_X1 U21545 ( .A1(n18600), .A2(n18453), .ZN(n18425) );
  AOI22_X1 U21546 ( .A1(n18637), .A2(n18449), .B1(n18631), .B2(n18425), .ZN(
        n18411) );
  INV_X1 U21547 ( .A(n18408), .ZN(n18409) );
  OAI221_X1 U21548 ( .B1(n18453), .B2(n18604), .C1(n18453), .C2(n18409), .A(
        n18602), .ZN(n18426) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18426), .B1(
        n18632), .B2(n18422), .ZN(n18410) );
  OAI211_X1 U21550 ( .C1(n18640), .C2(n18497), .A(n18411), .B(n18410), .ZN(
        P3_U2916) );
  AOI22_X1 U21551 ( .A1(n18643), .A2(n18422), .B1(n18641), .B2(n18425), .ZN(
        n18413) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18426), .B1(
        n18642), .B2(n18449), .ZN(n18412) );
  OAI211_X1 U21553 ( .C1(n18646), .C2(n18497), .A(n18413), .B(n18412), .ZN(
        P3_U2917) );
  AOI22_X1 U21554 ( .A1(n18552), .A2(n18422), .B1(n18648), .B2(n18425), .ZN(
        n18415) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18426), .B1(
        n18649), .B2(n18449), .ZN(n18414) );
  OAI211_X1 U21556 ( .C1(n18555), .C2(n18497), .A(n18415), .B(n18414), .ZN(
        P3_U2918) );
  AOI22_X1 U21557 ( .A1(n18581), .A2(n18449), .B1(n18654), .B2(n18425), .ZN(
        n18417) );
  INV_X1 U21558 ( .A(n18497), .ZN(n18486) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18426), .B1(
        n18656), .B2(n18486), .ZN(n18416) );
  OAI211_X1 U21560 ( .C1(n18584), .C2(n18429), .A(n18417), .B(n18416), .ZN(
        P3_U2919) );
  AOI22_X1 U21561 ( .A1(n18662), .A2(n18422), .B1(n18660), .B2(n18425), .ZN(
        n18419) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18426), .B1(
        n9625), .B2(n18486), .ZN(n18418) );
  OAI211_X1 U21563 ( .C1(n18666), .C2(n18447), .A(n18419), .B(n18418), .ZN(
        P3_U2920) );
  AOI22_X1 U21564 ( .A1(n18668), .A2(n18425), .B1(n18669), .B2(n18449), .ZN(
        n18421) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18426), .B1(
        n18670), .B2(n18486), .ZN(n18420) );
  OAI211_X1 U21566 ( .C1(n18673), .C2(n18429), .A(n18421), .B(n18420), .ZN(
        P3_U2921) );
  AOI22_X1 U21567 ( .A1(n18620), .A2(n18422), .B1(n18674), .B2(n18425), .ZN(
        n18424) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18426), .B1(
        n18676), .B2(n18486), .ZN(n18423) );
  OAI211_X1 U21569 ( .C1(n18623), .C2(n18447), .A(n18424), .B(n18423), .ZN(
        P3_U2922) );
  AOI22_X1 U21570 ( .A1(n18682), .A2(n18449), .B1(n18681), .B2(n18425), .ZN(
        n18428) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18426), .B1(
        n18684), .B2(n18486), .ZN(n18427) );
  OAI211_X1 U21572 ( .C1(n18690), .C2(n18429), .A(n18428), .B(n18427), .ZN(
        P3_U2923) );
  NAND2_X1 U21573 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18477), .ZN(
        n18520) );
  AND2_X1 U21574 ( .A1(n18600), .A2(n18477), .ZN(n18448) );
  AOI22_X1 U21575 ( .A1(n18637), .A2(n18465), .B1(n18631), .B2(n18448), .ZN(
        n18434) );
  NAND3_X1 U21576 ( .A1(n18432), .A2(n18431), .A3(n18430), .ZN(n18450) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18450), .B1(
        n18632), .B2(n18449), .ZN(n18433) );
  OAI211_X1 U21578 ( .C1(n18640), .C2(n18520), .A(n18434), .B(n18433), .ZN(
        P3_U2924) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18450), .B1(
        n18641), .B2(n18448), .ZN(n18436) );
  AOI22_X1 U21580 ( .A1(n18643), .A2(n18449), .B1(n18642), .B2(n18465), .ZN(
        n18435) );
  OAI211_X1 U21581 ( .C1(n18646), .C2(n18520), .A(n18436), .B(n18435), .ZN(
        P3_U2925) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18450), .B1(
        n18648), .B2(n18448), .ZN(n18438) );
  AOI22_X1 U21583 ( .A1(n18552), .A2(n18449), .B1(n18649), .B2(n18465), .ZN(
        n18437) );
  OAI211_X1 U21584 ( .C1(n18555), .C2(n18520), .A(n18438), .B(n18437), .ZN(
        P3_U2926) );
  AOI22_X1 U21585 ( .A1(n18581), .A2(n18465), .B1(n18654), .B2(n18448), .ZN(
        n18440) );
  INV_X1 U21586 ( .A(n18520), .ZN(n18513) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18450), .B1(
        n18656), .B2(n18513), .ZN(n18439) );
  OAI211_X1 U21588 ( .C1(n18584), .C2(n18447), .A(n18440), .B(n18439), .ZN(
        P3_U2927) );
  AOI22_X1 U21589 ( .A1(n18585), .A2(n18465), .B1(n18660), .B2(n18448), .ZN(
        n18442) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18450), .B1(
        n9625), .B2(n18513), .ZN(n18441) );
  OAI211_X1 U21591 ( .C1(n18588), .C2(n18447), .A(n18442), .B(n18441), .ZN(
        P3_U2928) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18450), .B1(
        n18668), .B2(n18448), .ZN(n18444) );
  AOI22_X1 U21593 ( .A1(n18590), .A2(n18449), .B1(n18670), .B2(n18513), .ZN(
        n18443) );
  OAI211_X1 U21594 ( .C1(n18593), .C2(n18474), .A(n18444), .B(n18443), .ZN(
        P3_U2929) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18450), .B1(
        n18674), .B2(n18448), .ZN(n18446) );
  AOI22_X1 U21596 ( .A1(n18676), .A2(n18513), .B1(n18675), .B2(n18465), .ZN(
        n18445) );
  OAI211_X1 U21597 ( .C1(n18679), .C2(n18447), .A(n18446), .B(n18445), .ZN(
        P3_U2930) );
  AOI22_X1 U21598 ( .A1(n18539), .A2(n18449), .B1(n18681), .B2(n18448), .ZN(
        n18452) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18450), .B1(
        n18684), .B2(n18513), .ZN(n18451) );
  OAI211_X1 U21600 ( .C1(n18543), .C2(n18474), .A(n18452), .B(n18451), .ZN(
        P3_U2931) );
  NAND2_X1 U21601 ( .A1(n18717), .A2(n18476), .ZN(n18532) );
  INV_X1 U21602 ( .A(n18532), .ZN(n18538) );
  NOR2_X1 U21603 ( .A1(n18513), .A2(n18538), .ZN(n18499) );
  NOR2_X1 U21604 ( .A1(n18752), .A2(n18499), .ZN(n18470) );
  AOI22_X1 U21605 ( .A1(n18632), .A2(n18465), .B1(n18631), .B2(n18470), .ZN(
        n18456) );
  INV_X1 U21606 ( .A(n18499), .ZN(n18454) );
  OAI221_X1 U21607 ( .B1(n18454), .B2(n18604), .C1(n18454), .C2(n18453), .A(
        n18602), .ZN(n18471) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18471), .B1(
        n18637), .B2(n18486), .ZN(n18455) );
  OAI211_X1 U21609 ( .C1(n18640), .C2(n18532), .A(n18456), .B(n18455), .ZN(
        P3_U2932) );
  AOI22_X1 U21610 ( .A1(n18643), .A2(n18465), .B1(n18641), .B2(n18470), .ZN(
        n18458) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18471), .B1(
        n18642), .B2(n18486), .ZN(n18457) );
  OAI211_X1 U21612 ( .C1(n18646), .C2(n18532), .A(n18458), .B(n18457), .ZN(
        P3_U2933) );
  AOI22_X1 U21613 ( .A1(n18648), .A2(n18470), .B1(n18649), .B2(n18486), .ZN(
        n18460) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18471), .B1(
        n18650), .B2(n18538), .ZN(n18459) );
  OAI211_X1 U21615 ( .C1(n18653), .C2(n18474), .A(n18460), .B(n18459), .ZN(
        P3_U2934) );
  AOI22_X1 U21616 ( .A1(n18655), .A2(n18465), .B1(n18654), .B2(n18470), .ZN(
        n18462) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18471), .B1(
        n18656), .B2(n18538), .ZN(n18461) );
  OAI211_X1 U21618 ( .C1(n18659), .C2(n18497), .A(n18462), .B(n18461), .ZN(
        P3_U2935) );
  AOI22_X1 U21619 ( .A1(n18662), .A2(n18465), .B1(n18660), .B2(n18470), .ZN(
        n18464) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18471), .B1(
        n9625), .B2(n18538), .ZN(n18463) );
  OAI211_X1 U21621 ( .C1(n18666), .C2(n18497), .A(n18464), .B(n18463), .ZN(
        P3_U2936) );
  AOI22_X1 U21622 ( .A1(n18590), .A2(n18465), .B1(n18668), .B2(n18470), .ZN(
        n18467) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18471), .B1(
        n18670), .B2(n18538), .ZN(n18466) );
  OAI211_X1 U21624 ( .C1(n18593), .C2(n18497), .A(n18467), .B(n18466), .ZN(
        P3_U2937) );
  AOI22_X1 U21625 ( .A1(n18675), .A2(n18486), .B1(n18674), .B2(n18470), .ZN(
        n18469) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18471), .B1(
        n18676), .B2(n18538), .ZN(n18468) );
  OAI211_X1 U21627 ( .C1(n18679), .C2(n18474), .A(n18469), .B(n18468), .ZN(
        P3_U2938) );
  AOI22_X1 U21628 ( .A1(n18682), .A2(n18486), .B1(n18681), .B2(n18470), .ZN(
        n18473) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18471), .B1(
        n18684), .B2(n18538), .ZN(n18472) );
  OAI211_X1 U21630 ( .C1(n18690), .C2(n18474), .A(n18473), .B(n18472), .ZN(
        P3_U2939) );
  NAND2_X1 U21631 ( .A1(n18476), .A2(n18475), .ZN(n18569) );
  INV_X1 U21632 ( .A(n18476), .ZN(n18498) );
  NOR2_X1 U21633 ( .A1(n18498), .A2(n18570), .ZN(n18493) );
  AOI22_X1 U21634 ( .A1(n18637), .A2(n18513), .B1(n18631), .B2(n18493), .ZN(
        n18479) );
  NOR2_X1 U21635 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18498), .ZN(
        n18521) );
  AOI22_X1 U21636 ( .A1(n18636), .A2(n18477), .B1(n18633), .B2(n18521), .ZN(
        n18494) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18494), .B1(
        n18632), .B2(n18486), .ZN(n18478) );
  OAI211_X1 U21638 ( .C1(n18640), .C2(n18569), .A(n18479), .B(n18478), .ZN(
        P3_U2940) );
  AOI22_X1 U21639 ( .A1(n18642), .A2(n18513), .B1(n18641), .B2(n18493), .ZN(
        n18481) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18494), .B1(
        n18643), .B2(n18486), .ZN(n18480) );
  OAI211_X1 U21641 ( .C1(n18646), .C2(n18569), .A(n18481), .B(n18480), .ZN(
        P3_U2941) );
  AOI22_X1 U21642 ( .A1(n18648), .A2(n18493), .B1(n18649), .B2(n18513), .ZN(
        n18483) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18494), .B1(
        n18552), .B2(n18486), .ZN(n18482) );
  OAI211_X1 U21644 ( .C1(n18555), .C2(n18569), .A(n18483), .B(n18482), .ZN(
        P3_U2942) );
  AOI22_X1 U21645 ( .A1(n18581), .A2(n18513), .B1(n18654), .B2(n18493), .ZN(
        n18485) );
  INV_X1 U21646 ( .A(n18569), .ZN(n18562) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18494), .B1(
        n18656), .B2(n18562), .ZN(n18484) );
  OAI211_X1 U21648 ( .C1(n18584), .C2(n18497), .A(n18485), .B(n18484), .ZN(
        P3_U2943) );
  AOI22_X1 U21649 ( .A1(n18662), .A2(n18486), .B1(n18660), .B2(n18493), .ZN(
        n18488) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18494), .B1(
        n9625), .B2(n18562), .ZN(n18487) );
  OAI211_X1 U21651 ( .C1(n18666), .C2(n18520), .A(n18488), .B(n18487), .ZN(
        P3_U2944) );
  AOI22_X1 U21652 ( .A1(n18668), .A2(n18493), .B1(n18669), .B2(n18513), .ZN(
        n18490) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18494), .B1(
        n18670), .B2(n18562), .ZN(n18489) );
  OAI211_X1 U21654 ( .C1(n18673), .C2(n18497), .A(n18490), .B(n18489), .ZN(
        P3_U2945) );
  AOI22_X1 U21655 ( .A1(n18675), .A2(n18513), .B1(n18674), .B2(n18493), .ZN(
        n18492) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18494), .B1(
        n18676), .B2(n18562), .ZN(n18491) );
  OAI211_X1 U21657 ( .C1(n18679), .C2(n18497), .A(n18492), .B(n18491), .ZN(
        P3_U2946) );
  AOI22_X1 U21658 ( .A1(n18682), .A2(n18513), .B1(n18681), .B2(n18493), .ZN(
        n18496) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18494), .B1(
        n18684), .B2(n18562), .ZN(n18495) );
  OAI211_X1 U21660 ( .C1(n18690), .C2(n18497), .A(n18496), .B(n18495), .ZN(
        P3_U2947) );
  NOR2_X1 U21661 ( .A1(n18714), .A2(n18498), .ZN(n18574) );
  NAND2_X1 U21662 ( .A1(n18574), .A2(n18713), .ZN(n18599) );
  NOR2_X1 U21663 ( .A1(n18562), .A2(n18589), .ZN(n18545) );
  NOR2_X1 U21664 ( .A1(n18752), .A2(n18545), .ZN(n18516) );
  AOI22_X1 U21665 ( .A1(n18632), .A2(n18513), .B1(n18631), .B2(n18516), .ZN(
        n18502) );
  OAI21_X1 U21666 ( .B1(n18499), .B2(n18544), .A(n18545), .ZN(n18500) );
  OAI211_X1 U21667 ( .C1(n18589), .C2(n18850), .A(n18547), .B(n18500), .ZN(
        n18517) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18517), .B1(
        n18637), .B2(n18538), .ZN(n18501) );
  OAI211_X1 U21669 ( .C1(n18640), .C2(n18599), .A(n18502), .B(n18501), .ZN(
        P3_U2948) );
  AOI22_X1 U21670 ( .A1(n18642), .A2(n18538), .B1(n18641), .B2(n18516), .ZN(
        n18504) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18517), .B1(
        n18643), .B2(n18513), .ZN(n18503) );
  OAI211_X1 U21672 ( .C1(n18646), .C2(n18599), .A(n18504), .B(n18503), .ZN(
        P3_U2949) );
  AOI22_X1 U21673 ( .A1(n18648), .A2(n18516), .B1(n18649), .B2(n18538), .ZN(
        n18506) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18517), .B1(
        n18650), .B2(n18589), .ZN(n18505) );
  OAI211_X1 U21675 ( .C1(n18653), .C2(n18520), .A(n18506), .B(n18505), .ZN(
        P3_U2950) );
  AOI22_X1 U21676 ( .A1(n18581), .A2(n18538), .B1(n18654), .B2(n18516), .ZN(
        n18508) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18517), .B1(
        n18656), .B2(n18589), .ZN(n18507) );
  OAI211_X1 U21678 ( .C1(n18584), .C2(n18520), .A(n18508), .B(n18507), .ZN(
        P3_U2951) );
  AOI22_X1 U21679 ( .A1(n18585), .A2(n18538), .B1(n18660), .B2(n18516), .ZN(
        n18510) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18517), .B1(
        n9625), .B2(n18589), .ZN(n18509) );
  OAI211_X1 U21681 ( .C1(n18588), .C2(n18520), .A(n18510), .B(n18509), .ZN(
        P3_U2952) );
  AOI22_X1 U21682 ( .A1(n18590), .A2(n18513), .B1(n18668), .B2(n18516), .ZN(
        n18512) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18517), .B1(
        n18670), .B2(n18589), .ZN(n18511) );
  OAI211_X1 U21684 ( .C1(n18593), .C2(n18532), .A(n18512), .B(n18511), .ZN(
        P3_U2953) );
  AOI22_X1 U21685 ( .A1(n18620), .A2(n18513), .B1(n18674), .B2(n18516), .ZN(
        n18515) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18517), .B1(
        n18676), .B2(n18589), .ZN(n18514) );
  OAI211_X1 U21687 ( .C1(n18623), .C2(n18532), .A(n18515), .B(n18514), .ZN(
        P3_U2954) );
  AOI22_X1 U21688 ( .A1(n18682), .A2(n18538), .B1(n18681), .B2(n18516), .ZN(
        n18519) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18517), .B1(
        n18684), .B2(n18589), .ZN(n18518) );
  OAI211_X1 U21690 ( .C1(n18690), .C2(n18520), .A(n18519), .B(n18518), .ZN(
        P3_U2955) );
  NAND2_X1 U21691 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18574), .ZN(
        n18629) );
  AND2_X1 U21692 ( .A1(n18600), .A2(n18574), .ZN(n18537) );
  AOI22_X1 U21693 ( .A1(n18632), .A2(n18538), .B1(n18631), .B2(n18537), .ZN(
        n18523) );
  AOI22_X1 U21694 ( .A1(n18636), .A2(n18521), .B1(n18633), .B2(n18574), .ZN(
        n18540) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18540), .B1(
        n18637), .B2(n18562), .ZN(n18522) );
  OAI211_X1 U21696 ( .C1(n18640), .C2(n18629), .A(n18523), .B(n18522), .ZN(
        P3_U2956) );
  AOI22_X1 U21697 ( .A1(n18643), .A2(n18538), .B1(n18641), .B2(n18537), .ZN(
        n18525) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18540), .B1(
        n18642), .B2(n18562), .ZN(n18524) );
  OAI211_X1 U21699 ( .C1(n18646), .C2(n18629), .A(n18525), .B(n18524), .ZN(
        P3_U2957) );
  AOI22_X1 U21700 ( .A1(n18648), .A2(n18537), .B1(n18649), .B2(n18562), .ZN(
        n18527) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18540), .B1(
        n18552), .B2(n18538), .ZN(n18526) );
  OAI211_X1 U21702 ( .C1(n18555), .C2(n18629), .A(n18527), .B(n18526), .ZN(
        P3_U2958) );
  AOI22_X1 U21703 ( .A1(n18655), .A2(n18538), .B1(n18654), .B2(n18537), .ZN(
        n18529) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18540), .B1(
        n18656), .B2(n18619), .ZN(n18528) );
  OAI211_X1 U21705 ( .C1(n18659), .C2(n18569), .A(n18529), .B(n18528), .ZN(
        P3_U2959) );
  AOI22_X1 U21706 ( .A1(n18585), .A2(n18562), .B1(n18660), .B2(n18537), .ZN(
        n18531) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18540), .B1(
        n9625), .B2(n18619), .ZN(n18530) );
  OAI211_X1 U21708 ( .C1(n18588), .C2(n18532), .A(n18531), .B(n18530), .ZN(
        P3_U2960) );
  AOI22_X1 U21709 ( .A1(n18590), .A2(n18538), .B1(n18668), .B2(n18537), .ZN(
        n18534) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18540), .B1(
        n18670), .B2(n18619), .ZN(n18533) );
  OAI211_X1 U21711 ( .C1(n18593), .C2(n18569), .A(n18534), .B(n18533), .ZN(
        P3_U2961) );
  AOI22_X1 U21712 ( .A1(n18620), .A2(n18538), .B1(n18674), .B2(n18537), .ZN(
        n18536) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18540), .B1(
        n18676), .B2(n18619), .ZN(n18535) );
  OAI211_X1 U21714 ( .C1(n18623), .C2(n18569), .A(n18536), .B(n18535), .ZN(
        P3_U2962) );
  AOI22_X1 U21715 ( .A1(n18539), .A2(n18538), .B1(n18681), .B2(n18537), .ZN(
        n18542) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18540), .B1(
        n18684), .B2(n18619), .ZN(n18541) );
  OAI211_X1 U21717 ( .C1(n18543), .C2(n18569), .A(n18542), .B(n18541), .ZN(
        P3_U2963) );
  NAND2_X1 U21718 ( .A1(n18717), .A2(n18573), .ZN(n18689) );
  INV_X1 U21719 ( .A(n18689), .ZN(n18661) );
  NOR2_X1 U21720 ( .A1(n18619), .A2(n18661), .ZN(n18601) );
  NOR2_X1 U21721 ( .A1(n18752), .A2(n18601), .ZN(n18565) );
  AOI22_X1 U21722 ( .A1(n18637), .A2(n18589), .B1(n18631), .B2(n18565), .ZN(
        n18549) );
  OAI21_X1 U21723 ( .B1(n18545), .B2(n18544), .A(n18601), .ZN(n18546) );
  OAI211_X1 U21724 ( .C1(n18661), .C2(n18850), .A(n18547), .B(n18546), .ZN(
        n18566) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18566), .B1(
        n18632), .B2(n18562), .ZN(n18548) );
  OAI211_X1 U21726 ( .C1(n18640), .C2(n18689), .A(n18549), .B(n18548), .ZN(
        P3_U2964) );
  AOI22_X1 U21727 ( .A1(n18643), .A2(n18562), .B1(n18641), .B2(n18565), .ZN(
        n18551) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18566), .B1(
        n18642), .B2(n18589), .ZN(n18550) );
  OAI211_X1 U21729 ( .C1(n18646), .C2(n18689), .A(n18551), .B(n18550), .ZN(
        P3_U2965) );
  AOI22_X1 U21730 ( .A1(n18552), .A2(n18562), .B1(n18648), .B2(n18565), .ZN(
        n18554) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18566), .B1(
        n18649), .B2(n18589), .ZN(n18553) );
  OAI211_X1 U21732 ( .C1(n18555), .C2(n18689), .A(n18554), .B(n18553), .ZN(
        P3_U2966) );
  AOI22_X1 U21733 ( .A1(n18655), .A2(n18562), .B1(n18654), .B2(n18565), .ZN(
        n18557) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18566), .B1(
        n18656), .B2(n18661), .ZN(n18556) );
  OAI211_X1 U21735 ( .C1(n18659), .C2(n18599), .A(n18557), .B(n18556), .ZN(
        P3_U2967) );
  AOI22_X1 U21736 ( .A1(n18662), .A2(n18562), .B1(n18660), .B2(n18565), .ZN(
        n18559) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18566), .B1(
        n9625), .B2(n18661), .ZN(n18558) );
  OAI211_X1 U21738 ( .C1(n18666), .C2(n18599), .A(n18559), .B(n18558), .ZN(
        P3_U2968) );
  AOI22_X1 U21739 ( .A1(n18590), .A2(n18562), .B1(n18668), .B2(n18565), .ZN(
        n18561) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18566), .B1(
        n18670), .B2(n18661), .ZN(n18560) );
  OAI211_X1 U21741 ( .C1(n18593), .C2(n18599), .A(n18561), .B(n18560), .ZN(
        P3_U2969) );
  AOI22_X1 U21742 ( .A1(n18620), .A2(n18562), .B1(n18674), .B2(n18565), .ZN(
        n18564) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18566), .B1(
        n18676), .B2(n18661), .ZN(n18563) );
  OAI211_X1 U21744 ( .C1(n18623), .C2(n18599), .A(n18564), .B(n18563), .ZN(
        P3_U2970) );
  AOI22_X1 U21745 ( .A1(n18682), .A2(n18589), .B1(n18681), .B2(n18565), .ZN(
        n18568) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18566), .B1(
        n18684), .B2(n18661), .ZN(n18567) );
  OAI211_X1 U21747 ( .C1(n18690), .C2(n18569), .A(n18568), .B(n18567), .ZN(
        P3_U2971) );
  NOR2_X1 U21748 ( .A1(n18571), .A2(n18570), .ZN(n18635) );
  AOI22_X1 U21749 ( .A1(n18637), .A2(n18619), .B1(n18631), .B2(n18635), .ZN(
        n18576) );
  AOI22_X1 U21750 ( .A1(n18636), .A2(n18574), .B1(n18573), .B2(n18572), .ZN(
        n18596) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18596), .B1(
        n18632), .B2(n18589), .ZN(n18575) );
  OAI211_X1 U21752 ( .C1(n18667), .C2(n18640), .A(n18576), .B(n18575), .ZN(
        P3_U2972) );
  AOI22_X1 U21753 ( .A1(n18643), .A2(n18589), .B1(n18641), .B2(n18635), .ZN(
        n18578) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18596), .B1(
        n18642), .B2(n18619), .ZN(n18577) );
  OAI211_X1 U21755 ( .C1(n18667), .C2(n18646), .A(n18578), .B(n18577), .ZN(
        P3_U2973) );
  AOI22_X1 U21756 ( .A1(n18648), .A2(n18635), .B1(n18649), .B2(n18619), .ZN(
        n18580) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18596), .B1(
        n18683), .B2(n18650), .ZN(n18579) );
  OAI211_X1 U21758 ( .C1(n18653), .C2(n18599), .A(n18580), .B(n18579), .ZN(
        P3_U2974) );
  AOI22_X1 U21759 ( .A1(n18581), .A2(n18619), .B1(n18654), .B2(n18635), .ZN(
        n18583) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18596), .B1(
        n18683), .B2(n18656), .ZN(n18582) );
  OAI211_X1 U21761 ( .C1(n18584), .C2(n18599), .A(n18583), .B(n18582), .ZN(
        P3_U2975) );
  AOI22_X1 U21762 ( .A1(n18585), .A2(n18619), .B1(n18660), .B2(n18635), .ZN(
        n18587) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18596), .B1(
        n18683), .B2(n9625), .ZN(n18586) );
  OAI211_X1 U21764 ( .C1(n18588), .C2(n18599), .A(n18587), .B(n18586), .ZN(
        P3_U2976) );
  AOI22_X1 U21765 ( .A1(n18590), .A2(n18589), .B1(n18668), .B2(n18635), .ZN(
        n18592) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18596), .B1(
        n18683), .B2(n18670), .ZN(n18591) );
  OAI211_X1 U21767 ( .C1(n18593), .C2(n18629), .A(n18592), .B(n18591), .ZN(
        P3_U2977) );
  AOI22_X1 U21768 ( .A1(n18675), .A2(n18619), .B1(n18674), .B2(n18635), .ZN(
        n18595) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18596), .B1(
        n18683), .B2(n18676), .ZN(n18594) );
  OAI211_X1 U21770 ( .C1(n18679), .C2(n18599), .A(n18595), .B(n18594), .ZN(
        P3_U2978) );
  AOI22_X1 U21771 ( .A1(n18682), .A2(n18619), .B1(n18681), .B2(n18635), .ZN(
        n18598) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18596), .B1(
        n18683), .B2(n18684), .ZN(n18597) );
  OAI211_X1 U21773 ( .C1(n18690), .C2(n18599), .A(n18598), .B(n18597), .ZN(
        P3_U2979) );
  AND2_X1 U21774 ( .A1(n18600), .A2(n18605), .ZN(n18624) );
  AOI22_X1 U21775 ( .A1(n18632), .A2(n18619), .B1(n18631), .B2(n18624), .ZN(
        n18607) );
  INV_X1 U21776 ( .A(n18601), .ZN(n18603) );
  OAI221_X1 U21777 ( .B1(n18605), .B2(n18604), .C1(n18605), .C2(n18603), .A(
        n18602), .ZN(n18626) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18626), .B1(
        n18637), .B2(n18661), .ZN(n18606) );
  OAI211_X1 U21779 ( .C1(n18610), .C2(n18640), .A(n18607), .B(n18606), .ZN(
        P3_U2980) );
  AOI22_X1 U21780 ( .A1(n18643), .A2(n18619), .B1(n18641), .B2(n18624), .ZN(
        n18609) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18626), .B1(
        n18642), .B2(n18661), .ZN(n18608) );
  OAI211_X1 U21782 ( .C1(n18610), .C2(n18646), .A(n18609), .B(n18608), .ZN(
        P3_U2981) );
  AOI22_X1 U21783 ( .A1(n18648), .A2(n18624), .B1(n18649), .B2(n18661), .ZN(
        n18612) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18650), .ZN(n18611) );
  OAI211_X1 U21785 ( .C1(n18653), .C2(n18629), .A(n18612), .B(n18611), .ZN(
        P3_U2982) );
  AOI22_X1 U21786 ( .A1(n18655), .A2(n18619), .B1(n18654), .B2(n18624), .ZN(
        n18614) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18656), .ZN(n18613) );
  OAI211_X1 U21788 ( .C1(n18659), .C2(n18689), .A(n18614), .B(n18613), .ZN(
        P3_U2983) );
  AOI22_X1 U21789 ( .A1(n18662), .A2(n18619), .B1(n18660), .B2(n18624), .ZN(
        n18616) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n9625), .ZN(n18615) );
  OAI211_X1 U21791 ( .C1(n18666), .C2(n18689), .A(n18616), .B(n18615), .ZN(
        P3_U2984) );
  AOI22_X1 U21792 ( .A1(n18668), .A2(n18624), .B1(n18669), .B2(n18661), .ZN(
        n18618) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18670), .ZN(n18617) );
  OAI211_X1 U21794 ( .C1(n18673), .C2(n18629), .A(n18618), .B(n18617), .ZN(
        P3_U2985) );
  AOI22_X1 U21795 ( .A1(n18620), .A2(n18619), .B1(n18674), .B2(n18624), .ZN(
        n18622) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18676), .ZN(n18621) );
  OAI211_X1 U21797 ( .C1(n18623), .C2(n18689), .A(n18622), .B(n18621), .ZN(
        P3_U2986) );
  AOI22_X1 U21798 ( .A1(n18682), .A2(n18661), .B1(n18681), .B2(n18624), .ZN(
        n18628) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n18684), .ZN(n18627) );
  OAI211_X1 U21800 ( .C1(n18690), .C2(n18629), .A(n18628), .B(n18627), .ZN(
        P3_U2987) );
  NOR2_X1 U21801 ( .A1(n18752), .A2(n18630), .ZN(n18680) );
  AOI22_X1 U21802 ( .A1(n18632), .A2(n18661), .B1(n18631), .B2(n18680), .ZN(
        n18639) );
  AOI22_X1 U21803 ( .A1(n18636), .A2(n18635), .B1(n18634), .B2(n18633), .ZN(
        n18686) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18686), .B1(
        n18683), .B2(n18637), .ZN(n18638) );
  OAI211_X1 U21805 ( .C1(n18647), .C2(n18640), .A(n18639), .B(n18638), .ZN(
        P3_U2988) );
  AOI22_X1 U21806 ( .A1(n18683), .A2(n18642), .B1(n18641), .B2(n18680), .ZN(
        n18645) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18686), .B1(
        n18643), .B2(n18661), .ZN(n18644) );
  OAI211_X1 U21808 ( .C1(n18647), .C2(n18646), .A(n18645), .B(n18644), .ZN(
        P3_U2989) );
  AOI22_X1 U21809 ( .A1(n18683), .A2(n18649), .B1(n18648), .B2(n18680), .ZN(
        n18652) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18650), .ZN(n18651) );
  OAI211_X1 U21811 ( .C1(n18653), .C2(n18689), .A(n18652), .B(n18651), .ZN(
        P3_U2990) );
  AOI22_X1 U21812 ( .A1(n18655), .A2(n18661), .B1(n18654), .B2(n18680), .ZN(
        n18658) );
  AOI22_X1 U21813 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18656), .ZN(n18657) );
  OAI211_X1 U21814 ( .C1(n18667), .C2(n18659), .A(n18658), .B(n18657), .ZN(
        P3_U2991) );
  AOI22_X1 U21815 ( .A1(n18662), .A2(n18661), .B1(n18660), .B2(n18680), .ZN(
        n18665) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n9625), .ZN(n18664) );
  OAI211_X1 U21817 ( .C1(n18667), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        P3_U2992) );
  AOI22_X1 U21818 ( .A1(n18683), .A2(n18669), .B1(n18668), .B2(n18680), .ZN(
        n18672) );
  AOI22_X1 U21819 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18670), .ZN(n18671) );
  OAI211_X1 U21820 ( .C1(n18673), .C2(n18689), .A(n18672), .B(n18671), .ZN(
        P3_U2993) );
  AOI22_X1 U21821 ( .A1(n18683), .A2(n18675), .B1(n18674), .B2(n18680), .ZN(
        n18678) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18676), .ZN(n18677) );
  OAI211_X1 U21823 ( .C1(n18679), .C2(n18689), .A(n18678), .B(n18677), .ZN(
        P3_U2994) );
  AOI22_X1 U21824 ( .A1(n18683), .A2(n18682), .B1(n18681), .B2(n18680), .ZN(
        n18688) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18684), .ZN(n18687) );
  OAI211_X1 U21826 ( .C1(n18690), .C2(n18689), .A(n18688), .B(n18687), .ZN(
        P3_U2995) );
  NOR2_X1 U21827 ( .A1(n18691), .A2(n15702), .ZN(n18693) );
  OAI222_X1 U21828 ( .A1(n18697), .A2(n18696), .B1(n18695), .B2(n18694), .C1(
        n18693), .C2(n18692), .ZN(n18890) );
  AOI21_X1 U21829 ( .B1(n18700), .B2(n18699), .A(n18698), .ZN(n18720) );
  AOI22_X1 U21830 ( .A1(n18865), .A2(n18701), .B1(n18704), .B2(n18712), .ZN(
        n18702) );
  OAI21_X1 U21831 ( .B1(n18703), .B2(n18720), .A(n18702), .ZN(n18855) );
  NOR2_X1 U21832 ( .A1(n18856), .A2(n18855), .ZN(n18707) );
  NOR2_X1 U21833 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18719), .ZN(
        n18705) );
  NOR2_X1 U21834 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18712), .ZN(
        n18709) );
  OAI22_X1 U21835 ( .A1(n18705), .A2(n18731), .B1(n18709), .B2(n18704), .ZN(
        n18852) );
  AOI21_X1 U21836 ( .B1(n18852), .B2(n18732), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18706) );
  AOI21_X1 U21837 ( .B1(n18732), .B2(n18707), .A(n18706), .ZN(n18736) );
  NAND2_X1 U21838 ( .A1(n17934), .A2(n18708), .ZN(n18711) );
  INV_X1 U21839 ( .A(n18709), .ZN(n18710) );
  AOI22_X1 U21840 ( .A1(n18870), .A2(n18711), .B1(n18873), .B2(n18710), .ZN(
        n18866) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18712), .B1(
        n18711), .B2(n18879), .ZN(n18715) );
  INV_X1 U21842 ( .A(n18715), .ZN(n18875) );
  NOR3_X1 U21843 ( .A1(n18714), .A2(n18713), .A3(n18875), .ZN(n18716) );
  OAI22_X1 U21844 ( .A1(n18866), .A2(n18716), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18715), .ZN(n18718) );
  NOR2_X1 U21845 ( .A1(n18719), .A2(n18865), .ZN(n18729) );
  OAI21_X1 U21846 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18725), .A(
        n18720), .ZN(n18728) );
  AOI211_X1 U21847 ( .C1(n18865), .C2(n18873), .A(n18722), .B(n18721), .ZN(
        n18727) );
  AOI211_X1 U21848 ( .C1(n18725), .C2(n18724), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18873), .ZN(n18726) );
  AOI211_X1 U21849 ( .C1(n18729), .C2(n18728), .A(n18727), .B(n18726), .ZN(
        n18730) );
  OAI21_X1 U21850 ( .B1(n18862), .B2(n18731), .A(n18730), .ZN(n18863) );
  AOI22_X1 U21851 ( .A1(n18742), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18863), .B2(n18732), .ZN(n18733) );
  OAI21_X1 U21852 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18733), .ZN(n18735) );
  OAI21_X1 U21853 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18737), .ZN(n18738) );
  AOI211_X1 U21854 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18742), .A(
        n18890), .B(n18741), .ZN(n18751) );
  INV_X1 U21855 ( .A(n18897), .ZN(n18743) );
  AOI22_X1 U21856 ( .A1(n18874), .A2(n18743), .B1(n18895), .B2(n18905), .ZN(
        n18744) );
  INV_X1 U21857 ( .A(n18744), .ZN(n18748) );
  OAI211_X1 U21858 ( .C1(n18746), .C2(n18745), .A(n18902), .B(n18751), .ZN(
        n18849) );
  NAND2_X1 U21859 ( .A1(n18895), .A2(n18905), .ZN(n18756) );
  NAND4_X1 U21860 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18895), .A4(n18910), .ZN(n18758) );
  OR3_X1 U21861 ( .A1(n18754), .A2(n18753), .A3(n18752), .ZN(n18755) );
  NAND4_X1 U21862 ( .A1(n18757), .A2(n18756), .A3(n18758), .A4(n18755), .ZN(
        P3_U2997) );
  AND4_X1 U21863 ( .A1(n18897), .A2(n18759), .A3(n18758), .A4(n18848), .ZN(
        P3_U2998) );
  INV_X1 U21864 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21075) );
  NOR2_X1 U21865 ( .A1(n21075), .A2(n18847), .ZN(P3_U2999) );
  AND2_X1 U21866 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18761), .ZN(
        P3_U3000) );
  AND2_X1 U21867 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18761), .ZN(
        P3_U3001) );
  AND2_X1 U21868 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18761), .ZN(
        P3_U3002) );
  AND2_X1 U21869 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18761), .ZN(
        P3_U3003) );
  AND2_X1 U21870 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18761), .ZN(
        P3_U3004) );
  AND2_X1 U21871 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18761), .ZN(
        P3_U3005) );
  AND2_X1 U21872 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18761), .ZN(
        P3_U3006) );
  AND2_X1 U21873 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18761), .ZN(
        P3_U3007) );
  AND2_X1 U21874 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18761), .ZN(
        P3_U3008) );
  AND2_X1 U21875 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18761), .ZN(
        P3_U3009) );
  AND2_X1 U21876 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18761), .ZN(
        P3_U3010) );
  AND2_X1 U21877 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18761), .ZN(
        P3_U3011) );
  AND2_X1 U21878 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18761), .ZN(
        P3_U3012) );
  AND2_X1 U21879 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18761), .ZN(
        P3_U3013) );
  AND2_X1 U21880 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18761), .ZN(
        P3_U3014) );
  AND2_X1 U21881 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18760), .ZN(
        P3_U3015) );
  AND2_X1 U21882 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18760), .ZN(
        P3_U3016) );
  AND2_X1 U21883 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18760), .ZN(
        P3_U3017) );
  INV_X1 U21884 ( .A(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21111) );
  NOR2_X1 U21885 ( .A1(n21111), .A2(n18847), .ZN(P3_U3018) );
  AND2_X1 U21886 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18760), .ZN(
        P3_U3019) );
  AND2_X1 U21887 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18760), .ZN(
        P3_U3020) );
  AND2_X1 U21888 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18760), .ZN(P3_U3021) );
  AND2_X1 U21889 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18760), .ZN(P3_U3022) );
  AND2_X1 U21890 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18760), .ZN(P3_U3023) );
  AND2_X1 U21891 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18760), .ZN(P3_U3024) );
  AND2_X1 U21892 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18760), .ZN(P3_U3025) );
  AND2_X1 U21893 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18761), .ZN(P3_U3026) );
  AND2_X1 U21894 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18761), .ZN(P3_U3027) );
  AND2_X1 U21895 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18761), .ZN(P3_U3028) );
  OAI21_X1 U21896 ( .B1(n19861), .B2(n18762), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18763) );
  INV_X1 U21897 ( .A(n18763), .ZN(n18765) );
  NAND2_X1 U21898 ( .A1(n18895), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18771) );
  AND2_X1 U21899 ( .A1(n18771), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18775) );
  AOI21_X1 U21900 ( .B1(NA), .B2(n18764), .A(n18776), .ZN(n18770) );
  OAI22_X1 U21901 ( .A1(n18843), .A2(n18765), .B1(n18775), .B2(n18770), .ZN(
        P3_U3029) );
  AND3_X1 U21902 ( .A1(n18776), .A2(P3_STATE_REG_1__SCAN_IN), .A3(HOLD), .ZN(
        n18766) );
  AOI221_X1 U21903 ( .B1(n18767), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19861), .C2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n18766), .ZN(n18769)
         );
  OAI211_X1 U21904 ( .C1(n18769), .C2(n18768), .A(n18771), .B(n18891), .ZN(
        P3_U3030) );
  INV_X1 U21905 ( .A(n18770), .ZN(n18774) );
  OAI222_X1 U21906 ( .A1(n18776), .A2(n19861), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n18771), .C2(NA), .ZN(n18772)
         );
  OAI211_X1 U21907 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n18772), .ZN(n18773) );
  OAI21_X1 U21908 ( .B1(n18775), .B2(n18774), .A(n18773), .ZN(P3_U3031) );
  OAI222_X1 U21909 ( .A1(n18881), .A2(n18830), .B1(n18777), .B2(n18843), .C1(
        n18778), .C2(n18826), .ZN(P3_U3032) );
  OAI222_X1 U21910 ( .A1(n18826), .A2(n18780), .B1(n18779), .B2(n18843), .C1(
        n18778), .C2(n18830), .ZN(P3_U3033) );
  INV_X1 U21911 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18782) );
  OAI222_X1 U21912 ( .A1(n18826), .A2(n18782), .B1(n18781), .B2(n18843), .C1(
        n18780), .C2(n18830), .ZN(P3_U3034) );
  OAI222_X1 U21913 ( .A1(n18826), .A2(n18784), .B1(n18783), .B2(n18843), .C1(
        n18782), .C2(n18830), .ZN(P3_U3035) );
  INV_X1 U21914 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18786) );
  OAI222_X1 U21915 ( .A1(n18826), .A2(n18786), .B1(n18785), .B2(n18843), .C1(
        n18784), .C2(n18830), .ZN(P3_U3036) );
  OAI222_X1 U21916 ( .A1(n18826), .A2(n18788), .B1(n18787), .B2(n18843), .C1(
        n18786), .C2(n18830), .ZN(P3_U3037) );
  INV_X1 U21917 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18790) );
  OAI222_X1 U21918 ( .A1(n18826), .A2(n18790), .B1(n18789), .B2(n18843), .C1(
        n18788), .C2(n18830), .ZN(P3_U3038) );
  OAI222_X1 U21919 ( .A1(n18826), .A2(n18792), .B1(n18791), .B2(n18843), .C1(
        n18790), .C2(n18830), .ZN(P3_U3039) );
  OAI222_X1 U21920 ( .A1(n18826), .A2(n18794), .B1(n18793), .B2(n18843), .C1(
        n18792), .C2(n18830), .ZN(P3_U3040) );
  OAI222_X1 U21921 ( .A1(n18826), .A2(n18796), .B1(n18795), .B2(n18843), .C1(
        n18794), .C2(n18830), .ZN(P3_U3041) );
  INV_X1 U21922 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18798) );
  OAI222_X1 U21923 ( .A1(n18826), .A2(n18798), .B1(n18797), .B2(n18843), .C1(
        n18796), .C2(n18830), .ZN(P3_U3042) );
  OAI222_X1 U21924 ( .A1(n18826), .A2(n18800), .B1(n18799), .B2(n18843), .C1(
        n18798), .C2(n18830), .ZN(P3_U3043) );
  OAI222_X1 U21925 ( .A1(n18826), .A2(n18803), .B1(n18801), .B2(n18843), .C1(
        n18800), .C2(n18836), .ZN(P3_U3044) );
  OAI222_X1 U21926 ( .A1(n18803), .A2(n18830), .B1(n18802), .B2(n18843), .C1(
        n18804), .C2(n18826), .ZN(P3_U3045) );
  OAI222_X1 U21927 ( .A1(n18826), .A2(n18805), .B1(n21118), .B2(n18843), .C1(
        n18804), .C2(n18836), .ZN(P3_U3046) );
  OAI222_X1 U21928 ( .A1(n18826), .A2(n18808), .B1(n18806), .B2(n18843), .C1(
        n18805), .C2(n18836), .ZN(P3_U3047) );
  OAI222_X1 U21929 ( .A1(n18808), .A2(n18830), .B1(n18807), .B2(n18843), .C1(
        n18809), .C2(n18826), .ZN(P3_U3048) );
  OAI222_X1 U21930 ( .A1(n18826), .A2(n18811), .B1(n18810), .B2(n18843), .C1(
        n18809), .C2(n18836), .ZN(P3_U3049) );
  OAI222_X1 U21931 ( .A1(n18826), .A2(n18814), .B1(n18812), .B2(n18843), .C1(
        n18811), .C2(n18836), .ZN(P3_U3050) );
  INV_X1 U21932 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20950) );
  OAI222_X1 U21933 ( .A1(n18814), .A2(n18830), .B1(n18813), .B2(n18843), .C1(
        n20950), .C2(n18826), .ZN(P3_U3051) );
  INV_X1 U21934 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18816) );
  OAI222_X1 U21935 ( .A1(n20950), .A2(n18830), .B1(n18815), .B2(n18843), .C1(
        n18816), .C2(n18826), .ZN(P3_U3052) );
  OAI222_X1 U21936 ( .A1(n18826), .A2(n18818), .B1(n18817), .B2(n18843), .C1(
        n18816), .C2(n18836), .ZN(P3_U3053) );
  OAI222_X1 U21937 ( .A1(n18826), .A2(n18820), .B1(n18819), .B2(n18843), .C1(
        n18818), .C2(n18830), .ZN(P3_U3054) );
  OAI222_X1 U21938 ( .A1(n18826), .A2(n18822), .B1(n18821), .B2(n18843), .C1(
        n18820), .C2(n18836), .ZN(P3_U3055) );
  OAI222_X1 U21939 ( .A1(n18826), .A2(n18824), .B1(n18823), .B2(n18843), .C1(
        n18822), .C2(n18830), .ZN(P3_U3056) );
  OAI222_X1 U21940 ( .A1(n18826), .A2(n18827), .B1(n18825), .B2(n18843), .C1(
        n18824), .C2(n18830), .ZN(P3_U3057) );
  OAI222_X1 U21941 ( .A1(n18826), .A2(n21059), .B1(n18828), .B2(n18843), .C1(
        n18827), .C2(n18830), .ZN(P3_U3058) );
  OAI222_X1 U21942 ( .A1(n21059), .A2(n18830), .B1(n18829), .B2(n18843), .C1(
        n18831), .C2(n18826), .ZN(P3_U3059) );
  OAI222_X1 U21943 ( .A1(n18826), .A2(n18835), .B1(n18832), .B2(n18843), .C1(
        n18831), .C2(n18836), .ZN(P3_U3060) );
  OAI222_X1 U21944 ( .A1(n18836), .A2(n18835), .B1(n18834), .B2(n18843), .C1(
        n18833), .C2(n18826), .ZN(P3_U3061) );
  INV_X1 U21945 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18837) );
  AOI22_X1 U21946 ( .A1(n18843), .A2(n18838), .B1(n18837), .B2(n18908), .ZN(
        P3_U3274) );
  INV_X1 U21947 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21107) );
  INV_X1 U21948 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18839) );
  AOI22_X1 U21949 ( .A1(n18843), .A2(n21107), .B1(n18839), .B2(n18908), .ZN(
        P3_U3275) );
  INV_X1 U21950 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18840) );
  AOI22_X1 U21951 ( .A1(n18843), .A2(n18841), .B1(n18840), .B2(n18908), .ZN(
        P3_U3276) );
  INV_X1 U21952 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18886) );
  INV_X1 U21953 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18842) );
  AOI22_X1 U21954 ( .A1(n18843), .A2(n18886), .B1(n18842), .B2(n18908), .ZN(
        P3_U3277) );
  OAI21_X1 U21955 ( .B1(n18847), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18845), 
        .ZN(n18844) );
  INV_X1 U21956 ( .A(n18844), .ZN(P3_U3280) );
  OAI21_X1 U21957 ( .B1(n18847), .B2(n18846), .A(n18845), .ZN(P3_U3281) );
  OAI221_X1 U21958 ( .B1(n18850), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18850), 
        .C2(n18849), .A(n18848), .ZN(P3_U3282) );
  NOR2_X1 U21959 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18851), .ZN(
        n18853) );
  AOI22_X1 U21960 ( .A1(n18874), .A2(n18854), .B1(n18853), .B2(n18852), .ZN(
        n18858) );
  AOI21_X1 U21961 ( .B1(n18911), .B2(n18855), .A(n18880), .ZN(n18857) );
  OAI22_X1 U21962 ( .A1(n18880), .A2(n18858), .B1(n18857), .B2(n18856), .ZN(
        P3_U3285) );
  NOR2_X1 U21963 ( .A1(n18859), .A2(n18876), .ZN(n18868) );
  AOI22_X1 U21964 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18861), .B2(n18860), .ZN(
        n18867) );
  AOI222_X1 U21965 ( .A1(n18863), .A2(n18911), .B1(n18868), .B2(n18867), .C1(
        n18874), .C2(n18862), .ZN(n18864) );
  AOI22_X1 U21966 ( .A1(n18880), .A2(n18865), .B1(n18864), .B2(n18877), .ZN(
        P3_U3288) );
  INV_X1 U21967 ( .A(n18866), .ZN(n18871) );
  INV_X1 U21968 ( .A(n18867), .ZN(n18869) );
  AOI222_X1 U21969 ( .A1(n18871), .A2(n18911), .B1(n18874), .B2(n18870), .C1(
        n18869), .C2(n18868), .ZN(n18872) );
  AOI22_X1 U21970 ( .A1(n18880), .A2(n18873), .B1(n18872), .B2(n18877), .ZN(
        P3_U3289) );
  AOI222_X1 U21971 ( .A1(n18876), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18911), 
        .B2(n18875), .C1(n18879), .C2(n18874), .ZN(n18878) );
  AOI22_X1 U21972 ( .A1(n18880), .A2(n18879), .B1(n18878), .B2(n18877), .ZN(
        P3_U3290) );
  AOI21_X1 U21973 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18882) );
  AOI22_X1 U21974 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18882), .B2(n18881), .ZN(n18884) );
  AOI22_X1 U21975 ( .A1(n18887), .A2(n18884), .B1(n21107), .B2(n18883), .ZN(
        P3_U3292) );
  OAI21_X1 U21976 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18887), .ZN(n18885) );
  OAI21_X1 U21977 ( .B1(n18887), .B2(n18886), .A(n18885), .ZN(P3_U3293) );
  INV_X1 U21978 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18888) );
  AOI22_X1 U21979 ( .A1(n18843), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18888), 
        .B2(n18908), .ZN(P3_U3294) );
  MUX2_X1 U21980 ( .A(P3_MORE_REG_SCAN_IN), .B(n18890), .S(n18889), .Z(
        P3_U3295) );
  AOI21_X1 U21981 ( .B1(n18893), .B2(n18892), .A(n18891), .ZN(n18894) );
  INV_X1 U21982 ( .A(n18894), .ZN(n18896) );
  AOI211_X1 U21983 ( .C1(n18912), .C2(n18896), .A(n18895), .B(n18910), .ZN(
        n18899) );
  OAI21_X1 U21984 ( .B1(n18899), .B2(n18898), .A(n18897), .ZN(n18907) );
  OAI21_X1 U21985 ( .B1(n18902), .B2(n18901), .A(n18900), .ZN(n18903) );
  AOI21_X1 U21986 ( .B1(n18905), .B2(n18904), .A(n18903), .ZN(n18906) );
  MUX2_X1 U21987 ( .A(n18907), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18906), 
        .Z(P3_U3296) );
  INV_X1 U21988 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18916) );
  INV_X1 U21989 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18909) );
  AOI22_X1 U21990 ( .A1(n18843), .A2(n18916), .B1(n18909), .B2(n18908), .ZN(
        P3_U3297) );
  AOI21_X1 U21991 ( .B1(n18911), .B2(n18910), .A(n18913), .ZN(n18917) );
  INV_X1 U21992 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18914) );
  AOI22_X1 U21993 ( .A1(n18917), .A2(n18914), .B1(n18913), .B2(n18912), .ZN(
        P3_U3298) );
  AOI21_X1 U21994 ( .B1(n18917), .B2(n18916), .A(n18915), .ZN(P3_U3299) );
  INV_X1 U21995 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19852) );
  INV_X1 U21996 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18918) );
  NAND2_X1 U21997 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19872), .ZN(n19860) );
  NAND2_X1 U21998 ( .A1(n19852), .A2(n19851), .ZN(n19856) );
  OAI21_X1 U21999 ( .B1(n19852), .B2(n19860), .A(n19856), .ZN(n19937) );
  OAI21_X1 U22000 ( .B1(n19852), .B2(n18918), .A(n19850), .ZN(P2_U2815) );
  INV_X1 U22001 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20973) );
  OAI22_X1 U22002 ( .A1(n18920), .A2(n20973), .B1(n13085), .B2(n18919), .ZN(
        P2_U2816) );
  NAND2_X1 U22003 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19852), .ZN(n20005) );
  AOI21_X1 U22004 ( .B1(n19852), .B2(n19872), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18921) );
  AOI22_X1 U22005 ( .A1(n19916), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18921), 
        .B2(n20005), .ZN(P2_U2817) );
  OAI21_X1 U22006 ( .B1(n19866), .B2(BS16), .A(n19937), .ZN(n19935) );
  OAI21_X1 U22007 ( .B1(n19937), .B2(n18922), .A(n19935), .ZN(P2_U2818) );
  NOR4_X1 U22008 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18926) );
  NOR4_X1 U22009 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18925) );
  NOR4_X1 U22010 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18924) );
  NOR4_X1 U22011 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18923) );
  NAND4_X1 U22012 ( .A1(n18926), .A2(n18925), .A3(n18924), .A4(n18923), .ZN(
        n18932) );
  NOR4_X1 U22013 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18930) );
  AOI211_X1 U22014 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18929) );
  NOR4_X1 U22015 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18928) );
  NOR4_X1 U22016 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18927) );
  NAND4_X1 U22017 ( .A1(n18930), .A2(n18929), .A3(n18928), .A4(n18927), .ZN(
        n18931) );
  NOR2_X1 U22018 ( .A1(n18932), .A2(n18931), .ZN(n18939) );
  INV_X1 U22019 ( .A(n18939), .ZN(n18938) );
  NOR2_X1 U22020 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18938), .ZN(n18933) );
  INV_X1 U22021 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19933) );
  AOI22_X1 U22022 ( .A1(n18933), .A2(n10242), .B1(n18938), .B2(n19933), .ZN(
        P2_U2820) );
  OR3_X1 U22023 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18937) );
  INV_X1 U22024 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U22025 ( .A1(n18933), .A2(n18937), .B1(n18938), .B2(n19931), .ZN(
        P2_U2821) );
  INV_X1 U22026 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19936) );
  NAND2_X1 U22027 ( .A1(n18933), .A2(n19936), .ZN(n18936) );
  OAI21_X1 U22028 ( .B1(n10242), .B2(n19874), .A(n18939), .ZN(n18934) );
  OAI21_X1 U22029 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18939), .A(n18934), 
        .ZN(n18935) );
  OAI221_X1 U22030 ( .B1(n18936), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18936), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18935), .ZN(P2_U2822) );
  INV_X1 U22031 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19929) );
  OAI221_X1 U22032 ( .B1(n18939), .B2(n19929), .C1(n18938), .C2(n18937), .A(
        n18936), .ZN(P2_U2823) );
  OAI22_X1 U22033 ( .A1(n18940), .A2(n19149), .B1(n19906), .B2(n19142), .ZN(
        n18944) );
  OAI22_X1 U22034 ( .A1(n19115), .A2(n18942), .B1(n18941), .B2(n19139), .ZN(
        n18943) );
  AOI211_X1 U22035 ( .C1(n18945), .C2(n19151), .A(n18944), .B(n18943), .ZN(
        n18950) );
  OAI211_X1 U22036 ( .C1(n18948), .C2(n18947), .A(n19123), .B(n18946), .ZN(
        n18949) );
  OAI211_X1 U22037 ( .C1(n19144), .C2(n18951), .A(n18950), .B(n18949), .ZN(
        P2_U2834) );
  AOI22_X1 U22038 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19146), .B1(n19089), 
        .B2(n18952), .ZN(n18961) );
  AOI22_X1 U22039 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19127), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19130), .ZN(n18960) );
  AOI22_X1 U22040 ( .A1(n18954), .A2(n19151), .B1(n18953), .B2(n19098), .ZN(
        n18959) );
  OAI211_X1 U22041 ( .C1(n18957), .C2(n18956), .A(n19123), .B(n18955), .ZN(
        n18958) );
  NAND4_X1 U22042 ( .A1(n18961), .A2(n18960), .A3(n18959), .A4(n18958), .ZN(
        P2_U2835) );
  OAI21_X1 U22043 ( .B1(n19903), .B2(n19142), .A(n19328), .ZN(n18965) );
  OAI22_X1 U22044 ( .A1(n18963), .A2(n19139), .B1(n18962), .B2(n19149), .ZN(
        n18964) );
  AOI211_X1 U22045 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19146), .A(n18965), .B(
        n18964), .ZN(n18972) );
  AOI22_X1 U22046 ( .A1(n18966), .A2(n19151), .B1(n10082), .B2(n19098), .ZN(
        n18971) );
  OAI211_X1 U22047 ( .C1(n18969), .C2(n18968), .A(n19123), .B(n18967), .ZN(
        n18970) );
  NAND3_X1 U22048 ( .A1(n18972), .A2(n18971), .A3(n18970), .ZN(P2_U2836) );
  AOI22_X1 U22049 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19127), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19146), .ZN(n18973) );
  OAI21_X1 U22050 ( .B1(n18974), .B2(n19149), .A(n18973), .ZN(n18975) );
  AOI211_X1 U22051 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19130), .A(n19291), 
        .B(n18975), .ZN(n18983) );
  AOI22_X1 U22052 ( .A1(n18977), .A2(n19151), .B1(n18976), .B2(n19098), .ZN(
        n18982) );
  OAI211_X1 U22053 ( .C1(n18980), .C2(n18979), .A(n19123), .B(n18978), .ZN(
        n18981) );
  NAND3_X1 U22054 ( .A1(n18983), .A2(n18982), .A3(n18981), .ZN(P2_U2837) );
  OAI21_X1 U22055 ( .B1(n19900), .B2(n19142), .A(n19328), .ZN(n18987) );
  OAI22_X1 U22056 ( .A1(n18985), .A2(n19139), .B1(n18984), .B2(n19149), .ZN(
        n18986) );
  AOI211_X1 U22057 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19146), .A(n18987), .B(
        n18986), .ZN(n18995) );
  AOI22_X1 U22058 ( .A1(n18989), .A2(n19098), .B1(n18988), .B2(n19151), .ZN(
        n18994) );
  OAI211_X1 U22059 ( .C1(n18992), .C2(n18991), .A(n19123), .B(n18990), .ZN(
        n18993) );
  NAND3_X1 U22060 ( .A1(n18995), .A2(n18994), .A3(n18993), .ZN(P2_U2838) );
  NAND2_X1 U22061 ( .A1(n9704), .A2(n18996), .ZN(n18997) );
  XNOR2_X1 U22062 ( .A(n18998), .B(n18997), .ZN(n19006) );
  OAI21_X1 U22063 ( .B1(n19898), .B2(n19142), .A(n19328), .ZN(n19002) );
  OAI22_X1 U22064 ( .A1(n19000), .A2(n19149), .B1(n18999), .B2(n19139), .ZN(
        n19001) );
  AOI211_X1 U22065 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19146), .A(n19002), .B(
        n19001), .ZN(n19005) );
  AOI22_X1 U22066 ( .A1(n19161), .A2(n19098), .B1(n19003), .B2(n19151), .ZN(
        n19004) );
  OAI211_X1 U22067 ( .C1(n19847), .C2(n19006), .A(n19005), .B(n19004), .ZN(
        P2_U2839) );
  OAI22_X1 U22068 ( .A1(n19008), .A2(n19139), .B1(n19007), .B2(n19149), .ZN(
        n19009) );
  AOI211_X1 U22069 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19130), .A(n19291), 
        .B(n19009), .ZN(n19017) );
  NOR2_X1 U22070 ( .A1(n9963), .A2(n19010), .ZN(n19011) );
  XNOR2_X1 U22071 ( .A(n19012), .B(n19011), .ZN(n19015) );
  OAI22_X1 U22072 ( .A1(n19013), .A2(n19121), .B1(n19168), .B2(n19144), .ZN(
        n19014) );
  AOI21_X1 U22073 ( .B1(n19015), .B2(n19123), .A(n19014), .ZN(n19016) );
  OAI211_X1 U22074 ( .C1(n19115), .C2(n10877), .A(n19017), .B(n19016), .ZN(
        P2_U2840) );
  NAND2_X1 U22075 ( .A1(n9704), .A2(n19018), .ZN(n19019) );
  XOR2_X1 U22076 ( .A(n19020), .B(n19019), .Z(n19027) );
  AOI22_X1 U22077 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19127), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19146), .ZN(n19021) );
  OAI21_X1 U22078 ( .B1(n19022), .B2(n19149), .A(n19021), .ZN(n19023) );
  AOI211_X1 U22079 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19130), .A(n19291), 
        .B(n19023), .ZN(n19026) );
  AOI22_X1 U22080 ( .A1(n19151), .A2(n19024), .B1(n19098), .B2(n19169), .ZN(
        n19025) );
  OAI211_X1 U22081 ( .C1(n19847), .C2(n19027), .A(n19026), .B(n19025), .ZN(
        P2_U2841) );
  OAI22_X1 U22082 ( .A1(n19115), .A2(n10870), .B1(n19028), .B2(n19149), .ZN(
        n19029) );
  AOI211_X1 U22083 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19130), .A(n19291), 
        .B(n19029), .ZN(n19037) );
  NOR2_X1 U22084 ( .A1(n9963), .A2(n19030), .ZN(n19031) );
  XNOR2_X1 U22085 ( .A(n19032), .B(n19031), .ZN(n19035) );
  OAI22_X1 U22086 ( .A1(n19121), .A2(n19033), .B1(n19144), .B2(n19173), .ZN(
        n19034) );
  AOI21_X1 U22087 ( .B1(n19035), .B2(n19123), .A(n19034), .ZN(n19036) );
  OAI211_X1 U22088 ( .C1(n19038), .C2(n19139), .A(n19037), .B(n19036), .ZN(
        P2_U2842) );
  NAND2_X1 U22089 ( .A1(n9704), .A2(n19039), .ZN(n19040) );
  XOR2_X1 U22090 ( .A(n19041), .B(n19040), .Z(n19048) );
  AOI22_X1 U22091 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19127), .B1(
        n19042), .B2(n19089), .ZN(n19043) );
  OAI211_X1 U22092 ( .C1(n19890), .C2(n19142), .A(n19043), .B(n19328), .ZN(
        n19044) );
  AOI21_X1 U22093 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n19146), .A(n19044), .ZN(
        n19047) );
  AOI22_X1 U22094 ( .A1(n19151), .A2(n19045), .B1(n19098), .B2(n19174), .ZN(
        n19046) );
  OAI211_X1 U22095 ( .C1(n19847), .C2(n19048), .A(n19047), .B(n19046), .ZN(
        P2_U2843) );
  NOR2_X1 U22096 ( .A1(n9963), .A2(n19049), .ZN(n19050) );
  XOR2_X1 U22097 ( .A(n19051), .B(n19050), .Z(n19058) );
  AOI22_X1 U22098 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19127), .B1(
        n19052), .B2(n19089), .ZN(n19053) );
  OAI211_X1 U22099 ( .C1(n19889), .C2(n19142), .A(n19053), .B(n19091), .ZN(
        n19056) );
  OAI22_X1 U22100 ( .A1(n19121), .A2(n19054), .B1(n19144), .B2(n19176), .ZN(
        n19055) );
  AOI211_X1 U22101 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19146), .A(n19056), .B(
        n19055), .ZN(n19057) );
  OAI21_X1 U22102 ( .B1(n19847), .B2(n19058), .A(n19057), .ZN(P2_U2844) );
  AOI22_X1 U22103 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(n19146), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19127), .ZN(n19059) );
  OAI21_X1 U22104 ( .B1(n19060), .B2(n19149), .A(n19059), .ZN(n19061) );
  AOI211_X1 U22105 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19130), .A(n19291), 
        .B(n19061), .ZN(n19067) );
  NAND2_X1 U22106 ( .A1(n9704), .A2(n19062), .ZN(n19063) );
  XNOR2_X1 U22107 ( .A(n19064), .B(n19063), .ZN(n19065) );
  AOI22_X1 U22108 ( .A1(n19123), .A2(n19065), .B1(n19098), .B2(n19177), .ZN(
        n19066) );
  OAI211_X1 U22109 ( .C1(n19121), .C2(n19068), .A(n19067), .B(n19066), .ZN(
        P2_U2845) );
  NOR2_X1 U22110 ( .A1(n9963), .A2(n19069), .ZN(n19070) );
  XOR2_X1 U22111 ( .A(n19071), .B(n19070), .Z(n19078) );
  AOI22_X1 U22112 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19127), .B1(
        n19089), .B2(n19072), .ZN(n19073) );
  OAI211_X1 U22113 ( .C1(n15253), .C2(n19142), .A(n19073), .B(n19091), .ZN(
        n19076) );
  OAI22_X1 U22114 ( .A1(n19121), .A2(n19074), .B1(n19144), .B2(n19181), .ZN(
        n19075) );
  AOI211_X1 U22115 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19146), .A(n19076), .B(
        n19075), .ZN(n19077) );
  OAI21_X1 U22116 ( .B1(n19847), .B2(n19078), .A(n19077), .ZN(P2_U2846) );
  NAND2_X1 U22117 ( .A1(n9704), .A2(n19079), .ZN(n19080) );
  XOR2_X1 U22118 ( .A(n19081), .B(n19080), .Z(n19088) );
  AOI22_X1 U22119 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19127), .B1(
        n19082), .B2(n19089), .ZN(n19083) );
  OAI211_X1 U22120 ( .C1(n19884), .C2(n19142), .A(n19083), .B(n19091), .ZN(
        n19084) );
  AOI21_X1 U22121 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19146), .A(n19084), .ZN(
        n19087) );
  AOI22_X1 U22122 ( .A1(n19151), .A2(n19085), .B1(n19098), .B2(n19182), .ZN(
        n19086) );
  OAI211_X1 U22123 ( .C1(n19847), .C2(n19088), .A(n19087), .B(n19086), .ZN(
        P2_U2847) );
  AOI22_X1 U22124 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19127), .B1(
        n19090), .B2(n19089), .ZN(n19092) );
  OAI211_X1 U22125 ( .C1(n19882), .C2(n19142), .A(n19092), .B(n19091), .ZN(
        n19093) );
  AOI21_X1 U22126 ( .B1(P2_EBX_REG_7__SCAN_IN), .B2(n19146), .A(n19093), .ZN(
        n19101) );
  NOR2_X1 U22127 ( .A1(n9963), .A2(n19094), .ZN(n19096) );
  XNOR2_X1 U22128 ( .A(n19096), .B(n19095), .ZN(n19099) );
  AOI22_X1 U22129 ( .A1(n19123), .A2(n19099), .B1(n19098), .B2(n19097), .ZN(
        n19100) );
  OAI211_X1 U22130 ( .C1(n19121), .C2(n19102), .A(n19101), .B(n19100), .ZN(
        P2_U2848) );
  OAI21_X1 U22131 ( .B1(n19880), .B2(n19142), .A(n19328), .ZN(n19106) );
  OAI22_X1 U22132 ( .A1(n19104), .A2(n19139), .B1(n19103), .B2(n19149), .ZN(
        n19105) );
  AOI211_X1 U22133 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19146), .A(n19106), .B(
        n19105), .ZN(n19113) );
  NAND2_X1 U22134 ( .A1(n9704), .A2(n19107), .ZN(n19108) );
  XNOR2_X1 U22135 ( .A(n19109), .B(n19108), .ZN(n19110) );
  AOI22_X1 U22136 ( .A1(n19151), .A2(n19111), .B1(n19123), .B2(n19110), .ZN(
        n19112) );
  OAI211_X1 U22137 ( .C1(n19144), .C2(n19188), .A(n19113), .B(n19112), .ZN(
        P2_U2849) );
  OAI22_X1 U22138 ( .A1(n19115), .A2(n10835), .B1(n19114), .B2(n19149), .ZN(
        n19116) );
  AOI211_X1 U22139 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19130), .A(n19291), .B(
        n19116), .ZN(n19126) );
  NOR2_X1 U22140 ( .A1(n9963), .A2(n19117), .ZN(n19118) );
  XNOR2_X1 U22141 ( .A(n19119), .B(n19118), .ZN(n19124) );
  OAI22_X1 U22142 ( .A1(n19121), .A2(n19120), .B1(n19144), .B2(n19196), .ZN(
        n19122) );
  AOI21_X1 U22143 ( .B1(n19124), .B2(n19123), .A(n19122), .ZN(n19125) );
  OAI211_X1 U22144 ( .C1(n9975), .C2(n19139), .A(n19126), .B(n19125), .ZN(
        P2_U2850) );
  AOI22_X1 U22145 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19127), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19146), .ZN(n19138) );
  OAI22_X1 U22146 ( .A1(n19128), .A2(n19149), .B1(n19144), .B2(n19329), .ZN(
        n19129) );
  AOI211_X1 U22147 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19130), .A(n19291), .B(
        n19129), .ZN(n19137) );
  INV_X1 U22148 ( .A(n19131), .ZN(n19192) );
  AOI22_X1 U22149 ( .A1(n19192), .A2(n19141), .B1(n19151), .B2(n19339), .ZN(
        n19136) );
  AND2_X1 U22150 ( .A1(n9704), .A2(n19132), .ZN(n19134) );
  AOI21_X1 U22151 ( .B1(n19289), .B2(n19134), .A(n19847), .ZN(n19133) );
  OAI21_X1 U22152 ( .B1(n19289), .B2(n19134), .A(n19133), .ZN(n19135) );
  NAND4_X1 U22153 ( .A1(n19138), .A2(n19137), .A3(n19136), .A4(n19135), .ZN(
        P2_U2851) );
  NAND2_X1 U22154 ( .A1(n19139), .A2(n19847), .ZN(n19140) );
  AOI22_X1 U22155 ( .A1(n19970), .A2(n19141), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19140), .ZN(n19153) );
  OAI22_X1 U22156 ( .A1(n19144), .A2(n19143), .B1(n10242), .B2(n19142), .ZN(
        n19145) );
  AOI21_X1 U22157 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19146), .A(n19145), .ZN(
        n19147) );
  OAI21_X1 U22158 ( .B1(n19149), .B2(n19148), .A(n19147), .ZN(n19150) );
  AOI21_X1 U22159 ( .B1(n19320), .B2(n19151), .A(n19150), .ZN(n19152) );
  NAND2_X1 U22160 ( .A1(n19153), .A2(n19152), .ZN(P2_U2855) );
  AOI22_X1 U22161 ( .A1(n19154), .A2(n19206), .B1(n19159), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19156) );
  AOI22_X1 U22162 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19205), .B1(n19160), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19155) );
  NAND2_X1 U22163 ( .A1(n19156), .A2(n19155), .ZN(P2_U2888) );
  AOI22_X1 U22164 ( .A1(n19158), .A2(n19157), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19205), .ZN(n19165) );
  AOI22_X1 U22165 ( .A1(n19160), .A2(BUF1_REG_16__SCAN_IN), .B1(n19159), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19164) );
  AOI22_X1 U22166 ( .A1(n19162), .A2(n19191), .B1(n19161), .B2(n19206), .ZN(
        n19163) );
  NAND3_X1 U22167 ( .A1(n19165), .A2(n19164), .A3(n19163), .ZN(P2_U2903) );
  INV_X1 U22168 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U22169 ( .A1(n19167), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19166), .ZN(n19288) );
  OAI222_X1 U22170 ( .A1(n19168), .A2(n19197), .B1(n19219), .B2(n19187), .C1(
        n19288), .C2(n19214), .ZN(P2_U2904) );
  INV_X1 U22171 ( .A(n19169), .ZN(n19172) );
  AOI22_X1 U22172 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19205), .B1(n19170), 
        .B2(n19189), .ZN(n19171) );
  OAI21_X1 U22173 ( .B1(n19197), .B2(n19172), .A(n19171), .ZN(P2_U2905) );
  INV_X1 U22174 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19223) );
  OAI222_X1 U22175 ( .A1(n19173), .A2(n19197), .B1(n19223), .B2(n19187), .C1(
        n19214), .C2(n19283), .ZN(P2_U2906) );
  INV_X1 U22176 ( .A(n19174), .ZN(n19175) );
  INV_X1 U22177 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19225) );
  OAI222_X1 U22178 ( .A1(n19175), .A2(n19197), .B1(n19225), .B2(n19187), .C1(
        n19214), .C2(n19281), .ZN(P2_U2907) );
  INV_X1 U22179 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19227) );
  OAI222_X1 U22180 ( .A1(n19176), .A2(n19197), .B1(n19227), .B2(n19187), .C1(
        n19214), .C2(n19279), .ZN(P2_U2908) );
  INV_X1 U22181 ( .A(n19177), .ZN(n19180) );
  AOI22_X1 U22182 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19205), .B1(n19178), 
        .B2(n19189), .ZN(n19179) );
  OAI21_X1 U22183 ( .B1(n19197), .B2(n19180), .A(n19179), .ZN(P2_U2909) );
  INV_X1 U22184 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19231) );
  OAI222_X1 U22185 ( .A1(n19181), .A2(n19197), .B1(n19231), .B2(n19187), .C1(
        n19214), .C2(n19277), .ZN(P2_U2910) );
  INV_X1 U22186 ( .A(n19182), .ZN(n19185) );
  AOI22_X1 U22187 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19205), .B1(n19183), .B2(
        n19189), .ZN(n19184) );
  OAI21_X1 U22188 ( .B1(n19197), .B2(n19185), .A(n19184), .ZN(P2_U2911) );
  INV_X1 U22189 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19235) );
  OAI222_X1 U22190 ( .A1(n19186), .A2(n19197), .B1(n19235), .B2(n19187), .C1(
        n19214), .C2(n19275), .ZN(P2_U2912) );
  INV_X1 U22191 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20965) );
  OAI222_X1 U22192 ( .A1(n19188), .A2(n19197), .B1(n20965), .B2(n19187), .C1(
        n19214), .C2(n19273), .ZN(P2_U2913) );
  INV_X1 U22193 ( .A(n19271), .ZN(n19190) );
  AOI22_X1 U22194 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19205), .B1(n19190), .B2(
        n19189), .ZN(n19195) );
  NAND3_X1 U22195 ( .A1(n19193), .A2(n19192), .A3(n19191), .ZN(n19194) );
  OAI211_X1 U22196 ( .C1(n19197), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        P2_U2914) );
  AOI22_X1 U22197 ( .A1(n19206), .A2(n19198), .B1(n19205), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19204) );
  AOI21_X1 U22198 ( .B1(n19201), .B2(n19200), .A(n19199), .ZN(n19202) );
  OR2_X1 U22199 ( .A1(n19202), .A2(n19210), .ZN(n19203) );
  OAI211_X1 U22200 ( .C1(n19358), .C2(n19214), .A(n19204), .B(n19203), .ZN(
        P2_U2916) );
  AOI22_X1 U22201 ( .A1(n19206), .A2(n19965), .B1(n19205), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19213) );
  AOI21_X1 U22202 ( .B1(n19209), .B2(n19208), .A(n19207), .ZN(n19211) );
  OR2_X1 U22203 ( .A1(n19211), .A2(n19210), .ZN(n19212) );
  OAI211_X1 U22204 ( .C1(n19349), .C2(n19214), .A(n19213), .B(n19212), .ZN(
        P2_U2918) );
  NOR2_X1 U22205 ( .A1(n19216), .A2(n19215), .ZN(P2_U2920) );
  AOI22_X1 U22206 ( .A1(n9637), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19218) );
  OAI21_X1 U22207 ( .B1(n19219), .B2(n19249), .A(n19218), .ZN(P2_U2936) );
  AOI22_X1 U22208 ( .A1(n9637), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19220) );
  OAI21_X1 U22209 ( .B1(n19221), .B2(n19249), .A(n19220), .ZN(P2_U2937) );
  AOI22_X1 U22210 ( .A1(n9637), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19222) );
  OAI21_X1 U22211 ( .B1(n19223), .B2(n19249), .A(n19222), .ZN(P2_U2938) );
  AOI22_X1 U22212 ( .A1(n9637), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19224) );
  OAI21_X1 U22213 ( .B1(n19225), .B2(n19249), .A(n19224), .ZN(P2_U2939) );
  AOI22_X1 U22214 ( .A1(n9637), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19226) );
  OAI21_X1 U22215 ( .B1(n19227), .B2(n19249), .A(n19226), .ZN(P2_U2940) );
  AOI22_X1 U22216 ( .A1(n9637), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19228) );
  OAI21_X1 U22217 ( .B1(n19229), .B2(n19249), .A(n19228), .ZN(P2_U2941) );
  AOI22_X1 U22218 ( .A1(n9637), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19230) );
  OAI21_X1 U22219 ( .B1(n19231), .B2(n19249), .A(n19230), .ZN(P2_U2942) );
  AOI22_X1 U22220 ( .A1(n9637), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19232) );
  OAI21_X1 U22221 ( .B1(n19233), .B2(n19249), .A(n19232), .ZN(P2_U2943) );
  AOI22_X1 U22222 ( .A1(n9637), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19234) );
  OAI21_X1 U22223 ( .B1(n19235), .B2(n19249), .A(n19234), .ZN(P2_U2944) );
  AOI22_X1 U22224 ( .A1(n9637), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19236) );
  OAI21_X1 U22225 ( .B1(n20965), .B2(n19249), .A(n19236), .ZN(P2_U2945) );
  INV_X1 U22226 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19238) );
  AOI22_X1 U22227 ( .A1(n9637), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19237) );
  OAI21_X1 U22228 ( .B1(n19238), .B2(n19249), .A(n19237), .ZN(P2_U2946) );
  INV_X1 U22229 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19240) );
  AOI22_X1 U22230 ( .A1(n9637), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19239) );
  OAI21_X1 U22231 ( .B1(n19240), .B2(n19249), .A(n19239), .ZN(P2_U2947) );
  INV_X1 U22232 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19242) );
  AOI22_X1 U22233 ( .A1(n9637), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19241) );
  OAI21_X1 U22234 ( .B1(n19242), .B2(n19249), .A(n19241), .ZN(P2_U2948) );
  INV_X1 U22235 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19244) );
  AOI22_X1 U22236 ( .A1(n9637), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19243) );
  OAI21_X1 U22237 ( .B1(n19244), .B2(n19249), .A(n19243), .ZN(P2_U2949) );
  INV_X1 U22238 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19246) );
  AOI22_X1 U22239 ( .A1(n9637), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19245) );
  OAI21_X1 U22240 ( .B1(n19246), .B2(n19249), .A(n19245), .ZN(P2_U2950) );
  INV_X1 U22241 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19250) );
  AOI22_X1 U22242 ( .A1(n9637), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19247), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19248) );
  OAI21_X1 U22243 ( .B1(n19250), .B2(n19249), .A(n19248), .ZN(P2_U2951) );
  AOI22_X1 U22244 ( .A1(n19285), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n19251) );
  OAI21_X1 U22245 ( .B1(n19349), .B2(n19287), .A(n19251), .ZN(P2_U2953) );
  INV_X1 U22246 ( .A(n19252), .ZN(n19353) );
  AOI22_X1 U22247 ( .A1(n13523), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19284), .ZN(n19253) );
  OAI21_X1 U22248 ( .B1(n19353), .B2(n19287), .A(n19253), .ZN(P2_U2954) );
  AOI22_X1 U22249 ( .A1(n13523), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n19254) );
  OAI21_X1 U22250 ( .B1(n19358), .B2(n19287), .A(n19254), .ZN(P2_U2955) );
  INV_X1 U22251 ( .A(n19255), .ZN(n19365) );
  AOI22_X1 U22252 ( .A1(n13523), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19284), .ZN(n19256) );
  OAI21_X1 U22253 ( .B1(n19365), .B2(n19287), .A(n19256), .ZN(P2_U2956) );
  AOI22_X1 U22254 ( .A1(n13523), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n19257) );
  OAI21_X1 U22255 ( .B1(n19271), .B2(n19287), .A(n19257), .ZN(P2_U2957) );
  AOI22_X1 U22256 ( .A1(n13523), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19284), .ZN(n19258) );
  OAI21_X1 U22257 ( .B1(n19273), .B2(n19287), .A(n19258), .ZN(P2_U2958) );
  AOI22_X1 U22258 ( .A1(n13523), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n19259) );
  OAI21_X1 U22259 ( .B1(n19275), .B2(n19287), .A(n19259), .ZN(P2_U2959) );
  AOI22_X1 U22260 ( .A1(n13523), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19284), .ZN(n19260) );
  OAI21_X1 U22261 ( .B1(n19277), .B2(n19287), .A(n19260), .ZN(P2_U2961) );
  AOI22_X1 U22262 ( .A1(n13523), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19284), .ZN(n19261) );
  OAI21_X1 U22263 ( .B1(n19279), .B2(n19287), .A(n19261), .ZN(P2_U2963) );
  AOI22_X1 U22264 ( .A1(n13523), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19284), .ZN(n19262) );
  OAI21_X1 U22265 ( .B1(n19281), .B2(n19287), .A(n19262), .ZN(P2_U2964) );
  AOI22_X1 U22266 ( .A1(n19285), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19284), .ZN(n19263) );
  OAI21_X1 U22267 ( .B1(n19283), .B2(n19287), .A(n19263), .ZN(P2_U2965) );
  AOI22_X1 U22268 ( .A1(n19285), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n19264) );
  OAI21_X1 U22269 ( .B1(n19265), .B2(n19287), .A(n19264), .ZN(P2_U2967) );
  AOI22_X1 U22270 ( .A1(n19285), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n19266) );
  OAI21_X1 U22271 ( .B1(n19349), .B2(n19287), .A(n19266), .ZN(P2_U2968) );
  AOI22_X1 U22272 ( .A1(n19285), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19284), .ZN(n19267) );
  OAI21_X1 U22273 ( .B1(n19353), .B2(n19287), .A(n19267), .ZN(P2_U2969) );
  AOI22_X1 U22274 ( .A1(n19285), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19284), .ZN(n19268) );
  OAI21_X1 U22275 ( .B1(n19358), .B2(n19287), .A(n19268), .ZN(P2_U2970) );
  AOI22_X1 U22276 ( .A1(n19285), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19284), .ZN(n19269) );
  OAI21_X1 U22277 ( .B1(n19365), .B2(n19287), .A(n19269), .ZN(P2_U2971) );
  AOI22_X1 U22278 ( .A1(n19285), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n19270) );
  OAI21_X1 U22279 ( .B1(n19271), .B2(n19287), .A(n19270), .ZN(P2_U2972) );
  AOI22_X1 U22280 ( .A1(n19285), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n19272) );
  OAI21_X1 U22281 ( .B1(n19273), .B2(n19287), .A(n19272), .ZN(P2_U2973) );
  AOI22_X1 U22282 ( .A1(n19285), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n19274) );
  OAI21_X1 U22283 ( .B1(n19275), .B2(n19287), .A(n19274), .ZN(P2_U2974) );
  AOI22_X1 U22284 ( .A1(n19285), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n19276) );
  OAI21_X1 U22285 ( .B1(n19277), .B2(n19287), .A(n19276), .ZN(P2_U2976) );
  AOI22_X1 U22286 ( .A1(n19285), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n19278) );
  OAI21_X1 U22287 ( .B1(n19279), .B2(n19287), .A(n19278), .ZN(P2_U2978) );
  AOI22_X1 U22288 ( .A1(n19285), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19284), .ZN(n19280) );
  OAI21_X1 U22289 ( .B1(n19281), .B2(n19287), .A(n19280), .ZN(P2_U2979) );
  AOI22_X1 U22290 ( .A1(n19285), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n19282) );
  OAI21_X1 U22291 ( .B1(n19283), .B2(n19287), .A(n19282), .ZN(P2_U2980) );
  AOI22_X1 U22292 ( .A1(n19285), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19284), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n19286) );
  OAI21_X1 U22293 ( .B1(n19288), .B2(n19287), .A(n19286), .ZN(P2_U2982) );
  AOI22_X1 U22294 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19291), .B1(n19290), 
        .B2(n19289), .ZN(n19300) );
  XOR2_X1 U22295 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n19292), .Z(
        n19293) );
  XNOR2_X1 U22296 ( .A(n19294), .B(n19293), .ZN(n19342) );
  XNOR2_X1 U22297 ( .A(n19296), .B(n19295), .ZN(n19332) );
  OAI22_X1 U22298 ( .A1(n19342), .A2(n19323), .B1(n19297), .B2(n19332), .ZN(
        n19298) );
  AOI21_X1 U22299 ( .B1(n19319), .B2(n19339), .A(n19298), .ZN(n19299) );
  OAI211_X1 U22300 ( .C1(n19301), .C2(n19312), .A(n19300), .B(n19299), .ZN(
        P2_U3010) );
  OAI22_X1 U22301 ( .A1(n19304), .A2(n19303), .B1(n19302), .B2(n19323), .ZN(
        n19307) );
  NOR2_X1 U22302 ( .A1(n10289), .A2(n19305), .ZN(n19306) );
  AOI211_X1 U22303 ( .C1(n19308), .C2(n19318), .A(n19307), .B(n19306), .ZN(
        n19310) );
  OAI211_X1 U22304 ( .C1(n19312), .C2(n19311), .A(n19310), .B(n19309), .ZN(
        P2_U3012) );
  OAI21_X1 U22305 ( .B1(n19314), .B2(n19313), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19327) );
  INV_X1 U22306 ( .A(n19315), .ZN(n19317) );
  AOI21_X1 U22307 ( .B1(n19318), .B2(n19317), .A(n19316), .ZN(n19322) );
  NAND2_X1 U22308 ( .A1(n19320), .A2(n19319), .ZN(n19321) );
  OAI211_X1 U22309 ( .C1(n19324), .C2(n19323), .A(n19322), .B(n19321), .ZN(
        n19325) );
  INV_X1 U22310 ( .A(n19325), .ZN(n19326) );
  NAND2_X1 U22311 ( .A1(n19327), .A2(n19326), .ZN(P2_U3014) );
  INV_X1 U22312 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19877) );
  NOR2_X1 U22313 ( .A1(n19877), .A2(n19328), .ZN(n19334) );
  OAI22_X1 U22314 ( .A1(n19332), .A2(n19331), .B1(n19330), .B2(n19329), .ZN(
        n19333) );
  AOI211_X1 U22315 ( .C1(n19336), .C2(n19335), .A(n19334), .B(n19333), .ZN(
        n19341) );
  AOI22_X1 U22316 ( .A1(n19339), .A2(n19338), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19337), .ZN(n19340) );
  OAI211_X1 U22317 ( .C1(n19343), .C2(n19342), .A(n19341), .B(n19340), .ZN(
        P2_U3042) );
  AOI22_X1 U22318 ( .A1(n19837), .A2(n19695), .B1(n19781), .B2(n19373), .ZN(
        n19345) );
  AOI22_X1 U22319 ( .A1(n19782), .A2(n19374), .B1(n19387), .B2(n19790), .ZN(
        n19344) );
  OAI211_X1 U22320 ( .C1(n19378), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P2_U3048) );
  AOI22_X1 U22321 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19361), .ZN(n19347) );
  NOR2_X2 U22322 ( .A1(n19348), .A2(n19363), .ZN(n19794) );
  AOI22_X1 U22323 ( .A1(n19837), .A2(n19796), .B1(n19373), .B2(n19794), .ZN(
        n19351) );
  NOR2_X2 U22324 ( .A1(n19349), .A2(n19601), .ZN(n19795) );
  AOI22_X2 U22325 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19361), .ZN(n19801) );
  INV_X1 U22326 ( .A(n19801), .ZN(n19750) );
  AOI22_X1 U22327 ( .A1(n19795), .A2(n19374), .B1(n19387), .B2(n19750), .ZN(
        n19350) );
  OAI211_X1 U22328 ( .C1(n19378), .C2(n10362), .A(n19351), .B(n19350), .ZN(
        P2_U3049) );
  AOI22_X2 U22329 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19361), .ZN(n19807) );
  INV_X1 U22330 ( .A(n19807), .ZN(n19753) );
  AND2_X1 U22331 ( .A1(n10205), .A2(n19352), .ZN(n19802) );
  AOI22_X1 U22332 ( .A1(n19753), .A2(n19837), .B1(n19373), .B2(n19802), .ZN(
        n19357) );
  NOR2_X2 U22333 ( .A1(n19353), .A2(n19601), .ZN(n19803) );
  OAI22_X2 U22334 ( .A1(n19355), .A2(n19368), .B1(n19354), .B2(n19366), .ZN(
        n19804) );
  AOI22_X1 U22335 ( .A1(n19803), .A2(n19374), .B1(n19387), .B2(n19804), .ZN(
        n19356) );
  OAI211_X1 U22336 ( .C1(n19378), .C2(n12773), .A(n19357), .B(n19356), .ZN(
        P2_U3050) );
  AOI22_X1 U22337 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19361), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19362), .ZN(n19813) );
  INV_X1 U22338 ( .A(n19813), .ZN(n19757) );
  NOR2_X2 U22339 ( .A1(n10204), .A2(n19363), .ZN(n19808) );
  AOI22_X1 U22340 ( .A1(n19757), .A2(n19837), .B1(n19373), .B2(n19808), .ZN(
        n19360) );
  NOR2_X2 U22341 ( .A1(n19358), .A2(n19601), .ZN(n19809) );
  OAI22_X2 U22342 ( .A1(n15111), .A2(n19368), .B1(n15109), .B2(n19366), .ZN(
        n19810) );
  AOI22_X1 U22343 ( .A1(n19809), .A2(n19374), .B1(n19387), .B2(n19810), .ZN(
        n19359) );
  OAI211_X1 U22344 ( .C1(n19378), .C2(n12758), .A(n19360), .B(n19359), .ZN(
        P2_U3051) );
  AOI22_X1 U22345 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19362), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19361), .ZN(n19819) );
  INV_X1 U22346 ( .A(n19819), .ZN(n19760) );
  AOI22_X1 U22347 ( .A1(n19760), .A2(n19837), .B1(n19373), .B2(n19814), .ZN(
        n19371) );
  NOR2_X2 U22348 ( .A1(n19365), .A2(n19601), .ZN(n19815) );
  OAI22_X2 U22349 ( .A1(n19369), .A2(n19368), .B1(n19367), .B2(n19366), .ZN(
        n19816) );
  AOI22_X1 U22350 ( .A1(n19815), .A2(n19374), .B1(n19387), .B2(n19816), .ZN(
        n19370) );
  OAI211_X1 U22351 ( .C1(n19378), .C2(n12780), .A(n19371), .B(n19370), .ZN(
        P2_U3052) );
  AOI22_X1 U22352 ( .A1(n19770), .A2(n19837), .B1(n19832), .B2(n19373), .ZN(
        n19376) );
  AOI22_X1 U22353 ( .A1(n19834), .A2(n19374), .B1(n19387), .B2(n19836), .ZN(
        n19375) );
  OAI211_X1 U22354 ( .C1(n19378), .C2(n19377), .A(n19376), .B(n19375), .ZN(
        P2_U3055) );
  AOI22_X1 U22355 ( .A1(n19395), .A2(n19782), .B1(n19781), .B2(n19394), .ZN(
        n19380) );
  AOI22_X1 U22356 ( .A1(n19426), .A2(n19790), .B1(n19387), .B2(n19695), .ZN(
        n19379) );
  OAI211_X1 U22357 ( .C1(n19382), .C2(n19381), .A(n19380), .B(n19379), .ZN(
        P2_U3056) );
  AOI22_X1 U22358 ( .A1(n19395), .A2(n19795), .B1(n19394), .B2(n19794), .ZN(
        n19384) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19396), .B1(
        n19387), .B2(n19796), .ZN(n19383) );
  OAI211_X1 U22360 ( .C1(n19801), .C2(n19423), .A(n19384), .B(n19383), .ZN(
        P2_U3057) );
  INV_X1 U22361 ( .A(n19387), .ZN(n19399) );
  AOI22_X1 U22362 ( .A1(n19395), .A2(n19803), .B1(n19394), .B2(n19802), .ZN(
        n19386) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19396), .B1(
        n19426), .B2(n19804), .ZN(n19385) );
  OAI211_X1 U22364 ( .C1(n19807), .C2(n19399), .A(n19386), .B(n19385), .ZN(
        P2_U3058) );
  INV_X1 U22365 ( .A(n19810), .ZN(n19668) );
  AOI22_X1 U22366 ( .A1(n19395), .A2(n19809), .B1(n19394), .B2(n19808), .ZN(
        n19389) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19396), .B1(
        n19387), .B2(n19757), .ZN(n19388) );
  OAI211_X1 U22368 ( .C1(n19668), .C2(n19423), .A(n19389), .B(n19388), .ZN(
        P2_U3059) );
  AOI22_X1 U22369 ( .A1(n19395), .A2(n19815), .B1(n19394), .B2(n19814), .ZN(
        n19391) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19396), .B1(
        n19426), .B2(n19816), .ZN(n19390) );
  OAI211_X1 U22371 ( .C1(n19819), .C2(n19399), .A(n19391), .B(n19390), .ZN(
        P2_U3060) );
  AOI22_X1 U22372 ( .A1(n19395), .A2(n19821), .B1(n19394), .B2(n19820), .ZN(
        n19393) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19396), .B1(
        n19426), .B2(n19822), .ZN(n19392) );
  OAI211_X1 U22374 ( .C1(n19825), .C2(n19399), .A(n19393), .B(n19392), .ZN(
        P2_U3061) );
  AOI22_X1 U22375 ( .A1(n19395), .A2(n19827), .B1(n19394), .B2(n19826), .ZN(
        n19398) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19396), .B1(
        n19426), .B2(n19828), .ZN(n19397) );
  OAI211_X1 U22377 ( .C1(n19831), .C2(n19399), .A(n19398), .B(n19397), .ZN(
        P2_U3062) );
  INV_X1 U22378 ( .A(n19404), .ZN(n19401) );
  NAND2_X1 U22379 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19431), .ZN(
        n19438) );
  NOR2_X1 U22380 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19438), .ZN(
        n19424) );
  OAI21_X1 U22381 ( .B1(n19401), .B2(n19424), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19403) );
  INV_X1 U22382 ( .A(n19632), .ZN(n19402) );
  NAND2_X1 U22383 ( .A1(n19402), .A2(n19431), .ZN(n19405) );
  NAND2_X1 U22384 ( .A1(n19403), .A2(n19405), .ZN(n19425) );
  AOI22_X1 U22385 ( .A1(n19425), .A2(n19782), .B1(n19781), .B2(n19424), .ZN(
        n19410) );
  AOI21_X1 U22386 ( .B1(n19404), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19408) );
  OAI21_X1 U22387 ( .B1(n19450), .B2(n19426), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19406) );
  NAND3_X1 U22388 ( .A1(n19406), .A2(n19938), .A3(n19405), .ZN(n19407) );
  OAI211_X1 U22389 ( .C1(n19424), .C2(n19408), .A(n19407), .B(n19788), .ZN(
        n19427) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19427), .B1(
        n19426), .B2(n19695), .ZN(n19409) );
  OAI211_X1 U22391 ( .C1(n19698), .C2(n19460), .A(n19410), .B(n19409), .ZN(
        P2_U3064) );
  AOI22_X1 U22392 ( .A1(n19425), .A2(n19795), .B1(n19794), .B2(n19424), .ZN(
        n19412) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19427), .B1(
        n19426), .B2(n19796), .ZN(n19411) );
  OAI211_X1 U22394 ( .C1(n19801), .C2(n19460), .A(n19412), .B(n19411), .ZN(
        P2_U3065) );
  AOI22_X1 U22395 ( .A1(n19425), .A2(n19803), .B1(n19802), .B2(n19424), .ZN(
        n19414) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19427), .B1(
        n19450), .B2(n19804), .ZN(n19413) );
  OAI211_X1 U22397 ( .C1(n19807), .C2(n19423), .A(n19414), .B(n19413), .ZN(
        P2_U3066) );
  AOI22_X1 U22398 ( .A1(n19425), .A2(n19809), .B1(n19808), .B2(n19424), .ZN(
        n19416) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19427), .B1(
        n19450), .B2(n19810), .ZN(n19415) );
  OAI211_X1 U22400 ( .C1(n19813), .C2(n19423), .A(n19416), .B(n19415), .ZN(
        P2_U3067) );
  INV_X1 U22401 ( .A(n19816), .ZN(n19650) );
  AOI22_X1 U22402 ( .A1(n19425), .A2(n19815), .B1(n9731), .B2(n19424), .ZN(
        n19418) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19427), .B1(
        n19426), .B2(n19760), .ZN(n19417) );
  OAI211_X1 U22404 ( .C1(n19650), .C2(n19460), .A(n19418), .B(n19417), .ZN(
        P2_U3068) );
  AOI22_X1 U22405 ( .A1(n19425), .A2(n19821), .B1(n19820), .B2(n19424), .ZN(
        n19420) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19427), .B1(
        n19426), .B2(n19763), .ZN(n19419) );
  OAI211_X1 U22407 ( .C1(n19710), .C2(n19460), .A(n19420), .B(n19419), .ZN(
        P2_U3069) );
  AOI22_X1 U22408 ( .A1(n19425), .A2(n19827), .B1(n19826), .B2(n19424), .ZN(
        n19422) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19427), .B1(
        n19450), .B2(n19828), .ZN(n19421) );
  OAI211_X1 U22410 ( .C1(n19831), .C2(n19423), .A(n19422), .B(n19421), .ZN(
        P2_U3070) );
  INV_X1 U22411 ( .A(n19836), .ZN(n19681) );
  AOI22_X1 U22412 ( .A1(n19425), .A2(n19834), .B1(n19832), .B2(n19424), .ZN(
        n19429) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19427), .B1(
        n19426), .B2(n19770), .ZN(n19428) );
  OAI211_X1 U22414 ( .C1(n19681), .C2(n19460), .A(n19429), .B(n19428), .ZN(
        P2_U3071) );
  NAND2_X1 U22415 ( .A1(n19548), .A2(n19430), .ZN(n19480) );
  AND2_X1 U22416 ( .A1(n19537), .A2(n19431), .ZN(n19455) );
  AOI22_X1 U22417 ( .A1(n19450), .A2(n19695), .B1(n19781), .B2(n19455), .ZN(
        n19441) );
  OAI21_X1 U22418 ( .B1(n19542), .B2(n19939), .A(n19938), .ZN(n19439) );
  INV_X1 U22419 ( .A(n19438), .ZN(n19434) );
  INV_X1 U22420 ( .A(n19455), .ZN(n19432) );
  OAI211_X1 U22421 ( .C1(n19435), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19989), 
        .B(n19432), .ZN(n19433) );
  OAI211_X1 U22422 ( .C1(n19439), .C2(n19434), .A(n19788), .B(n19433), .ZN(
        n19457) );
  INV_X1 U22423 ( .A(n19435), .ZN(n19436) );
  OAI21_X1 U22424 ( .B1(n19436), .B2(n19455), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19437) );
  OAI21_X1 U22425 ( .B1(n19439), .B2(n19438), .A(n19437), .ZN(n19456) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19457), .B1(
        n19782), .B2(n19456), .ZN(n19440) );
  OAI211_X1 U22427 ( .C1(n19698), .C2(n19480), .A(n19441), .B(n19440), .ZN(
        P2_U3072) );
  AOI22_X1 U22428 ( .A1(n19450), .A2(n19796), .B1(n19455), .B2(n19794), .ZN(
        n19443) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19457), .B1(
        n19795), .B2(n19456), .ZN(n19442) );
  OAI211_X1 U22430 ( .C1(n19801), .C2(n19480), .A(n19443), .B(n19442), .ZN(
        P2_U3073) );
  AOI22_X1 U22431 ( .A1(n19804), .A2(n19490), .B1(n19455), .B2(n19802), .ZN(
        n19445) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19457), .B1(
        n19803), .B2(n19456), .ZN(n19444) );
  OAI211_X1 U22433 ( .C1(n19807), .C2(n19460), .A(n19445), .B(n19444), .ZN(
        P2_U3074) );
  AOI22_X1 U22434 ( .A1(n19757), .A2(n19450), .B1(n19455), .B2(n19808), .ZN(
        n19447) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19457), .B1(
        n19809), .B2(n19456), .ZN(n19446) );
  OAI211_X1 U22436 ( .C1(n19668), .C2(n19480), .A(n19447), .B(n19446), .ZN(
        P2_U3075) );
  AOI22_X1 U22437 ( .A1(n19816), .A2(n19490), .B1(n19455), .B2(n19814), .ZN(
        n19449) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19457), .B1(
        n19815), .B2(n19456), .ZN(n19448) );
  OAI211_X1 U22439 ( .C1(n19819), .C2(n19460), .A(n19449), .B(n19448), .ZN(
        P2_U3076) );
  AOI22_X1 U22440 ( .A1(n19763), .A2(n19450), .B1(n19820), .B2(n19455), .ZN(
        n19452) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19457), .B1(
        n19821), .B2(n19456), .ZN(n19451) );
  OAI211_X1 U22442 ( .C1(n19710), .C2(n19480), .A(n19452), .B(n19451), .ZN(
        P2_U3077) );
  AOI22_X1 U22443 ( .A1(n19490), .A2(n19828), .B1(n19826), .B2(n19455), .ZN(
        n19454) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19457), .B1(
        n19827), .B2(n19456), .ZN(n19453) );
  OAI211_X1 U22445 ( .C1(n19831), .C2(n19460), .A(n19454), .B(n19453), .ZN(
        P2_U3078) );
  AOI22_X1 U22446 ( .A1(n19836), .A2(n19490), .B1(n19832), .B2(n19455), .ZN(
        n19459) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19457), .B1(
        n19834), .B2(n19456), .ZN(n19458) );
  OAI211_X1 U22448 ( .C1(n19842), .C2(n19460), .A(n19459), .B(n19458), .ZN(
        P2_U3079) );
  NOR2_X1 U22449 ( .A1(n19684), .A2(n19461), .ZN(n19489) );
  AOI22_X1 U22450 ( .A1(n19490), .A2(n19695), .B1(n19781), .B2(n19489), .ZN(
        n19475) );
  OAI21_X1 U22451 ( .B1(n19490), .B2(n19511), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19462) );
  NAND2_X1 U22452 ( .A1(n19462), .A2(n19938), .ZN(n19473) );
  INV_X1 U22453 ( .A(n19463), .ZN(n19465) );
  NAND2_X1 U22454 ( .A1(n19465), .A2(n19464), .ZN(n19690) );
  NOR2_X1 U22455 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19690), .ZN(
        n19468) );
  INV_X1 U22456 ( .A(n19489), .ZN(n19466) );
  OAI211_X1 U22457 ( .C1(n19469), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19989), 
        .B(n19466), .ZN(n19467) );
  OAI211_X1 U22458 ( .C1(n19473), .C2(n19468), .A(n19788), .B(n19467), .ZN(
        n19492) );
  INV_X1 U22459 ( .A(n19468), .ZN(n19472) );
  INV_X1 U22460 ( .A(n19469), .ZN(n19470) );
  OAI21_X1 U22461 ( .B1(n19470), .B2(n19489), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19471) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19492), .B1(
        n19782), .B2(n19491), .ZN(n19474) );
  OAI211_X1 U22463 ( .C1(n19698), .C2(n19495), .A(n19475), .B(n19474), .ZN(
        P2_U3080) );
  AOI22_X1 U22464 ( .A1(n19490), .A2(n19796), .B1(n19489), .B2(n19794), .ZN(
        n19477) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19492), .B1(
        n19795), .B2(n19491), .ZN(n19476) );
  OAI211_X1 U22466 ( .C1(n19801), .C2(n19495), .A(n19477), .B(n19476), .ZN(
        P2_U3081) );
  AOI22_X1 U22467 ( .A1(n19804), .A2(n19511), .B1(n19802), .B2(n19489), .ZN(
        n19479) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19492), .B1(
        n19803), .B2(n19491), .ZN(n19478) );
  OAI211_X1 U22469 ( .C1(n19807), .C2(n19480), .A(n19479), .B(n19478), .ZN(
        P2_U3082) );
  AOI22_X1 U22470 ( .A1(n19490), .A2(n19757), .B1(n19489), .B2(n19808), .ZN(
        n19482) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19492), .B1(
        n19809), .B2(n19491), .ZN(n19481) );
  OAI211_X1 U22472 ( .C1(n19668), .C2(n19495), .A(n19482), .B(n19481), .ZN(
        P2_U3083) );
  AOI22_X1 U22473 ( .A1(n19490), .A2(n19760), .B1(n9731), .B2(n19489), .ZN(
        n19484) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19492), .B1(
        n19815), .B2(n19491), .ZN(n19483) );
  OAI211_X1 U22475 ( .C1(n19650), .C2(n19495), .A(n19484), .B(n19483), .ZN(
        P2_U3084) );
  AOI22_X1 U22476 ( .A1(n19763), .A2(n19490), .B1(n19820), .B2(n19489), .ZN(
        n19486) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19492), .B1(
        n19821), .B2(n19491), .ZN(n19485) );
  OAI211_X1 U22478 ( .C1(n19710), .C2(n19495), .A(n19486), .B(n19485), .ZN(
        P2_U3085) );
  INV_X1 U22479 ( .A(n19831), .ZN(n19766) );
  AOI22_X1 U22480 ( .A1(n19490), .A2(n19766), .B1(n19826), .B2(n19489), .ZN(
        n19488) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19492), .B1(
        n19827), .B2(n19491), .ZN(n19487) );
  OAI211_X1 U22482 ( .C1(n19529), .C2(n19495), .A(n19488), .B(n19487), .ZN(
        P2_U3086) );
  AOI22_X1 U22483 ( .A1(n19490), .A2(n19770), .B1(n19832), .B2(n19489), .ZN(
        n19494) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19492), .B1(
        n19834), .B2(n19491), .ZN(n19493) );
  OAI211_X1 U22485 ( .C1(n19681), .C2(n19495), .A(n19494), .B(n19493), .ZN(
        P2_U3087) );
  INV_X1 U22486 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19498) );
  AOI22_X1 U22487 ( .A1(n19532), .A2(n19750), .B1(n19510), .B2(n19794), .ZN(
        n19497) );
  AOI22_X1 U22488 ( .A1(n19795), .A2(n19512), .B1(n19511), .B2(n19796), .ZN(
        n19496) );
  OAI211_X1 U22489 ( .C1(n19515), .C2(n19498), .A(n19497), .B(n19496), .ZN(
        P2_U3089) );
  INV_X1 U22490 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19501) );
  AOI22_X1 U22491 ( .A1(n19511), .A2(n19753), .B1(n19510), .B2(n19802), .ZN(
        n19500) );
  AOI22_X1 U22492 ( .A1(n19803), .A2(n19512), .B1(n19532), .B2(n19804), .ZN(
        n19499) );
  OAI211_X1 U22493 ( .C1(n19515), .C2(n19501), .A(n19500), .B(n19499), .ZN(
        P2_U3090) );
  AOI22_X1 U22494 ( .A1(n19757), .A2(n19511), .B1(n19510), .B2(n19808), .ZN(
        n19503) );
  AOI22_X1 U22495 ( .A1(n19809), .A2(n19512), .B1(n19532), .B2(n19810), .ZN(
        n19502) );
  OAI211_X1 U22496 ( .C1(n19515), .C2(n10416), .A(n19503), .B(n19502), .ZN(
        P2_U3091) );
  AOI22_X1 U22497 ( .A1(n19532), .A2(n19816), .B1(n19510), .B2(n19814), .ZN(
        n19505) );
  AOI22_X1 U22498 ( .A1(n19815), .A2(n19512), .B1(n19511), .B2(n19760), .ZN(
        n19504) );
  OAI211_X1 U22499 ( .C1(n19515), .C2(n12840), .A(n19505), .B(n19504), .ZN(
        P2_U3092) );
  AOI22_X1 U22500 ( .A1(n19763), .A2(n19511), .B1(n19820), .B2(n19510), .ZN(
        n19507) );
  AOI22_X1 U22501 ( .A1(n19821), .A2(n19512), .B1(n19532), .B2(n19822), .ZN(
        n19506) );
  OAI211_X1 U22502 ( .C1(n19515), .C2(n10448), .A(n19507), .B(n19506), .ZN(
        P2_U3093) );
  AOI22_X1 U22503 ( .A1(n19766), .A2(n19511), .B1(n19826), .B2(n19510), .ZN(
        n19509) );
  AOI22_X1 U22504 ( .A1(n19827), .A2(n19512), .B1(n19532), .B2(n19828), .ZN(
        n19508) );
  OAI211_X1 U22505 ( .C1(n19515), .C2(n12872), .A(n19509), .B(n19508), .ZN(
        P2_U3094) );
  AOI22_X1 U22506 ( .A1(n19511), .A2(n19770), .B1(n19832), .B2(n19510), .ZN(
        n19514) );
  AOI22_X1 U22507 ( .A1(n19834), .A2(n19512), .B1(n19532), .B2(n19836), .ZN(
        n19513) );
  OAI211_X1 U22508 ( .C1(n19515), .C2(n13426), .A(n19514), .B(n19513), .ZN(
        P2_U3095) );
  AOI22_X1 U22509 ( .A1(n19531), .A2(n19795), .B1(n19794), .B2(n19530), .ZN(
        n19517) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19796), .ZN(n19516) );
  OAI211_X1 U22511 ( .C1(n19801), .C2(n19563), .A(n19517), .B(n19516), .ZN(
        P2_U3097) );
  AOI22_X1 U22512 ( .A1(n19531), .A2(n19803), .B1(n19802), .B2(n19530), .ZN(
        n19519) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19533), .B1(
        n19565), .B2(n19804), .ZN(n19518) );
  OAI211_X1 U22514 ( .C1(n19807), .C2(n19520), .A(n19519), .B(n19518), .ZN(
        P2_U3098) );
  AOI22_X1 U22515 ( .A1(n19531), .A2(n19809), .B1(n19808), .B2(n19530), .ZN(
        n19522) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19757), .ZN(n19521) );
  OAI211_X1 U22517 ( .C1(n19668), .C2(n19563), .A(n19522), .B(n19521), .ZN(
        P2_U3099) );
  AOI22_X1 U22518 ( .A1(n19531), .A2(n19815), .B1(n9731), .B2(n19530), .ZN(
        n19524) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19760), .ZN(n19523) );
  OAI211_X1 U22520 ( .C1(n19650), .C2(n19563), .A(n19524), .B(n19523), .ZN(
        P2_U3100) );
  AOI22_X1 U22521 ( .A1(n19531), .A2(n19821), .B1(n19820), .B2(n19530), .ZN(
        n19526) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19763), .ZN(n19525) );
  OAI211_X1 U22523 ( .C1(n19710), .C2(n19563), .A(n19526), .B(n19525), .ZN(
        P2_U3101) );
  AOI22_X1 U22524 ( .A1(n19531), .A2(n19827), .B1(n19826), .B2(n19530), .ZN(
        n19528) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19766), .ZN(n19527) );
  OAI211_X1 U22526 ( .C1(n19529), .C2(n19563), .A(n19528), .B(n19527), .ZN(
        P2_U3102) );
  AOI22_X1 U22527 ( .A1(n19531), .A2(n19834), .B1(n19832), .B2(n19530), .ZN(
        n19535) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19770), .ZN(n19534) );
  OAI211_X1 U22529 ( .C1(n19681), .C2(n19563), .A(n19535), .B(n19534), .ZN(
        P2_U3103) );
  NAND2_X1 U22530 ( .A1(n19537), .A2(n19536), .ZN(n19545) );
  INV_X1 U22531 ( .A(n19545), .ZN(n19573) );
  NOR3_X1 U22532 ( .A1(n19538), .A2(n19573), .A3(n19777), .ZN(n19541) );
  INV_X1 U22533 ( .A(n19544), .ZN(n19539) );
  AOI21_X1 U22534 ( .B1(n19986), .B2(n19539), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19540) );
  AOI22_X1 U22535 ( .A1(n19564), .A2(n19782), .B1(n19781), .B2(n19573), .ZN(
        n19550) );
  INV_X1 U22536 ( .A(n19541), .ZN(n19547) );
  OR2_X1 U22537 ( .A1(n19543), .A2(n19542), .ZN(n19944) );
  AOI22_X1 U22538 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19545), .B1(n19544), 
        .B2(n19944), .ZN(n19546) );
  NAND3_X1 U22539 ( .A1(n19547), .A2(n19546), .A3(n19788), .ZN(n19566) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19566), .B1(
        n19588), .B2(n19790), .ZN(n19549) );
  OAI211_X1 U22541 ( .C1(n19793), .C2(n19563), .A(n19550), .B(n19549), .ZN(
        P2_U3104) );
  AOI22_X1 U22542 ( .A1(n19564), .A2(n19795), .B1(n19573), .B2(n19794), .ZN(
        n19552) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19796), .ZN(n19551) );
  OAI211_X1 U22544 ( .C1(n19801), .C2(n19598), .A(n19552), .B(n19551), .ZN(
        P2_U3105) );
  AOI22_X1 U22545 ( .A1(n19564), .A2(n19803), .B1(n19573), .B2(n19802), .ZN(
        n19554) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19566), .B1(
        n19588), .B2(n19804), .ZN(n19553) );
  OAI211_X1 U22547 ( .C1(n19807), .C2(n19563), .A(n19554), .B(n19553), .ZN(
        P2_U3106) );
  AOI22_X1 U22548 ( .A1(n19564), .A2(n19809), .B1(n19573), .B2(n19808), .ZN(
        n19556) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19566), .B1(
        n19588), .B2(n19810), .ZN(n19555) );
  OAI211_X1 U22550 ( .C1(n19813), .C2(n19563), .A(n19556), .B(n19555), .ZN(
        P2_U3107) );
  AOI22_X1 U22551 ( .A1(n19564), .A2(n19815), .B1(n19573), .B2(n19814), .ZN(
        n19558) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19566), .B1(
        n19588), .B2(n19816), .ZN(n19557) );
  OAI211_X1 U22553 ( .C1(n19819), .C2(n19563), .A(n19558), .B(n19557), .ZN(
        P2_U3108) );
  AOI22_X1 U22554 ( .A1(n19564), .A2(n19821), .B1(n19820), .B2(n19573), .ZN(
        n19560) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19763), .ZN(n19559) );
  OAI211_X1 U22556 ( .C1(n19710), .C2(n19598), .A(n19560), .B(n19559), .ZN(
        P2_U3109) );
  AOI22_X1 U22557 ( .A1(n19564), .A2(n19827), .B1(n19826), .B2(n19573), .ZN(
        n19562) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19566), .B1(
        n19588), .B2(n19828), .ZN(n19561) );
  OAI211_X1 U22559 ( .C1(n19831), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3110) );
  AOI22_X1 U22560 ( .A1(n19564), .A2(n19834), .B1(n19832), .B2(n19573), .ZN(
        n19568) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19566), .B1(
        n19565), .B2(n19770), .ZN(n19567) );
  OAI211_X1 U22562 ( .C1(n19681), .C2(n19598), .A(n19568), .B(n19567), .ZN(
        P2_U3111) );
  NOR2_X1 U22563 ( .A1(n19684), .A2(n19633), .ZN(n19593) );
  AOI22_X1 U22564 ( .A1(n19617), .A2(n19790), .B1(n19781), .B2(n19593), .ZN(
        n19579) );
  NOR3_X1 U22565 ( .A1(n19617), .A2(n19588), .A3(n19989), .ZN(n19570) );
  NOR2_X1 U22566 ( .A1(n19570), .A2(n19941), .ZN(n19577) );
  NOR2_X1 U22567 ( .A1(n19577), .A2(n19573), .ZN(n19571) );
  AOI211_X1 U22568 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n10553), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19571), .ZN(n19572) );
  NOR2_X1 U22569 ( .A1(n19573), .A2(n19593), .ZN(n19576) );
  INV_X1 U22570 ( .A(n10553), .ZN(n19574) );
  OAI21_X1 U22571 ( .B1(n19574), .B2(n19593), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19575) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19595), .B1(
        n19782), .B2(n19594), .ZN(n19578) );
  OAI211_X1 U22573 ( .C1(n19793), .C2(n19598), .A(n19579), .B(n19578), .ZN(
        P2_U3112) );
  AOI22_X1 U22574 ( .A1(n19588), .A2(n19796), .B1(n19794), .B2(n19593), .ZN(
        n19581) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19795), .ZN(n19580) );
  OAI211_X1 U22576 ( .C1(n19801), .C2(n19629), .A(n19581), .B(n19580), .ZN(
        P2_U3113) );
  AOI22_X1 U22577 ( .A1(n19617), .A2(n19804), .B1(n19802), .B2(n19593), .ZN(
        n19583) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19803), .ZN(n19582) );
  OAI211_X1 U22579 ( .C1(n19807), .C2(n19598), .A(n19583), .B(n19582), .ZN(
        P2_U3114) );
  AOI22_X1 U22580 ( .A1(n19617), .A2(n19810), .B1(n19808), .B2(n19593), .ZN(
        n19585) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19809), .ZN(n19584) );
  OAI211_X1 U22582 ( .C1(n19813), .C2(n19598), .A(n19585), .B(n19584), .ZN(
        P2_U3115) );
  AOI22_X1 U22583 ( .A1(n19617), .A2(n19816), .B1(n9731), .B2(n19593), .ZN(
        n19587) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19815), .ZN(n19586) );
  OAI211_X1 U22585 ( .C1(n19819), .C2(n19598), .A(n19587), .B(n19586), .ZN(
        P2_U3116) );
  AOI22_X1 U22586 ( .A1(n19763), .A2(n19588), .B1(n19820), .B2(n19593), .ZN(
        n19590) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19821), .ZN(n19589) );
  OAI211_X1 U22588 ( .C1(n19710), .C2(n19629), .A(n19590), .B(n19589), .ZN(
        P2_U3117) );
  AOI22_X1 U22589 ( .A1(n19617), .A2(n19828), .B1(n19826), .B2(n19593), .ZN(
        n19592) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19827), .ZN(n19591) );
  OAI211_X1 U22591 ( .C1(n19831), .C2(n19598), .A(n19592), .B(n19591), .ZN(
        P2_U3118) );
  AOI22_X1 U22592 ( .A1(n19617), .A2(n19836), .B1(n19832), .B2(n19593), .ZN(
        n19597) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19595), .B1(
        n19594), .B2(n19834), .ZN(n19596) );
  OAI211_X1 U22594 ( .C1(n19842), .C2(n19598), .A(n19597), .B(n19596), .ZN(
        P2_U3119) );
  NOR2_X1 U22595 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19633), .ZN(
        n19604) );
  NAND2_X1 U22596 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19604), .ZN(
        n19634) );
  INV_X1 U22597 ( .A(n19634), .ZN(n19624) );
  AOI22_X1 U22598 ( .A1(n19790), .A2(n19651), .B1(n19781), .B2(n19624), .ZN(
        n19610) );
  OAI21_X1 U22599 ( .B1(n19722), .B2(n19600), .A(n19938), .ZN(n19608) );
  INV_X1 U22600 ( .A(n10540), .ZN(n19605) );
  OAI21_X1 U22601 ( .B1(n19605), .B2(n19777), .A(n19986), .ZN(n19602) );
  AOI21_X1 U22602 ( .B1(n19602), .B2(n19634), .A(n19601), .ZN(n19603) );
  OAI21_X1 U22603 ( .B1(n19608), .B2(n19604), .A(n19603), .ZN(n19626) );
  INV_X1 U22604 ( .A(n19604), .ZN(n19607) );
  OAI21_X1 U22605 ( .B1(n19605), .B2(n19624), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19606) );
  OAI21_X1 U22606 ( .B1(n19608), .B2(n19607), .A(n19606), .ZN(n19625) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19626), .B1(
        n19782), .B2(n19625), .ZN(n19609) );
  OAI211_X1 U22608 ( .C1(n19793), .C2(n19629), .A(n19610), .B(n19609), .ZN(
        P2_U3120) );
  AOI22_X1 U22609 ( .A1(n19617), .A2(n19796), .B1(n19794), .B2(n19624), .ZN(
        n19612) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19626), .B1(
        n19795), .B2(n19625), .ZN(n19611) );
  OAI211_X1 U22611 ( .C1(n19801), .C2(n19661), .A(n19612), .B(n19611), .ZN(
        P2_U3121) );
  AOI22_X1 U22612 ( .A1(n19804), .A2(n19651), .B1(n19802), .B2(n19624), .ZN(
        n19614) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19626), .B1(
        n19803), .B2(n19625), .ZN(n19613) );
  OAI211_X1 U22614 ( .C1(n19807), .C2(n19629), .A(n19614), .B(n19613), .ZN(
        P2_U3122) );
  AOI22_X1 U22615 ( .A1(n19810), .A2(n19651), .B1(n19808), .B2(n19624), .ZN(
        n19616) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19626), .B1(
        n19809), .B2(n19625), .ZN(n19615) );
  OAI211_X1 U22617 ( .C1(n19813), .C2(n19629), .A(n19616), .B(n19615), .ZN(
        P2_U3123) );
  AOI22_X1 U22618 ( .A1(n19617), .A2(n19760), .B1(n9731), .B2(n19624), .ZN(
        n19619) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19626), .B1(
        n19815), .B2(n19625), .ZN(n19618) );
  OAI211_X1 U22620 ( .C1(n19650), .C2(n19661), .A(n19619), .B(n19618), .ZN(
        P2_U3124) );
  AOI22_X1 U22621 ( .A1(n19822), .A2(n19651), .B1(n19820), .B2(n19624), .ZN(
        n19621) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19626), .B1(
        n19821), .B2(n19625), .ZN(n19620) );
  OAI211_X1 U22623 ( .C1(n19825), .C2(n19629), .A(n19621), .B(n19620), .ZN(
        P2_U3125) );
  AOI22_X1 U22624 ( .A1(n19651), .A2(n19828), .B1(n19826), .B2(n19624), .ZN(
        n19623) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19626), .B1(
        n19827), .B2(n19625), .ZN(n19622) );
  OAI211_X1 U22626 ( .C1(n19831), .C2(n19629), .A(n19623), .B(n19622), .ZN(
        P2_U3126) );
  AOI22_X1 U22627 ( .A1(n19836), .A2(n19651), .B1(n19832), .B2(n19624), .ZN(
        n19628) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19626), .B1(
        n19834), .B2(n19625), .ZN(n19627) );
  OAI211_X1 U22629 ( .C1(n19842), .C2(n19629), .A(n19628), .B(n19627), .ZN(
        P2_U3127) );
  NOR3_X2 U22630 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10498), .A3(
        n19633), .ZN(n19656) );
  OAI21_X1 U22631 ( .B1(n10443), .B2(n19656), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19631) );
  OAI21_X1 U22632 ( .B1(n19633), .B2(n19632), .A(n19631), .ZN(n19657) );
  AOI22_X1 U22633 ( .A1(n19657), .A2(n19782), .B1(n19781), .B2(n19656), .ZN(
        n19641) );
  OAI21_X1 U22634 ( .B1(n19677), .B2(n19651), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19635) );
  AOI21_X1 U22635 ( .B1(n19635), .B2(n19634), .A(n19989), .ZN(n19639) );
  NAND3_X1 U22636 ( .A1(n10443), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19950), 
        .ZN(n19637) );
  INV_X1 U22637 ( .A(n19656), .ZN(n19636) );
  NAND2_X1 U22638 ( .A1(n19637), .A2(n19636), .ZN(n19638) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19658), .B1(
        n19651), .B2(n19695), .ZN(n19640) );
  OAI211_X1 U22640 ( .C1(n19698), .C2(n19671), .A(n19641), .B(n19640), .ZN(
        P2_U3128) );
  AOI22_X1 U22641 ( .A1(n19657), .A2(n19795), .B1(n19794), .B2(n19656), .ZN(
        n19643) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19658), .B1(
        n19651), .B2(n19796), .ZN(n19642) );
  OAI211_X1 U22643 ( .C1(n19801), .C2(n19671), .A(n19643), .B(n19642), .ZN(
        P2_U3129) );
  AOI22_X1 U22644 ( .A1(n19657), .A2(n19803), .B1(n19802), .B2(n19656), .ZN(
        n19645) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19658), .B1(
        n19677), .B2(n19804), .ZN(n19644) );
  OAI211_X1 U22646 ( .C1(n19807), .C2(n19661), .A(n19645), .B(n19644), .ZN(
        P2_U3130) );
  AOI22_X1 U22647 ( .A1(n19657), .A2(n19809), .B1(n19808), .B2(n19656), .ZN(
        n19647) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19658), .B1(
        n19677), .B2(n19810), .ZN(n19646) );
  OAI211_X1 U22649 ( .C1(n19813), .C2(n19661), .A(n19647), .B(n19646), .ZN(
        P2_U3131) );
  AOI22_X1 U22650 ( .A1(n19657), .A2(n19815), .B1(n9731), .B2(n19656), .ZN(
        n19649) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19658), .B1(
        n19651), .B2(n19760), .ZN(n19648) );
  OAI211_X1 U22652 ( .C1(n19650), .C2(n19671), .A(n19649), .B(n19648), .ZN(
        P2_U3132) );
  AOI22_X1 U22653 ( .A1(n19657), .A2(n19821), .B1(n19820), .B2(n19656), .ZN(
        n19653) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19658), .B1(
        n19651), .B2(n19763), .ZN(n19652) );
  OAI211_X1 U22655 ( .C1(n19710), .C2(n19671), .A(n19653), .B(n19652), .ZN(
        P2_U3133) );
  AOI22_X1 U22656 ( .A1(n19657), .A2(n19827), .B1(n19826), .B2(n19656), .ZN(
        n19655) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19658), .B1(
        n19677), .B2(n19828), .ZN(n19654) );
  OAI211_X1 U22658 ( .C1(n19831), .C2(n19661), .A(n19655), .B(n19654), .ZN(
        P2_U3134) );
  AOI22_X1 U22659 ( .A1(n19657), .A2(n19834), .B1(n19832), .B2(n19656), .ZN(
        n19660) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19658), .B1(
        n19677), .B2(n19836), .ZN(n19659) );
  OAI211_X1 U22661 ( .C1(n19842), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P2_U3135) );
  AOI22_X1 U22662 ( .A1(n19676), .A2(n19795), .B1(n19675), .B2(n19794), .ZN(
        n19663) );
  INV_X1 U22663 ( .A(n19674), .ZN(n19678) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19796), .ZN(n19662) );
  OAI211_X1 U22665 ( .C1(n19801), .C2(n19718), .A(n19663), .B(n19662), .ZN(
        P2_U3137) );
  AOI22_X1 U22666 ( .A1(n19803), .A2(n19676), .B1(n19675), .B2(n19802), .ZN(
        n19665) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19678), .B1(
        n19707), .B2(n19804), .ZN(n19664) );
  OAI211_X1 U22668 ( .C1(n19807), .C2(n19671), .A(n19665), .B(n19664), .ZN(
        P2_U3138) );
  AOI22_X1 U22669 ( .A1(n19676), .A2(n19809), .B1(n19675), .B2(n19808), .ZN(
        n19667) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19757), .ZN(n19666) );
  OAI211_X1 U22671 ( .C1(n19668), .C2(n19718), .A(n19667), .B(n19666), .ZN(
        P2_U3139) );
  AOI22_X1 U22672 ( .A1(n19815), .A2(n19676), .B1(n19675), .B2(n19814), .ZN(
        n19670) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19678), .B1(
        n19707), .B2(n19816), .ZN(n19669) );
  OAI211_X1 U22674 ( .C1(n19819), .C2(n19671), .A(n19670), .B(n19669), .ZN(
        P2_U3140) );
  AOI22_X1 U22675 ( .A1(n19827), .A2(n19676), .B1(n19675), .B2(n19826), .ZN(
        n19673) );
  AOI22_X1 U22676 ( .A1(n19707), .A2(n19828), .B1(n19677), .B2(n19766), .ZN(
        n19672) );
  OAI211_X1 U22677 ( .C1(n19674), .C2(n13062), .A(n19673), .B(n19672), .ZN(
        P2_U3142) );
  AOI22_X1 U22678 ( .A1(n19676), .A2(n19834), .B1(n19832), .B2(n19675), .ZN(
        n19680) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19678), .B1(
        n19677), .B2(n19770), .ZN(n19679) );
  OAI211_X1 U22680 ( .C1(n19681), .C2(n19718), .A(n19680), .B(n19679), .ZN(
        P2_U3143) );
  INV_X1 U22681 ( .A(n19683), .ZN(n19688) );
  INV_X1 U22682 ( .A(n19692), .ZN(n19686) );
  INV_X1 U22683 ( .A(n19719), .ZN(n19685) );
  NOR2_X1 U22684 ( .A1(n19685), .A2(n19684), .ZN(n19713) );
  OAI21_X1 U22685 ( .B1(n19686), .B2(n19713), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19687) );
  OAI21_X1 U22686 ( .B1(n19688), .B2(n19690), .A(n19687), .ZN(n19714) );
  AOI22_X1 U22687 ( .A1(n19714), .A2(n19782), .B1(n19781), .B2(n19713), .ZN(
        n19697) );
  OAI21_X1 U22688 ( .B1(n19707), .B2(n19730), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19689) );
  OAI21_X1 U22689 ( .B1(n19690), .B2(n12752), .A(n19689), .ZN(n19694) );
  INV_X1 U22690 ( .A(n19713), .ZN(n19691) );
  OAI211_X1 U22691 ( .C1(n19692), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19989), 
        .B(n19691), .ZN(n19693) );
  NAND3_X1 U22692 ( .A1(n19694), .A2(n19788), .A3(n19693), .ZN(n19715) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19715), .B1(
        n19707), .B2(n19695), .ZN(n19696) );
  OAI211_X1 U22694 ( .C1(n19698), .C2(n19749), .A(n19697), .B(n19696), .ZN(
        P2_U3144) );
  AOI22_X1 U22695 ( .A1(n19714), .A2(n19795), .B1(n19794), .B2(n19713), .ZN(
        n19700) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19715), .B1(
        n19707), .B2(n19796), .ZN(n19699) );
  OAI211_X1 U22697 ( .C1(n19801), .C2(n19749), .A(n19700), .B(n19699), .ZN(
        P2_U3145) );
  AOI22_X1 U22698 ( .A1(n19714), .A2(n19803), .B1(n19802), .B2(n19713), .ZN(
        n19702) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19715), .B1(
        n19730), .B2(n19804), .ZN(n19701) );
  OAI211_X1 U22700 ( .C1(n19807), .C2(n19718), .A(n19702), .B(n19701), .ZN(
        P2_U3146) );
  AOI22_X1 U22701 ( .A1(n19714), .A2(n19809), .B1(n19808), .B2(n19713), .ZN(
        n19704) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19715), .B1(
        n19730), .B2(n19810), .ZN(n19703) );
  OAI211_X1 U22703 ( .C1(n19813), .C2(n19718), .A(n19704), .B(n19703), .ZN(
        P2_U3147) );
  AOI22_X1 U22704 ( .A1(n19714), .A2(n19815), .B1(n9731), .B2(n19713), .ZN(
        n19706) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19715), .B1(
        n19730), .B2(n19816), .ZN(n19705) );
  OAI211_X1 U22706 ( .C1(n19819), .C2(n19718), .A(n19706), .B(n19705), .ZN(
        P2_U3148) );
  AOI22_X1 U22707 ( .A1(n19714), .A2(n19821), .B1(n19820), .B2(n19713), .ZN(
        n19709) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19715), .B1(
        n19707), .B2(n19763), .ZN(n19708) );
  OAI211_X1 U22709 ( .C1(n19710), .C2(n19749), .A(n19709), .B(n19708), .ZN(
        P2_U3149) );
  AOI22_X1 U22710 ( .A1(n19714), .A2(n19827), .B1(n19826), .B2(n19713), .ZN(
        n19712) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19715), .B1(
        n19730), .B2(n19828), .ZN(n19711) );
  OAI211_X1 U22712 ( .C1(n19831), .C2(n19718), .A(n19712), .B(n19711), .ZN(
        P2_U3150) );
  AOI22_X1 U22713 ( .A1(n19714), .A2(n19834), .B1(n19832), .B2(n19713), .ZN(
        n19717) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19715), .B1(
        n19730), .B2(n19836), .ZN(n19716) );
  OAI211_X1 U22715 ( .C1(n19842), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3151) );
  NAND2_X1 U22716 ( .A1(n19719), .A2(n10498), .ZN(n19725) );
  INV_X1 U22717 ( .A(n10550), .ZN(n19720) );
  NOR2_X1 U22718 ( .A1(n19973), .A2(n19725), .ZN(n19744) );
  NOR3_X1 U22719 ( .A1(n19720), .A2(n19744), .A3(n19777), .ZN(n19724) );
  AOI211_X2 U22720 ( .C1(n19725), .C2(n19777), .A(n19721), .B(n19724), .ZN(
        n19745) );
  AOI22_X1 U22721 ( .A1(n19745), .A2(n19782), .B1(n19781), .B2(n19744), .ZN(
        n19729) );
  INV_X1 U22722 ( .A(n19722), .ZN(n19784) );
  NAND2_X1 U22723 ( .A1(n19784), .A2(n19723), .ZN(n19726) );
  AOI21_X1 U22724 ( .B1(n19726), .B2(n19725), .A(n19724), .ZN(n19727) );
  OAI211_X1 U22725 ( .C1(n19744), .C2(n19950), .A(n19727), .B(n19788), .ZN(
        n19746) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19746), .B1(
        n19771), .B2(n19790), .ZN(n19728) );
  OAI211_X1 U22727 ( .C1(n19793), .C2(n19749), .A(n19729), .B(n19728), .ZN(
        P2_U3152) );
  INV_X1 U22728 ( .A(n19771), .ZN(n19733) );
  AOI22_X1 U22729 ( .A1(n19745), .A2(n19795), .B1(n19794), .B2(n19744), .ZN(
        n19732) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19746), .B1(
        n19730), .B2(n19796), .ZN(n19731) );
  OAI211_X1 U22731 ( .C1(n19801), .C2(n19733), .A(n19732), .B(n19731), .ZN(
        P2_U3153) );
  AOI22_X1 U22732 ( .A1(n19745), .A2(n19803), .B1(n19802), .B2(n19744), .ZN(
        n19735) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19746), .B1(
        n19771), .B2(n19804), .ZN(n19734) );
  OAI211_X1 U22734 ( .C1(n19807), .C2(n19749), .A(n19735), .B(n19734), .ZN(
        P2_U3154) );
  AOI22_X1 U22735 ( .A1(n19745), .A2(n19809), .B1(n19808), .B2(n19744), .ZN(
        n19737) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19746), .B1(
        n19771), .B2(n19810), .ZN(n19736) );
  OAI211_X1 U22737 ( .C1(n19813), .C2(n19749), .A(n19737), .B(n19736), .ZN(
        P2_U3155) );
  AOI22_X1 U22738 ( .A1(n19745), .A2(n19815), .B1(n9731), .B2(n19744), .ZN(
        n19739) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19746), .B1(
        n19771), .B2(n19816), .ZN(n19738) );
  OAI211_X1 U22740 ( .C1(n19819), .C2(n19749), .A(n19739), .B(n19738), .ZN(
        P2_U3156) );
  AOI22_X1 U22741 ( .A1(n19745), .A2(n19821), .B1(n19820), .B2(n19744), .ZN(
        n19741) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19746), .B1(
        n19771), .B2(n19822), .ZN(n19740) );
  OAI211_X1 U22743 ( .C1(n19825), .C2(n19749), .A(n19741), .B(n19740), .ZN(
        P2_U3157) );
  AOI22_X1 U22744 ( .A1(n19745), .A2(n19827), .B1(n19826), .B2(n19744), .ZN(
        n19743) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19746), .B1(
        n19771), .B2(n19828), .ZN(n19742) );
  OAI211_X1 U22746 ( .C1(n19831), .C2(n19749), .A(n19743), .B(n19742), .ZN(
        P2_U3158) );
  AOI22_X1 U22747 ( .A1(n19745), .A2(n19834), .B1(n19832), .B2(n19744), .ZN(
        n19748) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19746), .B1(
        n19771), .B2(n19836), .ZN(n19747) );
  OAI211_X1 U22749 ( .C1(n19842), .C2(n19749), .A(n19748), .B(n19747), .ZN(
        P2_U3159) );
  AOI22_X1 U22750 ( .A1(n19771), .A2(n19796), .B1(n19769), .B2(n19794), .ZN(
        n19752) );
  AOI22_X1 U22751 ( .A1(n19795), .A2(n19772), .B1(n19797), .B2(n19750), .ZN(
        n19751) );
  OAI211_X1 U22752 ( .C1(n19775), .C2(n10363), .A(n19752), .B(n19751), .ZN(
        P2_U3161) );
  AOI22_X1 U22753 ( .A1(n19753), .A2(n19771), .B1(n19769), .B2(n19802), .ZN(
        n19755) );
  AOI22_X1 U22754 ( .A1(n19803), .A2(n19772), .B1(n19797), .B2(n19804), .ZN(
        n19754) );
  OAI211_X1 U22755 ( .C1(n19775), .C2(n19756), .A(n19755), .B(n19754), .ZN(
        P2_U3162) );
  AOI22_X1 U22756 ( .A1(n19757), .A2(n19771), .B1(n19769), .B2(n19808), .ZN(
        n19759) );
  AOI22_X1 U22757 ( .A1(n19809), .A2(n19772), .B1(n19797), .B2(n19810), .ZN(
        n19758) );
  OAI211_X1 U22758 ( .C1(n19775), .C2(n10409), .A(n19759), .B(n19758), .ZN(
        P2_U3163) );
  AOI22_X1 U22759 ( .A1(n19760), .A2(n19771), .B1(n19769), .B2(n19814), .ZN(
        n19762) );
  AOI22_X1 U22760 ( .A1(n19815), .A2(n19772), .B1(n19797), .B2(n19816), .ZN(
        n19761) );
  OAI211_X1 U22761 ( .C1(n19775), .C2(n12849), .A(n19762), .B(n19761), .ZN(
        P2_U3164) );
  AOI22_X1 U22762 ( .A1(n19763), .A2(n19771), .B1(n19820), .B2(n19769), .ZN(
        n19765) );
  AOI22_X1 U22763 ( .A1(n19821), .A2(n19772), .B1(n19797), .B2(n19822), .ZN(
        n19764) );
  OAI211_X1 U22764 ( .C1(n19775), .C2(n10453), .A(n19765), .B(n19764), .ZN(
        P2_U3165) );
  AOI22_X1 U22765 ( .A1(n19766), .A2(n19771), .B1(n19769), .B2(n19826), .ZN(
        n19768) );
  AOI22_X1 U22766 ( .A1(n19827), .A2(n19772), .B1(n19797), .B2(n19828), .ZN(
        n19767) );
  OAI211_X1 U22767 ( .C1(n19775), .C2(n12881), .A(n19768), .B(n19767), .ZN(
        P2_U3166) );
  AOI22_X1 U22768 ( .A1(n19797), .A2(n19836), .B1(n19832), .B2(n19769), .ZN(
        n19774) );
  AOI22_X1 U22769 ( .A1(n19834), .A2(n19772), .B1(n19771), .B2(n19770), .ZN(
        n19773) );
  OAI211_X1 U22770 ( .C1(n19775), .C2(n11129), .A(n19774), .B(n19773), .ZN(
        P2_U3167) );
  INV_X1 U22771 ( .A(n19776), .ZN(n19778) );
  NOR3_X1 U22772 ( .A1(n19778), .A2(n19833), .A3(n19777), .ZN(n19785) );
  INV_X1 U22773 ( .A(n19786), .ZN(n19779) );
  AOI21_X1 U22774 ( .B1(n19986), .B2(n19779), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19780) );
  NOR2_X1 U22775 ( .A1(n19785), .A2(n19780), .ZN(n19835) );
  AOI22_X1 U22776 ( .A1(n19835), .A2(n19782), .B1(n19833), .B2(n19781), .ZN(
        n19792) );
  NAND2_X1 U22777 ( .A1(n19784), .A2(n19783), .ZN(n19787) );
  AOI21_X1 U22778 ( .B1(n19787), .B2(n19786), .A(n19785), .ZN(n19789) );
  OAI211_X1 U22779 ( .C1(n19833), .C2(n19950), .A(n19789), .B(n19788), .ZN(
        n19838) );
  AOI22_X1 U22780 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19838), .B1(
        n19837), .B2(n19790), .ZN(n19791) );
  OAI211_X1 U22781 ( .C1(n19793), .C2(n19841), .A(n19792), .B(n19791), .ZN(
        P2_U3168) );
  AOI22_X1 U22782 ( .A1(n19835), .A2(n19795), .B1(n19833), .B2(n19794), .ZN(
        n19799) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19838), .B1(
        n19797), .B2(n19796), .ZN(n19798) );
  OAI211_X1 U22784 ( .C1(n19801), .C2(n19800), .A(n19799), .B(n19798), .ZN(
        P2_U3169) );
  AOI22_X1 U22785 ( .A1(n19835), .A2(n19803), .B1(n19833), .B2(n19802), .ZN(
        n19806) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19838), .B1(
        n19837), .B2(n19804), .ZN(n19805) );
  OAI211_X1 U22787 ( .C1(n19807), .C2(n19841), .A(n19806), .B(n19805), .ZN(
        P2_U3170) );
  AOI22_X1 U22788 ( .A1(n19835), .A2(n19809), .B1(n19833), .B2(n19808), .ZN(
        n19812) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19838), .B1(
        n19837), .B2(n19810), .ZN(n19811) );
  OAI211_X1 U22790 ( .C1(n19813), .C2(n19841), .A(n19812), .B(n19811), .ZN(
        P2_U3171) );
  AOI22_X1 U22791 ( .A1(n19835), .A2(n19815), .B1(n19833), .B2(n19814), .ZN(
        n19818) );
  AOI22_X1 U22792 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19838), .B1(
        n19837), .B2(n19816), .ZN(n19817) );
  OAI211_X1 U22793 ( .C1(n19819), .C2(n19841), .A(n19818), .B(n19817), .ZN(
        P2_U3172) );
  AOI22_X1 U22794 ( .A1(n19835), .A2(n19821), .B1(n19833), .B2(n19820), .ZN(
        n19824) );
  AOI22_X1 U22795 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19838), .B1(
        n19837), .B2(n19822), .ZN(n19823) );
  OAI211_X1 U22796 ( .C1(n19825), .C2(n19841), .A(n19824), .B(n19823), .ZN(
        P2_U3173) );
  AOI22_X1 U22797 ( .A1(n19835), .A2(n19827), .B1(n19833), .B2(n19826), .ZN(
        n19830) );
  AOI22_X1 U22798 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19838), .B1(
        n19837), .B2(n19828), .ZN(n19829) );
  OAI211_X1 U22799 ( .C1(n19831), .C2(n19841), .A(n19830), .B(n19829), .ZN(
        P2_U3174) );
  AOI22_X1 U22800 ( .A1(n19835), .A2(n19834), .B1(n19833), .B2(n19832), .ZN(
        n19840) );
  AOI22_X1 U22801 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19838), .B1(
        n19837), .B2(n19836), .ZN(n19839) );
  OAI211_X1 U22802 ( .C1(n19842), .C2(n19841), .A(n19840), .B(n19839), .ZN(
        P2_U3175) );
  AOI21_X1 U22803 ( .B1(n19940), .B2(n19844), .A(n19843), .ZN(n19848) );
  NOR2_X1 U22804 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13085), .ZN(n19845) );
  OAI211_X1 U22805 ( .C1(n19849), .C2(n19845), .A(n19864), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19846) );
  OAI211_X1 U22806 ( .C1(n19849), .C2(n19848), .A(n19847), .B(n19846), .ZN(
        P2_U3177) );
  AND2_X1 U22807 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19850), .ZN(
        P2_U3179) );
  AND2_X1 U22808 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19850), .ZN(
        P2_U3180) );
  AND2_X1 U22809 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19850), .ZN(
        P2_U3181) );
  AND2_X1 U22810 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19850), .ZN(
        P2_U3182) );
  AND2_X1 U22811 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19850), .ZN(
        P2_U3183) );
  AND2_X1 U22812 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19850), .ZN(
        P2_U3184) );
  AND2_X1 U22813 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19850), .ZN(
        P2_U3185) );
  AND2_X1 U22814 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19850), .ZN(
        P2_U3186) );
  AND2_X1 U22815 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19850), .ZN(
        P2_U3187) );
  AND2_X1 U22816 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19850), .ZN(
        P2_U3188) );
  AND2_X1 U22817 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19850), .ZN(
        P2_U3189) );
  AND2_X1 U22818 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19850), .ZN(
        P2_U3190) );
  AND2_X1 U22819 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19850), .ZN(
        P2_U3191) );
  AND2_X1 U22820 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19850), .ZN(
        P2_U3192) );
  AND2_X1 U22821 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19850), .ZN(
        P2_U3193) );
  AND2_X1 U22822 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19850), .ZN(
        P2_U3194) );
  AND2_X1 U22823 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19850), .ZN(
        P2_U3195) );
  AND2_X1 U22824 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19850), .ZN(
        P2_U3196) );
  AND2_X1 U22825 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19850), .ZN(
        P2_U3197) );
  AND2_X1 U22826 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19850), .ZN(
        P2_U3198) );
  AND2_X1 U22827 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19850), .ZN(
        P2_U3199) );
  AND2_X1 U22828 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19850), .ZN(
        P2_U3200) );
  AND2_X1 U22829 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19850), .ZN(P2_U3201) );
  AND2_X1 U22830 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19850), .ZN(P2_U3202) );
  AND2_X1 U22831 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19850), .ZN(P2_U3203) );
  AND2_X1 U22832 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19850), .ZN(P2_U3204) );
  AND2_X1 U22833 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19850), .ZN(P2_U3205) );
  AND2_X1 U22834 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19850), .ZN(P2_U3206) );
  AND2_X1 U22835 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19850), .ZN(P2_U3207) );
  AND2_X1 U22836 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19850), .ZN(P2_U3208) );
  NOR2_X1 U22837 ( .A1(n19851), .A2(n19993), .ZN(n19865) );
  INV_X1 U22838 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20003) );
  OR3_X1 U22839 ( .A1(n19865), .A2(n20003), .A3(n19852), .ZN(n19854) );
  AOI211_X1 U22840 ( .C1(n19861), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19866), .B(n19916), .ZN(n19853) );
  INV_X1 U22841 ( .A(NA), .ZN(n20852) );
  NOR2_X1 U22842 ( .A1(n20852), .A2(n19856), .ZN(n19871) );
  AOI211_X1 U22843 ( .C1(n19872), .C2(n19854), .A(n19853), .B(n19871), .ZN(
        n19855) );
  INV_X1 U22844 ( .A(n19855), .ZN(P2_U3209) );
  AOI21_X1 U22845 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19861), .A(n19872), 
        .ZN(n19862) );
  NOR2_X1 U22846 ( .A1(n20003), .A2(n19862), .ZN(n19857) );
  AOI21_X1 U22847 ( .B1(n19857), .B2(n19856), .A(n19865), .ZN(n19859) );
  OAI211_X1 U22848 ( .C1(n19861), .C2(n19860), .A(n19859), .B(n19858), .ZN(
        P2_U3210) );
  AOI21_X1 U22849 ( .B1(n19864), .B2(n19863), .A(n19862), .ZN(n19870) );
  AOI22_X1 U22850 ( .A1(n20003), .A2(n19866), .B1(n20852), .B2(n19865), .ZN(
        n19867) );
  INV_X1 U22851 ( .A(n19867), .ZN(n19868) );
  OAI211_X1 U22852 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19868), .ZN(n19869) );
  OAI21_X1 U22853 ( .B1(n19871), .B2(n19870), .A(n19869), .ZN(P2_U3211) );
  NAND2_X1 U22854 ( .A1(n19916), .A2(n19872), .ZN(n19927) );
  CLKBUF_X1 U22855 ( .A(n19927), .Z(n19923) );
  OAI222_X1 U22856 ( .A1(n19924), .A2(n19874), .B1(n19873), .B2(n19916), .C1(
        n10267), .C2(n19923), .ZN(P2_U3212) );
  OAI222_X1 U22857 ( .A1(n19924), .A2(n10267), .B1(n19875), .B2(n19916), .C1(
        n13921), .C2(n19923), .ZN(P2_U3213) );
  OAI222_X1 U22858 ( .A1(n19924), .A2(n13921), .B1(n19876), .B2(n19916), .C1(
        n19877), .C2(n19923), .ZN(P2_U3214) );
  OAI222_X1 U22859 ( .A1(n19923), .A2(n10832), .B1(n19878), .B2(n19916), .C1(
        n19877), .C2(n19924), .ZN(P2_U3215) );
  OAI222_X1 U22860 ( .A1(n19927), .A2(n19880), .B1(n19879), .B2(n19916), .C1(
        n10832), .C2(n19924), .ZN(P2_U3216) );
  OAI222_X1 U22861 ( .A1(n19927), .A2(n19882), .B1(n19881), .B2(n19916), .C1(
        n19880), .C2(n19924), .ZN(P2_U3217) );
  OAI222_X1 U22862 ( .A1(n19927), .A2(n19884), .B1(n19883), .B2(n19916), .C1(
        n19882), .C2(n19924), .ZN(P2_U3218) );
  OAI222_X1 U22863 ( .A1(n19927), .A2(n15253), .B1(n19885), .B2(n19916), .C1(
        n19884), .C2(n19924), .ZN(P2_U3219) );
  INV_X1 U22864 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19887) );
  OAI222_X1 U22865 ( .A1(n19927), .A2(n19887), .B1(n19886), .B2(n19916), .C1(
        n15253), .C2(n19924), .ZN(P2_U3220) );
  OAI222_X1 U22866 ( .A1(n19923), .A2(n19889), .B1(n19888), .B2(n19916), .C1(
        n19887), .C2(n19924), .ZN(P2_U3221) );
  OAI222_X1 U22867 ( .A1(n19923), .A2(n19890), .B1(n20959), .B2(n19916), .C1(
        n19889), .C2(n19924), .ZN(P2_U3222) );
  OAI222_X1 U22868 ( .A1(n19923), .A2(n19892), .B1(n19891), .B2(n19916), .C1(
        n19890), .C2(n19924), .ZN(P2_U3223) );
  INV_X1 U22869 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19894) );
  OAI222_X1 U22870 ( .A1(n19923), .A2(n19894), .B1(n19893), .B2(n19916), .C1(
        n19892), .C2(n19924), .ZN(P2_U3224) );
  OAI222_X1 U22871 ( .A1(n19923), .A2(n19896), .B1(n19895), .B2(n19916), .C1(
        n19894), .C2(n19924), .ZN(P2_U3225) );
  OAI222_X1 U22872 ( .A1(n19923), .A2(n19898), .B1(n19897), .B2(n19916), .C1(
        n19896), .C2(n19924), .ZN(P2_U3226) );
  OAI222_X1 U22873 ( .A1(n19927), .A2(n19900), .B1(n19899), .B2(n19916), .C1(
        n19898), .C2(n19924), .ZN(P2_U3227) );
  OAI222_X1 U22874 ( .A1(n19927), .A2(n10886), .B1(n19901), .B2(n19916), .C1(
        n19900), .C2(n19924), .ZN(P2_U3228) );
  OAI222_X1 U22875 ( .A1(n19927), .A2(n19903), .B1(n19902), .B2(n19916), .C1(
        n10886), .C2(n19924), .ZN(P2_U3229) );
  OAI222_X1 U22876 ( .A1(n19927), .A2(n15218), .B1(n19904), .B2(n19916), .C1(
        n19903), .C2(n19924), .ZN(P2_U3230) );
  OAI222_X1 U22877 ( .A1(n19927), .A2(n19906), .B1(n19905), .B2(n19916), .C1(
        n15218), .C2(n19924), .ZN(P2_U3231) );
  OAI222_X1 U22878 ( .A1(n19927), .A2(n10902), .B1(n19907), .B2(n19916), .C1(
        n19906), .C2(n19924), .ZN(P2_U3232) );
  INV_X1 U22879 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19909) );
  OAI222_X1 U22880 ( .A1(n19923), .A2(n19909), .B1(n19908), .B2(n19916), .C1(
        n10902), .C2(n19924), .ZN(P2_U3233) );
  OAI222_X1 U22881 ( .A1(n19923), .A2(n19911), .B1(n19910), .B2(n19916), .C1(
        n19909), .C2(n19924), .ZN(P2_U3234) );
  OAI222_X1 U22882 ( .A1(n19923), .A2(n19913), .B1(n19912), .B2(n19916), .C1(
        n19911), .C2(n19924), .ZN(P2_U3235) );
  OAI222_X1 U22883 ( .A1(n19923), .A2(n15162), .B1(n19914), .B2(n19916), .C1(
        n19913), .C2(n19924), .ZN(P2_U3236) );
  OAI222_X1 U22884 ( .A1(n19923), .A2(n19918), .B1(n19915), .B2(n19916), .C1(
        n15162), .C2(n19924), .ZN(P2_U3237) );
  OAI222_X1 U22885 ( .A1(n19924), .A2(n19918), .B1(n19917), .B2(n19916), .C1(
        n19919), .C2(n19923), .ZN(P2_U3238) );
  OAI222_X1 U22886 ( .A1(n19923), .A2(n19921), .B1(n19920), .B2(n19916), .C1(
        n19919), .C2(n19924), .ZN(P2_U3239) );
  OAI222_X1 U22887 ( .A1(n19923), .A2(n19925), .B1(n19922), .B2(n19916), .C1(
        n19921), .C2(n19924), .ZN(P2_U3240) );
  OAI222_X1 U22888 ( .A1(n19927), .A2(n10955), .B1(n19926), .B2(n19916), .C1(
        n19925), .C2(n19924), .ZN(P2_U3241) );
  INV_X1 U22889 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19928) );
  AOI22_X1 U22890 ( .A1(n19916), .A2(n19929), .B1(n19928), .B2(n20005), .ZN(
        P2_U3585) );
  MUX2_X1 U22891 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19916), .Z(P2_U3586) );
  INV_X1 U22892 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19930) );
  AOI22_X1 U22893 ( .A1(n19916), .A2(n19931), .B1(n19930), .B2(n20005), .ZN(
        P2_U3587) );
  INV_X1 U22894 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U22895 ( .A1(n19916), .A2(n19933), .B1(n19932), .B2(n20005), .ZN(
        P2_U3588) );
  OAI21_X1 U22896 ( .B1(n19937), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19935), 
        .ZN(n19934) );
  INV_X1 U22897 ( .A(n19934), .ZN(P2_U3591) );
  OAI21_X1 U22898 ( .B1(n19937), .B2(n19936), .A(n19935), .ZN(P2_U3592) );
  NAND2_X1 U22899 ( .A1(n19938), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19962) );
  NOR2_X1 U22900 ( .A1(n19939), .A2(n19962), .ZN(n19952) );
  OR2_X1 U22901 ( .A1(n19963), .A2(n19989), .ZN(n19943) );
  NOR2_X1 U22902 ( .A1(n19941), .A2(n19940), .ZN(n19942) );
  NAND2_X1 U22903 ( .A1(n19943), .A2(n19942), .ZN(n19954) );
  OR2_X1 U22904 ( .A1(n19952), .A2(n19954), .ZN(n19948) );
  OAI22_X1 U22905 ( .A1(n19945), .A2(n19950), .B1(n19944), .B2(n19989), .ZN(
        n19946) );
  AOI21_X1 U22906 ( .B1(n19948), .B2(n19947), .A(n19946), .ZN(n19949) );
  AOI22_X1 U22907 ( .A1(n19974), .A2(n12752), .B1(n19949), .B2(n19971), .ZN(
        P2_U3602) );
  NOR2_X1 U22908 ( .A1(n19951), .A2(n19950), .ZN(n19953) );
  AOI211_X1 U22909 ( .C1(n19955), .C2(n19954), .A(n19953), .B(n19952), .ZN(
        n19956) );
  AOI22_X1 U22910 ( .A1(n19974), .A2(n19957), .B1(n19956), .B2(n19971), .ZN(
        P2_U3603) );
  INV_X1 U22911 ( .A(n19969), .ZN(n19959) );
  OR3_X1 U22912 ( .A1(n19960), .A2(n19959), .A3(n19958), .ZN(n19961) );
  OAI21_X1 U22913 ( .B1(n19963), .B2(n19962), .A(n19961), .ZN(n19964) );
  AOI21_X1 U22914 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19965), .A(n19964), 
        .ZN(n19966) );
  AOI22_X1 U22915 ( .A1(n19974), .A2(n10498), .B1(n19966), .B2(n19971), .ZN(
        P2_U3604) );
  AOI211_X1 U22916 ( .C1(n19970), .C2(n19969), .A(n19968), .B(n19967), .ZN(
        n19972) );
  AOI22_X1 U22917 ( .A1(n19974), .A2(n19973), .B1(n19972), .B2(n19971), .ZN(
        P2_U3605) );
  INV_X1 U22918 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19975) );
  AOI22_X1 U22919 ( .A1(n19916), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19975), 
        .B2(n20005), .ZN(P2_U3608) );
  INV_X1 U22920 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19985) );
  INV_X1 U22921 ( .A(n19976), .ZN(n19980) );
  AOI22_X1 U22922 ( .A1(n19980), .A2(n19979), .B1(n19978), .B2(n19977), .ZN(
        n19983) );
  NOR2_X1 U22923 ( .A1(n19981), .A2(n19984), .ZN(n19982) );
  AOI22_X1 U22924 ( .A1(n19985), .A2(n19984), .B1(n19983), .B2(n19982), .ZN(
        P2_U3609) );
  NAND2_X1 U22925 ( .A1(n9637), .A2(n19993), .ZN(n19990) );
  NAND2_X1 U22926 ( .A1(n19987), .A2(n19986), .ZN(n19988) );
  NAND4_X1 U22927 ( .A1(n19991), .A2(n19990), .A3(n19989), .A4(n19988), .ZN(
        n20004) );
  AOI21_X1 U22928 ( .B1(n19993), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19992), 
        .ZN(n20001) );
  AOI21_X1 U22929 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19995), .A(n19994), 
        .ZN(n19999) );
  NOR3_X1 U22930 ( .A1(n19996), .A2(n19995), .A3(n13085), .ZN(n19998) );
  MUX2_X1 U22931 ( .A(n19999), .B(n19998), .S(n19997), .Z(n20000) );
  OAI21_X1 U22932 ( .B1(n20001), .B2(n20000), .A(n20004), .ZN(n20002) );
  OAI21_X1 U22933 ( .B1(n20004), .B2(n20003), .A(n20002), .ZN(P2_U3610) );
  INV_X1 U22934 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20006) );
  AOI22_X1 U22935 ( .A1(n19916), .A2(n20007), .B1(n20006), .B2(n20005), .ZN(
        P2_U3611) );
  OAI21_X1 U22936 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20008), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20855) );
  NOR2_X2 U22937 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20008), .ZN(n20942) );
  OAI21_X1 U22938 ( .B1(n20855), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20893), .ZN(
        n20009) );
  INV_X1 U22939 ( .A(n20009), .ZN(P1_U2802) );
  OAI21_X1 U22940 ( .B1(n20011), .B2(n20010), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20012) );
  OAI21_X1 U22941 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20013), .A(n20012), 
        .ZN(P1_U2803) );
  NOR2_X1 U22942 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20015) );
  OAI21_X1 U22943 ( .B1(n20015), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20893), .ZN(
        n20014) );
  OAI21_X1 U22944 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20893), .A(n20014), 
        .ZN(P1_U2804) );
  NAND2_X1 U22945 ( .A1(n20855), .A2(n20928), .ZN(n20917) );
  INV_X1 U22946 ( .A(n20917), .ZN(n20921) );
  OAI21_X1 U22947 ( .B1(BS16), .B2(n20015), .A(n20921), .ZN(n20919) );
  OAI21_X1 U22948 ( .B1(n20921), .B2(n20418), .A(n20919), .ZN(P1_U2805) );
  OAI21_X1 U22949 ( .B1(n20018), .B2(n20017), .A(n20016), .ZN(P1_U2806) );
  NOR4_X1 U22950 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20022) );
  NOR4_X1 U22951 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20021) );
  NOR4_X1 U22952 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20020) );
  NOR4_X1 U22953 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20019) );
  NAND4_X1 U22954 ( .A1(n20022), .A2(n20021), .A3(n20020), .A4(n20019), .ZN(
        n20028) );
  NOR4_X1 U22955 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20026) );
  AOI211_X1 U22956 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_9__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20025) );
  NOR4_X1 U22957 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20024) );
  NOR4_X1 U22958 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20023) );
  NAND4_X1 U22959 ( .A1(n20026), .A2(n20025), .A3(n20024), .A4(n20023), .ZN(
        n20027) );
  NOR2_X1 U22960 ( .A1(n20028), .A2(n20027), .ZN(n20927) );
  INV_X1 U22961 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20914) );
  NOR3_X1 U22962 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20030) );
  OAI21_X1 U22963 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20030), .A(n20927), .ZN(
        n20029) );
  OAI21_X1 U22964 ( .B1(n20927), .B2(n20914), .A(n20029), .ZN(P1_U2807) );
  INV_X1 U22965 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20920) );
  AOI21_X1 U22966 ( .B1(n20243), .B2(n20920), .A(n20030), .ZN(n20031) );
  INV_X1 U22967 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20911) );
  INV_X1 U22968 ( .A(n20927), .ZN(n20923) );
  AOI22_X1 U22969 ( .A1(n20927), .A2(n20031), .B1(n20911), .B2(n20923), .ZN(
        P1_U2808) );
  OAI21_X1 U22970 ( .B1(n20033), .B2(n20032), .A(n20100), .ZN(n20048) );
  OAI22_X1 U22971 ( .A1(n20048), .A2(n20867), .B1(n20035), .B2(n20034), .ZN(
        n20036) );
  AOI211_X1 U22972 ( .C1(n20095), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20209), .B(n20036), .ZN(n20043) );
  NAND4_X1 U22973 ( .A1(n20090), .A2(n20072), .A3(P1_REIP_REG_6__SCAN_IN), 
        .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n20039) );
  INV_X1 U22974 ( .A(n20037), .ZN(n20038) );
  OAI22_X1 U22975 ( .A1(n20039), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20088), 
        .B2(n20038), .ZN(n20040) );
  AOI21_X1 U22976 ( .B1(n20052), .B2(n20041), .A(n20040), .ZN(n20042) );
  OAI211_X1 U22977 ( .C1(n20044), .C2(n20101), .A(n20043), .B(n20042), .ZN(
        P1_U2833) );
  NAND2_X1 U22978 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20046) );
  AOI21_X1 U22979 ( .B1(n20103), .B2(P1_EBX_REG_6__SCAN_IN), .A(n20209), .ZN(
        n20045) );
  OAI211_X1 U22980 ( .C1(n20088), .C2(n20047), .A(n20046), .B(n20045), .ZN(
        n20050) );
  INV_X1 U22981 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20865) );
  OAI211_X1 U22982 ( .C1(n20072), .C2(n20071), .A(P1_REIP_REG_5__SCAN_IN), .B(
        n20092), .ZN(n20059) );
  AOI21_X1 U22983 ( .B1(n20865), .B2(n20059), .A(n20048), .ZN(n20049) );
  AOI211_X1 U22984 ( .C1(n20052), .C2(n20051), .A(n20050), .B(n20049), .ZN(
        n20053) );
  OAI21_X1 U22985 ( .B1(n20054), .B2(n20101), .A(n20053), .ZN(P1_U2834) );
  INV_X1 U22986 ( .A(n20109), .ZN(n20085) );
  INV_X1 U22987 ( .A(n20110), .ZN(n20057) );
  NAND2_X1 U22988 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n20056) );
  AOI21_X1 U22989 ( .B1(n20103), .B2(P1_EBX_REG_5__SCAN_IN), .A(n20209), .ZN(
        n20055) );
  OAI211_X1 U22990 ( .C1(n20057), .C2(n20088), .A(n20056), .B(n20055), .ZN(
        n20058) );
  AOI21_X1 U22991 ( .B1(n20113), .B2(n20085), .A(n20058), .ZN(n20062) );
  AND2_X1 U22992 ( .A1(n20090), .A2(n20072), .ZN(n20060) );
  OAI21_X1 U22993 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20060), .A(n20059), .ZN(
        n20061) );
  OAI211_X1 U22994 ( .C1(n20101), .C2(n20063), .A(n20062), .B(n20061), .ZN(
        P1_U2835) );
  AOI21_X1 U22995 ( .B1(n20103), .B2(P1_EBX_REG_4__SCAN_IN), .A(n20209), .ZN(
        n20064) );
  OAI21_X1 U22996 ( .B1(n20065), .B2(n20088), .A(n20064), .ZN(n20068) );
  NOR2_X1 U22997 ( .A1(n20102), .A2(n20066), .ZN(n20067) );
  AOI211_X1 U22998 ( .C1(n20104), .C2(n20069), .A(n20068), .B(n20067), .ZN(
        n20076) );
  OAI21_X1 U22999 ( .B1(n20071), .B2(n20070), .A(n20862), .ZN(n20074) );
  OAI21_X1 U23000 ( .B1(n20072), .B2(n20071), .A(n20092), .ZN(n20073) );
  AOI22_X1 U23001 ( .A1(n20085), .A2(n20188), .B1(n20074), .B2(n20073), .ZN(
        n20075) );
  OAI211_X1 U23002 ( .C1(n20192), .C2(n20101), .A(n20076), .B(n20075), .ZN(
        P1_U2836) );
  AOI22_X1 U23003 ( .A1(n20077), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_EBX_REG_2__SCAN_IN), .B2(n20103), .ZN(n20087) );
  AOI22_X1 U23004 ( .A1(n20265), .A2(n20104), .B1(n20079), .B2(n20078), .ZN(
        n20081) );
  NAND2_X1 U23005 ( .A1(n20095), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n20080) );
  OAI211_X1 U23006 ( .C1(n20101), .C2(n20082), .A(n20081), .B(n20080), .ZN(
        n20083) );
  AOI21_X1 U23007 ( .B1(n20085), .B2(n20084), .A(n20083), .ZN(n20086) );
  OAI211_X1 U23008 ( .C1(n20088), .C2(n20227), .A(n20087), .B(n20086), .ZN(
        P1_U2838) );
  AOI22_X1 U23009 ( .A1(n20089), .A2(n20099), .B1(n20103), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n20097) );
  AOI22_X1 U23010 ( .A1(n20728), .A2(n20104), .B1(n20090), .B2(n20243), .ZN(
        n20091) );
  OAI21_X1 U23011 ( .B1(n20092), .B2(n20243), .A(n20091), .ZN(n20094) );
  NOR2_X1 U23012 ( .A1(n20101), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20093) );
  AOI211_X1 U23013 ( .C1(n20095), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n20094), .B(n20093), .ZN(n20096) );
  OAI211_X1 U23014 ( .C1(n20109), .C2(n20203), .A(n20097), .B(n20096), .ZN(
        P1_U2839) );
  AOI22_X1 U23015 ( .A1(n20100), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n20099), 
        .B2(n20098), .ZN(n20107) );
  NAND2_X1 U23016 ( .A1(n20102), .A2(n20101), .ZN(n20105) );
  INV_X1 U23017 ( .A(n11556), .ZN(n20379) );
  AOI222_X1 U23018 ( .A1(n20105), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20104), .B2(n20379), .C1(P1_EBX_REG_0__SCAN_IN), .C2(n20103), .ZN(
        n20106) );
  OAI211_X1 U23019 ( .C1(n20109), .C2(n20108), .A(n20107), .B(n20106), .ZN(
        P1_U2840) );
  AOI22_X1 U23020 ( .A1(n20113), .A2(n20112), .B1(n20111), .B2(n20110), .ZN(
        n20114) );
  OAI21_X1 U23021 ( .B1(n20116), .B2(n20115), .A(n20114), .ZN(P1_U2867) );
  AOI22_X1 U23022 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20117) );
  OAI21_X1 U23023 ( .B1(n13625), .B2(n20143), .A(n20117), .ZN(P1_U2921) );
  AOI22_X1 U23024 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20118) );
  OAI21_X1 U23025 ( .B1(n14639), .B2(n20143), .A(n20118), .ZN(P1_U2922) );
  AOI22_X1 U23026 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20119) );
  OAI21_X1 U23027 ( .B1(n14640), .B2(n20143), .A(n20119), .ZN(P1_U2923) );
  AOI22_X1 U23028 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n20121), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20120), .ZN(n20122) );
  OAI21_X1 U23029 ( .B1(n21055), .B2(n20123), .A(n20122), .ZN(P1_U2924) );
  AOI22_X1 U23030 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20124) );
  OAI21_X1 U23031 ( .B1(n14646), .B2(n20143), .A(n20124), .ZN(P1_U2925) );
  AOI22_X1 U23032 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20125) );
  OAI21_X1 U23033 ( .B1(n14226), .B2(n20143), .A(n20125), .ZN(P1_U2926) );
  AOI22_X1 U23034 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20126) );
  OAI21_X1 U23035 ( .B1(n14190), .B2(n20143), .A(n20126), .ZN(P1_U2927) );
  AOI22_X1 U23036 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20127) );
  OAI21_X1 U23037 ( .B1(n14082), .B2(n20143), .A(n20127), .ZN(P1_U2928) );
  AOI22_X1 U23038 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20128) );
  OAI21_X1 U23039 ( .B1(n11707), .B2(n20143), .A(n20128), .ZN(P1_U2929) );
  AOI22_X1 U23040 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20129) );
  OAI21_X1 U23041 ( .B1(n14069), .B2(n20143), .A(n20129), .ZN(P1_U2930) );
  AOI22_X1 U23042 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20130) );
  OAI21_X1 U23043 ( .B1(n20131), .B2(n20143), .A(n20130), .ZN(P1_U2931) );
  AOI22_X1 U23044 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20132) );
  OAI21_X1 U23045 ( .B1(n20133), .B2(n20143), .A(n20132), .ZN(P1_U2932) );
  AOI22_X1 U23046 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20134) );
  OAI21_X1 U23047 ( .B1(n20135), .B2(n20143), .A(n20134), .ZN(P1_U2933) );
  AOI22_X1 U23048 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20136) );
  OAI21_X1 U23049 ( .B1(n20137), .B2(n20143), .A(n20136), .ZN(P1_U2934) );
  AOI22_X1 U23050 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20139) );
  OAI21_X1 U23051 ( .B1(n20140), .B2(n20143), .A(n20139), .ZN(P1_U2935) );
  AOI22_X1 U23052 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20141), .B1(n20138), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20142) );
  OAI21_X1 U23053 ( .B1(n20144), .B2(n20143), .A(n20142), .ZN(P1_U2936) );
  AOI22_X1 U23054 ( .A1(n20181), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20151), .ZN(n20147) );
  INV_X1 U23055 ( .A(n20145), .ZN(n20146) );
  NAND2_X1 U23056 ( .A1(n20166), .A2(n20146), .ZN(n20168) );
  NAND2_X1 U23057 ( .A1(n20147), .A2(n20168), .ZN(P1_U2945) );
  AOI22_X1 U23058 ( .A1(n20181), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20151), .ZN(n20150) );
  INV_X1 U23059 ( .A(n20148), .ZN(n20149) );
  NAND2_X1 U23060 ( .A1(n20166), .A2(n20149), .ZN(n20170) );
  NAND2_X1 U23061 ( .A1(n20150), .A2(n20170), .ZN(P1_U2946) );
  AOI22_X1 U23062 ( .A1(n20181), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20151), .ZN(n20154) );
  INV_X1 U23063 ( .A(n20152), .ZN(n20153) );
  NAND2_X1 U23064 ( .A1(n20166), .A2(n20153), .ZN(n20172) );
  NAND2_X1 U23065 ( .A1(n20154), .A2(n20172), .ZN(P1_U2947) );
  AOI22_X1 U23066 ( .A1(n20181), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20176), .ZN(n20157) );
  INV_X1 U23067 ( .A(n20155), .ZN(n20156) );
  NAND2_X1 U23068 ( .A1(n20166), .A2(n20156), .ZN(n20174) );
  NAND2_X1 U23069 ( .A1(n20157), .A2(n20174), .ZN(P1_U2948) );
  AOI22_X1 U23070 ( .A1(n20181), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20176), .ZN(n20160) );
  INV_X1 U23071 ( .A(n20158), .ZN(n20159) );
  NAND2_X1 U23072 ( .A1(n20166), .A2(n20159), .ZN(n20177) );
  NAND2_X1 U23073 ( .A1(n20160), .A2(n20177), .ZN(P1_U2949) );
  AOI22_X1 U23074 ( .A1(n20181), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20176), .ZN(n20163) );
  INV_X1 U23075 ( .A(n20161), .ZN(n20162) );
  NAND2_X1 U23076 ( .A1(n20166), .A2(n20162), .ZN(n20179) );
  NAND2_X1 U23077 ( .A1(n20163), .A2(n20179), .ZN(P1_U2950) );
  AOI22_X1 U23078 ( .A1(n20181), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20176), .ZN(n20167) );
  INV_X1 U23079 ( .A(n20164), .ZN(n20165) );
  NAND2_X1 U23080 ( .A1(n20166), .A2(n20165), .ZN(n20182) );
  NAND2_X1 U23081 ( .A1(n20167), .A2(n20182), .ZN(P1_U2951) );
  AOI22_X1 U23082 ( .A1(n20181), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20176), .ZN(n20169) );
  NAND2_X1 U23083 ( .A1(n20169), .A2(n20168), .ZN(P1_U2960) );
  AOI22_X1 U23084 ( .A1(n20181), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20176), .ZN(n20171) );
  NAND2_X1 U23085 ( .A1(n20171), .A2(n20170), .ZN(P1_U2961) );
  AOI22_X1 U23086 ( .A1(n20181), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20176), .ZN(n20173) );
  NAND2_X1 U23087 ( .A1(n20173), .A2(n20172), .ZN(P1_U2962) );
  AOI22_X1 U23088 ( .A1(n20181), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20151), .ZN(n20175) );
  NAND2_X1 U23089 ( .A1(n20175), .A2(n20174), .ZN(P1_U2963) );
  AOI22_X1 U23090 ( .A1(n20181), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20176), .ZN(n20178) );
  NAND2_X1 U23091 ( .A1(n20178), .A2(n20177), .ZN(P1_U2964) );
  AOI22_X1 U23092 ( .A1(n20181), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20151), .ZN(n20180) );
  NAND2_X1 U23093 ( .A1(n20180), .A2(n20179), .ZN(P1_U2965) );
  AOI22_X1 U23094 ( .A1(n20181), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20151), .ZN(n20183) );
  NAND2_X1 U23095 ( .A1(n20183), .A2(n20182), .ZN(P1_U2966) );
  AOI22_X1 U23096 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20191) );
  OAI21_X1 U23097 ( .B1(n20186), .B2(n20185), .A(n20184), .ZN(n20187) );
  INV_X1 U23098 ( .A(n20187), .ZN(n20207) );
  AOI22_X1 U23099 ( .A1(n20207), .A2(n20200), .B1(n20189), .B2(n20188), .ZN(
        n20190) );
  OAI211_X1 U23100 ( .C1(n20193), .C2(n20192), .A(n20191), .B(n20190), .ZN(
        P1_U2995) );
  AOI22_X1 U23101 ( .A1(n20194), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20209), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20202) );
  OAI21_X1 U23102 ( .B1(n20196), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20195), .ZN(n20197) );
  INV_X1 U23103 ( .A(n20197), .ZN(n20250) );
  INV_X1 U23104 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20198) );
  AOI22_X1 U23105 ( .A1(n20250), .A2(n20200), .B1(n20199), .B2(n20198), .ZN(
        n20201) );
  OAI211_X1 U23106 ( .C1(n20258), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        P1_U2998) );
  AOI21_X1 U23107 ( .B1(n20206), .B2(n20205), .A(n20204), .ZN(n20221) );
  AOI222_X1 U23108 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20209), .B1(n20235), 
        .B2(n20208), .C1(n20249), .C2(n20207), .ZN(n20212) );
  OAI211_X1 U23109 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20216), .B(n20210), .ZN(n20211) );
  OAI211_X1 U23110 ( .C1(n20221), .C2(n20213), .A(n20212), .B(n20211), .ZN(
        P1_U3027) );
  AOI22_X1 U23111 ( .A1(n20209), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20235), 
        .B2(n20214), .ZN(n20219) );
  INV_X1 U23112 ( .A(n20215), .ZN(n20217) );
  AOI22_X1 U23113 ( .A1(n20217), .A2(n20249), .B1(n20220), .B2(n20216), .ZN(
        n20218) );
  OAI211_X1 U23114 ( .C1(n20221), .C2(n20220), .A(n20219), .B(n20218), .ZN(
        P1_U3028) );
  NAND2_X1 U23115 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20222), .ZN(
        n20239) );
  NOR3_X1 U23116 ( .A1(n20223), .A2(n20254), .A3(n20229), .ZN(n20225) );
  AOI211_X1 U23117 ( .C1(n20254), .C2(n20226), .A(n20225), .B(n20224), .ZN(
        n20237) );
  INV_X1 U23118 ( .A(n20227), .ZN(n20234) );
  OAI22_X1 U23119 ( .A1(n20229), .A2(n20228), .B1(n20078), .B2(n20244), .ZN(
        n20233) );
  NOR2_X1 U23120 ( .A1(n20231), .A2(n20230), .ZN(n20232) );
  AOI211_X1 U23121 ( .C1(n20235), .C2(n20234), .A(n20233), .B(n20232), .ZN(
        n20236) );
  OAI221_X1 U23122 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20239), .C1(
        n20238), .C2(n20237), .A(n20236), .ZN(P1_U3029) );
  INV_X1 U23123 ( .A(n20240), .ZN(n20241) );
  NOR3_X1 U23124 ( .A1(n20242), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20241), .ZN(n20248) );
  OAI22_X1 U23125 ( .A1(n20246), .A2(n20245), .B1(n20244), .B2(n20243), .ZN(
        n20247) );
  AOI211_X1 U23126 ( .C1(n20250), .C2(n20249), .A(n20248), .B(n20247), .ZN(
        n20251) );
  OAI221_X1 U23127 ( .B1(n20254), .B2(n20253), .C1(n20254), .C2(n20252), .A(
        n20251), .ZN(P1_U3030) );
  AND2_X1 U23128 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20255), .ZN(
        P1_U3032) );
  INV_X1 U23129 ( .A(n13980), .ZN(n20259) );
  NAND2_X1 U23130 ( .A1(n20338), .A2(n12353), .ZN(n20414) );
  OR2_X1 U23131 ( .A1(n12353), .A2(n20338), .ZN(n20372) );
  AOI22_X1 U23132 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9623), .B1(DATAI_24_), 
        .B2(n9622), .ZN(n20742) );
  NAND2_X1 U23133 ( .A1(n20590), .A2(n20537), .ZN(n20377) );
  OR2_X1 U23134 ( .A1(n20662), .A2(n20377), .ZN(n20307) );
  OR2_X1 U23135 ( .A1(n20261), .A2(n20289), .ZN(n20663) );
  OAI22_X1 U23136 ( .A1(n20837), .A2(n20742), .B1(n20307), .B2(n20663), .ZN(
        n20262) );
  INV_X1 U23137 ( .A(n20262), .ZN(n20274) );
  INV_X1 U23138 ( .A(n20591), .ZN(n20263) );
  NOR2_X1 U23139 ( .A1(n20538), .A2(n20263), .ZN(n20270) );
  NAND2_X1 U23140 ( .A1(n20269), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20729) );
  AND2_X1 U23141 ( .A1(n20421), .A2(n20729), .ZN(n20593) );
  NAND2_X1 U23142 ( .A1(n20337), .A2(n20837), .ZN(n20264) );
  AOI21_X1 U23143 ( .B1(n20264), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20782), 
        .ZN(n20268) );
  NAND2_X1 U23144 ( .A1(n9650), .A2(n14906), .ZN(n20271) );
  AOI22_X1 U23145 ( .A1(n20268), .A2(n20271), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20307), .ZN(n20266) );
  OAI211_X1 U23146 ( .C1(n20270), .C2(n20780), .A(n20593), .B(n20266), .ZN(
        n20311) );
  NOR2_X2 U23147 ( .A1(n20267), .A2(n20317), .ZN(n20784) );
  INV_X1 U23148 ( .A(n20268), .ZN(n20272) );
  OR2_X1 U23149 ( .A1(n20269), .A2(n20780), .ZN(n20595) );
  INV_X1 U23150 ( .A(n20270), .ZN(n20417) );
  OAI22_X1 U23151 ( .A1(n20272), .A2(n20271), .B1(n20595), .B2(n20417), .ZN(
        n20310) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20311), .B1(
        n20784), .B2(n20310), .ZN(n20273) );
  OAI211_X1 U23153 ( .C1(n20795), .C2(n20337), .A(n20274), .B(n20273), .ZN(
        P1_U3033) );
  AOI22_X1 U23154 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9623), .B1(DATAI_25_), 
        .B2(n9622), .ZN(n20746) );
  OAI22_X1 U23155 ( .A1(n20837), .A2(n20746), .B1(n20307), .B2(n20600), .ZN(
        n20276) );
  INV_X1 U23156 ( .A(n20276), .ZN(n20279) );
  NOR2_X2 U23157 ( .A1(n20277), .A2(n20317), .ZN(n20797) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20311), .B1(
        n20797), .B2(n20310), .ZN(n20278) );
  OAI211_X1 U23159 ( .C1(n20801), .C2(n20337), .A(n20279), .B(n20278), .ZN(
        P1_U3034) );
  AOI22_X1 U23160 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9623), .B1(DATAI_26_), 
        .B2(n9622), .ZN(n20750) );
  OR2_X1 U23161 ( .A1(n20280), .A2(n20289), .ZN(n20679) );
  OAI22_X1 U23162 ( .A1(n20837), .A2(n20750), .B1(n20307), .B2(n20679), .ZN(
        n20281) );
  INV_X1 U23163 ( .A(n20281), .ZN(n20284) );
  NOR2_X2 U23164 ( .A1(n20282), .A2(n20317), .ZN(n20803) );
  AOI22_X1 U23165 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20311), .B1(
        n20803), .B2(n20310), .ZN(n20283) );
  OAI211_X1 U23166 ( .C1(n20807), .C2(n20337), .A(n20284), .B(n20283), .ZN(
        P1_U3035) );
  AOI22_X1 U23167 ( .A1(DATAI_19_), .A2(n9622), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9623), .ZN(n20813) );
  OAI22_X1 U23168 ( .A1(n20837), .A2(n20754), .B1(n20307), .B2(n20607), .ZN(
        n20285) );
  INV_X1 U23169 ( .A(n20285), .ZN(n20288) );
  NOR2_X2 U23170 ( .A1(n20286), .A2(n20317), .ZN(n20809) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20311), .B1(
        n20809), .B2(n20310), .ZN(n20287) );
  OAI211_X1 U23172 ( .C1(n20813), .C2(n20337), .A(n20288), .B(n20287), .ZN(
        P1_U3036) );
  AOI22_X1 U23173 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9623), .B1(DATAI_28_), 
        .B2(n9622), .ZN(n20758) );
  OR2_X1 U23174 ( .A1(n20290), .A2(n20289), .ZN(n20686) );
  OAI22_X1 U23175 ( .A1(n20837), .A2(n20758), .B1(n20307), .B2(n20686), .ZN(
        n20291) );
  INV_X1 U23176 ( .A(n20291), .ZN(n20294) );
  NOR2_X2 U23177 ( .A1(n20292), .A2(n20317), .ZN(n21142) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20311), .B1(
        n21142), .B2(n20310), .ZN(n20293) );
  OAI211_X1 U23179 ( .C1(n21149), .C2(n20337), .A(n20294), .B(n20293), .ZN(
        P1_U3037) );
  AOI22_X1 U23180 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9623), .B1(DATAI_29_), 
        .B2(n9622), .ZN(n20762) );
  OAI22_X1 U23181 ( .A1(n20837), .A2(n20762), .B1(n20307), .B2(n20614), .ZN(
        n20296) );
  INV_X1 U23182 ( .A(n20296), .ZN(n20299) );
  NOR2_X2 U23183 ( .A1(n20297), .A2(n20317), .ZN(n20817) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20311), .B1(
        n20817), .B2(n20310), .ZN(n20298) );
  OAI211_X1 U23185 ( .C1(n20821), .C2(n20337), .A(n20299), .B(n20298), .ZN(
        P1_U3038) );
  AOI22_X1 U23186 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9623), .B1(DATAI_30_), 
        .B2(n9622), .ZN(n20766) );
  OAI22_X1 U23187 ( .A1(n20837), .A2(n20766), .B1(n20307), .B2(n20618), .ZN(
        n20300) );
  INV_X1 U23188 ( .A(n20300), .ZN(n20303) );
  NOR2_X2 U23189 ( .A1(n20301), .A2(n20317), .ZN(n20823) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20311), .B1(
        n20823), .B2(n20310), .ZN(n20302) );
  OAI211_X1 U23191 ( .C1(n20827), .C2(n20337), .A(n20303), .B(n20302), .ZN(
        P1_U3039) );
  AOI22_X1 U23192 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9623), .B1(DATAI_23_), 
        .B2(n9622), .ZN(n20838) );
  OAI22_X1 U23193 ( .A1(n20837), .A2(n20774), .B1(n20307), .B2(n20622), .ZN(
        n20308) );
  INV_X1 U23194 ( .A(n20308), .ZN(n20313) );
  NOR2_X2 U23195 ( .A1(n20309), .A2(n20317), .ZN(n20831) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20311), .B1(
        n20831), .B2(n20310), .ZN(n20312) );
  OAI211_X1 U23197 ( .C1(n20838), .C2(n20337), .A(n20313), .B(n20312), .ZN(
        P1_U3040) );
  INV_X1 U23198 ( .A(n12353), .ZN(n20339) );
  INV_X1 U23199 ( .A(n20700), .ZN(n20314) );
  INV_X1 U23200 ( .A(n20315), .ZN(n20702) );
  NOR3_X2 U23201 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20701), .A3(
        n20377), .ZN(n21139) );
  AOI21_X1 U23202 ( .B1(n9650), .B2(n20702), .A(n21139), .ZN(n20319) );
  INV_X1 U23203 ( .A(n20377), .ZN(n20374) );
  NAND2_X1 U23204 ( .A1(n20374), .A2(n20779), .ZN(n20316) );
  OAI22_X1 U23205 ( .A1(n20319), .A2(n20782), .B1(n20316), .B2(n20780), .ZN(
        n21141) );
  AOI22_X1 U23206 ( .A1(n20784), .A2(n21141), .B1(n20783), .B2(n21139), .ZN(
        n20323) );
  INV_X1 U23207 ( .A(n20316), .ZN(n20321) );
  INV_X1 U23208 ( .A(n20373), .ZN(n20318) );
  NOR2_X1 U23209 ( .A1(n20318), .A2(n20782), .ZN(n20382) );
  INV_X1 U23210 ( .A(n20666), .ZN(n20705) );
  OAI21_X1 U23211 ( .B1(n20382), .B2(n20705), .A(n20319), .ZN(n20320) );
  OAI211_X1 U23212 ( .C1(n20791), .C2(n20321), .A(n20789), .B(n20320), .ZN(
        n21145) );
  INV_X1 U23213 ( .A(n20337), .ZN(n21144) );
  INV_X1 U23214 ( .A(n20742), .ZN(n20792) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n20792), .ZN(n20322) );
  OAI211_X1 U23216 ( .C1(n20795), .C2(n21148), .A(n20323), .B(n20322), .ZN(
        P1_U3041) );
  AOI22_X1 U23217 ( .A1(n20797), .A2(n21141), .B1(n20796), .B2(n21139), .ZN(
        n20325) );
  INV_X1 U23218 ( .A(n21148), .ZN(n20334) );
  INV_X1 U23219 ( .A(n20801), .ZN(n20743) );
  AOI22_X1 U23220 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21145), .B1(
        n20334), .B2(n20743), .ZN(n20324) );
  OAI211_X1 U23221 ( .C1(n20746), .C2(n20337), .A(n20325), .B(n20324), .ZN(
        P1_U3042) );
  AOI22_X1 U23222 ( .A1(n20803), .A2(n21141), .B1(n20802), .B2(n21139), .ZN(
        n20327) );
  INV_X1 U23223 ( .A(n20750), .ZN(n20804) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n20804), .ZN(n20326) );
  OAI211_X1 U23225 ( .C1(n20807), .C2(n21148), .A(n20327), .B(n20326), .ZN(
        P1_U3043) );
  AOI22_X1 U23226 ( .A1(n20809), .A2(n21141), .B1(n20808), .B2(n21139), .ZN(
        n20329) );
  INV_X1 U23227 ( .A(n20813), .ZN(n20751) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21145), .B1(
        n20334), .B2(n20751), .ZN(n20328) );
  OAI211_X1 U23229 ( .C1(n20754), .C2(n20337), .A(n20329), .B(n20328), .ZN(
        P1_U3044) );
  AOI22_X1 U23230 ( .A1(n20817), .A2(n21141), .B1(n20816), .B2(n21139), .ZN(
        n20331) );
  INV_X1 U23231 ( .A(n20762), .ZN(n20818) );
  AOI22_X1 U23232 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n20818), .ZN(n20330) );
  OAI211_X1 U23233 ( .C1(n20821), .C2(n21148), .A(n20331), .B(n20330), .ZN(
        P1_U3046) );
  AOI22_X1 U23234 ( .A1(n20823), .A2(n21141), .B1(n20822), .B2(n21139), .ZN(
        n20333) );
  INV_X1 U23235 ( .A(n20827), .ZN(n20763) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21145), .B1(
        n20334), .B2(n20763), .ZN(n20332) );
  OAI211_X1 U23237 ( .C1(n20766), .C2(n20337), .A(n20333), .B(n20332), .ZN(
        P1_U3047) );
  AOI22_X1 U23238 ( .A1(n20831), .A2(n21141), .B1(n20828), .B2(n21139), .ZN(
        n20336) );
  INV_X1 U23239 ( .A(n20838), .ZN(n20769) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21145), .B1(
        n20334), .B2(n20769), .ZN(n20335) );
  OAI211_X1 U23241 ( .C1(n20774), .C2(n20337), .A(n20336), .B(n20335), .ZN(
        P1_U3048) );
  OR3_X1 U23242 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20779), .A3(
        n20377), .ZN(n20366) );
  OAI22_X1 U23243 ( .A1(n20413), .A2(n20795), .B1(n20663), .B2(n20366), .ZN(
        n20340) );
  INV_X1 U23244 ( .A(n20340), .ZN(n20347) );
  NAND3_X1 U23245 ( .A1(n21148), .A2(n20413), .A3(n20791), .ZN(n20341) );
  NAND2_X1 U23246 ( .A1(n20341), .A2(n20666), .ZN(n20343) );
  NAND2_X1 U23247 ( .A1(n9650), .A2(n20728), .ZN(n20344) );
  AOI22_X1 U23248 ( .A1(n20343), .A2(n20344), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20366), .ZN(n20342) );
  OR2_X1 U23249 ( .A1(n20591), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20476) );
  NAND2_X1 U23250 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20476), .ZN(n20473) );
  NAND3_X1 U23251 ( .A1(n20593), .A2(n20342), .A3(n20473), .ZN(n20369) );
  INV_X1 U23252 ( .A(n20343), .ZN(n20345) );
  OAI22_X1 U23253 ( .A1(n20345), .A2(n20344), .B1(n20595), .B2(n20476), .ZN(
        n20368) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20369), .B1(
        n20784), .B2(n20368), .ZN(n20346) );
  OAI211_X1 U23255 ( .C1(n20742), .C2(n21148), .A(n20347), .B(n20346), .ZN(
        P1_U3049) );
  OAI22_X1 U23256 ( .A1(n20413), .A2(n20801), .B1(n20366), .B2(n20600), .ZN(
        n20348) );
  INV_X1 U23257 ( .A(n20348), .ZN(n20350) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20369), .B1(
        n20797), .B2(n20368), .ZN(n20349) );
  OAI211_X1 U23259 ( .C1(n20746), .C2(n21148), .A(n20350), .B(n20349), .ZN(
        P1_U3050) );
  OAI22_X1 U23260 ( .A1(n20413), .A2(n20807), .B1(n20679), .B2(n20366), .ZN(
        n20351) );
  INV_X1 U23261 ( .A(n20351), .ZN(n20353) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20369), .B1(
        n20803), .B2(n20368), .ZN(n20352) );
  OAI211_X1 U23263 ( .C1(n20750), .C2(n21148), .A(n20353), .B(n20352), .ZN(
        P1_U3051) );
  OAI22_X1 U23264 ( .A1(n21148), .A2(n20754), .B1(n20607), .B2(n20366), .ZN(
        n20354) );
  INV_X1 U23265 ( .A(n20354), .ZN(n20356) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20369), .B1(
        n20809), .B2(n20368), .ZN(n20355) );
  OAI211_X1 U23267 ( .C1(n20813), .C2(n20413), .A(n20356), .B(n20355), .ZN(
        P1_U3052) );
  OAI22_X1 U23268 ( .A1(n21148), .A2(n20758), .B1(n20366), .B2(n20686), .ZN(
        n20357) );
  INV_X1 U23269 ( .A(n20357), .ZN(n20359) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20369), .B1(
        n21142), .B2(n20368), .ZN(n20358) );
  OAI211_X1 U23271 ( .C1(n21149), .C2(n20413), .A(n20359), .B(n20358), .ZN(
        P1_U3053) );
  OAI22_X1 U23272 ( .A1(n20413), .A2(n20821), .B1(n20614), .B2(n20366), .ZN(
        n20360) );
  INV_X1 U23273 ( .A(n20360), .ZN(n20362) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20369), .B1(
        n20817), .B2(n20368), .ZN(n20361) );
  OAI211_X1 U23275 ( .C1(n20762), .C2(n21148), .A(n20362), .B(n20361), .ZN(
        P1_U3054) );
  OAI22_X1 U23276 ( .A1(n20413), .A2(n20827), .B1(n20366), .B2(n20618), .ZN(
        n20363) );
  INV_X1 U23277 ( .A(n20363), .ZN(n20365) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20369), .B1(
        n20823), .B2(n20368), .ZN(n20364) );
  OAI211_X1 U23279 ( .C1(n20766), .C2(n21148), .A(n20365), .B(n20364), .ZN(
        P1_U3055) );
  OAI22_X1 U23280 ( .A1(n21148), .A2(n20774), .B1(n20622), .B2(n20366), .ZN(
        n20367) );
  INV_X1 U23281 ( .A(n20367), .ZN(n20371) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20369), .B1(
        n20831), .B2(n20368), .ZN(n20370) );
  OAI211_X1 U23283 ( .C1(n20838), .C2(n20413), .A(n20371), .B(n20370), .ZN(
        P1_U3056) );
  NAND2_X1 U23284 ( .A1(n20375), .A2(n20374), .ZN(n20407) );
  OAI22_X1 U23285 ( .A1(n20423), .A2(n20795), .B1(n20663), .B2(n20407), .ZN(
        n20376) );
  INV_X1 U23286 ( .A(n20376), .ZN(n20388) );
  NOR2_X1 U23287 ( .A1(n20779), .A2(n20377), .ZN(n20383) );
  AND2_X1 U23288 ( .A1(n20379), .A2(n20378), .ZN(n20776) );
  INV_X1 U23289 ( .A(n20407), .ZN(n20380) );
  AOI21_X1 U23290 ( .B1(n9650), .B2(n20776), .A(n20380), .ZN(n20386) );
  OAI21_X1 U23291 ( .B1(n20382), .B2(n20787), .A(n20386), .ZN(n20381) );
  OAI211_X1 U23292 ( .C1(n20791), .C2(n20383), .A(n20789), .B(n20381), .ZN(
        n20410) );
  NOR2_X1 U23293 ( .A1(n20382), .A2(n20787), .ZN(n20385) );
  INV_X1 U23294 ( .A(n20383), .ZN(n20384) );
  OAI22_X1 U23295 ( .A1(n20386), .A2(n20385), .B1(n20780), .B2(n20384), .ZN(
        n20409) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20410), .B1(
        n20784), .B2(n20409), .ZN(n20387) );
  OAI211_X1 U23297 ( .C1(n20742), .C2(n20413), .A(n20388), .B(n20387), .ZN(
        P1_U3057) );
  OAI22_X1 U23298 ( .A1(n20423), .A2(n20801), .B1(n20407), .B2(n20600), .ZN(
        n20389) );
  INV_X1 U23299 ( .A(n20389), .ZN(n20391) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20410), .B1(
        n20797), .B2(n20409), .ZN(n20390) );
  OAI211_X1 U23301 ( .C1(n20746), .C2(n20413), .A(n20391), .B(n20390), .ZN(
        P1_U3058) );
  OAI22_X1 U23302 ( .A1(n20413), .A2(n20750), .B1(n20679), .B2(n20407), .ZN(
        n20392) );
  INV_X1 U23303 ( .A(n20392), .ZN(n20394) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20410), .B1(
        n20803), .B2(n20409), .ZN(n20393) );
  OAI211_X1 U23305 ( .C1(n20807), .C2(n20423), .A(n20394), .B(n20393), .ZN(
        P1_U3059) );
  OAI22_X1 U23306 ( .A1(n20423), .A2(n20813), .B1(n20607), .B2(n20407), .ZN(
        n20395) );
  INV_X1 U23307 ( .A(n20395), .ZN(n20397) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20410), .B1(
        n20809), .B2(n20409), .ZN(n20396) );
  OAI211_X1 U23309 ( .C1(n20754), .C2(n20413), .A(n20397), .B(n20396), .ZN(
        P1_U3060) );
  OAI22_X1 U23310 ( .A1(n20413), .A2(n20758), .B1(n20686), .B2(n20407), .ZN(
        n20398) );
  INV_X1 U23311 ( .A(n20398), .ZN(n20400) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20410), .B1(
        n21142), .B2(n20409), .ZN(n20399) );
  OAI211_X1 U23313 ( .C1(n21149), .C2(n20423), .A(n20400), .B(n20399), .ZN(
        P1_U3061) );
  OAI22_X1 U23314 ( .A1(n20413), .A2(n20762), .B1(n20614), .B2(n20407), .ZN(
        n20401) );
  INV_X1 U23315 ( .A(n20401), .ZN(n20403) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20410), .B1(
        n20817), .B2(n20409), .ZN(n20402) );
  OAI211_X1 U23317 ( .C1(n20821), .C2(n20423), .A(n20403), .B(n20402), .ZN(
        P1_U3062) );
  OAI22_X1 U23318 ( .A1(n20423), .A2(n20827), .B1(n20407), .B2(n20618), .ZN(
        n20404) );
  INV_X1 U23319 ( .A(n20404), .ZN(n20406) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20410), .B1(
        n20823), .B2(n20409), .ZN(n20405) );
  OAI211_X1 U23321 ( .C1(n20766), .C2(n20413), .A(n20406), .B(n20405), .ZN(
        P1_U3063) );
  OAI22_X1 U23322 ( .A1(n20423), .A2(n20838), .B1(n20622), .B2(n20407), .ZN(
        n20408) );
  INV_X1 U23323 ( .A(n20408), .ZN(n20412) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20410), .B1(
        n20831), .B2(n20409), .ZN(n20411) );
  OAI211_X1 U23325 ( .C1(n20774), .C2(n20413), .A(n20412), .B(n20411), .ZN(
        P1_U3064) );
  NOR2_X1 U23326 ( .A1(n13698), .A2(n20415), .ZN(n20508) );
  NAND3_X1 U23327 ( .A1(n20508), .A2(n20791), .A3(n14906), .ZN(n20416) );
  OAI21_X1 U23328 ( .B1(n20729), .B2(n20417), .A(n20416), .ZN(n20438) );
  AOI22_X1 U23329 ( .A1(n20784), .A2(n20438), .B1(n20783), .B2(n10070), .ZN(
        n20425) );
  AOI21_X1 U23330 ( .B1(n20423), .B2(n20468), .A(n20418), .ZN(n20419) );
  AOI21_X1 U23331 ( .B1(n20508), .B2(n14906), .A(n20419), .ZN(n20420) );
  NOR2_X1 U23332 ( .A1(n20420), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20422) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20792), .ZN(n20424) );
  OAI211_X1 U23334 ( .C1(n20795), .C2(n20468), .A(n20425), .B(n20424), .ZN(
        P1_U3065) );
  AOI22_X1 U23335 ( .A1(n20797), .A2(n20438), .B1(n20796), .B2(n10070), .ZN(
        n20427) );
  INV_X1 U23336 ( .A(n20746), .ZN(n20798) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20798), .ZN(n20426) );
  OAI211_X1 U23338 ( .C1(n20801), .C2(n20468), .A(n20427), .B(n20426), .ZN(
        P1_U3066) );
  AOI22_X1 U23339 ( .A1(n20803), .A2(n20438), .B1(n20802), .B2(n10070), .ZN(
        n20429) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20804), .ZN(n20428) );
  OAI211_X1 U23341 ( .C1(n20807), .C2(n20468), .A(n20429), .B(n20428), .ZN(
        P1_U3067) );
  AOI22_X1 U23342 ( .A1(n20809), .A2(n20438), .B1(n20808), .B2(n10070), .ZN(
        n20431) );
  INV_X1 U23343 ( .A(n20754), .ZN(n20810) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20810), .ZN(n20430) );
  OAI211_X1 U23345 ( .C1(n20813), .C2(n20468), .A(n20431), .B(n20430), .ZN(
        P1_U3068) );
  AOI22_X1 U23346 ( .A1(n21142), .A2(n20438), .B1(n21140), .B2(n10070), .ZN(
        n20433) );
  INV_X1 U23347 ( .A(n20758), .ZN(n21143) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n21143), .ZN(n20432) );
  OAI211_X1 U23349 ( .C1(n21149), .C2(n20468), .A(n20433), .B(n20432), .ZN(
        P1_U3069) );
  AOI22_X1 U23350 ( .A1(n20817), .A2(n20438), .B1(n20816), .B2(n10070), .ZN(
        n20435) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20818), .ZN(n20434) );
  OAI211_X1 U23352 ( .C1(n20821), .C2(n20468), .A(n20435), .B(n20434), .ZN(
        P1_U3070) );
  AOI22_X1 U23353 ( .A1(n20823), .A2(n20438), .B1(n20822), .B2(n10070), .ZN(
        n20437) );
  INV_X1 U23354 ( .A(n20766), .ZN(n20824) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20824), .ZN(n20436) );
  OAI211_X1 U23356 ( .C1(n20827), .C2(n20468), .A(n20437), .B(n20436), .ZN(
        P1_U3071) );
  AOI22_X1 U23357 ( .A1(n20831), .A2(n20438), .B1(n20828), .B2(n10070), .ZN(
        n20442) );
  INV_X1 U23358 ( .A(n20774), .ZN(n20832) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20440), .B1(
        n20439), .B2(n20832), .ZN(n20441) );
  OAI211_X1 U23360 ( .C1(n20838), .C2(n20468), .A(n20442), .B(n20441), .ZN(
        P1_U3072) );
  NOR2_X1 U23361 ( .A1(n20470), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20446) );
  INV_X1 U23362 ( .A(n20446), .ZN(n20443) );
  NOR2_X1 U23363 ( .A1(n20701), .A2(n20443), .ZN(n20462) );
  AOI21_X1 U23364 ( .B1(n20508), .B2(n20702), .A(n20462), .ZN(n20444) );
  OAI22_X1 U23365 ( .A1(n20444), .A2(n20782), .B1(n20443), .B2(n20780), .ZN(
        n20463) );
  AOI22_X1 U23366 ( .A1(n20784), .A2(n20463), .B1(n20783), .B2(n20462), .ZN(
        n20448) );
  NOR2_X1 U23367 ( .A1(n20506), .A2(n20782), .ZN(n20511) );
  OAI21_X1 U23368 ( .B1(n20511), .B2(n20705), .A(n20444), .ZN(n20445) );
  OAI211_X1 U23369 ( .C1(n20791), .C2(n20446), .A(n20789), .B(n20445), .ZN(
        n20465) );
  INV_X1 U23370 ( .A(n20500), .ZN(n20464) );
  INV_X1 U23371 ( .A(n20795), .ZN(n20739) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20739), .ZN(n20447) );
  OAI211_X1 U23373 ( .C1(n20742), .C2(n20468), .A(n20448), .B(n20447), .ZN(
        P1_U3073) );
  AOI22_X1 U23374 ( .A1(n20797), .A2(n20463), .B1(n20796), .B2(n20462), .ZN(
        n20450) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20743), .ZN(n20449) );
  OAI211_X1 U23376 ( .C1(n20746), .C2(n20468), .A(n20450), .B(n20449), .ZN(
        P1_U3074) );
  AOI22_X1 U23377 ( .A1(n20803), .A2(n20463), .B1(n20802), .B2(n20462), .ZN(
        n20452) );
  INV_X1 U23378 ( .A(n20468), .ZN(n20459) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20465), .B1(
        n20459), .B2(n20804), .ZN(n20451) );
  OAI211_X1 U23380 ( .C1(n20807), .C2(n20500), .A(n20452), .B(n20451), .ZN(
        P1_U3075) );
  AOI22_X1 U23381 ( .A1(n20809), .A2(n20463), .B1(n20808), .B2(n20462), .ZN(
        n20454) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20751), .ZN(n20453) );
  OAI211_X1 U23383 ( .C1(n20754), .C2(n20468), .A(n20454), .B(n20453), .ZN(
        P1_U3076) );
  AOI22_X1 U23384 ( .A1(n21142), .A2(n20463), .B1(n21140), .B2(n20462), .ZN(
        n20456) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20465), .B1(
        n20459), .B2(n21143), .ZN(n20455) );
  OAI211_X1 U23386 ( .C1(n21149), .C2(n20500), .A(n20456), .B(n20455), .ZN(
        P1_U3077) );
  AOI22_X1 U23387 ( .A1(n20817), .A2(n20463), .B1(n20816), .B2(n20462), .ZN(
        n20458) );
  INV_X1 U23388 ( .A(n20821), .ZN(n20759) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20759), .ZN(n20457) );
  OAI211_X1 U23390 ( .C1(n20762), .C2(n20468), .A(n20458), .B(n20457), .ZN(
        P1_U3078) );
  AOI22_X1 U23391 ( .A1(n20823), .A2(n20463), .B1(n20822), .B2(n20462), .ZN(
        n20461) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20465), .B1(
        n20459), .B2(n20824), .ZN(n20460) );
  OAI211_X1 U23393 ( .C1(n20827), .C2(n20500), .A(n20461), .B(n20460), .ZN(
        P1_U3079) );
  AOI22_X1 U23394 ( .A1(n20831), .A2(n20463), .B1(n20828), .B2(n20462), .ZN(
        n20467) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20769), .ZN(n20466) );
  OAI211_X1 U23396 ( .C1(n20774), .C2(n20468), .A(n20467), .B(n20466), .ZN(
        P1_U3080) );
  NOR2_X1 U23397 ( .A1(n20779), .A2(n20470), .ZN(n20513) );
  INV_X1 U23398 ( .A(n20513), .ZN(n20509) );
  OR2_X1 U23399 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20509), .ZN(
        n20499) );
  OAI22_X1 U23400 ( .A1(n20500), .A2(n20742), .B1(n20499), .B2(n20663), .ZN(
        n20471) );
  INV_X1 U23401 ( .A(n20471), .ZN(n20480) );
  NAND3_X1 U23402 ( .A1(n20535), .A2(n20500), .A3(n20791), .ZN(n20472) );
  NAND2_X1 U23403 ( .A1(n20472), .A2(n20666), .ZN(n20475) );
  NAND2_X1 U23404 ( .A1(n20508), .A2(n20728), .ZN(n20477) );
  AOI22_X1 U23405 ( .A1(n20475), .A2(n20477), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20499), .ZN(n20474) );
  NAND3_X1 U23406 ( .A1(n20737), .A2(n20474), .A3(n20473), .ZN(n20503) );
  INV_X1 U23407 ( .A(n20475), .ZN(n20478) );
  OAI22_X1 U23408 ( .A1(n20478), .A2(n20477), .B1(n20476), .B2(n20729), .ZN(
        n20502) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20503), .B1(
        n20784), .B2(n20502), .ZN(n20479) );
  OAI211_X1 U23410 ( .C1(n20795), .C2(n20535), .A(n20480), .B(n20479), .ZN(
        P1_U3081) );
  OAI22_X1 U23411 ( .A1(n20500), .A2(n20746), .B1(n20600), .B2(n20499), .ZN(
        n20481) );
  INV_X1 U23412 ( .A(n20481), .ZN(n20483) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20503), .B1(
        n20797), .B2(n20502), .ZN(n20482) );
  OAI211_X1 U23414 ( .C1(n20801), .C2(n20535), .A(n20483), .B(n20482), .ZN(
        P1_U3082) );
  OAI22_X1 U23415 ( .A1(n20535), .A2(n20807), .B1(n20679), .B2(n20499), .ZN(
        n20484) );
  INV_X1 U23416 ( .A(n20484), .ZN(n20486) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20503), .B1(
        n20803), .B2(n20502), .ZN(n20485) );
  OAI211_X1 U23418 ( .C1(n20750), .C2(n20500), .A(n20486), .B(n20485), .ZN(
        P1_U3083) );
  OAI22_X1 U23419 ( .A1(n20500), .A2(n20754), .B1(n20499), .B2(n20607), .ZN(
        n20487) );
  INV_X1 U23420 ( .A(n20487), .ZN(n20489) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20503), .B1(
        n20809), .B2(n20502), .ZN(n20488) );
  OAI211_X1 U23422 ( .C1(n20813), .C2(n20535), .A(n20489), .B(n20488), .ZN(
        P1_U3084) );
  OAI22_X1 U23423 ( .A1(n20500), .A2(n20758), .B1(n20499), .B2(n20686), .ZN(
        n20490) );
  INV_X1 U23424 ( .A(n20490), .ZN(n20492) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20503), .B1(
        n21142), .B2(n20502), .ZN(n20491) );
  OAI211_X1 U23426 ( .C1(n21149), .C2(n20535), .A(n20492), .B(n20491), .ZN(
        P1_U3085) );
  OAI22_X1 U23427 ( .A1(n20535), .A2(n20821), .B1(n20614), .B2(n20499), .ZN(
        n20493) );
  INV_X1 U23428 ( .A(n20493), .ZN(n20495) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20503), .B1(
        n20817), .B2(n20502), .ZN(n20494) );
  OAI211_X1 U23430 ( .C1(n20762), .C2(n20500), .A(n20495), .B(n20494), .ZN(
        P1_U3086) );
  OAI22_X1 U23431 ( .A1(n20500), .A2(n20766), .B1(n20618), .B2(n20499), .ZN(
        n20496) );
  INV_X1 U23432 ( .A(n20496), .ZN(n20498) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20503), .B1(
        n20823), .B2(n20502), .ZN(n20497) );
  OAI211_X1 U23434 ( .C1(n20827), .C2(n20535), .A(n20498), .B(n20497), .ZN(
        P1_U3087) );
  OAI22_X1 U23435 ( .A1(n20500), .A2(n20774), .B1(n20499), .B2(n20622), .ZN(
        n20501) );
  INV_X1 U23436 ( .A(n20501), .ZN(n20505) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20503), .B1(
        n20831), .B2(n20502), .ZN(n20504) );
  OAI211_X1 U23438 ( .C1(n20838), .C2(n20535), .A(n20505), .B(n20504), .ZN(
        P1_U3088) );
  NAND2_X1 U23439 ( .A1(n20506), .A2(n20630), .ZN(n20529) );
  INV_X1 U23440 ( .A(n20507), .ZN(n20530) );
  AOI21_X1 U23441 ( .B1(n20508), .B2(n20776), .A(n20530), .ZN(n20510) );
  OAI22_X1 U23442 ( .A1(n20510), .A2(n20782), .B1(n20509), .B2(n20780), .ZN(
        n20531) );
  AOI22_X1 U23443 ( .A1(n20784), .A2(n20531), .B1(n20530), .B2(n20783), .ZN(
        n20515) );
  OAI21_X1 U23444 ( .B1(n20787), .B2(n20511), .A(n20510), .ZN(n20512) );
  OAI211_X1 U23445 ( .C1(n20791), .C2(n20513), .A(n20789), .B(n20512), .ZN(
        n20532) );
  INV_X1 U23446 ( .A(n20535), .ZN(n20526) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20532), .B1(
        n20526), .B2(n20792), .ZN(n20514) );
  OAI211_X1 U23448 ( .C1(n20795), .C2(n20529), .A(n20515), .B(n20514), .ZN(
        P1_U3089) );
  AOI22_X1 U23449 ( .A1(n20797), .A2(n20531), .B1(n20530), .B2(n20796), .ZN(
        n20517) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20532), .B1(
        n20526), .B2(n20798), .ZN(n20516) );
  OAI211_X1 U23451 ( .C1(n20801), .C2(n20529), .A(n20517), .B(n20516), .ZN(
        P1_U3090) );
  AOI22_X1 U23452 ( .A1(n20803), .A2(n20531), .B1(n20530), .B2(n20802), .ZN(
        n20519) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20532), .B1(
        n20526), .B2(n20804), .ZN(n20518) );
  OAI211_X1 U23454 ( .C1(n20807), .C2(n20529), .A(n20519), .B(n20518), .ZN(
        P1_U3091) );
  AOI22_X1 U23455 ( .A1(n20809), .A2(n20531), .B1(n20530), .B2(n20808), .ZN(
        n20521) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20532), .B1(
        n20558), .B2(n20751), .ZN(n20520) );
  OAI211_X1 U23457 ( .C1(n20754), .C2(n20535), .A(n20521), .B(n20520), .ZN(
        P1_U3092) );
  AOI22_X1 U23458 ( .A1(n21142), .A2(n20531), .B1(n20530), .B2(n21140), .ZN(
        n20523) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20532), .B1(
        n20526), .B2(n21143), .ZN(n20522) );
  OAI211_X1 U23460 ( .C1(n21149), .C2(n20529), .A(n20523), .B(n20522), .ZN(
        P1_U3093) );
  AOI22_X1 U23461 ( .A1(n20817), .A2(n20531), .B1(n20530), .B2(n20816), .ZN(
        n20525) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20532), .B1(
        n20526), .B2(n20818), .ZN(n20524) );
  OAI211_X1 U23463 ( .C1(n20821), .C2(n20529), .A(n20525), .B(n20524), .ZN(
        P1_U3094) );
  AOI22_X1 U23464 ( .A1(n20823), .A2(n20531), .B1(n20530), .B2(n20822), .ZN(
        n20528) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20532), .B1(
        n20526), .B2(n20824), .ZN(n20527) );
  OAI211_X1 U23466 ( .C1(n20827), .C2(n20529), .A(n20528), .B(n20527), .ZN(
        P1_U3095) );
  AOI22_X1 U23467 ( .A1(n20831), .A2(n20531), .B1(n20530), .B2(n20828), .ZN(
        n20534) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20532), .B1(
        n20558), .B2(n20769), .ZN(n20533) );
  OAI211_X1 U23469 ( .C1(n20774), .C2(n20535), .A(n20534), .B(n20533), .ZN(
        P1_U3096) );
  NAND2_X1 U23470 ( .A1(n20536), .A2(n13698), .ZN(n20589) );
  INV_X1 U23471 ( .A(n20589), .ZN(n20634) );
  NAND2_X1 U23472 ( .A1(n20537), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20632) );
  AOI21_X1 U23473 ( .B1(n20634), .B2(n14906), .A(n10077), .ZN(n20540) );
  NAND2_X1 U23474 ( .A1(n20538), .A2(n20591), .ZN(n20672) );
  OAI22_X1 U23475 ( .A1(n20540), .A2(n20782), .B1(n20595), .B2(n20672), .ZN(
        n20557) );
  AOI22_X1 U23476 ( .A1(n20784), .A2(n20557), .B1(n10077), .B2(n20783), .ZN(
        n20544) );
  INV_X1 U23477 ( .A(n20586), .ZN(n20539) );
  OAI21_X1 U23478 ( .B1(n20539), .B2(n20558), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20541) );
  NAND2_X1 U23479 ( .A1(n20541), .A2(n20540), .ZN(n20542) );
  OAI211_X1 U23480 ( .C1(n10077), .C2(n20671), .A(n20593), .B(n20542), .ZN(
        n20559) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20792), .ZN(n20543) );
  OAI211_X1 U23482 ( .C1(n20795), .C2(n20586), .A(n20544), .B(n20543), .ZN(
        P1_U3097) );
  AOI22_X1 U23483 ( .A1(n20797), .A2(n20557), .B1(n10077), .B2(n20796), .ZN(
        n20546) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20798), .ZN(n20545) );
  OAI211_X1 U23485 ( .C1(n20801), .C2(n20586), .A(n20546), .B(n20545), .ZN(
        P1_U3098) );
  AOI22_X1 U23486 ( .A1(n20803), .A2(n20557), .B1(n10077), .B2(n20802), .ZN(
        n20548) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20804), .ZN(n20547) );
  OAI211_X1 U23488 ( .C1(n20807), .C2(n20586), .A(n20548), .B(n20547), .ZN(
        P1_U3099) );
  AOI22_X1 U23489 ( .A1(n20809), .A2(n20557), .B1(n10077), .B2(n20808), .ZN(
        n20550) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20810), .ZN(n20549) );
  OAI211_X1 U23491 ( .C1(n20813), .C2(n20586), .A(n20550), .B(n20549), .ZN(
        P1_U3100) );
  AOI22_X1 U23492 ( .A1(n21142), .A2(n20557), .B1(n10077), .B2(n21140), .ZN(
        n20552) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n21143), .ZN(n20551) );
  OAI211_X1 U23494 ( .C1(n21149), .C2(n20586), .A(n20552), .B(n20551), .ZN(
        P1_U3101) );
  AOI22_X1 U23495 ( .A1(n20817), .A2(n20557), .B1(n10077), .B2(n20816), .ZN(
        n20554) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20818), .ZN(n20553) );
  OAI211_X1 U23497 ( .C1(n20821), .C2(n20586), .A(n20554), .B(n20553), .ZN(
        P1_U3102) );
  AOI22_X1 U23498 ( .A1(n20823), .A2(n20557), .B1(n10077), .B2(n20822), .ZN(
        n20556) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20824), .ZN(n20555) );
  OAI211_X1 U23500 ( .C1(n20827), .C2(n20586), .A(n20556), .B(n20555), .ZN(
        P1_U3103) );
  AOI22_X1 U23501 ( .A1(n20831), .A2(n20557), .B1(n10077), .B2(n20828), .ZN(
        n20561) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20559), .B1(
        n20558), .B2(n20832), .ZN(n20560) );
  OAI211_X1 U23503 ( .C1(n20838), .C2(n20586), .A(n20561), .B(n20560), .ZN(
        P1_U3104) );
  NOR2_X1 U23504 ( .A1(n20632), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20565) );
  INV_X1 U23505 ( .A(n20565), .ZN(n20562) );
  NOR2_X1 U23506 ( .A1(n20701), .A2(n20562), .ZN(n20580) );
  AOI21_X1 U23507 ( .B1(n20634), .B2(n20702), .A(n20580), .ZN(n20563) );
  OAI22_X1 U23508 ( .A1(n20563), .A2(n20782), .B1(n20562), .B2(n20780), .ZN(
        n20581) );
  AOI22_X1 U23509 ( .A1(n20784), .A2(n20581), .B1(n20783), .B2(n20580), .ZN(
        n20567) );
  NOR2_X1 U23510 ( .A1(n20631), .A2(n20782), .ZN(n20637) );
  OAI21_X1 U23511 ( .B1(n20637), .B2(n20705), .A(n20563), .ZN(n20564) );
  OAI211_X1 U23512 ( .C1(n20791), .C2(n20565), .A(n20789), .B(n20564), .ZN(
        n20583) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20739), .ZN(n20566) );
  OAI211_X1 U23514 ( .C1(n20742), .C2(n20586), .A(n20567), .B(n20566), .ZN(
        P1_U3105) );
  AOI22_X1 U23515 ( .A1(n20797), .A2(n20581), .B1(n20796), .B2(n20580), .ZN(
        n20569) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20743), .ZN(n20568) );
  OAI211_X1 U23517 ( .C1(n20746), .C2(n20586), .A(n20569), .B(n20568), .ZN(
        P1_U3106) );
  AOI22_X1 U23518 ( .A1(n20803), .A2(n20581), .B1(n20802), .B2(n20580), .ZN(
        n20571) );
  INV_X1 U23519 ( .A(n20807), .ZN(n20747) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20747), .ZN(n20570) );
  OAI211_X1 U23521 ( .C1(n20750), .C2(n20586), .A(n20571), .B(n20570), .ZN(
        P1_U3107) );
  AOI22_X1 U23522 ( .A1(n20809), .A2(n20581), .B1(n20808), .B2(n20580), .ZN(
        n20573) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20751), .ZN(n20572) );
  OAI211_X1 U23524 ( .C1(n20754), .C2(n20586), .A(n20573), .B(n20572), .ZN(
        P1_U3108) );
  AOI22_X1 U23525 ( .A1(n21142), .A2(n20581), .B1(n21140), .B2(n20580), .ZN(
        n20575) );
  INV_X1 U23526 ( .A(n21149), .ZN(n20755) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20755), .ZN(n20574) );
  OAI211_X1 U23528 ( .C1(n20758), .C2(n20586), .A(n20575), .B(n20574), .ZN(
        P1_U3109) );
  AOI22_X1 U23529 ( .A1(n20817), .A2(n20581), .B1(n20816), .B2(n20580), .ZN(
        n20577) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20759), .ZN(n20576) );
  OAI211_X1 U23531 ( .C1(n20762), .C2(n20586), .A(n20577), .B(n20576), .ZN(
        P1_U3110) );
  AOI22_X1 U23532 ( .A1(n20823), .A2(n20581), .B1(n20822), .B2(n20580), .ZN(
        n20579) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20763), .ZN(n20578) );
  OAI211_X1 U23534 ( .C1(n20766), .C2(n20586), .A(n20579), .B(n20578), .ZN(
        P1_U3111) );
  AOI22_X1 U23535 ( .A1(n20831), .A2(n20581), .B1(n20828), .B2(n20580), .ZN(
        n20585) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20583), .B1(
        n20582), .B2(n20769), .ZN(n20584) );
  OAI211_X1 U23537 ( .C1(n20774), .C2(n20586), .A(n20585), .B(n20584), .ZN(
        P1_U3112) );
  NOR2_X1 U23538 ( .A1(n20779), .A2(n20632), .ZN(n20639) );
  INV_X1 U23539 ( .A(n20639), .ZN(n20635) );
  OR2_X1 U23540 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20635), .ZN(
        n20623) );
  OAI22_X1 U23541 ( .A1(n20624), .A2(n20742), .B1(n20663), .B2(n20623), .ZN(
        n20587) );
  INV_X1 U23542 ( .A(n20587), .ZN(n20599) );
  NAND3_X1 U23543 ( .A1(n20648), .A2(n20624), .A3(n20791), .ZN(n20588) );
  NAND2_X1 U23544 ( .A1(n20588), .A2(n20666), .ZN(n20594) );
  OR2_X1 U23545 ( .A1(n20589), .A2(n14906), .ZN(n20596) );
  AOI22_X1 U23546 ( .A1(n20594), .A2(n20596), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20623), .ZN(n20592) );
  OR2_X1 U23547 ( .A1(n20591), .A2(n20590), .ZN(n20730) );
  NAND2_X1 U23548 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20730), .ZN(n20736) );
  NAND3_X1 U23549 ( .A1(n20593), .A2(n20592), .A3(n20736), .ZN(n20627) );
  INV_X1 U23550 ( .A(n20594), .ZN(n20597) );
  OAI22_X1 U23551 ( .A1(n20597), .A2(n20596), .B1(n20595), .B2(n20730), .ZN(
        n20626) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20627), .B1(
        n20784), .B2(n20626), .ZN(n20598) );
  OAI211_X1 U23553 ( .C1(n20795), .C2(n20648), .A(n20599), .B(n20598), .ZN(
        P1_U3113) );
  OAI22_X1 U23554 ( .A1(n20648), .A2(n20801), .B1(n20623), .B2(n20600), .ZN(
        n20601) );
  INV_X1 U23555 ( .A(n20601), .ZN(n20603) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20627), .B1(
        n20797), .B2(n20626), .ZN(n20602) );
  OAI211_X1 U23557 ( .C1(n20746), .C2(n20624), .A(n20603), .B(n20602), .ZN(
        P1_U3114) );
  OAI22_X1 U23558 ( .A1(n20624), .A2(n20750), .B1(n20623), .B2(n20679), .ZN(
        n20604) );
  INV_X1 U23559 ( .A(n20604), .ZN(n20606) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20627), .B1(
        n20803), .B2(n20626), .ZN(n20605) );
  OAI211_X1 U23561 ( .C1(n20807), .C2(n20648), .A(n20606), .B(n20605), .ZN(
        P1_U3115) );
  OAI22_X1 U23562 ( .A1(n20624), .A2(n20754), .B1(n20623), .B2(n20607), .ZN(
        n20608) );
  INV_X1 U23563 ( .A(n20608), .ZN(n20610) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20627), .B1(
        n20809), .B2(n20626), .ZN(n20609) );
  OAI211_X1 U23565 ( .C1(n20813), .C2(n20648), .A(n20610), .B(n20609), .ZN(
        P1_U3116) );
  OAI22_X1 U23566 ( .A1(n20648), .A2(n21149), .B1(n20623), .B2(n20686), .ZN(
        n20611) );
  INV_X1 U23567 ( .A(n20611), .ZN(n20613) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20627), .B1(
        n21142), .B2(n20626), .ZN(n20612) );
  OAI211_X1 U23569 ( .C1(n20758), .C2(n20624), .A(n20613), .B(n20612), .ZN(
        P1_U3117) );
  OAI22_X1 U23570 ( .A1(n20624), .A2(n20762), .B1(n20623), .B2(n20614), .ZN(
        n20615) );
  INV_X1 U23571 ( .A(n20615), .ZN(n20617) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20627), .B1(
        n20817), .B2(n20626), .ZN(n20616) );
  OAI211_X1 U23573 ( .C1(n20821), .C2(n20648), .A(n20617), .B(n20616), .ZN(
        P1_U3118) );
  OAI22_X1 U23574 ( .A1(n20648), .A2(n20827), .B1(n20623), .B2(n20618), .ZN(
        n20619) );
  INV_X1 U23575 ( .A(n20619), .ZN(n20621) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20627), .B1(
        n20823), .B2(n20626), .ZN(n20620) );
  OAI211_X1 U23577 ( .C1(n20766), .C2(n20624), .A(n20621), .B(n20620), .ZN(
        P1_U3119) );
  OAI22_X1 U23578 ( .A1(n20624), .A2(n20774), .B1(n20623), .B2(n20622), .ZN(
        n20625) );
  INV_X1 U23579 ( .A(n20625), .ZN(n20629) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20627), .B1(
        n20831), .B2(n20626), .ZN(n20628) );
  OAI211_X1 U23581 ( .C1(n20838), .C2(n20648), .A(n20629), .B(n20628), .ZN(
        P1_U3120) );
  NOR2_X1 U23582 ( .A1(n20633), .A2(n20632), .ZN(n20655) );
  AOI21_X1 U23583 ( .B1(n20634), .B2(n20776), .A(n20655), .ZN(n20636) );
  OAI22_X1 U23584 ( .A1(n20636), .A2(n20782), .B1(n20635), .B2(n20780), .ZN(
        n20656) );
  AOI22_X1 U23585 ( .A1(n20784), .A2(n20656), .B1(n20783), .B2(n20655), .ZN(
        n20641) );
  OAI21_X1 U23586 ( .B1(n20787), .B2(n20637), .A(n20636), .ZN(n20638) );
  OAI211_X1 U23587 ( .C1(n20791), .C2(n20639), .A(n20789), .B(n20638), .ZN(
        n20658) );
  INV_X1 U23588 ( .A(n20648), .ZN(n20657) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20792), .ZN(n20640) );
  OAI211_X1 U23590 ( .C1(n20795), .C2(n20699), .A(n20641), .B(n20640), .ZN(
        P1_U3121) );
  AOI22_X1 U23591 ( .A1(n20797), .A2(n20656), .B1(n20796), .B2(n20655), .ZN(
        n20643) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20798), .ZN(n20642) );
  OAI211_X1 U23593 ( .C1(n20801), .C2(n20699), .A(n20643), .B(n20642), .ZN(
        P1_U3122) );
  AOI22_X1 U23594 ( .A1(n20803), .A2(n20656), .B1(n20802), .B2(n20655), .ZN(
        n20645) );
  INV_X1 U23595 ( .A(n20699), .ZN(n20665) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20658), .B1(
        n20665), .B2(n20747), .ZN(n20644) );
  OAI211_X1 U23597 ( .C1(n20750), .C2(n20648), .A(n20645), .B(n20644), .ZN(
        P1_U3123) );
  AOI22_X1 U23598 ( .A1(n20809), .A2(n20656), .B1(n20808), .B2(n20655), .ZN(
        n20647) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20658), .B1(
        n20665), .B2(n20751), .ZN(n20646) );
  OAI211_X1 U23600 ( .C1(n20754), .C2(n20648), .A(n20647), .B(n20646), .ZN(
        P1_U3124) );
  AOI22_X1 U23601 ( .A1(n21142), .A2(n20656), .B1(n21140), .B2(n20655), .ZN(
        n20650) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n21143), .ZN(n20649) );
  OAI211_X1 U23603 ( .C1(n21149), .C2(n20699), .A(n20650), .B(n20649), .ZN(
        P1_U3125) );
  AOI22_X1 U23604 ( .A1(n20817), .A2(n20656), .B1(n20816), .B2(n20655), .ZN(
        n20652) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20818), .ZN(n20651) );
  OAI211_X1 U23606 ( .C1(n20821), .C2(n20699), .A(n20652), .B(n20651), .ZN(
        P1_U3126) );
  AOI22_X1 U23607 ( .A1(n20823), .A2(n20656), .B1(n20822), .B2(n20655), .ZN(
        n20654) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20824), .ZN(n20653) );
  OAI211_X1 U23609 ( .C1(n20827), .C2(n20699), .A(n20654), .B(n20653), .ZN(
        P1_U3127) );
  AOI22_X1 U23610 ( .A1(n20831), .A2(n20656), .B1(n20828), .B2(n20655), .ZN(
        n20660) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20658), .B1(
        n20657), .B2(n20832), .ZN(n20659) );
  OAI211_X1 U23612 ( .C1(n20838), .C2(n20699), .A(n20660), .B(n20659), .ZN(
        P1_U3128) );
  OR2_X1 U23613 ( .A1(n20662), .A2(n20778), .ZN(n20685) );
  NOR2_X1 U23614 ( .A1(n20663), .A2(n20685), .ZN(n20664) );
  AOI21_X1 U23615 ( .B1(n20724), .B2(n20739), .A(n20664), .ZN(n20676) );
  INV_X1 U23616 ( .A(n20685), .ZN(n20694) );
  NOR3_X1 U23617 ( .A1(n20665), .A2(n20724), .A3(n20782), .ZN(n20667) );
  NOR2_X1 U23618 ( .A1(n20667), .A2(n20705), .ZN(n20674) );
  INV_X1 U23619 ( .A(n20674), .ZN(n20669) );
  NOR2_X1 U23620 ( .A1(n13698), .A2(n20668), .ZN(n20777) );
  NAND2_X1 U23621 ( .A1(n20777), .A2(n14906), .ZN(n20673) );
  AOI22_X1 U23622 ( .A1(n20669), .A2(n20673), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20672), .ZN(n20670) );
  OAI211_X1 U23623 ( .C1(n20694), .C2(n20671), .A(n20737), .B(n20670), .ZN(
        n20696) );
  OAI22_X1 U23624 ( .A1(n20674), .A2(n20673), .B1(n20672), .B2(n20729), .ZN(
        n20695) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20696), .B1(
        n20784), .B2(n20695), .ZN(n20675) );
  OAI211_X1 U23626 ( .C1(n20742), .C2(n20699), .A(n20676), .B(n20675), .ZN(
        P1_U3129) );
  AOI22_X1 U23627 ( .A1(n20724), .A2(n20743), .B1(n20796), .B2(n20694), .ZN(
        n20678) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20696), .B1(
        n20797), .B2(n20695), .ZN(n20677) );
  OAI211_X1 U23629 ( .C1(n20746), .C2(n20699), .A(n20678), .B(n20677), .ZN(
        P1_U3130) );
  NOR2_X1 U23630 ( .A1(n20679), .A2(n20685), .ZN(n20680) );
  AOI21_X1 U23631 ( .B1(n20724), .B2(n20747), .A(n20680), .ZN(n20682) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20696), .B1(
        n20803), .B2(n20695), .ZN(n20681) );
  OAI211_X1 U23633 ( .C1(n20750), .C2(n20699), .A(n20682), .B(n20681), .ZN(
        P1_U3131) );
  AOI22_X1 U23634 ( .A1(n20724), .A2(n20751), .B1(n20808), .B2(n20694), .ZN(
        n20684) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20696), .B1(
        n20809), .B2(n20695), .ZN(n20683) );
  OAI211_X1 U23636 ( .C1(n20754), .C2(n20699), .A(n20684), .B(n20683), .ZN(
        P1_U3132) );
  NOR2_X1 U23637 ( .A1(n20686), .A2(n20685), .ZN(n20687) );
  AOI21_X1 U23638 ( .B1(n20724), .B2(n20755), .A(n20687), .ZN(n20689) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20696), .B1(
        n21142), .B2(n20695), .ZN(n20688) );
  OAI211_X1 U23640 ( .C1(n20758), .C2(n20699), .A(n20689), .B(n20688), .ZN(
        P1_U3133) );
  AOI22_X1 U23641 ( .A1(n20724), .A2(n20759), .B1(n20816), .B2(n20694), .ZN(
        n20691) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20696), .B1(
        n20817), .B2(n20695), .ZN(n20690) );
  OAI211_X1 U23643 ( .C1(n20762), .C2(n20699), .A(n20691), .B(n20690), .ZN(
        P1_U3134) );
  AOI22_X1 U23644 ( .A1(n20724), .A2(n20763), .B1(n20822), .B2(n20694), .ZN(
        n20693) );
  AOI22_X1 U23645 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20696), .B1(
        n20823), .B2(n20695), .ZN(n20692) );
  OAI211_X1 U23646 ( .C1(n20766), .C2(n20699), .A(n20693), .B(n20692), .ZN(
        P1_U3135) );
  AOI22_X1 U23647 ( .A1(n20724), .A2(n20769), .B1(n20828), .B2(n20694), .ZN(
        n20698) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20696), .B1(
        n20831), .B2(n20695), .ZN(n20697) );
  OAI211_X1 U23649 ( .C1(n20774), .C2(n20699), .A(n20698), .B(n20697), .ZN(
        P1_U3136) );
  NOR3_X2 U23650 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20701), .A3(
        n20778), .ZN(n20722) );
  AOI21_X1 U23651 ( .B1(n20777), .B2(n20702), .A(n20722), .ZN(n20704) );
  NOR2_X1 U23652 ( .A1(n20778), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20707) );
  INV_X1 U23653 ( .A(n20707), .ZN(n20703) );
  OAI22_X1 U23654 ( .A1(n20704), .A2(n20782), .B1(n20703), .B2(n20780), .ZN(
        n20723) );
  AOI22_X1 U23655 ( .A1(n20784), .A2(n20723), .B1(n20783), .B2(n20722), .ZN(
        n20709) );
  NOR2_X1 U23656 ( .A1(n20732), .A2(n20782), .ZN(n20786) );
  OAI21_X1 U23657 ( .B1(n20786), .B2(n20705), .A(n20704), .ZN(n20706) );
  OAI211_X1 U23658 ( .C1(n20791), .C2(n20707), .A(n20789), .B(n20706), .ZN(
        n20725) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20792), .ZN(n20708) );
  OAI211_X1 U23660 ( .C1(n20795), .C2(n20773), .A(n20709), .B(n20708), .ZN(
        P1_U3137) );
  AOI22_X1 U23661 ( .A1(n20797), .A2(n20723), .B1(n20796), .B2(n20722), .ZN(
        n20711) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20798), .ZN(n20710) );
  OAI211_X1 U23663 ( .C1(n20801), .C2(n20773), .A(n20711), .B(n20710), .ZN(
        P1_U3138) );
  AOI22_X1 U23664 ( .A1(n20803), .A2(n20723), .B1(n20802), .B2(n20722), .ZN(
        n20713) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20804), .ZN(n20712) );
  OAI211_X1 U23666 ( .C1(n20807), .C2(n20773), .A(n20713), .B(n20712), .ZN(
        P1_U3139) );
  AOI22_X1 U23667 ( .A1(n20809), .A2(n20723), .B1(n20808), .B2(n20722), .ZN(
        n20715) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20810), .ZN(n20714) );
  OAI211_X1 U23669 ( .C1(n20813), .C2(n20773), .A(n20715), .B(n20714), .ZN(
        P1_U3140) );
  AOI22_X1 U23670 ( .A1(n21142), .A2(n20723), .B1(n21140), .B2(n20722), .ZN(
        n20717) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n21143), .ZN(n20716) );
  OAI211_X1 U23672 ( .C1(n21149), .C2(n20773), .A(n20717), .B(n20716), .ZN(
        P1_U3141) );
  AOI22_X1 U23673 ( .A1(n20817), .A2(n20723), .B1(n20816), .B2(n20722), .ZN(
        n20719) );
  AOI22_X1 U23674 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20818), .ZN(n20718) );
  OAI211_X1 U23675 ( .C1(n20821), .C2(n20773), .A(n20719), .B(n20718), .ZN(
        P1_U3142) );
  AOI22_X1 U23676 ( .A1(n20823), .A2(n20723), .B1(n20822), .B2(n20722), .ZN(
        n20721) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20824), .ZN(n20720) );
  OAI211_X1 U23678 ( .C1(n20827), .C2(n20773), .A(n20721), .B(n20720), .ZN(
        P1_U3143) );
  AOI22_X1 U23679 ( .A1(n20831), .A2(n20723), .B1(n20828), .B2(n20722), .ZN(
        n20727) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20725), .B1(
        n20724), .B2(n20832), .ZN(n20726) );
  OAI211_X1 U23681 ( .C1(n20838), .C2(n20773), .A(n20727), .B(n20726), .ZN(
        P1_U3144) );
  NAND2_X1 U23682 ( .A1(n20777), .A2(n20728), .ZN(n20734) );
  OAI22_X1 U23683 ( .A1(n20734), .A2(n20782), .B1(n20730), .B2(n20729), .ZN(
        n20768) );
  NOR3_X2 U23684 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20779), .A3(
        n20778), .ZN(n20767) );
  AOI22_X1 U23685 ( .A1(n20784), .A2(n20768), .B1(n20783), .B2(n20767), .ZN(
        n20741) );
  INV_X1 U23686 ( .A(n20773), .ZN(n20733) );
  OAI21_X1 U23687 ( .B1(n20733), .B2(n20833), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20735) );
  AOI21_X1 U23688 ( .B1(n20735), .B2(n20734), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20738) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20739), .ZN(n20740) );
  OAI211_X1 U23690 ( .C1(n20742), .C2(n20773), .A(n20741), .B(n20740), .ZN(
        P1_U3145) );
  AOI22_X1 U23691 ( .A1(n20797), .A2(n20768), .B1(n20796), .B2(n20767), .ZN(
        n20745) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20743), .ZN(n20744) );
  OAI211_X1 U23693 ( .C1(n20746), .C2(n20773), .A(n20745), .B(n20744), .ZN(
        P1_U3146) );
  AOI22_X1 U23694 ( .A1(n20803), .A2(n20768), .B1(n20802), .B2(n20767), .ZN(
        n20749) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20747), .ZN(n20748) );
  OAI211_X1 U23696 ( .C1(n20750), .C2(n20773), .A(n20749), .B(n20748), .ZN(
        P1_U3147) );
  AOI22_X1 U23697 ( .A1(n20809), .A2(n20768), .B1(n20808), .B2(n20767), .ZN(
        n20753) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20751), .ZN(n20752) );
  OAI211_X1 U23699 ( .C1(n20754), .C2(n20773), .A(n20753), .B(n20752), .ZN(
        P1_U3148) );
  AOI22_X1 U23700 ( .A1(n21142), .A2(n20768), .B1(n21140), .B2(n20767), .ZN(
        n20757) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20755), .ZN(n20756) );
  OAI211_X1 U23702 ( .C1(n20758), .C2(n20773), .A(n20757), .B(n20756), .ZN(
        P1_U3149) );
  AOI22_X1 U23703 ( .A1(n20817), .A2(n20768), .B1(n20816), .B2(n20767), .ZN(
        n20761) );
  AOI22_X1 U23704 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20759), .ZN(n20760) );
  OAI211_X1 U23705 ( .C1(n20762), .C2(n20773), .A(n20761), .B(n20760), .ZN(
        P1_U3150) );
  AOI22_X1 U23706 ( .A1(n20823), .A2(n20768), .B1(n20822), .B2(n20767), .ZN(
        n20765) );
  AOI22_X1 U23707 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20763), .ZN(n20764) );
  OAI211_X1 U23708 ( .C1(n20766), .C2(n20773), .A(n20765), .B(n20764), .ZN(
        P1_U3151) );
  AOI22_X1 U23709 ( .A1(n20831), .A2(n20768), .B1(n20828), .B2(n20767), .ZN(
        n20772) );
  AOI22_X1 U23710 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20770), .B1(
        n20833), .B2(n20769), .ZN(n20771) );
  OAI211_X1 U23711 ( .C1(n20774), .C2(n20773), .A(n20772), .B(n20771), .ZN(
        P1_U3152) );
  INV_X1 U23712 ( .A(n20775), .ZN(n20829) );
  AOI21_X1 U23713 ( .B1(n20777), .B2(n20776), .A(n20829), .ZN(n20785) );
  NOR2_X1 U23714 ( .A1(n20779), .A2(n20778), .ZN(n20790) );
  INV_X1 U23715 ( .A(n20790), .ZN(n20781) );
  OAI22_X1 U23716 ( .A1(n20785), .A2(n20782), .B1(n20781), .B2(n20780), .ZN(
        n20830) );
  AOI22_X1 U23717 ( .A1(n20784), .A2(n20830), .B1(n20829), .B2(n20783), .ZN(
        n20794) );
  OAI21_X1 U23718 ( .B1(n20787), .B2(n20786), .A(n20785), .ZN(n20788) );
  OAI211_X1 U23719 ( .C1(n20791), .C2(n20790), .A(n20789), .B(n20788), .ZN(
        n20834) );
  AOI22_X1 U23720 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n20792), .ZN(n20793) );
  OAI211_X1 U23721 ( .C1(n20795), .C2(n20837), .A(n20794), .B(n20793), .ZN(
        P1_U3153) );
  AOI22_X1 U23722 ( .A1(n20797), .A2(n20830), .B1(n20829), .B2(n20796), .ZN(
        n20800) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n20798), .ZN(n20799) );
  OAI211_X1 U23724 ( .C1(n20801), .C2(n20837), .A(n20800), .B(n20799), .ZN(
        P1_U3154) );
  AOI22_X1 U23725 ( .A1(n20803), .A2(n20830), .B1(n20829), .B2(n20802), .ZN(
        n20806) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n20804), .ZN(n20805) );
  OAI211_X1 U23727 ( .C1(n20807), .C2(n20837), .A(n20806), .B(n20805), .ZN(
        P1_U3155) );
  AOI22_X1 U23728 ( .A1(n20809), .A2(n20830), .B1(n20829), .B2(n20808), .ZN(
        n20812) );
  AOI22_X1 U23729 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n20810), .ZN(n20811) );
  OAI211_X1 U23730 ( .C1(n20813), .C2(n20837), .A(n20812), .B(n20811), .ZN(
        P1_U3156) );
  AOI22_X1 U23731 ( .A1(n21142), .A2(n20830), .B1(n20829), .B2(n21140), .ZN(
        n20815) );
  AOI22_X1 U23732 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n21143), .ZN(n20814) );
  OAI211_X1 U23733 ( .C1(n21149), .C2(n20837), .A(n20815), .B(n20814), .ZN(
        P1_U3157) );
  AOI22_X1 U23734 ( .A1(n20817), .A2(n20830), .B1(n20829), .B2(n20816), .ZN(
        n20820) );
  AOI22_X1 U23735 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n20818), .ZN(n20819) );
  OAI211_X1 U23736 ( .C1(n20821), .C2(n20837), .A(n20820), .B(n20819), .ZN(
        P1_U3158) );
  AOI22_X1 U23737 ( .A1(n20823), .A2(n20830), .B1(n20829), .B2(n20822), .ZN(
        n20826) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n20824), .ZN(n20825) );
  OAI211_X1 U23739 ( .C1(n20827), .C2(n20837), .A(n20826), .B(n20825), .ZN(
        P1_U3159) );
  AOI22_X1 U23740 ( .A1(n20831), .A2(n20830), .B1(n20829), .B2(n20828), .ZN(
        n20836) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20834), .B1(
        n20833), .B2(n20832), .ZN(n20835) );
  OAI211_X1 U23742 ( .C1(n20838), .C2(n20837), .A(n20836), .B(n20835), .ZN(
        P1_U3160) );
  NAND2_X1 U23743 ( .A1(n20840), .A2(n20839), .ZN(P1_U3163) );
  AND2_X1 U23744 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20917), .ZN(
        P1_U3164) );
  AND2_X1 U23745 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20917), .ZN(
        P1_U3165) );
  AND2_X1 U23746 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20917), .ZN(
        P1_U3166) );
  AND2_X1 U23747 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20917), .ZN(
        P1_U3167) );
  AND2_X1 U23748 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20917), .ZN(
        P1_U3168) );
  AND2_X1 U23749 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20917), .ZN(
        P1_U3169) );
  AND2_X1 U23750 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20917), .ZN(
        P1_U3170) );
  AND2_X1 U23751 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20917), .ZN(
        P1_U3171) );
  AND2_X1 U23752 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20917), .ZN(
        P1_U3172) );
  AND2_X1 U23753 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20917), .ZN(
        P1_U3173) );
  AND2_X1 U23754 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20917), .ZN(
        P1_U3174) );
  AND2_X1 U23755 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20917), .ZN(
        P1_U3175) );
  AND2_X1 U23756 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20917), .ZN(
        P1_U3176) );
  AND2_X1 U23757 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20917), .ZN(
        P1_U3177) );
  AND2_X1 U23758 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20917), .ZN(
        P1_U3178) );
  AND2_X1 U23759 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20917), .ZN(
        P1_U3179) );
  AND2_X1 U23760 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20917), .ZN(
        P1_U3180) );
  AND2_X1 U23761 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20917), .ZN(
        P1_U3181) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20917), .ZN(
        P1_U3182) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20917), .ZN(
        P1_U3183) );
  AND2_X1 U23764 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20917), .ZN(
        P1_U3184) );
  AND2_X1 U23765 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20917), .ZN(
        P1_U3185) );
  INV_X1 U23766 ( .A(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20952) );
  NOR2_X1 U23767 ( .A1(n20921), .A2(n20952), .ZN(P1_U3186) );
  AND2_X1 U23768 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20917), .ZN(P1_U3187) );
  AND2_X1 U23769 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20917), .ZN(P1_U3188) );
  AND2_X1 U23770 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20917), .ZN(P1_U3189) );
  AND2_X1 U23771 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20917), .ZN(P1_U3190) );
  AND2_X1 U23772 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20917), .ZN(P1_U3191) );
  AND2_X1 U23773 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20917), .ZN(P1_U3192) );
  AND2_X1 U23774 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20917), .ZN(P1_U3193) );
  NAND2_X1 U23775 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20848), .ZN(n20851) );
  INV_X1 U23776 ( .A(n20851), .ZN(n20844) );
  NAND2_X1 U23777 ( .A1(n20852), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20847) );
  AOI22_X1 U23778 ( .A1(HOLD), .A2(n20842), .B1(n20847), .B2(n20841), .ZN(
        n20843) );
  OAI22_X1 U23779 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20844), .B1(n20942), 
        .B2(n20843), .ZN(P1_U3194) );
  INV_X1 U23780 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20845) );
  OAI21_X1 U23781 ( .B1(n20845), .B2(P1_STATE_REG_2__SCAN_IN), .A(HOLD), .ZN(
        n20846) );
  OAI21_X1 U23782 ( .B1(n20848), .B2(n20847), .A(n20846), .ZN(n20849) );
  INV_X1 U23783 ( .A(n20849), .ZN(n20856) );
  NAND3_X1 U23784 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20850), .A3(n20852), 
        .ZN(n20854) );
  OAI211_X1 U23785 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20852), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20851), .ZN(n20853) );
  OAI221_X1 U23786 ( .B1(n20856), .B2(n20855), .C1(n20856), .C2(n20854), .A(
        n20853), .ZN(P1_U3196) );
  NAND2_X1 U23787 ( .A1(n20942), .A2(n20857), .ZN(n20908) );
  NAND2_X1 U23788 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20942), .ZN(n20904) );
  OAI222_X1 U23789 ( .A1(n20908), .A2(n20078), .B1(n20858), .B2(n20942), .C1(
        n20243), .C2(n20904), .ZN(P1_U3197) );
  INV_X1 U23790 ( .A(n20904), .ZN(n20906) );
  INV_X1 U23791 ( .A(n20908), .ZN(n20902) );
  AOI222_X1 U23792 ( .A1(n20906), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20928), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20902), .ZN(n20859) );
  INV_X1 U23793 ( .A(n20859), .ZN(P1_U3198) );
  AOI222_X1 U23794 ( .A1(n20906), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20928), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20902), .ZN(n20860) );
  INV_X1 U23795 ( .A(n20860), .ZN(P1_U3199) );
  AOI22_X1 U23796 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20928), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20902), .ZN(n20861) );
  OAI21_X1 U23797 ( .B1(n20862), .B2(n20904), .A(n20861), .ZN(P1_U3200) );
  AOI22_X1 U23798 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20928), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20906), .ZN(n20863) );
  OAI21_X1 U23799 ( .B1(n20865), .B2(n20908), .A(n20863), .ZN(P1_U3201) );
  INV_X1 U23800 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20864) );
  OAI222_X1 U23801 ( .A1(n20904), .A2(n20865), .B1(n20864), .B2(n20942), .C1(
        n20867), .C2(n20908), .ZN(P1_U3202) );
  INV_X1 U23802 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20866) );
  OAI222_X1 U23803 ( .A1(n20904), .A2(n20867), .B1(n20866), .B2(n20942), .C1(
        n14095), .C2(n20908), .ZN(P1_U3203) );
  INV_X1 U23804 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20868) );
  OAI222_X1 U23805 ( .A1(n20908), .A2(n20870), .B1(n20868), .B2(n20942), .C1(
        n14095), .C2(n20904), .ZN(P1_U3204) );
  INV_X1 U23806 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20869) );
  INV_X1 U23807 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20871) );
  OAI222_X1 U23808 ( .A1(n20904), .A2(n20870), .B1(n20869), .B2(n20942), .C1(
        n20871), .C2(n20908), .ZN(P1_U3205) );
  INV_X1 U23809 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20872) );
  OAI222_X1 U23810 ( .A1(n20908), .A2(n20873), .B1(n20872), .B2(n20942), .C1(
        n20871), .C2(n20904), .ZN(P1_U3206) );
  AOI222_X1 U23811 ( .A1(n20906), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20928), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20902), .ZN(n20874) );
  INV_X1 U23812 ( .A(n20874), .ZN(P1_U3207) );
  AOI222_X1 U23813 ( .A1(n20906), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20928), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20902), .ZN(n20875) );
  INV_X1 U23814 ( .A(n20875), .ZN(P1_U3208) );
  AOI22_X1 U23815 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20928), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20902), .ZN(n20876) );
  OAI21_X1 U23816 ( .B1(n20877), .B2(n20904), .A(n20876), .ZN(P1_U3209) );
  AOI22_X1 U23817 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20893), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20906), .ZN(n20878) );
  OAI21_X1 U23818 ( .B1(n20880), .B2(n20908), .A(n20878), .ZN(P1_U3210) );
  AOI22_X1 U23819 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20893), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20902), .ZN(n20879) );
  OAI21_X1 U23820 ( .B1(n20880), .B2(n20904), .A(n20879), .ZN(P1_U3211) );
  AOI22_X1 U23821 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20893), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20906), .ZN(n20881) );
  OAI21_X1 U23822 ( .B1(n20883), .B2(n20908), .A(n20881), .ZN(P1_U3212) );
  INV_X1 U23823 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20882) );
  OAI222_X1 U23824 ( .A1(n20904), .A2(n20883), .B1(n20882), .B2(n20942), .C1(
        n20884), .C2(n20908), .ZN(P1_U3213) );
  INV_X1 U23825 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20885) );
  OAI222_X1 U23826 ( .A1(n20908), .A2(n20887), .B1(n20885), .B2(n20942), .C1(
        n20884), .C2(n20904), .ZN(P1_U3214) );
  AOI22_X1 U23827 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20893), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20902), .ZN(n20886) );
  OAI21_X1 U23828 ( .B1(n20887), .B2(n20904), .A(n20886), .ZN(P1_U3215) );
  AOI22_X1 U23829 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20893), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20906), .ZN(n20888) );
  OAI21_X1 U23830 ( .B1(n20890), .B2(n20908), .A(n20888), .ZN(P1_U3216) );
  INV_X1 U23831 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20889) );
  OAI222_X1 U23832 ( .A1(n20904), .A2(n20890), .B1(n20889), .B2(n20942), .C1(
        n20892), .C2(n20908), .ZN(P1_U3217) );
  AOI22_X1 U23833 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20893), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20902), .ZN(n20891) );
  OAI21_X1 U23834 ( .B1(n20892), .B2(n20904), .A(n20891), .ZN(P1_U3218) );
  AOI22_X1 U23835 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20893), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20906), .ZN(n20894) );
  OAI21_X1 U23836 ( .B1(n14704), .B2(n20908), .A(n20894), .ZN(P1_U3219) );
  INV_X1 U23837 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20895) );
  OAI222_X1 U23838 ( .A1(n20904), .A2(n14704), .B1(n20895), .B2(n20942), .C1(
        n20897), .C2(n20908), .ZN(P1_U3220) );
  AOI22_X1 U23839 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20902), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20928), .ZN(n20896) );
  OAI21_X1 U23840 ( .B1(n20897), .B2(n20904), .A(n20896), .ZN(P1_U3221) );
  INV_X1 U23841 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20900) );
  AOI22_X1 U23842 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20906), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20928), .ZN(n20898) );
  OAI21_X1 U23843 ( .B1(n20900), .B2(n20908), .A(n20898), .ZN(P1_U3222) );
  AOI22_X1 U23844 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20902), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20928), .ZN(n20899) );
  OAI21_X1 U23845 ( .B1(n20900), .B2(n20904), .A(n20899), .ZN(P1_U3223) );
  AOI22_X1 U23846 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20906), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20928), .ZN(n20901) );
  OAI21_X1 U23847 ( .B1(n20905), .B2(n20908), .A(n20901), .ZN(P1_U3224) );
  AOI22_X1 U23848 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20902), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20928), .ZN(n20903) );
  OAI21_X1 U23849 ( .B1(n20905), .B2(n20904), .A(n20903), .ZN(P1_U3225) );
  AOI22_X1 U23850 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20906), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20928), .ZN(n20907) );
  OAI21_X1 U23851 ( .B1(n20909), .B2(n20908), .A(n20907), .ZN(P1_U3226) );
  INV_X1 U23852 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20910) );
  AOI22_X1 U23853 ( .A1(n20942), .A2(n20911), .B1(n20910), .B2(n20928), .ZN(
        P1_U3458) );
  INV_X1 U23854 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20953) );
  INV_X1 U23855 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20912) );
  AOI22_X1 U23856 ( .A1(n20942), .A2(n20953), .B1(n20912), .B2(n20928), .ZN(
        P1_U3459) );
  INV_X1 U23857 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20913) );
  AOI22_X1 U23858 ( .A1(n20942), .A2(n20914), .B1(n20913), .B2(n20928), .ZN(
        P1_U3460) );
  INV_X1 U23859 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20926) );
  INV_X1 U23860 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20915) );
  AOI22_X1 U23861 ( .A1(n20942), .A2(n20926), .B1(n20915), .B2(n20928), .ZN(
        P1_U3461) );
  INV_X1 U23862 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20918) );
  INV_X1 U23863 ( .A(n20919), .ZN(n20916) );
  AOI21_X1 U23864 ( .B1(n20918), .B2(n20917), .A(n20916), .ZN(P1_U3464) );
  OAI21_X1 U23865 ( .B1(n20921), .B2(n20920), .A(n20919), .ZN(P1_U3465) );
  AOI21_X1 U23866 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20922) );
  AOI22_X1 U23867 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20922), .B2(n20243), .ZN(n20924) );
  AOI22_X1 U23868 ( .A1(n20927), .A2(n20924), .B1(n20953), .B2(n20923), .ZN(
        P1_U3481) );
  OAI21_X1 U23869 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20927), .ZN(n20925) );
  OAI21_X1 U23870 ( .B1(n20927), .B2(n20926), .A(n20925), .ZN(P1_U3482) );
  AOI22_X1 U23871 ( .A1(n20942), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20929), 
        .B2(n20928), .ZN(P1_U3483) );
  NAND2_X1 U23872 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20930), .ZN(n20933) );
  INV_X1 U23873 ( .A(n20931), .ZN(n20932) );
  OAI21_X1 U23874 ( .B1(n20934), .B2(n20933), .A(n20932), .ZN(n20941) );
  AOI211_X1 U23875 ( .C1(n20938), .C2(n20937), .A(n20936), .B(n20935), .ZN(
        n20940) );
  NAND2_X1 U23876 ( .A1(n20940), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20939) );
  OAI21_X1 U23877 ( .B1(n20941), .B2(n20940), .A(n20939), .ZN(P1_U3485) );
  MUX2_X1 U23878 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20942), .Z(P1_U3486) );
  OAI22_X1 U23879 ( .A1(n20945), .A2(keyinput96), .B1(n20944), .B2(keyinput88), 
        .ZN(n20943) );
  AOI221_X1 U23880 ( .B1(n20945), .B2(keyinput96), .C1(keyinput88), .C2(n20944), .A(n20943), .ZN(n20957) );
  OAI22_X1 U23881 ( .A1(n20947), .A2(keyinput80), .B1(n21061), .B2(keyinput119), .ZN(n20946) );
  AOI221_X1 U23882 ( .B1(n20947), .B2(keyinput80), .C1(keyinput119), .C2(
        n21061), .A(n20946), .ZN(n20956) );
  OAI22_X1 U23883 ( .A1(n20950), .A2(keyinput127), .B1(n20949), .B2(
        keyinput117), .ZN(n20948) );
  AOI221_X1 U23884 ( .B1(n20950), .B2(keyinput127), .C1(keyinput117), .C2(
        n20949), .A(n20948), .ZN(n20955) );
  OAI22_X1 U23885 ( .A1(n20953), .A2(keyinput108), .B1(n20952), .B2(
        keyinput120), .ZN(n20951) );
  AOI221_X1 U23886 ( .B1(n20953), .B2(keyinput108), .C1(keyinput120), .C2(
        n20952), .A(n20951), .ZN(n20954) );
  NAND4_X1 U23887 ( .A1(n20957), .A2(n20956), .A3(n20955), .A4(n20954), .ZN(
        n20992) );
  AOI22_X1 U23888 ( .A1(n21056), .A2(keyinput93), .B1(n21096), .B2(keyinput97), 
        .ZN(n20958) );
  OAI221_X1 U23889 ( .B1(n21056), .B2(keyinput93), .C1(n21096), .C2(keyinput97), .A(n20958), .ZN(n20962) );
  XOR2_X1 U23890 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B(keyinput68), .Z(
        n20961) );
  XNOR2_X1 U23891 ( .A(n20959), .B(keyinput112), .ZN(n20960) );
  OR3_X1 U23892 ( .A1(n20962), .A2(n20961), .A3(n20960), .ZN(n20969) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(keyinput66), 
        .B1(n21120), .B2(keyinput71), .ZN(n20963) );
  OAI221_X1 U23894 ( .B1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput66), 
        .C1(n21120), .C2(keyinput71), .A(n20963), .ZN(n20968) );
  AOI22_X1 U23895 ( .A1(n20966), .A2(keyinput74), .B1(keyinput79), .B2(n20965), 
        .ZN(n20964) );
  OAI221_X1 U23896 ( .B1(n20966), .B2(keyinput74), .C1(n20965), .C2(keyinput79), .A(n20964), .ZN(n20967) );
  OR3_X1 U23897 ( .A1(n20969), .A2(n20968), .A3(n20967), .ZN(n20991) );
  OAI22_X1 U23898 ( .A1(n9979), .A2(keyinput81), .B1(n15060), .B2(keyinput103), 
        .ZN(n20970) );
  AOI221_X1 U23899 ( .B1(n9979), .B2(keyinput81), .C1(keyinput103), .C2(n15060), .A(n20970), .ZN(n20978) );
  INV_X1 U23900 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21092) );
  OAI22_X1 U23901 ( .A1(n9976), .A2(keyinput126), .B1(n21092), .B2(keyinput76), 
        .ZN(n20971) );
  AOI221_X1 U23902 ( .B1(n9976), .B2(keyinput126), .C1(keyinput76), .C2(n21092), .A(n20971), .ZN(n20977) );
  OAI22_X1 U23903 ( .A1(n21126), .A2(keyinput99), .B1(n20973), .B2(keyinput110), .ZN(n20972) );
  AOI221_X1 U23904 ( .B1(n21126), .B2(keyinput99), .C1(keyinput110), .C2(
        n20973), .A(n20972), .ZN(n20976) );
  OAI22_X1 U23905 ( .A1(n21090), .A2(keyinput87), .B1(n21075), .B2(keyinput92), 
        .ZN(n20974) );
  AOI221_X1 U23906 ( .B1(n21090), .B2(keyinput87), .C1(keyinput92), .C2(n21075), .A(n20974), .ZN(n20975) );
  NAND4_X1 U23907 ( .A1(n20978), .A2(n20977), .A3(n20976), .A4(n20975), .ZN(
        n20990) );
  OAI22_X1 U23908 ( .A1(n21087), .A2(keyinput78), .B1(n21086), .B2(keyinput118), .ZN(n20979) );
  AOI221_X1 U23909 ( .B1(n21087), .B2(keyinput78), .C1(keyinput118), .C2(
        n21086), .A(n20979), .ZN(n20988) );
  INV_X1 U23910 ( .A(DATAI_26_), .ZN(n20981) );
  OAI22_X1 U23911 ( .A1(n20981), .A2(keyinput67), .B1(n21125), .B2(keyinput84), 
        .ZN(n20980) );
  AOI221_X1 U23912 ( .B1(n20981), .B2(keyinput67), .C1(keyinput84), .C2(n21125), .A(n20980), .ZN(n20987) );
  OAI22_X1 U23913 ( .A1(n21117), .A2(keyinput82), .B1(n20983), .B2(keyinput125), .ZN(n20982) );
  AOI221_X1 U23914 ( .B1(n21117), .B2(keyinput82), .C1(keyinput125), .C2(
        n20983), .A(n20982), .ZN(n20986) );
  INV_X1 U23915 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n21102) );
  OAI22_X1 U23916 ( .A1(n12752), .A2(keyinput109), .B1(n21102), .B2(
        keyinput111), .ZN(n20984) );
  AOI221_X1 U23917 ( .B1(n12752), .B2(keyinput109), .C1(keyinput111), .C2(
        n21102), .A(n20984), .ZN(n20985) );
  NAND4_X1 U23918 ( .A1(n20988), .A2(n20987), .A3(n20986), .A4(n20985), .ZN(
        n20989) );
  NOR4_X1 U23919 ( .A1(n20992), .A2(n20991), .A3(n20990), .A4(n20989), .ZN(
        n21138) );
  OAI22_X1 U23920 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(keyinput123), 
        .B1(keyinput73), .B2(P3_REIP_REG_28__SCAN_IN), .ZN(n20993) );
  AOI221_X1 U23921 ( .B1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput123), 
        .C1(P3_REIP_REG_28__SCAN_IN), .C2(keyinput73), .A(n20993), .ZN(n21000)
         );
  OAI22_X1 U23922 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(keyinput100), 
        .B1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput98), .ZN(n20994) );
  AOI221_X1 U23923 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput100), 
        .C1(keyinput98), .C2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A(n20994), .ZN(
        n20999) );
  OAI22_X1 U23924 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(keyinput107), .B1(
        keyinput121), .B2(P1_EBX_REG_4__SCAN_IN), .ZN(n20995) );
  AOI221_X1 U23925 ( .B1(P2_REIP_REG_30__SCAN_IN), .B2(keyinput107), .C1(
        P1_EBX_REG_4__SCAN_IN), .C2(keyinput121), .A(n20995), .ZN(n20998) );
  OAI22_X1 U23926 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput101), 
        .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput77), .ZN(n20996) );
  AOI221_X1 U23927 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput101), 
        .C1(keyinput77), .C2(P3_BYTEENABLE_REG_2__SCAN_IN), .A(n20996), .ZN(
        n20997) );
  NAND4_X1 U23928 ( .A1(n21000), .A2(n20999), .A3(n20998), .A4(n20997), .ZN(
        n21028) );
  OAI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(keyinput113), 
        .B1(keyinput95), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n21001) );
  AOI221_X1 U23930 ( .B1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B2(keyinput113), 
        .C1(P3_REIP_REG_12__SCAN_IN), .C2(keyinput95), .A(n21001), .ZN(n21008)
         );
  OAI22_X1 U23931 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(keyinput65), 
        .B1(P1_DATAO_REG_12__SCAN_IN), .B2(keyinput83), .ZN(n21002) );
  AOI221_X1 U23932 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput65), 
        .C1(keyinput83), .C2(P1_DATAO_REG_12__SCAN_IN), .A(n21002), .ZN(n21007) );
  OAI22_X1 U23933 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(keyinput86), .B1(
        P1_INSTQUEUE_REG_11__7__SCAN_IN), .B2(keyinput91), .ZN(n21003) );
  AOI221_X1 U23934 ( .B1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput86), 
        .C1(keyinput91), .C2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(n21003), 
        .ZN(n21006) );
  OAI22_X1 U23935 ( .A1(BUF1_REG_23__SCAN_IN), .A2(keyinput116), .B1(
        BUF2_REG_1__SCAN_IN), .B2(keyinput105), .ZN(n21004) );
  AOI221_X1 U23936 ( .B1(BUF1_REG_23__SCAN_IN), .B2(keyinput116), .C1(
        keyinput105), .C2(BUF2_REG_1__SCAN_IN), .A(n21004), .ZN(n21005) );
  NAND4_X1 U23937 ( .A1(n21008), .A2(n21007), .A3(n21006), .A4(n21005), .ZN(
        n21027) );
  OAI22_X1 U23938 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput115), 
        .B1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput102), .ZN(n21009)
         );
  AOI221_X1 U23939 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput115), 
        .C1(keyinput102), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(n21009), 
        .ZN(n21016) );
  OAI22_X1 U23940 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(keyinput114), .B1(
        keyinput106), .B2(READY2), .ZN(n21010) );
  AOI221_X1 U23941 ( .B1(P1_EBX_REG_0__SCAN_IN), .B2(keyinput114), .C1(READY2), 
        .C2(keyinput106), .A(n21010), .ZN(n21015) );
  OAI22_X1 U23942 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(keyinput124), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(keyinput90), .ZN(n21011) );
  AOI221_X1 U23943 ( .B1(P2_ADDRESS_REG_25__SCAN_IN), .B2(keyinput124), .C1(
        keyinput90), .C2(P3_ADDRESS_REG_14__SCAN_IN), .A(n21011), .ZN(n21014)
         );
  OAI22_X1 U23944 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(keyinput94), 
        .B1(P3_UWORD_REG_9__SCAN_IN), .B2(keyinput64), .ZN(n21012) );
  AOI221_X1 U23945 ( .B1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(keyinput94), 
        .C1(keyinput64), .C2(P3_UWORD_REG_9__SCAN_IN), .A(n21012), .ZN(n21013)
         );
  NAND4_X1 U23946 ( .A1(n21016), .A2(n21015), .A3(n21014), .A4(n21013), .ZN(
        n21026) );
  OAI22_X1 U23947 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(keyinput75), .B1(
        P3_INSTQUEUE_REG_15__0__SCAN_IN), .B2(keyinput122), .ZN(n21017) );
  AOI221_X1 U23948 ( .B1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(keyinput75), 
        .C1(keyinput122), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(n21017), 
        .ZN(n21024) );
  OAI22_X1 U23949 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(keyinput72), 
        .B1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B2(keyinput104), .ZN(n21018) );
  AOI221_X1 U23950 ( .B1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B2(keyinput72), 
        .C1(keyinput104), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(n21018), 
        .ZN(n21023) );
  OAI22_X1 U23951 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(keyinput89), .B1(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput69), .ZN(n21019) );
  AOI221_X1 U23952 ( .B1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B2(keyinput89), 
        .C1(keyinput69), .C2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(n21019), 
        .ZN(n21022) );
  OAI22_X1 U23953 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(keyinput85), 
        .B1(P3_DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput70), .ZN(n21020) );
  AOI221_X1 U23954 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput85), 
        .C1(keyinput70), .C2(P3_DATAWIDTH_REG_12__SCAN_IN), .A(n21020), .ZN(
        n21021) );
  NAND4_X1 U23955 ( .A1(n21024), .A2(n21023), .A3(n21022), .A4(n21021), .ZN(
        n21025) );
  NOR4_X1 U23956 ( .A1(n21028), .A2(n21027), .A3(n21026), .A4(n21025), .ZN(
        n21137) );
  AOI22_X1 U23957 ( .A1(DATAI_26_), .A2(keyinput3), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput1), .ZN(n21029) );
  OAI221_X1 U23958 ( .B1(DATAI_26_), .B2(keyinput3), .C1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(keyinput1), .A(n21029), .ZN(
        n21036) );
  AOI22_X1 U23959 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(keyinput16), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput36), .ZN(n21030) );
  OAI221_X1 U23960 ( .B1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput16), 
        .C1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(keyinput36), .A(n21030), .ZN(
        n21035) );
  AOI22_X1 U23961 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(keyinput53), .B1(
        BUF1_REG_27__SCAN_IN), .B2(keyinput39), .ZN(n21031) );
  OAI221_X1 U23962 ( .B1(P2_UWORD_REG_9__SCAN_IN), .B2(keyinput53), .C1(
        BUF1_REG_27__SCAN_IN), .C2(keyinput39), .A(n21031), .ZN(n21034) );
  AOI22_X1 U23963 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput44), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput61), .ZN(n21032) );
  OAI221_X1 U23964 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput44), .C1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(keyinput61), .A(n21032), .ZN(
        n21033) );
  NOR4_X1 U23965 ( .A1(n21036), .A2(n21035), .A3(n21034), .A4(n21033), .ZN(
        n21070) );
  AOI22_X1 U23966 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(keyinput8), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput62), .ZN(n21037) );
  OAI221_X1 U23967 ( .B1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B2(keyinput8), 
        .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(keyinput62), .A(n21037), 
        .ZN(n21044) );
  AOI22_X1 U23968 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput10), 
        .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput24), .ZN(n21038)
         );
  OAI221_X1 U23969 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput10), 
        .C1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(keyinput24), .A(n21038), 
        .ZN(n21043) );
  AOI22_X1 U23970 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(keyinput56), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(keyinput43), .ZN(n21039) );
  OAI221_X1 U23971 ( .B1(P1_DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput56), .C1(
        P2_REIP_REG_30__SCAN_IN), .C2(keyinput43), .A(n21039), .ZN(n21042) );
  AOI22_X1 U23972 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(keyinput48), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(keyinput15), .ZN(n21040) );
  OAI221_X1 U23973 ( .B1(P2_ADDRESS_REG_10__SCAN_IN), .B2(keyinput48), .C1(
        P2_EAX_REG_6__SCAN_IN), .C2(keyinput15), .A(n21040), .ZN(n21041) );
  NOR4_X1 U23974 ( .A1(n21044), .A2(n21043), .A3(n21042), .A4(n21041), .ZN(
        n21069) );
  AOI22_X1 U23975 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(keyinput63), .B1(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput37), .ZN(n21045) );
  OAI221_X1 U23976 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(keyinput63), .C1(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(keyinput37), .A(n21045), .ZN(
        n21052) );
  AOI22_X1 U23977 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(keyinput50), .B1(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput2), .ZN(n21046) );
  OAI221_X1 U23978 ( .B1(P1_EBX_REG_0__SCAN_IN), .B2(keyinput50), .C1(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .C2(keyinput2), .A(n21046), .ZN(
        n21051) );
  AOI22_X1 U23979 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(keyinput46), .B1(
        P2_ADDRESS_REG_25__SCAN_IN), .B2(keyinput60), .ZN(n21047) );
  OAI221_X1 U23980 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(keyinput46), .C1(
        P2_ADDRESS_REG_25__SCAN_IN), .C2(keyinput60), .A(n21047), .ZN(n21050)
         );
  AOI22_X1 U23981 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(keyinput25), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(keyinput32), .ZN(n21048) );
  OAI221_X1 U23982 ( .B1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B2(keyinput25), 
        .C1(P2_EBX_REG_4__SCAN_IN), .C2(keyinput32), .A(n21048), .ZN(n21049)
         );
  NOR4_X1 U23983 ( .A1(n21052), .A2(n21051), .A3(n21050), .A4(n21049), .ZN(
        n21068) );
  AOI22_X1 U23984 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(keyinput31), .B1(
        P2_INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput4), .ZN(n21053) );
  OAI221_X1 U23985 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(keyinput31), .C1(
        P2_INSTQUEUE_REG_5__0__SCAN_IN), .C2(keyinput4), .A(n21053), .ZN(
        n21066) );
  AOI22_X1 U23986 ( .A1(n21056), .A2(keyinput29), .B1(keyinput19), .B2(n21055), 
        .ZN(n21054) );
  OAI221_X1 U23987 ( .B1(n21056), .B2(keyinput29), .C1(n21055), .C2(keyinput19), .A(n21054), .ZN(n21065) );
  AOI22_X1 U23988 ( .A1(n21059), .A2(keyinput9), .B1(n21058), .B2(keyinput59), 
        .ZN(n21057) );
  OAI221_X1 U23989 ( .B1(n21059), .B2(keyinput9), .C1(n21058), .C2(keyinput59), 
        .A(n21057), .ZN(n21064) );
  INV_X1 U23990 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n21062) );
  AOI22_X1 U23991 ( .A1(n21062), .A2(keyinput49), .B1(keyinput55), .B2(n21061), 
        .ZN(n21060) );
  OAI221_X1 U23992 ( .B1(n21062), .B2(keyinput49), .C1(n21061), .C2(keyinput55), .A(n21060), .ZN(n21063) );
  NOR4_X1 U23993 ( .A1(n21066), .A2(n21065), .A3(n21064), .A4(n21063), .ZN(
        n21067) );
  NAND4_X1 U23994 ( .A1(n21070), .A2(n21069), .A3(n21068), .A4(n21067), .ZN(
        n21136) );
  INV_X1 U23995 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21073) );
  AOI22_X1 U23996 ( .A1(n21073), .A2(keyinput22), .B1(keyinput40), .B2(n21072), 
        .ZN(n21071) );
  OAI221_X1 U23997 ( .B1(n21073), .B2(keyinput22), .C1(n21072), .C2(keyinput40), .A(n21071), .ZN(n21084) );
  AOI22_X1 U23998 ( .A1(n12752), .A2(keyinput45), .B1(keyinput28), .B2(n21075), 
        .ZN(n21074) );
  OAI221_X1 U23999 ( .B1(n12752), .B2(keyinput45), .C1(n21075), .C2(keyinput28), .A(n21074), .ZN(n21083) );
  AOI22_X1 U24000 ( .A1(n21077), .A2(keyinput11), .B1(n9979), .B2(keyinput17), 
        .ZN(n21076) );
  OAI221_X1 U24001 ( .B1(n21077), .B2(keyinput11), .C1(n9979), .C2(keyinput17), 
        .A(n21076), .ZN(n21082) );
  XOR2_X1 U24002 ( .A(n21078), .B(keyinput38), .Z(n21080) );
  XNOR2_X1 U24003 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B(keyinput34), .ZN(
        n21079) );
  NAND2_X1 U24004 ( .A1(n21080), .A2(n21079), .ZN(n21081) );
  NOR4_X1 U24005 ( .A1(n21084), .A2(n21083), .A3(n21082), .A4(n21081), .ZN(
        n21134) );
  AOI22_X1 U24006 ( .A1(n21087), .A2(keyinput14), .B1(keyinput54), .B2(n21086), 
        .ZN(n21085) );
  OAI221_X1 U24007 ( .B1(n21087), .B2(keyinput14), .C1(n21086), .C2(keyinput54), .A(n21085), .ZN(n21100) );
  AOI22_X1 U24008 ( .A1(n21090), .A2(keyinput23), .B1(n21089), .B2(keyinput5), 
        .ZN(n21088) );
  OAI221_X1 U24009 ( .B1(n21090), .B2(keyinput23), .C1(n21089), .C2(keyinput5), 
        .A(n21088), .ZN(n21099) );
  AOI22_X1 U24010 ( .A1(n21093), .A2(keyinput27), .B1(keyinput12), .B2(n21092), 
        .ZN(n21091) );
  OAI221_X1 U24011 ( .B1(n21093), .B2(keyinput27), .C1(n21092), .C2(keyinput12), .A(n21091), .ZN(n21098) );
  AOI22_X1 U24012 ( .A1(n21096), .A2(keyinput33), .B1(keyinput21), .B2(n21095), 
        .ZN(n21094) );
  OAI221_X1 U24013 ( .B1(n21096), .B2(keyinput33), .C1(n21095), .C2(keyinput21), .A(n21094), .ZN(n21097) );
  NOR4_X1 U24014 ( .A1(n21100), .A2(n21099), .A3(n21098), .A4(n21097), .ZN(
        n21133) );
  AOI22_X1 U24015 ( .A1(n21103), .A2(keyinput52), .B1(n21102), .B2(keyinput47), 
        .ZN(n21101) );
  OAI221_X1 U24016 ( .B1(n21103), .B2(keyinput52), .C1(n21102), .C2(keyinput47), .A(n21101), .ZN(n21115) );
  AOI22_X1 U24017 ( .A1(n21105), .A2(keyinput57), .B1(n9967), .B2(keyinput51), 
        .ZN(n21104) );
  OAI221_X1 U24018 ( .B1(n21105), .B2(keyinput57), .C1(n9967), .C2(keyinput51), 
        .A(n21104), .ZN(n21114) );
  AOI22_X1 U24019 ( .A1(n21108), .A2(keyinput41), .B1(keyinput13), .B2(n21107), 
        .ZN(n21106) );
  OAI221_X1 U24020 ( .B1(n21108), .B2(keyinput41), .C1(n21107), .C2(keyinput13), .A(n21106), .ZN(n21113) );
  AOI22_X1 U24021 ( .A1(n21111), .A2(keyinput6), .B1(n21110), .B2(keyinput58), 
        .ZN(n21109) );
  OAI221_X1 U24022 ( .B1(n21111), .B2(keyinput6), .C1(n21110), .C2(keyinput58), 
        .A(n21109), .ZN(n21112) );
  NOR4_X1 U24023 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21132) );
  AOI22_X1 U24024 ( .A1(n21118), .A2(keyinput26), .B1(n21117), .B2(keyinput18), 
        .ZN(n21116) );
  OAI221_X1 U24025 ( .B1(n21118), .B2(keyinput26), .C1(n21117), .C2(keyinput18), .A(n21116), .ZN(n21130) );
  INV_X1 U24026 ( .A(READY2), .ZN(n21121) );
  AOI22_X1 U24027 ( .A1(n21121), .A2(keyinput42), .B1(n21120), .B2(keyinput7), 
        .ZN(n21119) );
  OAI221_X1 U24028 ( .B1(n21121), .B2(keyinput42), .C1(n21120), .C2(keyinput7), 
        .A(n21119), .ZN(n21129) );
  AOI22_X1 U24029 ( .A1(n10373), .A2(keyinput30), .B1(keyinput0), .B2(n21123), 
        .ZN(n21122) );
  OAI221_X1 U24030 ( .B1(n10373), .B2(keyinput30), .C1(n21123), .C2(keyinput0), 
        .A(n21122), .ZN(n21128) );
  AOI22_X1 U24031 ( .A1(n21126), .A2(keyinput35), .B1(keyinput20), .B2(n21125), 
        .ZN(n21124) );
  OAI221_X1 U24032 ( .B1(n21126), .B2(keyinput35), .C1(n21125), .C2(keyinput20), .A(n21124), .ZN(n21127) );
  NOR4_X1 U24033 ( .A1(n21130), .A2(n21129), .A3(n21128), .A4(n21127), .ZN(
        n21131) );
  NAND4_X1 U24034 ( .A1(n21134), .A2(n21133), .A3(n21132), .A4(n21131), .ZN(
        n21135) );
  AOI211_X1 U24035 ( .C1(n21138), .C2(n21137), .A(n21136), .B(n21135), .ZN(
        n21151) );
  AOI22_X1 U24036 ( .A1(n21142), .A2(n21141), .B1(n21140), .B2(n21139), .ZN(
        n21147) );
  AOI22_X1 U24037 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21145), .B1(
        n21144), .B2(n21143), .ZN(n21146) );
  OAI211_X1 U24038 ( .C1(n21149), .C2(n21148), .A(n21147), .B(n21146), .ZN(
        n21150) );
  XOR2_X1 U24039 ( .A(n21151), .B(n21150), .Z(P1_U3045) );
  INV_X1 U12369 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10138) );
  OR2_X1 U13240 ( .A1(n10314), .A2(n10309), .ZN(n15566) );
  NAND2_X1 U11405 ( .A1(n11539), .A2(n11609), .ZN(n13980) );
  INV_X1 U11073 ( .A(n19291), .ZN(n19328) );
  CLKBUF_X1 U11104 ( .A(n12234), .Z(n11980) );
  CLKBUF_X1 U11116 ( .A(n17233), .Z(n9629) );
  XNOR2_X1 U11122 ( .A(n9759), .B(n11446), .ZN(n20378) );
  NAND2_X1 U11148 ( .A1(n11452), .A2(n11451), .ZN(n13970) );
  NAND2_X1 U11152 ( .A1(n14994), .A2(n12990), .ZN(n13012) );
  CLKBUF_X1 U11153 ( .A(n10442), .Z(n19538) );
  NAND2_X1 U11157 ( .A1(n9717), .A2(n10090), .ZN(n13892) );
  CLKBUF_X1 U11167 ( .A(n12939), .Z(n15017) );
  CLKBUF_X1 U11389 ( .A(n10294), .Z(n10295) );
  CLKBUF_X1 U11418 ( .A(n16557), .Z(n16563) );
  OR2_X1 U12199 ( .A1(n18281), .A2(n18295), .ZN(n21152) );
  CLKBUF_X1 U12268 ( .A(n18905), .Z(n17507) );
endmodule

