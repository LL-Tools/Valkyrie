

module b17_C_gen_AntiSAT_k_128_3 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164;

  NAND3_X1 U11079 ( .A1(n10184), .A2(n13884), .A3(n11921), .ZN(n13996) );
  AND2_X1 U11080 ( .A1(n12316), .A2(n12315), .ZN(n14596) );
  XNOR2_X1 U11081 ( .A(n12880), .B(n13425), .ZN(n13947) );
  INV_X1 U11082 ( .A(n19074), .ZN(n16733) );
  INV_X2 U11083 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11760) );
  OR2_X1 U11084 ( .A1(n10434), .A2(n10431), .ZN(n19789) );
  CLKBUF_X2 U11085 ( .A(n10416), .Z(n9639) );
  AND2_X2 U11086 ( .A1(n14499), .A2(n10275), .ZN(n11033) );
  OAI21_X1 U11087 ( .B1(n19321), .B2(n13307), .A(n13268), .ZN(n13314) );
  AND2_X1 U11088 ( .A1(n14503), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10644) );
  AND2_X1 U11089 ( .A1(n14503), .A2(n10275), .ZN(n14351) );
  AND2_X1 U11090 ( .A1(n9682), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10639) );
  AND2_X1 U11091 ( .A1(n14504), .A2(n10275), .ZN(n10659) );
  AND2_X1 U11092 ( .A1(n10451), .A2(n10275), .ZN(n14352) );
  CLKBUF_X2 U11093 ( .A(n12581), .Z(n17355) );
  CLKBUF_X2 U11094 ( .A(n17369), .Z(n17350) );
  CLKBUF_X2 U11095 ( .A(n11560), .Z(n12511) );
  INV_X1 U11096 ( .A(n17197), .ZN(n17388) );
  CLKBUF_X2 U11097 ( .A(n12698), .Z(n9652) );
  CLKBUF_X1 U11098 ( .A(n12719), .Z(n9650) );
  CLKBUF_X2 U11099 ( .A(n12602), .Z(n17369) );
  BUF_X1 U11100 ( .A(n12563), .Z(n17214) );
  INV_X1 U11101 ( .A(n17197), .ZN(n17367) );
  CLKBUF_X2 U11102 ( .A(n9692), .Z(n9685) );
  BUF_X1 U11103 ( .A(n11614), .Z(n15194) );
  NOR2_X1 U11104 ( .A1(n10330), .A2(n10844), .ZN(n10350) );
  INV_X1 U11105 ( .A(n13749), .ZN(n12869) );
  AND2_X1 U11106 ( .A1(n11458), .A2(n11459), .ZN(n9669) );
  OAI22_X2 U11107 ( .A1(n16629), .A2(n13764), .B1(n21140), .B2(n13763), .ZN(
        n20824) );
  NAND2_X2 U11108 ( .A1(n20344), .A2(n14260), .ZN(n13764) );
  INV_X1 U11110 ( .A(n21163), .ZN(n9636) );
  CLKBUF_X2 U11112 ( .A(n11551), .Z(n9690) );
  INV_X1 U11113 ( .A(n12198), .ZN(n11553) );
  AND4_X1 U11114 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11514) );
  AND2_X1 U11115 ( .A1(n14500), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10654) );
  AND2_X1 U11116 ( .A1(n13803), .A2(n10417), .ZN(n10410) );
  INV_X1 U11117 ( .A(n12585), .ZN(n12541) );
  INV_X1 U11118 ( .A(n13817), .ZN(n10184) );
  XNOR2_X1 U11119 ( .A(n11781), .B(n11782), .ZN(n13755) );
  NAND2_X1 U11120 ( .A1(n10725), .A2(n14554), .ZN(n10724) );
  AND3_X1 U11121 ( .A1(n10942), .A2(n20152), .A3(n13434), .ZN(n10329) );
  NOR2_X1 U11122 ( .A1(n9639), .A2(n10415), .ZN(n19566) );
  NAND2_X1 U11123 ( .A1(n18363), .A2(n18872), .ZN(n18248) );
  NAND3_X1 U11124 ( .A1(n16171), .A2(n12370), .A3(n10151), .ZN(n9911) );
  INV_X1 U11125 ( .A(n13900), .ZN(n11635) );
  INV_X1 U11126 ( .A(n14552), .ZN(n11295) );
  OR2_X1 U11127 ( .A1(n11308), .A2(n11307), .ZN(n16350) );
  OR2_X1 U11128 ( .A1(n15410), .A2(n15409), .ZN(n15412) );
  OAI21_X1 U11129 ( .B1(n16350), .B2(n10536), .A(n15732), .ZN(n15587) );
  AOI21_X1 U11130 ( .B1(n10067), .B2(n9846), .A(n9845), .ZN(n15573) );
  INV_X1 U11131 ( .A(n17083), .ZN(n9975) );
  INV_X1 U11132 ( .A(n18436), .ZN(n17447) );
  AOI21_X1 U11133 ( .B1(n16022), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9864), .ZN(n12675) );
  NOR2_X2 U11134 ( .A1(n13908), .A2(n13907), .ZN(n20229) );
  OR2_X1 U11135 ( .A1(n11298), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11305) );
  AND2_X1 U11136 ( .A1(n13437), .A2(n9823), .ZN(n13433) );
  NAND2_X1 U11137 ( .A1(n10405), .A2(n10407), .ZN(n10412) );
  AND2_X1 U11138 ( .A1(n10861), .A2(n16538), .ZN(n11201) );
  INV_X1 U11139 ( .A(n18416), .ZN(n17600) );
  INV_X1 U11140 ( .A(n17911), .ZN(n17927) );
  INV_X1 U11141 ( .A(n18062), .ZN(n18071) );
  AOI22_X1 U11142 ( .A1(n12677), .A2(n12676), .B1(n16021), .B2(n12675), .ZN(
        n16582) );
  INV_X1 U11143 ( .A(n20229), .ZN(n20244) );
  INV_X2 U11144 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19097) );
  AOI211_X1 U11145 ( .C1(n15823), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15822), .B(n15821), .ZN(n15824) );
  AND2_X1 U11146 ( .A1(n11602), .A2(n10219), .ZN(n9637) );
  AND4_X1 U11147 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n9638) );
  AND2_X1 U11148 ( .A1(n13669), .A2(n11359), .ZN(n11713) );
  NAND3_X2 U11149 ( .A1(n9911), .A2(n9909), .A3(n9717), .ZN(n10149) );
  AND4_X4 U11150 ( .A1(n11515), .A2(n9721), .A3(n11514), .A4(n11513), .ZN(
        n13013) );
  AOI21_X2 U11151 ( .B1(n13947), .B2(n13895), .A(n12881), .ZN(n13793) );
  XNOR2_X1 U11152 ( .A(n10408), .B(n10409), .ZN(n10416) );
  INV_X2 U11153 ( .A(n10258), .ZN(n9640) );
  INV_X1 U11154 ( .A(n10258), .ZN(n9641) );
  INV_X1 U11155 ( .A(n9640), .ZN(n9642) );
  INV_X1 U11156 ( .A(n9640), .ZN(n9643) );
  INV_X1 U11157 ( .A(n9640), .ZN(n9644) );
  INV_X1 U11158 ( .A(n9640), .ZN(n9645) );
  INV_X1 U11159 ( .A(n9641), .ZN(n9646) );
  INV_X1 U11160 ( .A(n9641), .ZN(n9647) );
  AND2_X2 U11161 ( .A1(n9802), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10258) );
  NOR3_X1 U11162 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n12540), .ZN(n9648) );
  NAND2_X2 U11163 ( .A1(n10316), .A2(n10315), .ZN(n10325) );
  NOR2_X2 U11164 ( .A1(n19176), .A2(n19177), .ZN(n19175) );
  NOR2_X1 U11165 ( .A1(n12539), .A2(n18884), .ZN(n9649) );
  NOR2_X2 U11166 ( .A1(n12815), .A2(n18385), .ZN(n18075) );
  NOR2_X2 U11167 ( .A1(n12494), .A2(n10146), .ZN(n14529) );
  NOR2_X1 U11168 ( .A1(n12539), .A2(n18888), .ZN(n12719) );
  AND2_X2 U11170 ( .A1(n10441), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10507) );
  BUF_X1 U11171 ( .A(n12698), .Z(n9651) );
  NOR2_X1 U11172 ( .A1(n18884), .A2(n12542), .ZN(n12698) );
  NAND2_X1 U11173 ( .A1(n14707), .A2(n9658), .ZN(n14651) );
  AND2_X1 U11174 ( .A1(n14707), .A2(n10185), .ZN(n14650) );
  NAND2_X1 U11175 ( .A1(n10155), .A2(n14991), .ZN(n10154) );
  AND2_X1 U11176 ( .A1(n12404), .A2(n10159), .ZN(n10158) );
  AND2_X1 U11177 ( .A1(n10032), .A2(n10031), .ZN(n16324) );
  AND2_X1 U11178 ( .A1(n9869), .A2(n9868), .ZN(n17754) );
  OR2_X1 U11179 ( .A1(n16339), .A2(n19288), .ZN(n10032) );
  NOR2_X1 U11180 ( .A1(n16340), .A2(n16341), .ZN(n16339) );
  INV_X4 U11181 ( .A(n14933), .ZN(n16146) );
  INV_X1 U11182 ( .A(n10579), .ZN(n10515) );
  OAI21_X1 U11183 ( .B1(n13916), .B2(n12338), .A(n12329), .ZN(n12352) );
  NOR2_X1 U11184 ( .A1(n15579), .A2(n15304), .ZN(n15303) );
  NAND2_X1 U11185 ( .A1(n13398), .A2(n13397), .ZN(n13432) );
  INV_X1 U11186 ( .A(n13803), .ZN(n13399) );
  NAND2_X1 U11189 ( .A1(n20270), .A2(n14843), .ZN(n20265) );
  NAND3_X1 U11190 ( .A1(n17992), .A2(n17978), .A3(n9722), .ZN(n17964) );
  OR2_X1 U11191 ( .A1(n16080), .A2(n12921), .ZN(n16081) );
  INV_X2 U11192 ( .A(n18249), .ZN(n18852) );
  NAND2_X1 U11193 ( .A1(n19074), .A2(n18345), .ZN(n18249) );
  INV_X2 U11194 ( .A(n18894), .ZN(n18864) );
  NOR2_X1 U11195 ( .A1(n11652), .A2(n11651), .ZN(n11686) );
  INV_X2 U11196 ( .A(n18897), .ZN(n18872) );
  AOI22_X1 U11197 ( .A1(n10927), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16539), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10362) );
  INV_X4 U11198 ( .A(n17955), .ZN(n17978) );
  NAND2_X1 U11199 ( .A1(n12886), .A2(n12874), .ZN(n12927) );
  NAND2_X1 U11200 ( .A1(n11618), .A2(n11617), .ZN(n11634) );
  MUX2_X1 U11201 ( .A(n11616), .B(n13018), .S(n13749), .Z(n11617) );
  NAND2_X1 U11202 ( .A1(n17447), .A2(n17444), .ZN(n12790) );
  INV_X2 U11203 ( .A(n13013), .ZN(n11682) );
  NAND2_X1 U11204 ( .A1(n10269), .A2(n10270), .ZN(n10328) );
  INV_X2 U11205 ( .A(n10939), .ZN(n19474) );
  NAND2_X1 U11206 ( .A1(n12571), .A2(n12572), .ZN(n9867) );
  INV_X1 U11207 ( .A(n10537), .ZN(n9653) );
  AND4_X1 U11208 ( .A1(n11453), .A2(n11452), .A3(n11451), .A4(n11450), .ZN(
        n11459) );
  NAND4_X1 U11209 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11615) );
  BUF_X2 U11210 ( .A(n11553), .Z(n12124) );
  AND4_X1 U11211 ( .A1(n10296), .A2(n10295), .A3(n10294), .A4(n10293), .ZN(
        n10303) );
  BUF_X2 U11212 ( .A(n12584), .Z(n17393) );
  BUF_X4 U11213 ( .A(n12697), .Z(n17395) );
  CLKBUF_X2 U11214 ( .A(n11703), .Z(n11690) );
  BUF_X2 U11215 ( .A(n11529), .Z(n11491) );
  BUF_X2 U11216 ( .A(n11558), .Z(n11575) );
  CLKBUF_X2 U11217 ( .A(n11713), .Z(n9687) );
  CLKBUF_X2 U11218 ( .A(n10442), .Z(n14499) );
  AND2_X4 U11219 ( .A1(n10220), .A2(n14333), .ZN(n14500) );
  INV_X4 U11220 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11350) );
  NAND2_X1 U11221 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12540) );
  AND2_X1 U11222 ( .A1(n9894), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9891) );
  OAI21_X1 U11223 ( .B1(n15556), .B2(n16524), .A(n12865), .ZN(n9998) );
  AND2_X1 U11224 ( .A1(n12494), .A2(n10022), .ZN(n14527) );
  AOI21_X1 U11225 ( .B1(n14592), .B2(n16519), .A(n9837), .ZN(n9836) );
  AOI21_X1 U11226 ( .B1(n14911), .B2(n20344), .A(n14910), .ZN(n14912) );
  AND2_X1 U11227 ( .A1(n10193), .A2(n10191), .ZN(n14251) );
  AND2_X1 U11228 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  AOI211_X1 U11229 ( .C1(n14655), .C2(P1_REIP_REG_26__SCAN_IN), .A(n14654), 
        .B(n14653), .ZN(n14656) );
  NOR2_X2 U11230 ( .A1(n15584), .A2(n15732), .ZN(n15578) );
  XNOR2_X1 U11231 ( .A(n15549), .B(n15548), .ZN(n15701) );
  INV_X1 U11232 ( .A(n10191), .ZN(n12527) );
  INV_X1 U11233 ( .A(n15391), .ZN(n9809) );
  NAND2_X1 U11234 ( .A1(n12489), .A2(n14924), .ZN(n13016) );
  NAND2_X1 U11235 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15713) );
  INV_X1 U11236 ( .A(n14651), .ZN(n14629) );
  OAI21_X1 U11237 ( .B1(n15835), .B2(n10060), .A(n10058), .ZN(n15668) );
  NAND2_X1 U11238 ( .A1(n9918), .A2(n16391), .ZN(n15835) );
  CLKBUF_X1 U11239 ( .A(n15573), .Z(n15597) );
  CLKBUF_X1 U11240 ( .A(n14732), .Z(n14733) );
  AND2_X1 U11241 ( .A1(n10207), .A2(n9817), .ZN(n9814) );
  NAND2_X1 U11242 ( .A1(n10153), .A2(n10158), .ZN(n14992) );
  NAND2_X1 U11243 ( .A1(n9902), .A2(n10154), .ZN(n9901) );
  NAND2_X1 U11244 ( .A1(n10067), .A2(n10064), .ZN(n9918) );
  NAND2_X1 U11245 ( .A1(n14750), .A2(n9780), .ZN(n14732) );
  INV_X1 U11246 ( .A(n14749), .ZN(n14750) );
  OR2_X1 U11247 ( .A1(n14414), .A2(n14413), .ZN(n10207) );
  AND2_X1 U11248 ( .A1(n10012), .A2(n10203), .ZN(n9959) );
  AND2_X1 U11249 ( .A1(n11186), .A2(n11192), .ZN(n10166) );
  XNOR2_X1 U11250 ( .A(n14566), .B(n14565), .ZN(n15382) );
  NAND2_X1 U11251 ( .A1(n10140), .A2(n10137), .ZN(n10136) );
  AND2_X1 U11252 ( .A1(n11193), .A2(n10161), .ZN(n10160) );
  NAND2_X1 U11253 ( .A1(n9865), .A2(n17955), .ZN(n16592) );
  AND2_X1 U11254 ( .A1(n14159), .A2(n10137), .ZN(n9917) );
  AND2_X1 U11255 ( .A1(n10158), .A2(n9783), .ZN(n9900) );
  XNOR2_X1 U11256 ( .A(n10695), .B(n14218), .ZN(n14159) );
  NAND2_X1 U11257 ( .A1(n9915), .A2(n10625), .ZN(n14158) );
  NAND2_X1 U11258 ( .A1(n9992), .A2(n9991), .ZN(n17725) );
  AND2_X1 U11259 ( .A1(n9910), .A2(n16158), .ZN(n9909) );
  NAND2_X1 U11260 ( .A1(n9989), .A2(n9996), .ZN(n9994) );
  AND2_X1 U11261 ( .A1(n16134), .A2(n16138), .ZN(n12401) );
  NOR2_X1 U11262 ( .A1(n16157), .A2(n10152), .ZN(n10151) );
  AOI21_X1 U11263 ( .B1(n19332), .B2(n19305), .A(n10081), .ZN(n15274) );
  NAND2_X1 U11264 ( .A1(n11174), .A2(n16506), .ZN(n16445) );
  NAND2_X1 U11265 ( .A1(n11169), .A2(n11168), .ZN(n13874) );
  AND2_X1 U11266 ( .A1(n15008), .A2(n12399), .ZN(n16134) );
  OAI21_X1 U11267 ( .B1(n15035), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15008), .ZN(n15019) );
  AND2_X1 U11268 ( .A1(n11175), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11183) );
  NAND2_X1 U11269 ( .A1(n9841), .A2(n10627), .ZN(n10689) );
  NAND2_X1 U11270 ( .A1(n11902), .A2(n11901), .ZN(n13884) );
  NOR2_X1 U11271 ( .A1(n17772), .A2(n18139), .ZN(n9868) );
  NAND2_X1 U11272 ( .A1(n14933), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15008) );
  NOR2_X1 U11273 ( .A1(n14933), .A2(n9779), .ZN(n15017) );
  AND2_X2 U11274 ( .A1(n13697), .A2(n11841), .ZN(n9672) );
  NAND2_X1 U11275 ( .A1(n11889), .A2(n11888), .ZN(n13818) );
  NOR2_X1 U11276 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17766), .ZN(
        n17765) );
  XNOR2_X1 U11277 ( .A(n12324), .B(n11893), .ZN(n12384) );
  AND2_X1 U11278 ( .A1(n15803), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15792) );
  AND2_X1 U11279 ( .A1(n10616), .A2(n10615), .ZN(n10627) );
  NAND2_X1 U11280 ( .A1(n11890), .A2(n11891), .ZN(n12371) );
  OR3_X1 U11281 ( .A1(n10686), .A2(n10685), .A3(n10684), .ZN(n10687) );
  AND2_X1 U11282 ( .A1(n13836), .A2(n9757), .ZN(n14190) );
  OAI21_X1 U11283 ( .B1(n13916), .B2(n11997), .A(n11840), .ZN(n13773) );
  OR2_X1 U11284 ( .A1(n16182), .A2(n13040), .ZN(n15055) );
  NAND2_X1 U11285 ( .A1(n11833), .A2(n11842), .ZN(n13916) );
  XNOR2_X1 U11286 ( .A(n11842), .B(n11843), .ZN(n12354) );
  NAND2_X1 U11287 ( .A1(n11761), .A2(n12097), .ZN(n11781) );
  OR2_X1 U11288 ( .A1(n14634), .A2(n14254), .ZN(n14256) );
  NAND2_X1 U11289 ( .A1(n11809), .A2(n13691), .ZN(n11842) );
  CLKBUF_X1 U11290 ( .A(n12330), .Z(n13690) );
  XNOR2_X1 U11291 ( .A(n13433), .B(n13432), .ZN(n20103) );
  AND2_X1 U11292 ( .A1(n11759), .A2(n11832), .ZN(n12330) );
  AND2_X1 U11293 ( .A1(n10411), .A2(n9928), .ZN(n19855) );
  AND2_X1 U11294 ( .A1(n9738), .A2(n13435), .ZN(n9799) );
  NAND2_X1 U11295 ( .A1(n9839), .A2(n9838), .ZN(n10581) );
  AND2_X1 U11296 ( .A1(n9857), .A2(n19439), .ZN(n10596) );
  AND2_X1 U11297 ( .A1(n10410), .A2(n9639), .ZN(n19885) );
  NAND2_X1 U11298 ( .A1(n9898), .A2(n11808), .ZN(n13691) );
  NOR2_X1 U11299 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17922), .ZN(
        n17876) );
  OR2_X1 U11300 ( .A1(n10432), .A2(n10433), .ZN(n19454) );
  AND2_X1 U11301 ( .A1(n10030), .A2(n19257), .ZN(n15319) );
  NOR2_X1 U11302 ( .A1(n15856), .A2(n10065), .ZN(n10064) );
  CLKBUF_X1 U11303 ( .A(n12477), .Z(n16118) );
  AND2_X1 U11304 ( .A1(n9803), .A2(n10120), .ZN(n13438) );
  CLKBUF_X1 U11305 ( .A(n12479), .Z(n16117) );
  NOR2_X1 U11306 ( .A1(n13443), .A2(n10002), .ZN(n13561) );
  NOR2_X1 U11307 ( .A1(n15217), .A2(n13811), .ZN(n20828) );
  NOR2_X1 U11308 ( .A1(n15217), .A2(n13734), .ZN(n20834) );
  NOR2_X1 U11309 ( .A1(n15217), .A2(n13744), .ZN(n20816) );
  INV_X1 U11310 ( .A(n16390), .ZN(n10065) );
  NOR2_X1 U11311 ( .A1(n15217), .A2(n13739), .ZN(n20803) );
  NOR2_X1 U11312 ( .A1(n15217), .A2(n13831), .ZN(n20849) );
  NOR2_X1 U11313 ( .A1(n15217), .A2(n13887), .ZN(n20855) );
  NAND2_X1 U11314 ( .A1(n11667), .A2(n11666), .ZN(n11786) );
  NOR2_X1 U11315 ( .A1(n13990), .A2(n19453), .ZN(n19333) );
  NAND2_X1 U11316 ( .A1(n10175), .A2(n9734), .ZN(n11754) );
  AND2_X1 U11317 ( .A1(n15977), .A2(n15976), .ZN(n15988) );
  INV_X1 U11318 ( .A(n13702), .ZN(n11751) );
  NAND2_X2 U11319 ( .A1(n20270), .A2(n11567), .ZN(n14842) );
  OR2_X1 U11320 ( .A1(n9664), .A2(n12652), .ZN(n9663) );
  AOI22_X1 U11321 ( .A1(n18853), .A2(n18852), .B1(n18857), .B2(n15969), .ZN(
        n18861) );
  XNOR2_X1 U11322 ( .A(n11773), .B(n11774), .ZN(n20431) );
  OAI21_X1 U11323 ( .B1(n19136), .B2(n19125), .A(n19257), .ZN(n15977) );
  NAND2_X1 U11324 ( .A1(n11750), .A2(n11658), .ZN(n11667) );
  NOR2_X2 U11325 ( .A1(n14552), .A2(n19498), .ZN(n19485) );
  OR2_X1 U11326 ( .A1(n14781), .A2(n14782), .ZN(n16080) );
  NAND2_X1 U11327 ( .A1(n20477), .A2(n11654), .ZN(n11750) );
  NAND2_X1 U11328 ( .A1(n18007), .A2(n12648), .ZN(n12651) );
  XNOR2_X1 U11329 ( .A(n13304), .B(n13302), .ZN(n10409) );
  OAI211_X1 U11330 ( .C1(n13924), .C2(n12321), .A(n11665), .B(n11664), .ZN(
        n11666) );
  NAND2_X1 U11331 ( .A1(n11775), .A2(n20865), .ZN(n11723) );
  NOR2_X1 U11332 ( .A1(n13448), .A2(n13444), .ZN(n10003) );
  OR2_X1 U11333 ( .A1(n11787), .A2(n11350), .ZN(n11791) );
  OR2_X1 U11334 ( .A1(n11787), .A2(n9887), .ZN(n11665) );
  CLKBUF_X1 U11335 ( .A(n11662), .Z(n11787) );
  NAND2_X1 U11336 ( .A1(n10391), .A2(n10390), .ZN(n10393) );
  XNOR2_X1 U11337 ( .A(n10381), .B(n10380), .ZN(n10404) );
  NAND2_X1 U11338 ( .A1(n10363), .A2(n10362), .ZN(n10380) );
  INV_X1 U11339 ( .A(n9670), .ZN(n11656) );
  NAND2_X1 U11340 ( .A1(n10386), .A2(n10385), .ZN(n13302) );
  OAI21_X1 U11341 ( .B1(n10384), .B2(n9720), .A(n10379), .ZN(n10407) );
  NAND2_X1 U11342 ( .A1(n10398), .A2(n10397), .ZN(n10868) );
  AND2_X1 U11343 ( .A1(n10389), .A2(n10388), .ZN(n10390) );
  OR2_X1 U11344 ( .A1(n10384), .A2(n14333), .ZN(n10386) );
  AOI21_X1 U11345 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(n10379) );
  AND2_X1 U11346 ( .A1(n10372), .A2(n10371), .ZN(n10374) );
  NOR2_X1 U11347 ( .A1(n10618), .A2(n10617), .ZN(n10621) );
  OR2_X2 U11348 ( .A1(n17638), .A2(n18917), .ZN(n17706) );
  OR2_X1 U11349 ( .A1(n14517), .A2(n19115), .ZN(n10373) );
  OAI21_X1 U11350 ( .B1(n12460), .B2(n12993), .A(n13012), .ZN(n11626) );
  NAND2_X1 U11351 ( .A1(n9889), .A2(n13895), .ZN(n11620) );
  AND2_X1 U11352 ( .A1(n9946), .A2(n13080), .ZN(n10359) );
  INV_X1 U11353 ( .A(n14517), .ZN(n14562) );
  CLKBUF_X1 U11354 ( .A(n12460), .Z(n9686) );
  NOR2_X1 U11355 ( .A1(n16405), .A2(n13073), .ZN(n19227) );
  AND4_X1 U11356 ( .A1(n11650), .A2(n11645), .A3(n13017), .A4(n20955), .ZN(
        n11633) );
  AND2_X1 U11357 ( .A1(n10338), .A2(n10337), .ZN(n11151) );
  NOR2_X1 U11358 ( .A1(n11632), .A2(n13356), .ZN(n11649) );
  NAND2_X1 U11359 ( .A1(n18055), .A2(n12636), .ZN(n18042) );
  OR2_X1 U11360 ( .A1(n10945), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10167) );
  NAND2_X1 U11361 ( .A1(n13029), .A2(n11631), .ZN(n13356) );
  NAND2_X1 U11362 ( .A1(n13269), .A2(n10537), .ZN(n13291) );
  CLKBUF_X1 U11363 ( .A(n11627), .Z(n11628) );
  NAND2_X1 U11364 ( .A1(n11793), .A2(n11792), .ZN(n12280) );
  NAND3_X1 U11365 ( .A1(n12775), .A2(n12774), .A3(n12773), .ZN(n17444) );
  INV_X2 U11366 ( .A(U212), .ZN(n16660) );
  OR2_X2 U11367 ( .A1(n16661), .A2(n16605), .ZN(n16663) );
  BUF_X2 U11368 ( .A(n9653), .Z(n14552) );
  XNOR2_X1 U11369 ( .A(n17593), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18067) );
  CLKBUF_X1 U11370 ( .A(n10325), .Z(n11330) );
  INV_X1 U11371 ( .A(n10328), .ZN(n13269) );
  CLKBUF_X1 U11372 ( .A(n10328), .Z(n13434) );
  INV_X1 U11373 ( .A(n13326), .ZN(n9654) );
  NAND3_X1 U11374 ( .A1(n11682), .A2(n13900), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12301) );
  OR2_X1 U11375 ( .A1(n11719), .A2(n11718), .ZN(n12342) );
  OR2_X1 U11376 ( .A1(n11682), .A2(n20865), .ZN(n11793) );
  NAND2_X1 U11377 ( .A1(n9638), .A2(n9723), .ZN(n11630) );
  AND2_X1 U11378 ( .A1(n9669), .A2(n11615), .ZN(n11627) );
  OR2_X1 U11379 ( .A1(n11702), .A2(n11701), .ZN(n12389) );
  NAND2_X2 U11380 ( .A1(n10198), .A2(n11544), .ZN(n13749) );
  CLKBUF_X1 U11381 ( .A(n11615), .Z(n13357) );
  NOR2_X2 U11382 ( .A1(n12704), .A2(n12703), .ZN(n19074) );
  NAND2_X2 U11383 ( .A1(n11458), .A2(n11459), .ZN(n11624) );
  AND3_X1 U11384 ( .A1(n11490), .A2(n11489), .A3(n9661), .ZN(n11496) );
  AND4_X1 U11385 ( .A1(n12570), .A2(n10209), .A3(n12569), .A4(n12568), .ZN(
        n12571) );
  AND4_X1 U11386 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11544) );
  NAND2_X1 U11387 ( .A1(n10244), .A2(n10243), .ZN(n10537) );
  AND3_X1 U11388 ( .A1(n10216), .A2(n11534), .A3(n11533), .ZN(n10198) );
  AND4_X1 U11389 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11592) );
  NOR2_X1 U11390 ( .A1(n11478), .A2(n10218), .ZN(n11479) );
  NAND2_X1 U11391 ( .A1(n20344), .A2(n13718), .ZN(n13763) );
  AND4_X1 U11392 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11591) );
  AND4_X1 U11393 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11590) );
  AND4_X1 U11394 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  AND4_X1 U11395 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11612) );
  AND4_X1 U11396 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11480) );
  AND4_X1 U11397 ( .A1(n11457), .A2(n11456), .A3(n11455), .A4(n11454), .ZN(
        n11458) );
  AND3_X1 U11398 ( .A1(n11494), .A2(n11493), .A3(n11492), .ZN(n10215) );
  BUF_X2 U11399 ( .A(n12575), .Z(n17368) );
  BUF_X2 U11400 ( .A(n12575), .Z(n17385) );
  BUF_X2 U11401 ( .A(n12719), .Z(n17366) );
  NAND2_X2 U11402 ( .A1(n19083), .A2(n18954), .ZN(n19013) );
  INV_X2 U11403 ( .A(n12503), .ZN(n12173) );
  NAND2_X2 U11404 ( .A1(n19083), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19017) );
  AOI22_X1 U11405 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11562), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11451) );
  NAND2_X2 U11406 ( .A1(n20159), .A2(n20046), .ZN(n20089) );
  BUF_X2 U11407 ( .A(n10309), .Z(n10441) );
  OR2_X1 U11408 ( .A1(n12503), .A2(n20395), .ZN(n10200) );
  INV_X2 U11409 ( .A(n16702), .ZN(n16704) );
  INV_X2 U11410 ( .A(n16729), .ZN(n9655) );
  NAND2_X2 U11411 ( .A1(n13660), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12198) );
  INV_X1 U11412 ( .A(n18871), .ZN(n17096) );
  NOR2_X4 U11413 ( .A1(n18888), .A2(n12542), .ZN(n12697) );
  AND2_X2 U11414 ( .A1(n11358), .A2(n13659), .ZN(n11477) );
  AND2_X2 U11415 ( .A1(n13659), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13660) );
  AND2_X2 U11416 ( .A1(n13656), .A2(n11354), .ZN(n9671) );
  AND2_X2 U11417 ( .A1(n11347), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11360) );
  AND2_X1 U11418 ( .A1(n11350), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13669) );
  AND2_X2 U11419 ( .A1(n9887), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11358) );
  AND2_X2 U11420 ( .A1(n11353), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11359) );
  NAND2_X1 U11421 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12679), .ZN(
        n12543) );
  NAND2_X1 U11422 ( .A1(n12678), .A2(n19048), .ZN(n18884) );
  AND2_X1 U11423 ( .A1(n13594), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9802) );
  NAND2_X1 U11424 ( .A1(n9939), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12532) );
  AND2_X2 U11425 ( .A1(n10220), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10442) );
  NOR2_X1 U11426 ( .A1(n12679), .A2(n12540), .ZN(n18871) );
  INV_X1 U11427 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19048) );
  NOR2_X1 U11429 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9939) );
  AND2_X2 U11430 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13489) );
  INV_X2 U11431 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14333) );
  NOR2_X2 U11432 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10220) );
  INV_X1 U11433 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11587) );
  NOR2_X2 U11434 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13656) );
  AND2_X1 U11435 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11354) );
  AND2_X2 U11436 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13659) );
  NAND2_X1 U11437 ( .A1(n18040), .A2(n18354), .ZN(n9656) );
  NOR2_X2 U11438 ( .A1(n15552), .A2(n15279), .ZN(n15278) );
  INV_X2 U11439 ( .A(n14998), .ZN(n10157) );
  OR2_X1 U11440 ( .A1(n12339), .A2(n9654), .ZN(n12346) );
  XNOR2_X1 U11441 ( .A(n9657), .B(n15639), .ZN(n15800) );
  AND2_X1 U11442 ( .A1(n15637), .A2(n15636), .ZN(n9657) );
  NAND2_X2 U11443 ( .A1(n15685), .A2(n11194), .ZN(n15883) );
  NOR2_X4 U11444 ( .A1(n10843), .A2(n20152), .ZN(n10340) );
  NAND2_X2 U11445 ( .A1(n12992), .A2(n12493), .ZN(n12494) );
  AOI21_X1 U11446 ( .B1(n15407), .B2(n10207), .A(n9817), .ZN(n9816) );
  NAND2_X2 U11447 ( .A1(n9800), .A2(n9799), .ZN(n13542) );
  NAND2_X2 U11448 ( .A1(n10364), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10387) );
  AND2_X1 U11449 ( .A1(n10185), .A2(n14652), .ZN(n9658) );
  CLKBUF_X1 U11450 ( .A(n10184), .Z(n9659) );
  CLKBUF_X1 U11451 ( .A(n14750), .Z(n9660) );
  AND2_X1 U11452 ( .A1(n11487), .A2(n11488), .ZN(n9661) );
  NAND2_X1 U11453 ( .A1(n17993), .A2(n9665), .ZN(n9662) );
  AND2_X2 U11454 ( .A1(n9662), .A2(n9663), .ZN(n18276) );
  INV_X1 U11455 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9664) );
  AND2_X1 U11456 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U11457 ( .A1(n9667), .A2(n12645), .ZN(n9666) );
  NAND2_X1 U11458 ( .A1(n18024), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9667) );
  CLKBUF_X1 U11459 ( .A(n18040), .Z(n9668) );
  XNOR2_X2 U11460 ( .A(n9862), .B(n12643), .ZN(n18024) );
  NAND2_X2 U11461 ( .A1(n18030), .A2(n12641), .ZN(n9862) );
  NOR2_X1 U11462 ( .A1(n16592), .A2(n16578), .ZN(n12672) );
  NAND2_X2 U11463 ( .A1(n9728), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9670) );
  INV_X1 U11464 ( .A(n9671), .ZN(n11569) );
  NAND2_X2 U11465 ( .A1(n14161), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14160) );
  NAND2_X4 U11466 ( .A1(n10000), .A2(n10122), .ZN(n13803) );
  AOI21_X2 U11467 ( .B1(n10399), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10348), .ZN(n10381) );
  AND2_X2 U11468 ( .A1(n10579), .A2(n10580), .ZN(n11157) );
  INV_X1 U11469 ( .A(n9672), .ZN(n13696) );
  AND2_X1 U11470 ( .A1(n10041), .A2(n13659), .ZN(n11550) );
  NOR2_X2 U11471 ( .A1(n12714), .A2(n12713), .ZN(n18416) );
  OR2_X2 U11472 ( .A1(n15838), .A2(n11195), .ZN(n9999) );
  XNOR2_X2 U11473 ( .A(n10580), .B(n10515), .ZN(n13798) );
  NAND2_X2 U11474 ( .A1(n9947), .A2(n10459), .ZN(n10580) );
  AND2_X1 U11475 ( .A1(n13669), .A2(n11359), .ZN(n9673) );
  INV_X1 U11476 ( .A(n9687), .ZN(n9674) );
  AND2_X1 U11477 ( .A1(n11360), .A2(n11354), .ZN(n9675) );
  AOI21_X1 U11478 ( .B1(n11614), .B2(n11630), .A(n11613), .ZN(n11618) );
  AOI22_X2 U11479 ( .A1(n9725), .A2(n19438), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16456), .ZN(n15829) );
  AND2_X1 U11480 ( .A1(n11359), .A2(n10041), .ZN(n9677) );
  AND2_X1 U11481 ( .A1(n11359), .A2(n10041), .ZN(n9678) );
  AND2_X1 U11482 ( .A1(n11359), .A2(n10041), .ZN(n11560) );
  AND2_X1 U11483 ( .A1(n11359), .A2(n11354), .ZN(n9679) );
  AND2_X1 U11484 ( .A1(n11359), .A2(n11354), .ZN(n9680) );
  AND2_X1 U11485 ( .A1(n11359), .A2(n11354), .ZN(n11596) );
  AND2_X4 U11486 ( .A1(n11360), .A2(n11358), .ZN(n11545) );
  INV_X2 U11487 ( .A(n11615), .ZN(n12278) );
  AND2_X1 U11488 ( .A1(n11360), .A2(n11354), .ZN(n11551) );
  OR2_X2 U11489 ( .A1(n11626), .A2(n13011), .ZN(n9728) );
  NAND3_X2 U11490 ( .A1(n14950), .A2(n10148), .A3(n9905), .ZN(n12491) );
  XNOR2_X2 U11491 ( .A(n11157), .B(n10997), .ZN(n13872) );
  OAI21_X1 U11492 ( .B1(n14650), .B2(n14652), .A(n14651), .ZN(n14921) );
  XNOR2_X1 U11493 ( .A(n11786), .B(n20506), .ZN(n20618) );
  OR2_X2 U11494 ( .A1(n14651), .A2(n10192), .ZN(n10191) );
  INV_X2 U11495 ( .A(n14498), .ZN(n9681) );
  INV_X2 U11496 ( .A(n14498), .ZN(n9682) );
  INV_X2 U11497 ( .A(n14498), .ZN(n14461) );
  XNOR2_X2 U11498 ( .A(n9888), .B(n9670), .ZN(n20477) );
  AND2_X4 U11499 ( .A1(n14722), .A2(n14723), .ZN(n14707) );
  NAND2_X2 U11500 ( .A1(n11785), .A2(n11784), .ZN(n13697) );
  NAND3_X2 U11501 ( .A1(n9672), .A2(n13818), .A3(n9870), .ZN(n13817) );
  AND2_X1 U11502 ( .A1(n11360), .A2(n10041), .ZN(n9683) );
  INV_X1 U11503 ( .A(n11491), .ZN(n9684) );
  AND2_X1 U11504 ( .A1(n11360), .A2(n10041), .ZN(n11529) );
  AND2_X1 U11505 ( .A1(n11359), .A2(n11354), .ZN(n9692) );
  NOR2_X4 U11506 ( .A1(n13996), .A2(n14014), .ZN(n14013) );
  NOR2_X4 U11507 ( .A1(n11634), .A2(n10202), .ZN(n13002) );
  NOR2_X4 U11508 ( .A1(n14732), .A2(n14734), .ZN(n14722) );
  NAND3_X4 U11509 ( .A1(n11496), .A2(n11495), .A3(n10215), .ZN(n11567) );
  NOR2_X2 U11510 ( .A1(n13021), .A2(n12457), .ZN(n10027) );
  INV_X1 U11511 ( .A(n11575), .ZN(n9688) );
  AND2_X2 U11512 ( .A1(n11358), .A2(n11359), .ZN(n11558) );
  XNOR2_X2 U11513 ( .A(n11687), .B(n11686), .ZN(n11775) );
  OAI21_X1 U11514 ( .B1(n11667), .B2(n11666), .A(n11786), .ZN(n13657) );
  NAND2_X2 U11515 ( .A1(n13002), .A2(n9654), .ZN(n12449) );
  AND2_X1 U11516 ( .A1(n13669), .A2(n11359), .ZN(n9691) );
  AND2_X1 U11518 ( .A1(n14003), .A2(n10907), .ZN(n10021) );
  INV_X1 U11519 ( .A(n16408), .ZN(n10138) );
  XNOR2_X1 U11520 ( .A(n10869), .B(n10868), .ZN(n10866) );
  NAND2_X1 U11521 ( .A1(n10027), .A2(n11613), .ZN(n11621) );
  AOI21_X1 U11522 ( .B1(n10574), .B2(n10573), .A(n10572), .ZN(n10790) );
  INV_X1 U11523 ( .A(n10626), .ZN(n9841) );
  NOR2_X1 U11524 ( .A1(n10468), .A2(n9735), .ZN(n9914) );
  NAND2_X1 U11525 ( .A1(n10000), .A2(n9848), .ZN(n9855) );
  OAI22_X1 U11526 ( .A1(n10582), .A2(n10435), .B1(n10581), .B2(n10436), .ZN(
        n10437) );
  NAND2_X1 U11527 ( .A1(n10965), .A2(n10939), .ZN(n10335) );
  AOI21_X1 U11528 ( .B1(n18679), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12680), .ZN(n12686) );
  AND2_X1 U11529 ( .A1(n12797), .A2(n12796), .ZN(n12680) );
  OAI22_X1 U11530 ( .A1(n12678), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18906), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12685) );
  OR2_X1 U11531 ( .A1(n15194), .A2(n20865), .ZN(n12437) );
  INV_X1 U11532 ( .A(n14767), .ZN(n10180) );
  NAND2_X1 U11533 ( .A1(n11760), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12097) );
  INV_X1 U11534 ( .A(n13889), .ZN(n12434) );
  NOR2_X1 U11535 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13889) );
  INV_X1 U11536 ( .A(n12434), .ZN(n12523) );
  NOR2_X2 U11537 ( .A1(n11624), .A2(n11760), .ZN(n12052) );
  NAND2_X1 U11538 ( .A1(n12491), .A2(n15060), .ZN(n12488) );
  INV_X1 U11539 ( .A(n9906), .ZN(n9902) );
  NAND2_X1 U11540 ( .A1(n14998), .A2(n10154), .ZN(n9903) );
  INV_X1 U11541 ( .A(n14015), .ZN(n10051) );
  NOR2_X1 U11542 ( .A1(n10217), .A2(n11512), .ZN(n11513) );
  OAI21_X1 U11543 ( .B1(n11703), .B2(n11511), .A(n11510), .ZN(n11512) );
  INV_X1 U11544 ( .A(n12952), .ZN(n12961) );
  OAI21_X1 U11545 ( .B1(n11682), .B2(n11624), .A(n11567), .ZN(n11613) );
  OR2_X1 U11546 ( .A1(n12874), .A2(n11619), .ZN(n13029) );
  NOR2_X1 U11547 ( .A1(n10960), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10963) );
  INV_X1 U11548 ( .A(n14206), .ZN(n10130) );
  NAND2_X1 U11549 ( .A1(n10087), .A2(n13352), .ZN(n10086) );
  INV_X1 U11550 ( .A(n13284), .ZN(n10087) );
  AND2_X1 U11551 ( .A1(n13278), .A2(n14487), .ZN(n14450) );
  NAND2_X1 U11552 ( .A1(n11206), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15584) );
  AND2_X1 U11553 ( .A1(n9745), .A2(n10094), .ZN(n10093) );
  INV_X1 U11554 ( .A(n13708), .ZN(n10094) );
  AND4_X1 U11555 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n10535) );
  OAI21_X1 U11556 ( .B1(n14487), .B2(n11005), .A(n10687), .ZN(n11180) );
  NOR2_X1 U11557 ( .A1(n10552), .A2(n10549), .ZN(n10547) );
  NAND2_X1 U11558 ( .A1(n10547), .A2(n10546), .ZN(n10618) );
  NAND2_X1 U11559 ( .A1(n9852), .A2(n10000), .ZN(n10432) );
  AND2_X1 U11560 ( .A1(n10122), .A2(n19321), .ZN(n9852) );
  NAND2_X1 U11561 ( .A1(n10308), .A2(n10275), .ZN(n10316) );
  NAND2_X1 U11562 ( .A1(n10314), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10315) );
  NOR2_X1 U11563 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12679), .ZN(
        n12796) );
  NOR2_X1 U11564 ( .A1(n14075), .A2(n14074), .ZN(n15945) );
  NAND2_X1 U11565 ( .A1(n13326), .A2(n11630), .ZN(n12874) );
  OR2_X1 U11566 ( .A1(n14596), .A2(n20162), .ZN(n13328) );
  INV_X1 U11567 ( .A(n14533), .ZN(n10192) );
  INV_X1 U11568 ( .A(n12445), .ZN(n10194) );
  AND2_X1 U11569 ( .A1(n10810), .A2(n11200), .ZN(n11332) );
  INV_X1 U11570 ( .A(n14067), .ZN(n10020) );
  NAND2_X1 U11571 ( .A1(n13392), .A2(n13307), .ZN(n10120) );
  CLKBUF_X2 U11572 ( .A(n10984), .Z(n14577) );
  NAND2_X1 U11573 ( .A1(n13292), .A2(n10963), .ZN(n14579) );
  AND2_X1 U11574 ( .A1(n11257), .A2(n11256), .ZN(n14576) );
  NAND2_X1 U11575 ( .A1(n15397), .A2(n9809), .ZN(n9821) );
  AND2_X1 U11576 ( .A1(n15534), .A2(n15518), .ZN(n15520) );
  AND2_X1 U11577 ( .A1(n9653), .A2(n10332), .ZN(n13292) );
  NAND2_X1 U11578 ( .A1(n13433), .A2(n13432), .ZN(n9800) );
  INV_X1 U11579 ( .A(n13820), .ZN(n10898) );
  NAND2_X1 U11580 ( .A1(n10062), .A2(n16374), .ZN(n10061) );
  INV_X1 U11581 ( .A(n11277), .ZN(n10062) );
  NAND2_X1 U11582 ( .A1(n10136), .A2(n10069), .ZN(n10068) );
  INV_X1 U11583 ( .A(n15855), .ZN(n10069) );
  INV_X1 U11584 ( .A(n13277), .ZN(n19439) );
  OR2_X1 U11585 ( .A1(n20103), .A2(n20130), .ZN(n19757) );
  AND2_X1 U11586 ( .A1(n17753), .A2(n9774), .ZN(n9989) );
  NAND2_X1 U11587 ( .A1(n13277), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n9849) );
  CLKBUF_X1 U11588 ( .A(n11477), .Z(n12145) );
  INV_X1 U11589 ( .A(n11562), .ZN(n12503) );
  AOI21_X1 U11590 ( .B1(n10817), .B2(n10540), .A(n10539), .ZN(n10543) );
  INV_X1 U11591 ( .A(n15617), .ZN(n10143) );
  AOI21_X1 U11592 ( .B1(n10145), .B2(n15607), .A(n11294), .ZN(n10142) );
  AND2_X1 U11593 ( .A1(n10672), .A2(n10671), .ZN(n10690) );
  INV_X1 U11594 ( .A(n10981), .ZN(n11162) );
  NAND2_X1 U11595 ( .A1(n10222), .A2(n19097), .ZN(n10168) );
  NAND2_X1 U11596 ( .A1(n13291), .A2(n10939), .ZN(n10320) );
  NOR2_X1 U11597 ( .A1(n12637), .A2(n17581), .ZN(n12638) );
  NOR2_X1 U11598 ( .A1(n12815), .A2(n12816), .ZN(n12824) );
  NOR2_X1 U11599 ( .A1(n17600), .A2(n18448), .ZN(n12788) );
  NOR2_X1 U11600 ( .A1(n13900), .A2(n11623), .ZN(n13023) );
  NAND2_X1 U11601 ( .A1(n12869), .A2(n11622), .ZN(n11623) );
  NAND2_X1 U11602 ( .A1(n11523), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12215) );
  NOR2_X1 U11603 ( .A1(n14684), .A2(n10187), .ZN(n10186) );
  INV_X1 U11604 ( .A(n10188), .ZN(n10187) );
  NOR2_X1 U11605 ( .A1(n14696), .A2(n10189), .ZN(n10188) );
  INV_X1 U11606 ( .A(n14708), .ZN(n10189) );
  OR2_X1 U11607 ( .A1(n12184), .A2(n14710), .ZN(n12206) );
  INV_X1 U11608 ( .A(n14828), .ZN(n12038) );
  OAI211_X1 U11609 ( .C1(n14013), .C2(n9875), .A(n9871), .B(n9873), .ZN(n10183) );
  NAND2_X1 U11610 ( .A1(n9877), .A2(n9874), .ZN(n9873) );
  INV_X1 U11611 ( .A(n9877), .ZN(n9875) );
  INV_X1 U11612 ( .A(n14697), .ZN(n10054) );
  AND2_X1 U11613 ( .A1(n10056), .A2(n14724), .ZN(n10055) );
  INV_X1 U11614 ( .A(n14712), .ZN(n10056) );
  NAND2_X1 U11615 ( .A1(n10026), .A2(n16146), .ZN(n10156) );
  NAND2_X1 U11616 ( .A1(n16124), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10026) );
  NAND2_X1 U11617 ( .A1(n10157), .A2(n10156), .ZN(n10153) );
  NOR2_X1 U11618 ( .A1(n11891), .A2(n9908), .ZN(n9907) );
  INV_X1 U11619 ( .A(n11866), .ZN(n9908) );
  INV_X1 U11620 ( .A(n14009), .ZN(n10052) );
  INV_X1 U11621 ( .A(n12382), .ZN(n10152) );
  INV_X1 U11622 ( .A(n10177), .ZN(n10176) );
  OAI21_X1 U11623 ( .B1(n11722), .B2(n10178), .A(n11726), .ZN(n10177) );
  OR2_X1 U11624 ( .A1(n11741), .A2(n11740), .ZN(n12341) );
  INV_X1 U11625 ( .A(n11793), .ZN(n12325) );
  NOR2_X1 U11626 ( .A1(n11466), .A2(n11465), .ZN(n11482) );
  AOI21_X1 U11627 ( .B1(n11545), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n11470), .ZN(n11481) );
  OAI21_X1 U11628 ( .B1(n20958), .B2(n15188), .A(n15199), .ZN(n13720) );
  NAND2_X1 U11629 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20135), .ZN(
        n10795) );
  NOR2_X1 U11630 ( .A1(n11319), .A2(n11320), .ZN(n14548) );
  NOR2_X1 U11631 ( .A1(n10116), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10115) );
  OR2_X1 U11632 ( .A1(n10762), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10767) );
  OR2_X1 U11633 ( .A1(n9713), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10754) );
  AND2_X1 U11634 ( .A1(n10113), .A2(n9750), .ZN(n10112) );
  NOR2_X1 U11635 ( .A1(n10110), .A2(n10703), .ZN(n10109) );
  AND2_X1 U11636 ( .A1(n10621), .A2(n10620), .ZN(n10693) );
  AND2_X1 U11637 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10448), .ZN(
        n14358) );
  INV_X1 U11638 ( .A(n14450), .ZN(n14429) );
  NAND2_X1 U11639 ( .A1(n10280), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10281) );
  INV_X1 U11640 ( .A(n15416), .ZN(n10128) );
  NOR2_X1 U11641 ( .A1(n16418), .A2(n10040), .ZN(n10039) );
  INV_X1 U11642 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10040) );
  XNOR2_X1 U11643 ( .A(n10626), .B(n10627), .ZN(n11175) );
  NAND2_X1 U11644 ( .A1(n15573), .A2(n11301), .ZN(n11313) );
  NAND2_X1 U11645 ( .A1(n11300), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11301) );
  NOR2_X1 U11646 ( .A1(n15317), .A2(n10536), .ZN(n11323) );
  NAND2_X1 U11647 ( .A1(n15426), .A2(n15340), .ZN(n10016) );
  NOR2_X1 U11648 ( .A1(n15638), .A2(n15667), .ZN(n11274) );
  NOR2_X1 U11649 ( .A1(n10079), .A2(n10078), .ZN(n10077) );
  INV_X1 U11650 ( .A(n15637), .ZN(n10079) );
  INV_X1 U11651 ( .A(n15648), .ZN(n10078) );
  INV_X1 U11652 ( .A(n14579), .ZN(n11251) );
  NAND2_X1 U11653 ( .A1(n15877), .A2(n9835), .ZN(n15817) );
  INV_X1 U11654 ( .A(n11195), .ZN(n9835) );
  INV_X1 U11655 ( .A(n13085), .ZN(n10096) );
  NOR2_X1 U11656 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  INV_X1 U11657 ( .A(n13089), .ZN(n10007) );
  NOR2_X1 U11658 ( .A1(n15675), .A2(n15673), .ZN(n10141) );
  NOR2_X1 U11659 ( .A1(n13620), .A2(n10011), .ZN(n10010) );
  INV_X1 U11660 ( .A(n13545), .ZN(n10011) );
  INV_X1 U11661 ( .A(n11180), .ZN(n10688) );
  NAND2_X1 U11662 ( .A1(n14158), .A2(n14159), .ZN(n10697) );
  OR2_X1 U11663 ( .A1(n10384), .A2(n10275), .ZN(n10398) );
  AOI21_X1 U11664 ( .B1(n10399), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10403), .ZN(n10869) );
  OR2_X1 U11665 ( .A1(n10457), .A2(n10456), .ZN(n10993) );
  AND2_X1 U11666 ( .A1(n10333), .A2(n10196), .ZN(n10338) );
  AND2_X1 U11667 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13313) );
  NAND2_X1 U11668 ( .A1(n15374), .A2(n10417), .ZN(n10413) );
  NAND2_X1 U11669 ( .A1(n19439), .A2(n15374), .ZN(n10431) );
  INV_X1 U11670 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U11671 ( .A1(n9985), .A2(n17978), .ZN(n12664) );
  NOR2_X1 U11672 ( .A1(n9987), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9986) );
  NAND2_X1 U11673 ( .A1(n12656), .A2(n12657), .ZN(n9987) );
  AOI21_X1 U11674 ( .B1(n17565), .B2(n12623), .A(n17955), .ZN(n12649) );
  XNOR2_X1 U11675 ( .A(n17577), .B(n12638), .ZN(n12639) );
  XNOR2_X1 U11676 ( .A(n12824), .B(n17586), .ZN(n12825) );
  INV_X1 U11677 ( .A(n12788), .ZN(n12777) );
  NOR2_X1 U11678 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n17096), .ZN(
        n12575) );
  AND2_X1 U11679 ( .A1(n20198), .A2(n14268), .ZN(n14789) );
  INV_X1 U11680 ( .A(n20949), .ZN(n13903) );
  AND2_X1 U11681 ( .A1(n12941), .A2(n12940), .ZN(n14735) );
  AND2_X1 U11682 ( .A1(n12895), .A2(n12894), .ZN(n16302) );
  AOI21_X1 U11683 ( .B1(n12164), .B2(n12163), .A(n12162), .ZN(n14723) );
  NAND2_X1 U11684 ( .A1(n12371), .A2(n12052), .ZN(n11889) );
  INV_X1 U11685 ( .A(n12097), .ZN(n14531) );
  AND2_X1 U11686 ( .A1(n12446), .A2(n9741), .ZN(n14533) );
  OR2_X1 U11687 ( .A1(n14929), .A2(n12434), .ZN(n12238) );
  INV_X1 U11688 ( .A(n12494), .ZN(n10147) );
  NAND2_X1 U11689 ( .A1(n15035), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10148) );
  NOR2_X1 U11690 ( .A1(n11503), .A2(n11502), .ZN(n11515) );
  NAND2_X1 U11691 ( .A1(n16171), .A2(n12370), .ZN(n16166) );
  AND2_X1 U11692 ( .A1(n16015), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13373) );
  NOR2_X1 U11693 ( .A1(n9689), .A2(n20506), .ZN(n20589) );
  NAND2_X1 U11694 ( .A1(n13690), .A2(n13692), .ZN(n20587) );
  NOR2_X1 U11695 ( .A1(n20685), .A2(n15217), .ZN(n20769) );
  NAND2_X1 U11696 ( .A1(n20865), .A2(n13720), .ZN(n15217) );
  NOR2_X1 U11697 ( .A1(n14595), .A2(n14596), .ZN(n16004) );
  OR2_X1 U11698 ( .A1(n10792), .A2(n10791), .ZN(n10794) );
  NOR2_X1 U11699 ( .A1(n16324), .A2(n19288), .ZN(n15279) );
  NOR2_X1 U11700 ( .A1(n11298), .A2(n10116), .ZN(n11308) );
  AND2_X1 U11701 ( .A1(n11314), .A2(n14554), .ZN(n11303) );
  AND2_X1 U11702 ( .A1(n15250), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15247) );
  AND2_X1 U11703 ( .A1(n11337), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15265) );
  NAND2_X1 U11704 ( .A1(n10714), .A2(n13630), .ZN(n10725) );
  AOI22_X1 U11705 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n14567), .B2(n19097), .ZN(
        n15243) );
  OR2_X1 U11706 ( .A1(n11076), .A2(n11075), .ZN(n13641) );
  INV_X1 U11707 ( .A(n9796), .ZN(n9795) );
  OAI21_X1 U11708 ( .B1(n9809), .B2(n9797), .A(n14492), .ZN(n9796) );
  INV_X1 U11709 ( .A(n9818), .ZN(n9797) );
  NOR2_X1 U11710 ( .A1(n15483), .A2(n10099), .ZN(n11257) );
  OR3_X1 U11711 ( .A1(n15307), .A2(n10100), .A3(n10102), .ZN(n10099) );
  OAI211_X1 U11712 ( .C1(n9811), .C2(n9812), .A(n9810), .B(n14453), .ZN(n9808)
         );
  INV_X1 U11713 ( .A(n11242), .ZN(n10098) );
  OR2_X1 U11714 ( .A1(n13970), .A2(n13969), .ZN(n13971) );
  NOR2_X1 U11715 ( .A1(n13285), .A2(n9744), .ZN(n13429) );
  AND2_X1 U11716 ( .A1(n9781), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9935) );
  NOR2_X1 U11717 ( .A1(n14582), .A2(n11317), .ZN(n10173) );
  NOR2_X1 U11718 ( .A1(n9788), .A2(n9930), .ZN(n9929) );
  XNOR2_X1 U11719 ( .A(n11323), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11311) );
  AND2_X1 U11720 ( .A1(n9709), .A2(n15335), .ZN(n10097) );
  OR2_X1 U11721 ( .A1(n15331), .A2(n10536), .ZN(n15595) );
  OAI21_X1 U11722 ( .B1(n11284), .B2(n15617), .A(n15615), .ZN(n10145) );
  NAND2_X1 U11723 ( .A1(n10067), .A2(n9697), .ZN(n11285) );
  INV_X1 U11724 ( .A(n10077), .ZN(n10073) );
  INV_X1 U11725 ( .A(n11280), .ZN(n10072) );
  INV_X1 U11726 ( .A(n10075), .ZN(n10074) );
  NOR2_X1 U11727 ( .A1(n10774), .A2(n9751), .ZN(n10075) );
  NAND2_X1 U11728 ( .A1(n15647), .A2(n10077), .ZN(n10076) );
  INV_X1 U11729 ( .A(n14185), .ZN(n10019) );
  AND2_X1 U11730 ( .A1(n13987), .A2(n10088), .ZN(n15534) );
  AND2_X1 U11731 ( .A1(n10090), .A2(n10089), .ZN(n10088) );
  INV_X1 U11732 ( .A(n15531), .ZN(n10089) );
  NAND2_X1 U11733 ( .A1(n13836), .A2(n10021), .ZN(n14068) );
  AOI21_X1 U11734 ( .B1(n10059), .B2(n10061), .A(n15667), .ZN(n10058) );
  INV_X1 U11735 ( .A(n10061), .ZN(n10060) );
  INV_X1 U11736 ( .A(n10063), .ZN(n10059) );
  AND2_X1 U11737 ( .A1(n16374), .A2(n15834), .ZN(n10063) );
  OR2_X1 U11738 ( .A1(n10731), .A2(n16468), .ZN(n16391) );
  NAND2_X1 U11739 ( .A1(n9916), .A2(n10722), .ZN(n10070) );
  NAND2_X1 U11740 ( .A1(n9917), .A2(n14158), .ZN(n9916) );
  NOR2_X1 U11741 ( .A1(n13619), .A2(n10008), .ZN(n13556) );
  OAI21_X1 U11742 ( .B1(n10163), .B2(n10166), .A(n14160), .ZN(n10162) );
  AND2_X1 U11743 ( .A1(n11014), .A2(n11013), .ZN(n13284) );
  AOI21_X1 U11744 ( .B1(n9752), .B2(n13800), .A(n9923), .ZN(n9922) );
  NOR2_X1 U11745 ( .A1(n13863), .A2(n16522), .ZN(n9923) );
  NOR2_X1 U11746 ( .A1(n13800), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9924) );
  AND2_X1 U11747 ( .A1(n10990), .A2(n9754), .ZN(n10084) );
  INV_X1 U11748 ( .A(n13783), .ZN(n10085) );
  AND2_X1 U11749 ( .A1(n16539), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10376) );
  OAI21_X1 U11750 ( .B1(n13277), .B2(n13307), .A(n13276), .ZN(n13281) );
  NAND2_X1 U11751 ( .A1(n9825), .A2(n9824), .ZN(n9823) );
  INV_X1 U11752 ( .A(n13393), .ZN(n9824) );
  INV_X1 U11753 ( .A(n13438), .ZN(n9825) );
  NAND2_X1 U11754 ( .A1(n9851), .A2(n13277), .ZN(n9850) );
  AND2_X1 U11755 ( .A1(n9639), .A2(n10417), .ZN(n10418) );
  NOR2_X1 U11756 ( .A1(n9854), .A2(n9853), .ZN(n9857) );
  NOR2_X1 U11757 ( .A1(n20111), .A2(n20121), .ZN(n19755) );
  NOR2_X1 U11758 ( .A1(n15374), .A2(n19439), .ZN(n9928) );
  AND2_X1 U11759 ( .A1(n20111), .A2(n20099), .ZN(n19894) );
  AND2_X1 U11760 ( .A1(n9639), .A2(n19439), .ZN(n9927) );
  INV_X1 U11761 ( .A(n14487), .ZN(n10458) );
  NOR2_X1 U11762 ( .A1(n20103), .A2(n19713), .ZN(n19921) );
  INV_X1 U11763 ( .A(n19757), .ZN(n19895) );
  NAND2_X1 U11764 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19964), .ZN(n19498) );
  INV_X1 U11765 ( .A(n20107), .ZN(n19969) );
  INV_X1 U11766 ( .A(n19964), .ZN(n19889) );
  NAND2_X1 U11767 ( .A1(n10832), .A2(n10831), .ZN(n13488) );
  OR2_X1 U11768 ( .A1(n10830), .A2(n13223), .ZN(n10831) );
  AOI21_X1 U11769 ( .B1(n12799), .B2(n12801), .A(n12798), .ZN(n18856) );
  NAND2_X1 U11770 ( .A1(n9972), .A2(n9969), .ZN(n16762) );
  INV_X1 U11771 ( .A(n9970), .ZN(n9969) );
  OAI21_X1 U11772 ( .B1(n9975), .B2(n9971), .A(n9974), .ZN(n9970) );
  AOI21_X1 U11773 ( .B1(n17083), .B2(n17822), .A(n17803), .ZN(n9963) );
  INV_X1 U11774 ( .A(n19089), .ZN(n19067) );
  NOR2_X1 U11775 ( .A1(n14076), .A2(n15945), .ZN(n16038) );
  NOR3_X2 U11776 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18888), .ZN(n12582) );
  INV_X1 U11777 ( .A(n12776), .ZN(n17640) );
  AND2_X1 U11778 ( .A1(n17739), .A2(n9755), .ZN(n16567) );
  INV_X1 U11779 ( .A(n18276), .ZN(n17904) );
  INV_X1 U11780 ( .A(n17765), .ZN(n9869) );
  INV_X1 U11781 ( .A(n18142), .ZN(n17885) );
  NOR2_X1 U11782 ( .A1(n9863), .A2(n12658), .ZN(n17977) );
  NAND2_X1 U11783 ( .A1(n18276), .A2(n17955), .ZN(n9863) );
  NAND2_X1 U11784 ( .A1(n18005), .A2(n9731), .ZN(n9937) );
  INV_X1 U11785 ( .A(n18000), .ZN(n9936) );
  NAND2_X1 U11786 ( .A1(n18005), .A2(n12836), .ZN(n17999) );
  NAND2_X1 U11787 ( .A1(n18023), .A2(n12645), .ZN(n18008) );
  XNOR2_X1 U11788 ( .A(n12639), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18032) );
  INV_X1 U11789 ( .A(n18856), .ZN(n16710) );
  NOR2_X1 U11790 ( .A1(n18436), .A2(n12802), .ZN(n15961) );
  NAND2_X1 U11791 ( .A1(n13264), .A2(n13296), .ZN(n20949) );
  NAND2_X1 U11792 ( .A1(n12448), .A2(n12447), .ZN(n10193) );
  OR2_X1 U11793 ( .A1(n20338), .A2(n13517), .ZN(n20349) );
  NAND2_X1 U11794 ( .A1(n10044), .A2(n10042), .ZN(n15059) );
  OR2_X1 U11795 ( .A1(n14610), .A2(n10045), .ZN(n10044) );
  XNOR2_X1 U11796 ( .A(n14612), .B(n12899), .ZN(n10045) );
  NAND2_X1 U11797 ( .A1(n10025), .A2(n10024), .ZN(n14530) );
  NAND2_X1 U11798 ( .A1(n14527), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10025) );
  NAND2_X1 U11799 ( .A1(n14529), .A2(n14528), .ZN(n10024) );
  XNOR2_X1 U11800 ( .A(n12498), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15077) );
  NAND2_X1 U11801 ( .A1(n12497), .A2(n12496), .ZN(n12498) );
  CLKBUF_X1 U11802 ( .A(n13702), .Z(n20619) );
  NOR2_X1 U11803 ( .A1(n13916), .A2(n13690), .ZN(n20680) );
  INV_X1 U11804 ( .A(n20622), .ZN(n20643) );
  NAND2_X1 U11805 ( .A1(n11332), .A2(n11331), .ZN(n13124) );
  INV_X1 U11806 ( .A(n19320), .ZN(n19285) );
  AND2_X1 U11807 ( .A1(n9712), .A2(n12857), .ZN(n16338) );
  OR2_X1 U11808 ( .A1(n11060), .A2(n11059), .ZN(n13551) );
  INV_X1 U11809 ( .A(n15450), .ZN(n15434) );
  NAND2_X1 U11810 ( .A1(n15440), .A2(n10332), .ZN(n15450) );
  OAI211_X1 U11811 ( .C1(n15544), .C2(n15545), .A(n15546), .B(n15543), .ZN(
        n14558) );
  AND2_X1 U11812 ( .A1(n16453), .A2(n20117), .ZN(n19428) );
  INV_X1 U11813 ( .A(n16440), .ZN(n19432) );
  AND2_X1 U11814 ( .A1(n16453), .A2(n13245), .ZN(n16440) );
  NAND2_X1 U11815 ( .A1(n14591), .A2(n14590), .ZN(n9837) );
  NAND2_X1 U11816 ( .A1(n19332), .A2(n19436), .ZN(n14590) );
  NAND2_X1 U11817 ( .A1(n15382), .A2(n19440), .ZN(n14591) );
  XNOR2_X1 U11818 ( .A(n15542), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15703) );
  NAND2_X1 U11819 ( .A1(n9932), .A2(n12849), .ZN(n15556) );
  NAND2_X1 U11820 ( .A1(n9933), .A2(n11317), .ZN(n9932) );
  XNOR2_X1 U11821 ( .A(n9842), .B(n12855), .ZN(n15564) );
  NAND2_X1 U11822 ( .A1(n15713), .A2(n9843), .ZN(n9842) );
  NAND2_X1 U11823 ( .A1(n12852), .A2(n9844), .ZN(n9843) );
  INV_X1 U11824 ( .A(n15831), .ZN(n9858) );
  NAND2_X1 U11825 ( .A1(n9861), .A2(n9859), .ZN(n15831) );
  NOR2_X1 U11826 ( .A1(n16460), .A2(n9860), .ZN(n9859) );
  INV_X1 U11827 ( .A(n15815), .ZN(n9861) );
  AND2_X1 U11828 ( .A1(n15816), .A2(n16455), .ZN(n9860) );
  INV_X1 U11829 ( .A(n19440), .ZN(n16527) );
  OR2_X1 U11830 ( .A1(n13314), .A2(n13271), .ZN(n20130) );
  INV_X1 U11831 ( .A(n17126), .ZN(n17091) );
  INV_X1 U11832 ( .A(n17121), .ZN(n17095) );
  INV_X1 U11833 ( .A(n17127), .ZN(n17116) );
  AOI21_X1 U11834 ( .B1(n18248), .B2(n18149), .A(n9945), .ZN(n9944) );
  OAI21_X1 U11835 ( .B1(n18363), .B2(n18160), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9945) );
  AND2_X1 U11836 ( .A1(n9942), .A2(n18382), .ZN(n9941) );
  OAI21_X1 U11837 ( .B1(n18152), .B2(n18150), .A(n18151), .ZN(n9942) );
  AOI21_X1 U11838 ( .B1(n10589), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n10499), .ZN(n10462) );
  NAND2_X1 U11839 ( .A1(n10822), .A2(n10823), .ZN(n9830) );
  NAND2_X1 U11840 ( .A1(n13269), .A2(n9653), .ZN(n10354) );
  OAI21_X1 U11841 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n12678), .A(
        n12681), .ZN(n12682) );
  OR2_X1 U11842 ( .A1(n12685), .A2(n12686), .ZN(n12681) );
  AND2_X1 U11843 ( .A1(n13691), .A2(n11843), .ZN(n10028) );
  NOR2_X1 U11844 ( .A1(n12198), .A2(n11568), .ZN(n11570) );
  INV_X1 U11845 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11568) );
  NOR2_X1 U11846 ( .A1(n9878), .A2(n9874), .ZN(n9872) );
  AOI21_X1 U11847 ( .B1(n14778), .B2(n11978), .A(n11977), .ZN(n9878) );
  AND2_X1 U11848 ( .A1(n11977), .A2(n14778), .ZN(n9877) );
  INV_X1 U11849 ( .A(n14024), .ZN(n9874) );
  OR2_X1 U11850 ( .A1(n11881), .A2(n11880), .ZN(n12377) );
  OR2_X1 U11851 ( .A1(n11823), .A2(n11822), .ZN(n12364) );
  INV_X1 U11852 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U11853 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11539), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U11854 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11457) );
  OR2_X1 U11855 ( .A1(n13900), .A2(n20865), .ZN(n11792) );
  NAND2_X1 U11856 ( .A1(n10545), .A2(n10544), .ZN(n10570) );
  AND2_X1 U11857 ( .A1(n10112), .A2(n9759), .ZN(n10111) );
  AND4_X1 U11858 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10534) );
  NOR2_X1 U11859 ( .A1(n9724), .A2(n9913), .ZN(n9912) );
  OR2_X1 U11860 ( .A1(n10354), .A2(n10334), .ZN(n10336) );
  NAND2_X1 U11861 ( .A1(n10106), .A2(n10105), .ZN(n10549) );
  NAND2_X1 U11862 ( .A1(n14552), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10105) );
  NAND2_X1 U11863 ( .A1(n10802), .A2(n11295), .ZN(n10106) );
  NAND2_X1 U11864 ( .A1(n13291), .A2(n10837), .ZN(n10835) );
  AOI22_X1 U11865 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10264) );
  INV_X1 U11866 ( .A(n10354), .ZN(n10846) );
  NOR2_X1 U11867 ( .A1(n18441), .A2(n17447), .ZN(n12804) );
  OR2_X1 U11868 ( .A1(n12439), .A2(n14621), .ZN(n12441) );
  NOR2_X1 U11869 ( .A1(n14894), .A2(n10182), .ZN(n10181) );
  INV_X1 U11870 ( .A(n14833), .ZN(n10048) );
  NOR2_X1 U11871 ( .A1(n12198), .A2(n11501), .ZN(n11502) );
  INV_X1 U11872 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11501) );
  AND2_X1 U11873 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  NAND2_X1 U11874 ( .A1(n12869), .A2(n11630), .ZN(n12457) );
  INV_X1 U11875 ( .A(n12967), .ZN(n12946) );
  NOR2_X1 U11876 ( .A1(n11643), .A2(n13013), .ZN(n11632) );
  INV_X1 U11877 ( .A(n20477), .ZN(n11749) );
  INV_X1 U11878 ( .A(n11745), .ZN(n10179) );
  OR2_X1 U11879 ( .A1(n11807), .A2(n11806), .ZN(n12355) );
  INV_X1 U11880 ( .A(n12301), .ZN(n12307) );
  INV_X1 U11881 ( .A(n11620), .ZN(n13365) );
  NAND2_X1 U11882 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11535) );
  AND2_X1 U11883 ( .A1(n20728), .A2(n11661), .ZN(n13924) );
  NOR2_X1 U11884 ( .A1(n12301), .A2(n12338), .ZN(n12303) );
  AND2_X1 U11885 ( .A1(n12272), .A2(n12304), .ZN(n12450) );
  OR2_X1 U11886 ( .A1(n12305), .A2(n12271), .ZN(n12272) );
  OR2_X1 U11887 ( .A1(n10513), .A2(n10512), .ZN(n10981) );
  NAND2_X1 U11888 ( .A1(n11265), .A2(n11264), .ZN(n11319) );
  NAND2_X1 U11889 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  INV_X1 U11890 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10118) );
  NOR2_X1 U11891 ( .A1(n10732), .A2(n10114), .ZN(n10113) );
  INV_X1 U11892 ( .A(n10723), .ZN(n10114) );
  NAND2_X1 U11893 ( .A1(n10101), .A2(n15292), .ZN(n10100) );
  INV_X1 U11894 ( .A(n15484), .ZN(n10101) );
  INV_X1 U11895 ( .A(n10206), .ZN(n9817) );
  INV_X1 U11896 ( .A(n15439), .ZN(n14319) );
  AND2_X1 U11897 ( .A1(n14181), .A2(n14058), .ZN(n10131) );
  NAND3_X1 U11898 ( .A1(n10361), .A2(n10339), .A3(n10928), .ZN(n10364) );
  NOR2_X1 U11899 ( .A1(n11316), .A2(n11317), .ZN(n9952) );
  AND2_X1 U11900 ( .A1(n11312), .A2(n10132), .ZN(n9955) );
  AND2_X1 U11901 ( .A1(n10135), .A2(n11321), .ZN(n10132) );
  INV_X1 U11902 ( .A(n10133), .ZN(n9954) );
  AOI21_X1 U11903 ( .B1(n11321), .B2(n9782), .A(n10134), .ZN(n10133) );
  INV_X1 U11904 ( .A(n12850), .ZN(n10134) );
  NOR2_X1 U11905 ( .A1(n15661), .A2(n10035), .ZN(n10034) );
  AOI21_X1 U11906 ( .B1(n9922), .B2(n9924), .A(n9921), .ZN(n9920) );
  INV_X1 U11907 ( .A(n13870), .ZN(n9921) );
  NAND2_X1 U11908 ( .A1(n10866), .A2(n10119), .ZN(n10121) );
  INV_X1 U11909 ( .A(n10396), .ZN(n9804) );
  NOR2_X1 U11910 ( .A1(n15743), .A2(n15745), .ZN(n15719) );
  AND2_X1 U11911 ( .A1(n9736), .A2(n9697), .ZN(n9846) );
  INV_X1 U11912 ( .A(n10142), .ZN(n9845) );
  OR2_X1 U11913 ( .A1(n10172), .A2(n11231), .ZN(n10171) );
  NAND2_X1 U11914 ( .A1(n11197), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10172) );
  NOR2_X1 U11915 ( .A1(n14059), .A2(n10091), .ZN(n10090) );
  INV_X1 U11916 ( .A(n13988), .ZN(n10091) );
  AND2_X1 U11917 ( .A1(n16371), .A2(n16373), .ZN(n11277) );
  INV_X1 U11918 ( .A(n13963), .ZN(n10907) );
  INV_X1 U11919 ( .A(n13083), .ZN(n10095) );
  INV_X1 U11920 ( .A(n13553), .ZN(n10009) );
  AND2_X1 U11921 ( .A1(n14233), .A2(n11186), .ZN(n10163) );
  AND2_X1 U11922 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11189) );
  NAND2_X1 U11923 ( .A1(n9847), .A2(n19274), .ZN(n10695) );
  OR2_X1 U11924 ( .A1(n10613), .A2(n10612), .ZN(n11001) );
  NAND2_X1 U11925 ( .A1(n10458), .A2(n10993), .ZN(n10459) );
  OAI211_X1 U11926 ( .C1(n11150), .C2(n20152), .A(n10353), .B(n10352), .ZN(
        n10370) );
  NAND2_X1 U11927 ( .A1(n10368), .A2(n20152), .ZN(n10353) );
  NAND2_X1 U11928 ( .A1(n10169), .A2(n13592), .ZN(n10378) );
  NOR2_X1 U11929 ( .A1(n9834), .A2(n19470), .ZN(n9833) );
  AND2_X1 U11930 ( .A1(n10973), .A2(n10972), .ZN(n10979) );
  NOR2_X1 U11931 ( .A1(n10486), .A2(n10485), .ZN(n11159) );
  INV_X1 U11932 ( .A(n10393), .ZN(n13304) );
  AND3_X1 U11933 ( .A1(n10355), .A2(n10499), .A3(n13291), .ZN(n10935) );
  OR2_X1 U11934 ( .A1(n14429), .A2(n13300), .ZN(n13394) );
  NAND2_X1 U11935 ( .A1(n9840), .A2(n10411), .ZN(n10582) );
  INV_X1 U11936 ( .A(n10433), .ZN(n9840) );
  NAND2_X1 U11937 ( .A1(n10427), .A2(n15374), .ZN(n19815) );
  AND4_X1 U11938 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  NAND2_X1 U11939 ( .A1(n10301), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10302) );
  INV_X1 U11940 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10221) );
  NAND3_X1 U11941 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20107), .A3(n19964), 
        .ZN(n19452) );
  INV_X1 U11942 ( .A(n13221), .ZN(n13502) );
  NAND2_X1 U11944 ( .A1(n9976), .A2(n16773), .ZN(n9974) );
  INV_X1 U11945 ( .A(n17710), .ZN(n9971) );
  OR2_X1 U11947 ( .A1(n18884), .A2(n9866), .ZN(n14122) );
  NAND2_X1 U11948 ( .A1(n12533), .A2(n12679), .ZN(n9866) );
  NAND2_X1 U11949 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12539) );
  NAND2_X1 U11950 ( .A1(n12576), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12568) );
  NAND2_X1 U11951 ( .A1(n18871), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14110) );
  NAND2_X1 U11952 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12533), .ZN(
        n12542) );
  NOR2_X1 U11953 ( .A1(n17906), .A2(n9982), .ZN(n9981) );
  NAND2_X1 U11954 ( .A1(n18044), .A2(n12829), .ZN(n12830) );
  INV_X1 U11955 ( .A(n17593), .ZN(n12816) );
  XNOR2_X1 U11956 ( .A(n9867), .B(n17593), .ZN(n12635) );
  NOR2_X1 U11957 ( .A1(n19074), .A2(n12776), .ZN(n16730) );
  INV_X1 U11958 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20196) );
  OR2_X1 U11959 ( .A1(n20949), .A2(n13906), .ZN(n20198) );
  AND2_X1 U11960 ( .A1(n12920), .A2(n12919), .ZN(n16077) );
  AND3_X1 U11961 ( .A1(n11940), .A2(n11939), .A3(n11938), .ZN(n14014) );
  INV_X1 U11962 ( .A(n11630), .ZN(n11622) );
  NOR2_X1 U11963 ( .A1(n13696), .A2(n13814), .ZN(n13813) );
  OR2_X1 U11964 ( .A1(n14909), .A2(n12434), .ZN(n12259) );
  AOI21_X1 U11965 ( .B1(n12249), .B2(n12248), .A(n12247), .ZN(n14652) );
  AND2_X1 U11966 ( .A1(n14913), .A2(n12523), .ZN(n12247) );
  NAND2_X1 U11967 ( .A1(n11524), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12236) );
  AND2_X1 U11968 ( .A1(n12240), .A2(n10186), .ZN(n10185) );
  NOR2_X1 U11969 ( .A1(n14673), .A2(n14660), .ZN(n12240) );
  AND2_X1 U11970 ( .A1(n12187), .A2(n12186), .ZN(n14708) );
  INV_X1 U11971 ( .A(n12117), .ZN(n11521) );
  NAND2_X1 U11972 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n11520), .ZN(
        n12117) );
  INV_X1 U11973 ( .A(n12096), .ZN(n11520) );
  NAND2_X1 U11974 ( .A1(n12062), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12096) );
  CLKBUF_X1 U11975 ( .A(n14765), .Z(n14766) );
  NAND2_X1 U11976 ( .A1(n12018), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12039) );
  CLKBUF_X1 U11977 ( .A(n14828), .Z(n14829) );
  NOR2_X1 U11978 ( .A1(n11959), .A2(n15038), .ZN(n11993) );
  NAND2_X1 U11979 ( .A1(n11941), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11959) );
  NOR2_X1 U11980 ( .A1(n11936), .A2(n14792), .ZN(n11941) );
  NAND2_X1 U11981 ( .A1(n11917), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11936) );
  AND3_X1 U11982 ( .A1(n11920), .A2(n11919), .A3(n11918), .ZN(n13998) );
  CLKBUF_X1 U11983 ( .A(n13996), .Z(n13997) );
  NOR2_X1 U11984 ( .A1(n11894), .A2(n20196), .ZN(n11917) );
  INV_X1 U11985 ( .A(n11900), .ZN(n11901) );
  INV_X1 U11986 ( .A(n13814), .ZN(n9870) );
  INV_X1 U11987 ( .A(n11860), .ZN(n11884) );
  NAND2_X1 U11988 ( .A1(n11861), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11860) );
  NOR2_X1 U11989 ( .A1(n11834), .A2(n20235), .ZN(n11861) );
  INV_X1 U11990 ( .A(n11762), .ZN(n11835) );
  NAND2_X1 U11991 ( .A1(n11835), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11834) );
  NAND2_X1 U11992 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11762) );
  OAI21_X1 U11993 ( .B1(n13915), .B2(n12338), .A(n12334), .ZN(n20340) );
  XNOR2_X1 U11994 ( .A(n14612), .B(n14609), .ZN(n10043) );
  NAND2_X1 U11995 ( .A1(n9746), .A2(n14247), .ZN(n10146) );
  NOR2_X1 U11996 ( .A1(n12495), .A2(n10023), .ZN(n10022) );
  INV_X1 U11997 ( .A(n15087), .ZN(n10023) );
  NAND2_X1 U11998 ( .A1(n14665), .A2(n12966), .ZN(n14634) );
  AND2_X1 U11999 ( .A1(n14662), .A2(n14663), .ZN(n14665) );
  NAND2_X1 U12000 ( .A1(n14949), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14922) );
  AND2_X1 U12001 ( .A1(n14737), .A2(n9758), .ZN(n14687) );
  INV_X1 U12002 ( .A(n14688), .ZN(n10053) );
  NAND2_X1 U12003 ( .A1(n14737), .A2(n9743), .ZN(n14699) );
  AND4_X1 U12004 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n16206), .A4(n13047), .ZN(
        n13048) );
  NAND2_X1 U12005 ( .A1(n9899), .A2(n15035), .ZN(n14950) );
  NAND2_X1 U12006 ( .A1(n10153), .A2(n9900), .ZN(n9899) );
  NAND2_X1 U12007 ( .A1(n14737), .A2(n10055), .ZN(n14714) );
  INV_X1 U12008 ( .A(n10158), .ZN(n10155) );
  AND2_X1 U12009 ( .A1(n12938), .A2(n12937), .ZN(n14751) );
  INV_X1 U12010 ( .A(n12401), .ZN(n16125) );
  NOR3_X1 U12011 ( .A1(n16081), .A2(n14833), .A3(n10049), .ZN(n14826) );
  NOR2_X1 U12012 ( .A1(n16081), .A2(n14833), .ZN(n14832) );
  NAND2_X1 U12013 ( .A1(n9740), .A2(n10029), .ZN(n15009) );
  OR2_X1 U12014 ( .A1(n16146), .A2(n12403), .ZN(n15028) );
  OR2_X1 U12015 ( .A1(n16146), .A2(n12402), .ZN(n15026) );
  AND2_X1 U12016 ( .A1(n9727), .A2(n14210), .ZN(n10050) );
  AND2_X1 U12017 ( .A1(n16305), .A2(n9727), .ZN(n14211) );
  NAND2_X1 U12018 ( .A1(n16305), .A2(n9719), .ZN(n14016) );
  NAND2_X1 U12019 ( .A1(n16305), .A2(n12903), .ZN(n16290) );
  AND2_X1 U12020 ( .A1(n12902), .A2(n12901), .ZN(n16287) );
  AND2_X1 U12021 ( .A1(n16303), .A2(n16302), .ZN(n16305) );
  INV_X1 U12022 ( .A(n15175), .ZN(n16269) );
  AND2_X1 U12023 ( .A1(n12890), .A2(n10046), .ZN(n16303) );
  AND2_X1 U12024 ( .A1(n9716), .A2(n12889), .ZN(n10046) );
  AND2_X1 U12025 ( .A1(n12890), .A2(n12889), .ZN(n13774) );
  NOR2_X1 U12026 ( .A1(n13056), .A2(n13033), .ZN(n15170) );
  OAI21_X1 U12027 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11657), .A(
        n11656), .ZN(n11658) );
  NAND2_X1 U12028 ( .A1(n11753), .A2(n11752), .ZN(n12339) );
  INV_X1 U12029 ( .A(n13765), .ZN(n13750) );
  NAND2_X1 U12030 ( .A1(n13916), .A2(n13915), .ZN(n20485) );
  INV_X1 U12031 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20647) );
  NAND2_X1 U12032 ( .A1(n13688), .A2(n15191), .ZN(n20586) );
  AOI21_X1 U12033 ( .B1(n20647), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n15217), 
        .ZN(n20809) );
  INV_X1 U12034 ( .A(n20677), .ZN(n20802) );
  NAND2_X1 U12035 ( .A1(n10326), .A2(n10358), .ZN(n10333) );
  OAI21_X1 U12036 ( .B1(n10981), .B2(n10358), .A(n10107), .ZN(n10802) );
  NAND2_X1 U12037 ( .A1(n10358), .A2(n10815), .ZN(n10107) );
  AND2_X1 U12038 ( .A1(n10830), .A2(n10797), .ZN(n13579) );
  OR2_X1 U12039 ( .A1(n15333), .A2(n15608), .ZN(n10030) );
  AND2_X1 U12040 ( .A1(n10748), .A2(n10754), .ZN(n19191) );
  NAND2_X1 U12041 ( .A1(n10724), .A2(n10113), .ZN(n10743) );
  NAND2_X1 U12042 ( .A1(n10724), .A2(n10723), .ZN(n10733) );
  AND2_X1 U12043 ( .A1(n10700), .A2(n9700), .ZN(n10714) );
  NAND2_X1 U12044 ( .A1(n10700), .A2(n10109), .ZN(n10710) );
  OR2_X1 U12045 ( .A1(n11136), .A2(n11135), .ZN(n13961) );
  NOR2_X1 U12046 ( .A1(n9819), .A2(n15392), .ZN(n9818) );
  NAND2_X1 U12047 ( .A1(n14434), .A2(n9767), .ZN(n10123) );
  NOR3_X1 U12048 ( .A1(n15483), .A2(n15307), .A3(n15484), .ZN(n15306) );
  NAND2_X1 U12049 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  NAND2_X1 U12050 ( .A1(n14371), .A2(n10128), .ZN(n9822) );
  INV_X1 U12051 ( .A(n15422), .ZN(n10127) );
  NOR2_X1 U12052 ( .A1(n15423), .A2(n15422), .ZN(n15421) );
  CLKBUF_X1 U12053 ( .A(n14306), .Z(n14205) );
  NAND2_X1 U12054 ( .A1(n13987), .A2(n13988), .ZN(n14060) );
  AND3_X1 U12055 ( .A1(n11079), .A2(n11078), .A3(n11077), .ZN(n13085) );
  AND3_X1 U12056 ( .A1(n11048), .A2(n11047), .A3(n11046), .ZN(n13422) );
  OR2_X1 U12057 ( .A1(n19379), .A2(n13294), .ZN(n13990) );
  AND2_X1 U12058 ( .A1(n13222), .A2(n20151), .ZN(n19388) );
  INV_X1 U12059 ( .A(n13201), .ZN(n19453) );
  XNOR2_X1 U12060 ( .A(n13072), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14567) );
  NAND2_X1 U12061 ( .A1(n9953), .A2(n9950), .ZN(n14546) );
  NAND2_X1 U12062 ( .A1(n11313), .A2(n9951), .ZN(n9950) );
  AOI21_X1 U12063 ( .B1(n11313), .B2(n9955), .A(n9954), .ZN(n9953) );
  AND2_X1 U12064 ( .A1(n11312), .A2(n9952), .ZN(n9951) );
  AND2_X1 U12065 ( .A1(n15247), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15246) );
  NAND2_X1 U12066 ( .A1(n15247), .A2(n9708), .ZN(n15244) );
  AND2_X1 U12067 ( .A1(n15265), .A2(n9773), .ZN(n15250) );
  NAND2_X1 U12068 ( .A1(n15265), .A2(n9704), .ZN(n15251) );
  AND2_X1 U12069 ( .A1(n15265), .A2(n9764), .ZN(n15254) );
  AND2_X1 U12070 ( .A1(n15261), .A2(n10033), .ZN(n15264) );
  AND2_X1 U12071 ( .A1(n9701), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10033) );
  NAND2_X1 U12072 ( .A1(n15261), .A2(n9701), .ZN(n15262) );
  NAND2_X1 U12073 ( .A1(n15261), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15260) );
  NOR2_X1 U12074 ( .A1(n15258), .A2(n16381), .ZN(n15261) );
  AND2_X1 U12075 ( .A1(n13070), .A2(n9756), .ZN(n15259) );
  NAND2_X1 U12076 ( .A1(n13070), .A2(n9698), .ZN(n15256) );
  AND2_X1 U12077 ( .A1(n13070), .A2(n10039), .ZN(n15257) );
  NAND2_X1 U12078 ( .A1(n13070), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13069) );
  NOR2_X1 U12079 ( .A1(n13068), .A2(n16430), .ZN(n13070) );
  NAND2_X1 U12080 ( .A1(n13063), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13068) );
  NAND3_X1 U12081 ( .A1(n10038), .A2(n10036), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13067) );
  NOR2_X1 U12082 ( .A1(n16454), .A2(n10037), .ZN(n10036) );
  NOR2_X1 U12083 ( .A1(n13064), .A2(n13807), .ZN(n13066) );
  NOR2_X1 U12084 ( .A1(n10866), .A2(n10119), .ZN(n9805) );
  NAND2_X1 U12085 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13064) );
  INV_X1 U12086 ( .A(n10404), .ZN(n10414) );
  OR3_X1 U12087 ( .A1(n14551), .A2(n10536), .A3(n14584), .ZN(n15546) );
  INV_X1 U12088 ( .A(n12853), .ZN(n9844) );
  AND2_X1 U12089 ( .A1(n15719), .A2(n15720), .ZN(n15705) );
  XNOR2_X1 U12090 ( .A(n12852), .B(n12853), .ZN(n15570) );
  NOR2_X1 U12091 ( .A1(n11318), .A2(n9930), .ZN(n9931) );
  OR2_X1 U12092 ( .A1(n15769), .A2(n11238), .ZN(n15743) );
  OR2_X1 U12093 ( .A1(n15323), .A2(n15324), .ZN(n15483) );
  NAND2_X1 U12094 ( .A1(n10015), .A2(n10017), .ZN(n10014) );
  INV_X1 U12095 ( .A(n15322), .ZN(n10017) );
  INV_X1 U12096 ( .A(n10925), .ZN(n10015) );
  AND2_X1 U12097 ( .A1(n9935), .A2(n9787), .ZN(n9934) );
  INV_X1 U12098 ( .A(n10171), .ZN(n10170) );
  NAND2_X1 U12099 ( .A1(n11237), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15769) );
  NOR3_X1 U12100 ( .A1(n15448), .A2(n10925), .A3(n10018), .ZN(n15429) );
  NOR2_X1 U12101 ( .A1(n15652), .A2(n10171), .ZN(n11205) );
  AND2_X1 U12102 ( .A1(n15792), .A2(n11197), .ZN(n11237) );
  NOR2_X1 U12103 ( .A1(n15448), .A2(n10925), .ZN(n15427) );
  AND2_X1 U12104 ( .A1(n10772), .A2(n15802), .ZN(n15638) );
  NOR2_X1 U12105 ( .A1(n15817), .A2(n10959), .ZN(n15803) );
  AND2_X1 U12106 ( .A1(n11145), .A2(n11144), .ZN(n15531) );
  NAND2_X1 U12107 ( .A1(n13987), .A2(n10090), .ZN(n15532) );
  OR2_X1 U12108 ( .A1(n19165), .A2(n10764), .ZN(n15648) );
  NAND2_X1 U12109 ( .A1(n10093), .A2(n15844), .ZN(n10092) );
  AND2_X1 U12110 ( .A1(n13836), .A2(n10907), .ZN(n14004) );
  AND3_X1 U12111 ( .A1(n11110), .A2(n11109), .A3(n11108), .ZN(n13708) );
  CLKBUF_X1 U12112 ( .A(n13088), .Z(n13637) );
  NAND2_X1 U12113 ( .A1(n10697), .A2(n10139), .ZN(n15869) );
  INV_X1 U12114 ( .A(n15877), .ZN(n16478) );
  NAND2_X1 U12115 ( .A1(n10005), .A2(n10010), .ZN(n13554) );
  AOI21_X1 U12116 ( .B1(n14232), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10165), .ZN(n10164) );
  INV_X1 U12117 ( .A(n14233), .ZN(n10165) );
  NOR2_X1 U12118 ( .A1(n13619), .A2(n13620), .ZN(n13544) );
  AND2_X1 U12119 ( .A1(n19260), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15673) );
  NOR2_X1 U12120 ( .A1(n14218), .A2(n14219), .ZN(n16491) );
  NAND2_X1 U12121 ( .A1(n13846), .A2(n11006), .ZN(n14221) );
  NAND2_X1 U12122 ( .A1(n13531), .A2(n10003), .ZN(n10002) );
  INV_X1 U12123 ( .A(n10003), .ZN(n10001) );
  NAND2_X1 U12124 ( .A1(n11182), .A2(n11181), .ZN(n14161) );
  NAND2_X1 U12125 ( .A1(n16441), .A2(n16442), .ZN(n9915) );
  NAND2_X1 U12126 ( .A1(n10004), .A2(n10876), .ZN(n13449) );
  INV_X1 U12127 ( .A(n13443), .ZN(n10004) );
  INV_X1 U12128 ( .A(n15814), .ZN(n13877) );
  OR2_X1 U12129 ( .A1(n14579), .A2(n19115), .ZN(n10970) );
  OR2_X1 U12130 ( .A1(n10498), .A2(n10497), .ZN(n13242) );
  NAND2_X1 U12131 ( .A1(n13267), .A2(n19854), .ZN(n13391) );
  INV_X1 U12132 ( .A(n10340), .ZN(n11149) );
  NAND2_X1 U12133 ( .A1(n21164), .A2(n13316), .ZN(n13398) );
  AND2_X1 U12134 ( .A1(n13315), .A2(n13318), .ZN(n13316) );
  INV_X1 U12135 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16035) );
  INV_X1 U12136 ( .A(n19454), .ZN(n19461) );
  INV_X1 U12137 ( .A(n10432), .ZN(n9838) );
  INV_X1 U12138 ( .A(n10431), .ZN(n9839) );
  INV_X1 U12139 ( .A(n10581), .ZN(n19532) );
  INV_X1 U12140 ( .A(n10596), .ZN(n19659) );
  AND2_X1 U12141 ( .A1(n20103), .A2(n20130), .ZN(n19656) );
  INV_X1 U12142 ( .A(n19789), .ZN(n19783) );
  AND2_X1 U12143 ( .A1(n20111), .A2(n20121), .ZN(n19920) );
  INV_X1 U12144 ( .A(n19492), .ZN(n19494) );
  NOR2_X2 U12145 ( .A1(n19451), .A2(n19452), .ZN(n19493) );
  NOR2_X2 U12146 ( .A1(n19453), .A2(n19452), .ZN(n19492) );
  INV_X1 U12147 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19884) );
  OR2_X1 U12148 ( .A1(n13077), .A2(n19884), .ZN(n13508) );
  NOR3_X1 U12149 ( .A1(n16731), .A2(n16730), .A3(n18885), .ZN(n18855) );
  OAI21_X1 U12150 ( .B1(n16876), .B2(n9962), .A(n9976), .ZN(n9964) );
  INV_X1 U12151 ( .A(n9963), .ZN(n9962) );
  OR2_X1 U12152 ( .A1(n16876), .A2(n17822), .ZN(n9965) );
  NAND2_X1 U12153 ( .A1(n16734), .A2(n16737), .ZN(n17118) );
  AND2_X1 U12154 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n9983), .ZN(
        n12534) );
  NOR2_X1 U12155 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9983) );
  NOR3_X1 U12156 ( .A1(n16038), .A2(n17600), .A3(n16733), .ZN(n16039) );
  NOR2_X1 U12157 ( .A1(n17638), .A2(n17599), .ZN(n17618) );
  NOR2_X1 U12158 ( .A1(n18924), .A2(n16710), .ZN(n17639) );
  NAND2_X1 U12159 ( .A1(n17739), .A2(n9703), .ZN(n12810) );
  NOR2_X1 U12160 ( .A1(n17712), .A2(n9967), .ZN(n9966) );
  INV_X1 U12161 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U12162 ( .A1(n17739), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17711) );
  NOR2_X1 U12163 ( .A1(n17757), .A2(n17758), .ZN(n17739) );
  NAND2_X1 U12164 ( .A1(n17777), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17757) );
  NAND2_X1 U12165 ( .A1(n17818), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17795) );
  NOR2_X1 U12166 ( .A1(n17829), .A2(n17830), .ZN(n17818) );
  AND3_X1 U12167 ( .A1(n9981), .A2(n18013), .A3(n9979), .ZN(n17851) );
  AND2_X1 U12168 ( .A1(n9726), .A2(n9980), .ZN(n9979) );
  INV_X1 U12169 ( .A(n17868), .ZN(n9980) );
  OR2_X1 U12170 ( .A1(n17890), .A2(n12657), .ZN(n18142) );
  AOI21_X1 U12171 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17780), .A(
        n18798), .ZN(n17910) );
  AND2_X1 U12172 ( .A1(n9981), .A2(n18013), .ZN(n17925) );
  INV_X1 U12173 ( .A(n17979), .ZN(n17938) );
  NOR2_X1 U12174 ( .A1(n18021), .A2(n18020), .ZN(n18013) );
  INV_X1 U12175 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17097) );
  AND2_X1 U12176 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18047) );
  OR2_X1 U12177 ( .A1(n12674), .A2(n12673), .ZN(n9864) );
  NOR2_X1 U12178 ( .A1(n18087), .A2(n16578), .ZN(n16558) );
  INV_X1 U12179 ( .A(n17726), .ZN(n9865) );
  NAND2_X1 U12180 ( .A1(n9988), .A2(n9994), .ZN(n9992) );
  AND2_X1 U12181 ( .A1(n17955), .A2(n18083), .ZN(n9993) );
  NAND2_X1 U12182 ( .A1(n17824), .A2(n12668), .ZN(n17766) );
  AOI21_X1 U12183 ( .B1(n17864), .B2(n17764), .A(n12666), .ZN(n12667) );
  OR3_X2 U12184 ( .A1(n17811), .A2(n18151), .A3(n17790), .ZN(n17772) );
  NAND2_X1 U12185 ( .A1(n17984), .A2(n12842), .ZN(n17903) );
  NAND2_X1 U12186 ( .A1(n17903), .A2(n17896), .ZN(n17890) );
  INV_X1 U12187 ( .A(n12658), .ZN(n17954) );
  XNOR2_X1 U12188 ( .A(n12830), .B(n9938), .ZN(n18034) );
  INV_X1 U12189 ( .A(n12831), .ZN(n9938) );
  NAND2_X1 U12190 ( .A1(n18058), .A2(n12828), .ZN(n18045) );
  NAND2_X1 U12191 ( .A1(n18045), .A2(n18046), .ZN(n18044) );
  XNOR2_X1 U12192 ( .A(n12825), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18060) );
  XNOR2_X1 U12193 ( .A(n12635), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18057) );
  AOI211_X1 U12194 ( .C1(n12692), .C2(n12691), .A(n12801), .B(n12798), .ZN(
        n18853) );
  NOR2_X1 U12195 ( .A1(n12633), .A2(n12632), .ZN(n12815) );
  NAND2_X1 U12196 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n12678), .ZN(
        n18888) );
  NOR2_X1 U12197 ( .A1(n19088), .A2(n14074), .ZN(n18881) );
  NAND2_X1 U12198 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18875) );
  NOR2_X2 U12199 ( .A1(n18865), .A2(n18863), .ZN(n18885) );
  NOR2_X1 U12200 ( .A1(n12735), .A2(n12734), .ZN(n18427) );
  NOR2_X1 U12201 ( .A1(n12765), .A2(n12764), .ZN(n18432) );
  NOR2_X1 U12202 ( .A1(n12745), .A2(n12744), .ZN(n18436) );
  NOR2_X1 U12203 ( .A1(n12725), .A2(n12724), .ZN(n18448) );
  OAI21_X1 U12204 ( .B1(n15947), .B2(n17599), .A(n15946), .ZN(n18900) );
  NOR2_X1 U12205 ( .A1(n18929), .A2(n19086), .ZN(n19069) );
  INV_X1 U12206 ( .A(n19453), .ZN(n19451) );
  INV_X1 U12207 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16057) );
  OR2_X1 U12208 ( .A1(n13903), .A2(n13902), .ZN(n16102) );
  INV_X1 U12209 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14792) );
  AND2_X1 U12210 ( .A1(n20198), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20215) );
  NAND2_X1 U12211 ( .A1(n20949), .A2(n13905), .ZN(n20220) );
  INV_X1 U12212 ( .A(n20257), .ZN(n20243) );
  INV_X1 U12213 ( .A(n20215), .ZN(n20245) );
  INV_X1 U12214 ( .A(n20220), .ZN(n20248) );
  INV_X1 U12215 ( .A(n14251), .ZN(n14293) );
  INV_X1 U12216 ( .A(n14253), .ZN(n14851) );
  INV_X1 U12217 ( .A(n16122), .ZN(n14885) );
  NAND2_X2 U12218 ( .A1(n12466), .A2(n13373), .ZN(n16115) );
  OR2_X1 U12219 ( .A1(n13370), .A2(n12465), .ZN(n12466) );
  INV_X1 U12220 ( .A(n14902), .ZN(n14898) );
  NAND2_X1 U12221 ( .A1(n14903), .A2(n13511), .ZN(n14902) );
  AND2_X1 U12222 ( .A1(n13330), .A2(n13329), .ZN(n20274) );
  OAI21_X1 U12223 ( .B1(n14629), .B2(n9741), .A(n14630), .ZN(n14907) );
  NAND2_X1 U12224 ( .A1(n9876), .A2(n11977), .ZN(n14837) );
  INV_X1 U12225 ( .A(n14023), .ZN(n9876) );
  INV_X1 U12226 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15038) );
  INV_X1 U12227 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20235) );
  CLKBUF_X1 U12228 ( .A(n13755), .Z(n13756) );
  AND2_X2 U12229 ( .A1(n20810), .A2(n12262), .ZN(n20344) );
  OAI211_X1 U12230 ( .C1(n9895), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n9892), .B(n9890), .ZN(n15085) );
  NAND2_X1 U12231 ( .A1(n9895), .A2(n9891), .ZN(n9890) );
  NAND2_X1 U12232 ( .A1(n9909), .A2(n9911), .ZN(n14029) );
  NAND2_X1 U12233 ( .A1(n16164), .A2(n12382), .ZN(n16161) );
  OR2_X1 U12234 ( .A1(n20379), .A2(n15169), .ZN(n15175) );
  INV_X1 U12235 ( .A(n20352), .ZN(n20372) );
  INV_X1 U12236 ( .A(n16278), .ZN(n20375) );
  INV_X1 U12237 ( .A(n20802), .ZN(n20810) );
  INV_X1 U12238 ( .A(n12330), .ZN(n13915) );
  INV_X1 U12239 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20727) );
  INV_X1 U12240 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20386) );
  OR2_X1 U12241 ( .A1(n13687), .A2(n13686), .ZN(n20385) );
  INV_X1 U12243 ( .A(n20936), .ZN(n15199) );
  NOR2_X1 U12244 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20937) );
  NOR2_X2 U12245 ( .A1(n20485), .A2(n20764), .ZN(n20501) );
  OAI21_X1 U12246 ( .B1(n20528), .B2(n20512), .A(n20769), .ZN(n20530) );
  NOR2_X2 U12247 ( .A1(n20587), .A2(n20653), .ZN(n20581) );
  OAI211_X1 U12248 ( .C1(n20642), .C2(n20689), .A(n20688), .B(n20626), .ZN(
        n20644) );
  AND2_X1 U12249 ( .A1(n20680), .A2(n20654), .ZN(n20720) );
  NOR2_X1 U12250 ( .A1(n20807), .A2(n20616), .ZN(n20758) );
  INV_X1 U12251 ( .A(n20763), .ZN(n15240) );
  OAI211_X1 U12252 ( .C1(n20771), .C2(n20793), .A(n20770), .B(n20769), .ZN(
        n20795) );
  INV_X1 U12253 ( .A(n20447), .ZN(n20823) );
  INV_X1 U12254 ( .A(n20451), .ZN(n20829) );
  INV_X1 U12255 ( .A(n20455), .ZN(n20835) );
  INV_X1 U12256 ( .A(n20863), .ZN(n20843) );
  INV_X1 U12257 ( .A(n20846), .ZN(n20859) );
  INV_X1 U12258 ( .A(n20468), .ZN(n20857) );
  NOR2_X1 U12259 ( .A1(n20689), .A2(n14596), .ZN(n20936) );
  NAND2_X1 U12260 ( .A1(n10201), .A2(n10082), .ZN(n10081) );
  INV_X1 U12261 ( .A(n15272), .ZN(n10082) );
  AOI21_X1 U12262 ( .B1(n15279), .B2(n15552), .A(n19289), .ZN(n15280) );
  INV_X1 U12263 ( .A(n16326), .ZN(n10031) );
  INV_X1 U12264 ( .A(n10032), .ZN(n16325) );
  NAND2_X1 U12265 ( .A1(n11303), .A2(n11304), .ZN(n15317) );
  NOR2_X1 U12266 ( .A1(n15988), .A2(n19288), .ZN(n15333) );
  INV_X1 U12267 ( .A(n10030), .ZN(n15332) );
  AND2_X1 U12268 ( .A1(n13090), .A2(n13081), .ZN(n19317) );
  OR2_X1 U12269 ( .A1(n13092), .A2(n13091), .ZN(n19320) );
  NAND2_X1 U12270 ( .A1(n13836), .A2(n9742), .ZN(n14184) );
  OR2_X1 U12271 ( .A1(n11091), .A2(n11090), .ZN(n13644) );
  CLKBUF_X1 U12272 ( .A(n13972), .Z(n13643) );
  OR2_X1 U12273 ( .A1(n11027), .A2(n11026), .ZN(n13623) );
  CLKBUF_X1 U12274 ( .A(n13399), .Z(n16512) );
  XNOR2_X1 U12275 ( .A(n10083), .B(n14580), .ZN(n19332) );
  NAND2_X1 U12276 ( .A1(n14576), .A2(n14575), .ZN(n10083) );
  XNOR2_X1 U12277 ( .A(n14576), .B(n14575), .ZN(n15692) );
  XNOR2_X1 U12278 ( .A(n9798), .B(n14514), .ZN(n14526) );
  OAI21_X1 U12279 ( .B1(n15397), .B2(n9797), .A(n9795), .ZN(n9798) );
  NAND2_X1 U12280 ( .A1(n9821), .A2(n14486), .ZN(n9820) );
  NAND2_X1 U12281 ( .A1(n9821), .A2(n9818), .ZN(n15387) );
  NOR2_X1 U12282 ( .A1(n9811), .A2(n9812), .ZN(n15402) );
  AND2_X1 U12283 ( .A1(n15520), .A2(n9709), .ZN(n15336) );
  NAND2_X1 U12284 ( .A1(n15520), .A2(n9707), .ZN(n15768) );
  OR2_X1 U12285 ( .A1(n19379), .A2(n13293), .ZN(n15522) );
  NOR2_X1 U12286 ( .A1(n13285), .A2(n13284), .ZN(n13351) );
  AND2_X1 U12287 ( .A1(n19356), .A2(n15538), .ZN(n19351) );
  NAND2_X1 U12288 ( .A1(n9800), .A2(n13435), .ZN(n13441) );
  INV_X1 U12289 ( .A(n20130), .ZN(n19713) );
  INV_X1 U12290 ( .A(n19356), .ZN(n19381) );
  NAND2_X1 U12291 ( .A1(n13290), .A2(n16538), .ZN(n19379) );
  INV_X1 U12292 ( .A(n15538), .ZN(n19380) );
  NOR2_X1 U12293 ( .A1(n19388), .A2(n20146), .ZN(n19387) );
  BUF_X1 U12295 ( .A(n19387), .Z(n19416) );
  OR2_X1 U12296 ( .A1(n15838), .A2(n9711), .ZN(n15664) );
  INV_X1 U12297 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16430) );
  NAND2_X1 U12298 ( .A1(n13124), .A2(n11335), .ZN(n16453) );
  INV_X1 U12299 ( .A(n16453), .ZN(n19421) );
  INV_X1 U12300 ( .A(n19424), .ZN(n16450) );
  INV_X1 U12301 ( .A(n19428), .ZN(n15688) );
  AOI21_X1 U12302 ( .B1(n14582), .B2(n12849), .A(n15542), .ZN(n11333) );
  NAND2_X1 U12303 ( .A1(n11325), .A2(n16519), .ZN(n11326) );
  INV_X1 U12304 ( .A(n11343), .ZN(n11325) );
  INV_X1 U12305 ( .A(n11311), .ZN(n15577) );
  OAI21_X1 U12306 ( .B1(n11285), .B2(n15617), .A(n10144), .ZN(n15606) );
  INV_X1 U12307 ( .A(n10145), .ZN(n10144) );
  AND2_X1 U12308 ( .A1(n11285), .A2(n11284), .ZN(n15619) );
  OAI21_X1 U12309 ( .B1(n15647), .B2(n10074), .A(n10071), .ZN(n10789) );
  AOI21_X1 U12310 ( .B1(n10075), .B2(n10073), .A(n10072), .ZN(n10071) );
  NAND2_X1 U12311 ( .A1(n9925), .A2(n9751), .ZN(n15780) );
  NAND2_X1 U12312 ( .A1(n10076), .A2(n10080), .ZN(n9925) );
  NAND2_X1 U12313 ( .A1(n10076), .A2(n10075), .ZN(n15779) );
  NAND2_X1 U12314 ( .A1(n10057), .A2(n10061), .ZN(n10214) );
  NAND2_X1 U12315 ( .A1(n15835), .A2(n10063), .ZN(n10057) );
  NAND2_X1 U12316 ( .A1(n15835), .A2(n15834), .ZN(n16372) );
  NAND2_X1 U12317 ( .A1(n10067), .A2(n11267), .ZN(n16393) );
  OR2_X1 U12318 ( .A1(n10070), .A2(n10066), .ZN(n15858) );
  INV_X1 U12319 ( .A(n10136), .ZN(n10066) );
  OR2_X1 U12320 ( .A1(n10957), .A2(n16523), .ZN(n14219) );
  INV_X1 U12321 ( .A(n16524), .ZN(n19438) );
  OAI21_X1 U12322 ( .B1(n10548), .B2(n9924), .A(n9922), .ZN(n13871) );
  AND2_X1 U12323 ( .A1(n9771), .A2(n13111), .ZN(n13784) );
  NAND2_X1 U12324 ( .A1(n10548), .A2(n13863), .ZN(n13802) );
  NAND2_X1 U12325 ( .A1(n11201), .A2(n13583), .ZN(n15814) );
  OAI21_X2 U12326 ( .B1(n10407), .B2(n10406), .A(n10412), .ZN(n19321) );
  INV_X1 U12327 ( .A(n19436), .ZN(n16526) );
  INV_X1 U12328 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20135) );
  INV_X1 U12329 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20116) );
  AOI221_X1 U12330 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16535), .C1(n20140), .C2(
        n16535), .A(n19964), .ZN(n20133) );
  INV_X1 U12331 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16037) );
  INV_X1 U12332 ( .A(n20121), .ZN(n20099) );
  AND2_X1 U12333 ( .A1(n19656), .A2(n19822), .ZN(n19583) );
  NAND2_X1 U12334 ( .A1(n19693), .A2(n19822), .ZN(n19607) );
  OAI21_X1 U12335 ( .B1(n19602), .B2(n19601), .A(n19600), .ZN(n19620) );
  INV_X1 U12336 ( .A(n19638), .ZN(n19650) );
  AND2_X1 U12337 ( .A1(n19812), .A2(n19625), .ZN(n19719) );
  INV_X1 U12338 ( .A(n19743), .ZN(n19733) );
  NOR2_X2 U12339 ( .A1(n19757), .A2(n19756), .ZN(n19807) );
  INV_X1 U12340 ( .A(n19835), .ZN(n19844) );
  OAI21_X1 U12341 ( .B1(n19860), .B2(n19859), .A(n19858), .ZN(n19881) );
  INV_X1 U12342 ( .A(n19852), .ZN(n19880) );
  OAI21_X1 U12343 ( .B1(n19930), .B2(n19929), .A(n19928), .ZN(n19954) );
  INV_X1 U12344 ( .A(n19898), .ZN(n19974) );
  INV_X1 U12345 ( .A(n19906), .ZN(n19992) );
  INV_X1 U12346 ( .A(n20026), .ZN(n20005) );
  OAI22_X1 U12347 ( .A1(n19484), .A2(n19496), .B1(n19483), .B2(n19494), .ZN(
        n20004) );
  INV_X1 U12348 ( .A(n19948), .ZN(n20006) );
  INV_X1 U12349 ( .A(n19914), .ZN(n20013) );
  INV_X1 U12350 ( .A(n20001), .ZN(n20022) );
  NAND2_X1 U12351 ( .A1(n13488), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16544) );
  INV_X1 U12352 ( .A(n13508), .ZN(n16538) );
  INV_X1 U12353 ( .A(n19077), .ZN(n19088) );
  INV_X1 U12354 ( .A(n17639), .ZN(n17638) );
  INV_X1 U12355 ( .A(n9978), .ZN(n16772) );
  AND2_X1 U12356 ( .A1(n9978), .A2(n9977), .ZN(n16771) );
  OR2_X1 U12357 ( .A1(n16784), .A2(n9975), .ZN(n9978) );
  AND2_X1 U12358 ( .A1(n9965), .A2(n9976), .ZN(n16865) );
  NAND2_X1 U12359 ( .A1(n16876), .A2(n9976), .ZN(n9961) );
  NOR2_X1 U12360 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16956), .ZN(n16944) );
  INV_X1 U12361 ( .A(n17118), .ZN(n17106) );
  INV_X1 U12362 ( .A(n17130), .ZN(n17115) );
  NAND4_X1 U12363 ( .A1(n9655), .A2(n19067), .A3(n18933), .A4(n18922), .ZN(
        n17130) );
  NOR2_X1 U12364 ( .A1(n16910), .A2(n17276), .ZN(n17264) );
  NOR2_X1 U12365 ( .A1(n17418), .A2(n17417), .ZN(n17416) );
  INV_X1 U12366 ( .A(n17453), .ZN(n17449) );
  NOR2_X1 U12367 ( .A1(n17666), .A2(n17462), .ZN(n17458) );
  NOR2_X1 U12368 ( .A1(n17662), .A2(n17471), .ZN(n17467) );
  INV_X1 U12369 ( .A(n17476), .ZN(n17472) );
  NAND2_X1 U12370 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17472), .ZN(n17471) );
  NOR4_X1 U12371 ( .A1(n17517), .A2(n17654), .A3(n17652), .A4(n17443), .ZN(
        n17482) );
  NOR2_X1 U12372 ( .A1(n17648), .A2(n17505), .ZN(n17500) );
  NOR2_X1 U12373 ( .A1(n17707), .A2(n17525), .ZN(n17518) );
  NAND2_X1 U12374 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17518), .ZN(n17517) );
  NOR2_X1 U12375 ( .A1(n17523), .A2(n17522), .ZN(n17567) );
  NOR2_X1 U12376 ( .A1(n12601), .A2(n12600), .ZN(n17581) );
  INV_X1 U12377 ( .A(n17598), .ZN(n17585) );
  INV_X1 U12378 ( .A(n17595), .ZN(n17590) );
  AND2_X1 U12379 ( .A1(n17564), .A2(n17591), .ZN(n17598) );
  INV_X1 U12380 ( .A(n17563), .ZN(n17591) );
  NOR2_X1 U12381 ( .A1(n18893), .A2(n17563), .ZN(n17594) );
  CLKBUF_X1 U12382 ( .A(n17615), .Z(n17634) );
  CLKBUF_X1 U12383 ( .A(n17703), .Z(n17695) );
  NOR2_X1 U12384 ( .A1(n19074), .A2(n17695), .ZN(n17696) );
  OAI211_X1 U12385 ( .C1(n19074), .C2(n19075), .A(n17640), .B(n17639), .ZN(
        n17703) );
  NOR2_X1 U12387 ( .A1(n17795), .A2(n17796), .ZN(n17777) );
  NAND2_X1 U12388 ( .A1(n17876), .A2(n18269), .ZN(n17894) );
  NAND2_X1 U12389 ( .A1(n12654), .A2(n12653), .ZN(n17960) );
  NOR2_X2 U12390 ( .A1(n17565), .A2(n18079), .ZN(n17973) );
  NAND2_X1 U12391 ( .A1(n18013), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17994) );
  INV_X1 U12392 ( .A(n18076), .ZN(n18022) );
  NAND2_X1 U12393 ( .A1(n18047), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18021) );
  OAI21_X1 U12394 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19068), .A(n16713), 
        .ZN(n18076) );
  NAND2_X1 U12395 ( .A1(n9996), .A2(n9995), .ZN(n17744) );
  INV_X1 U12396 ( .A(n9994), .ZN(n17743) );
  AND2_X1 U12397 ( .A1(n17753), .A2(n9763), .ZN(n9995) );
  NOR2_X1 U12398 ( .A1(n18104), .A2(n15973), .ZN(n18152) );
  INV_X1 U12399 ( .A(n18105), .ZN(n18135) );
  NAND2_X1 U12400 ( .A1(n17954), .A2(n18276), .ZN(n18311) );
  INV_X1 U12401 ( .A(n9937), .ZN(n17998) );
  AND2_X1 U12402 ( .A1(n9656), .A2(n9715), .ZN(n18031) );
  INV_X1 U12403 ( .A(n18881), .ZN(n18363) );
  INV_X1 U12404 ( .A(n18359), .ZN(n18383) );
  INV_X1 U12405 ( .A(n18382), .ZN(n18399) );
  INV_X1 U12406 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19049) );
  NAND2_X1 U12407 ( .A1(n18952), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19084) );
  INV_X1 U12408 ( .A(n13718), .ZN(n14260) );
  CLKBUF_X1 U12409 ( .A(n16692), .Z(n16698) );
  NAND2_X1 U12410 ( .A1(n9883), .A2(n9882), .ZN(P1_U2843) );
  AOI22_X1 U12411 ( .A1(n12976), .A2(n12975), .B1(n14840), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12412 ( .A1(n14251), .A2(n12977), .ZN(n9883) );
  AOI21_X1 U12413 ( .B1(n16152), .B2(n14278), .A(n12528), .ZN(n12529) );
  NOR2_X1 U12414 ( .A1(n15059), .A2(n20352), .ZN(n15065) );
  AND2_X1 U12415 ( .A1(n13542), .A2(n9702), .ZN(n13552) );
  AOI21_X1 U12416 ( .B1(n15562), .B2(n16449), .A(n15561), .ZN(n15563) );
  OAI211_X1 U12417 ( .C1(n14593), .C2(n16524), .A(n9836), .B(n10208), .ZN(
        P2_U3015) );
  NAND2_X1 U12418 ( .A1(n15700), .A2(n9959), .ZN(n9958) );
  NOR2_X1 U12419 ( .A1(n15698), .A2(n15697), .ZN(n15700) );
  NAND2_X1 U12420 ( .A1(n9997), .A2(n10104), .ZN(P2_U3018) );
  INV_X1 U12421 ( .A(n9998), .ZN(n9997) );
  NAND2_X1 U12422 ( .A1(n9858), .A2(n9766), .ZN(n15823) );
  OR2_X1 U12423 ( .A1(n16777), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9960) );
  INV_X1 U12424 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17094) );
  AOI21_X1 U12425 ( .B1(n9943), .B2(n9941), .A(n9940), .ZN(n18154) );
  AND2_X1 U12426 ( .A1(n18359), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9940) );
  INV_X1 U12427 ( .A(n9690), .ZN(n11348) );
  NAND2_X1 U12428 ( .A1(n12038), .A2(n9762), .ZN(n14764) );
  NAND2_X1 U12429 ( .A1(n14707), .A2(n14708), .ZN(n14695) );
  INV_X1 U12430 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13807) );
  NAND2_X1 U12431 ( .A1(n14629), .A2(n9741), .ZN(n14630) );
  INV_X1 U12432 ( .A(n12576), .ZN(n17150) );
  NOR2_X1 U12433 ( .A1(n12533), .A2(n12532), .ZN(n12576) );
  OR3_X1 U12434 ( .A1(n16081), .A2(n10047), .A3(n16049), .ZN(n9693) );
  AND2_X1 U12435 ( .A1(n14707), .A2(n10186), .ZN(n14657) );
  INV_X2 U12436 ( .A(n9639), .ZN(n15374) );
  NAND2_X1 U12437 ( .A1(n13489), .A2(n14333), .ZN(n14498) );
  NAND2_X1 U12438 ( .A1(n15883), .A2(n9935), .ZN(n15652) );
  AND2_X1 U12439 ( .A1(n15578), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9694) );
  INV_X1 U12440 ( .A(n13064), .ZN(n10038) );
  AND4_X1 U12441 ( .A1(n10038), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9695) );
  OR3_X1 U12442 ( .A1(n15448), .A2(n10016), .A3(n10925), .ZN(n9696) );
  AND2_X1 U12443 ( .A1(n11275), .A2(n11274), .ZN(n9697) );
  INV_X1 U12444 ( .A(n9999), .ZN(n15837) );
  AND2_X1 U12445 ( .A1(n10039), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9698) );
  AND2_X1 U12446 ( .A1(n10109), .A2(n10108), .ZN(n9699) );
  NAND2_X1 U12447 ( .A1(n14776), .A2(n14778), .ZN(n14777) );
  AND2_X1 U12448 ( .A1(n9699), .A2(n13559), .ZN(n9700) );
  AND2_X1 U12449 ( .A1(n10034), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9701) );
  AND2_X1 U12450 ( .A1(n13541), .A2(n13543), .ZN(n9702) );
  AND2_X1 U12451 ( .A1(n9966), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9703) );
  AND2_X1 U12452 ( .A1(n9764), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9704) );
  AND2_X1 U12453 ( .A1(n10095), .A2(n10093), .ZN(n9705) );
  INV_X1 U12454 ( .A(n9801), .ZN(n14057) );
  NAND2_X2 U12455 ( .A1(n10292), .A2(n10291), .ZN(n19470) );
  AND2_X1 U12456 ( .A1(n9702), .A2(n13551), .ZN(n9706) );
  XOR2_X1 U12457 ( .A(n16760), .B(n12809), .Z(n17083) );
  AND2_X1 U12458 ( .A1(n10098), .A2(n15509), .ZN(n9707) );
  AND2_X1 U12459 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9708) );
  NAND2_X1 U12460 ( .A1(n13110), .A2(n13109), .ZN(n13111) );
  AND2_X1 U12461 ( .A1(n9707), .A2(n9778), .ZN(n9709) );
  AND2_X1 U12462 ( .A1(n9708), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9710) );
  OR2_X1 U12463 ( .A1(n11195), .A2(n9785), .ZN(n9711) );
  INV_X4 U12464 ( .A(n14110), .ZN(n12550) );
  OR2_X1 U12465 ( .A1(n15291), .A2(n12856), .ZN(n9712) );
  INV_X1 U12466 ( .A(n10899), .ZN(n10400) );
  INV_X2 U12467 ( .A(n10899), .ZN(n14561) );
  INV_X1 U12468 ( .A(n9975), .ZN(n9976) );
  NAND2_X1 U12469 ( .A1(n15883), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15838) );
  AND2_X1 U12470 ( .A1(n10364), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U12471 ( .A1(n10724), .A2(n10112), .ZN(n9713) );
  AND4_X1 U12472 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n10200), .ZN(
        n9714) );
  OR2_X1 U12473 ( .A1(n18042), .A2(n18041), .ZN(n9715) );
  NAND2_X1 U12474 ( .A1(n10697), .A2(n10696), .ZN(n14229) );
  INV_X2 U12475 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12679) );
  NOR2_X1 U12476 ( .A1(n15652), .A2(n15802), .ZN(n15631) );
  NAND2_X1 U12477 ( .A1(n11615), .A2(n13013), .ZN(n11619) );
  NOR2_X1 U12478 ( .A1(n13067), .A2(n16438), .ZN(n13063) );
  OR2_X1 U12479 ( .A1(n12892), .A2(n12891), .ZN(n9716) );
  OR2_X1 U12480 ( .A1(n12394), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9717) );
  OR2_X1 U12481 ( .A1(n17725), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9718) );
  CLKBUF_X3 U12482 ( .A(n10903), .Z(n11210) );
  NOR2_X1 U12483 ( .A1(n12539), .A2(n18877), .ZN(n12573) );
  AND2_X1 U12484 ( .A1(n10052), .A2(n12903), .ZN(n9719) );
  AND2_X1 U12485 ( .A1(n10899), .A2(n10222), .ZN(n9720) );
  AND3_X1 U12486 ( .A1(n11505), .A2(n11504), .A3(n9884), .ZN(n9721) );
  NAND2_X1 U12487 ( .A1(n12038), .A2(n12037), .ZN(n14821) );
  NAND2_X1 U12488 ( .A1(n15883), .A2(n9934), .ZN(n15598) );
  OAI21_X2 U12489 ( .B1(n10303), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10302), .ZN(n10939) );
  NAND2_X1 U12490 ( .A1(n14160), .A2(n11186), .ZN(n14232) );
  AND2_X1 U12491 ( .A1(n12652), .A2(n9664), .ZN(n9722) );
  AND4_X1 U12492 ( .A1(n11565), .A2(n11566), .A3(n11563), .A4(n11564), .ZN(
        n9723) );
  INV_X1 U12493 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20125) );
  AND2_X1 U12494 ( .A1(n19566), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9724) );
  AND2_X1 U12495 ( .A1(n15837), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9725) );
  AND2_X1 U12496 ( .A1(n17914), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9726) );
  AND2_X1 U12497 ( .A1(n9719), .A2(n10051), .ZN(n9727) );
  NAND2_X1 U12498 ( .A1(n13803), .A2(n19321), .ZN(n10434) );
  INV_X1 U12499 ( .A(n10434), .ZN(n10411) );
  AND2_X1 U12500 ( .A1(n15869), .A2(n10712), .ZN(n9729) );
  NAND2_X1 U12501 ( .A1(n12406), .A2(n15046), .ZN(n14949) );
  AND2_X1 U12502 ( .A1(n10271), .A2(n10273), .ZN(n9730) );
  INV_X1 U12503 ( .A(n10164), .ZN(n15680) );
  INV_X1 U12504 ( .A(n13444), .ZN(n10876) );
  NAND2_X1 U12505 ( .A1(n14707), .A2(n10188), .ZN(n10190) );
  INV_X1 U12506 ( .A(n12396), .ZN(n15035) );
  AND2_X1 U12507 ( .A1(n12836), .A2(n9936), .ZN(n9731) );
  AND2_X1 U12508 ( .A1(n10121), .A2(n13392), .ZN(n9732) );
  AND2_X1 U12509 ( .A1(n10197), .A2(n14027), .ZN(n9733) );
  NAND2_X1 U12510 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  OR2_X1 U12511 ( .A1(n15652), .A2(n10172), .ZN(n11199) );
  AND2_X1 U12512 ( .A1(n10176), .A2(n10179), .ZN(n9734) );
  NAND2_X1 U12513 ( .A1(n11187), .A2(n9957), .ZN(n11184) );
  INV_X1 U12514 ( .A(n11316), .ZN(n10135) );
  AND2_X1 U12515 ( .A1(n12853), .A2(n11318), .ZN(n11316) );
  NAND2_X1 U12516 ( .A1(n9856), .A2(n9855), .ZN(n9735) );
  INV_X1 U12517 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12533) );
  AND2_X1 U12518 ( .A1(n15607), .A2(n10143), .ZN(n9736) );
  INV_X1 U12519 ( .A(n10140), .ZN(n10139) );
  NAND2_X1 U12520 ( .A1(n10696), .A2(n10141), .ZN(n10140) );
  INV_X1 U12521 ( .A(n14122), .ZN(n12583) );
  AND2_X1 U12522 ( .A1(n13080), .A2(n10168), .ZN(n9737) );
  NAND2_X1 U12523 ( .A1(n14765), .A2(n16047), .ZN(n14749) );
  INV_X1 U12524 ( .A(n11774), .ZN(n10178) );
  OAI211_X1 U12525 ( .C1(n12301), .C2(n20391), .A(n11725), .B(n11724), .ZN(
        n11774) );
  NAND2_X1 U12526 ( .A1(n10123), .A2(n9806), .ZN(n15391) );
  NAND2_X1 U12527 ( .A1(n13438), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9738) );
  AND2_X1 U12528 ( .A1(n10138), .A2(n10712), .ZN(n10137) );
  OR2_X1 U12529 ( .A1(n12388), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16158) );
  INV_X1 U12530 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13594) );
  INV_X1 U12531 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16454) );
  AND2_X1 U12532 ( .A1(n17824), .A2(n17809), .ZN(n17811) );
  NAND2_X1 U12533 ( .A1(n11622), .A2(n13900), .ZN(n12886) );
  NAND2_X1 U12534 ( .A1(n15520), .A2(n15509), .ZN(n11243) );
  INV_X2 U12535 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12678) );
  NOR2_X1 U12536 ( .A1(n13083), .A2(n10092), .ZN(n15348) );
  AND2_X1 U12537 ( .A1(n15265), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15252) );
  NAND2_X1 U12538 ( .A1(n14057), .A2(n14058), .ZN(n14180) );
  NAND2_X1 U12539 ( .A1(n14306), .A2(n15445), .ZN(n15437) );
  NOR2_X1 U12540 ( .A1(n15437), .A2(n14319), .ZN(n15431) );
  AND2_X1 U12541 ( .A1(n15261), .A2(n10034), .ZN(n9739) );
  NAND2_X1 U12542 ( .A1(n14190), .A2(n14189), .ZN(n14188) );
  NAND2_X1 U12543 ( .A1(n10183), .A2(n14836), .ZN(n14835) );
  NAND2_X1 U12544 ( .A1(n16146), .A2(n12403), .ZN(n9740) );
  AND2_X1 U12545 ( .A1(n12260), .A2(n12259), .ZN(n9741) );
  AND2_X1 U12546 ( .A1(n10021), .A2(n10020), .ZN(n9742) );
  AND2_X1 U12547 ( .A1(n10055), .A2(n10054), .ZN(n9743) );
  AND2_X1 U12548 ( .A1(n14687), .A2(n14674), .ZN(n14662) );
  OR2_X1 U12549 ( .A1(n10086), .A2(n13422), .ZN(n9744) );
  INV_X1 U12550 ( .A(n10536), .ZN(n14550) );
  NOR2_X1 U12551 ( .A1(n13083), .A2(n13085), .ZN(n13084) );
  NAND2_X1 U12552 ( .A1(n9659), .A2(n13884), .ZN(n13883) );
  AND2_X1 U12553 ( .A1(n10096), .A2(n13627), .ZN(n9745) );
  INV_X1 U12554 ( .A(n10699), .ZN(n10110) );
  NAND2_X1 U12555 ( .A1(n10149), .A2(n14027), .ZN(n15045) );
  AND2_X1 U12556 ( .A1(n15348), .A2(n15349), .ZN(n13987) );
  AND2_X1 U12557 ( .A1(n15035), .A2(n15088), .ZN(n9746) );
  INV_X1 U12559 ( .A(n15243), .ZN(n19257) );
  NAND2_X1 U12560 ( .A1(n14057), .A2(n10131), .ZN(n14204) );
  XNOR2_X1 U12561 ( .A(n14023), .B(n11977), .ZN(n14776) );
  NAND2_X1 U12562 ( .A1(n14737), .A2(n14724), .ZN(n14711) );
  XNOR2_X1 U12563 ( .A(n14414), .B(n14410), .ZN(n15406) );
  INV_X1 U12564 ( .A(n14933), .ZN(n15046) );
  OR2_X1 U12565 ( .A1(n16081), .A2(n10047), .ZN(n9747) );
  NOR2_X1 U12566 ( .A1(n13837), .A2(n13838), .ZN(n13836) );
  AND2_X1 U12567 ( .A1(n10700), .A2(n9699), .ZN(n9748) );
  INV_X1 U12568 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9887) );
  NOR2_X1 U12569 ( .A1(n15421), .A2(n14371), .ZN(n9749) );
  OR2_X1 U12570 ( .A1(n11295), .A2(n10742), .ZN(n9750) );
  NOR3_X1 U12571 ( .A1(n15448), .A2(n10016), .A3(n10014), .ZN(n10013) );
  NAND2_X1 U12572 ( .A1(n10780), .A2(n11280), .ZN(n9751) );
  NOR2_X1 U12573 ( .A1(n15483), .A2(n15484), .ZN(n10103) );
  INV_X1 U12574 ( .A(n13543), .ZN(n13549) );
  OR2_X1 U12575 ( .A1(n11045), .A2(n11044), .ZN(n13543) );
  INV_X1 U12576 ( .A(n10774), .ZN(n10080) );
  AND2_X1 U12577 ( .A1(n11883), .A2(n11882), .ZN(n11891) );
  NAND2_X1 U12578 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  NAND2_X1 U12579 ( .A1(n13863), .A2(n16522), .ZN(n9752) );
  AND2_X1 U12580 ( .A1(n15035), .A2(n15087), .ZN(n9753) );
  AND2_X1 U12581 ( .A1(n10085), .A2(n13785), .ZN(n9754) );
  AND2_X1 U12582 ( .A1(n9703), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9755) );
  AND2_X1 U12583 ( .A1(n9698), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9756) );
  AND2_X1 U12584 ( .A1(n9742), .A2(n10019), .ZN(n9757) );
  AND2_X1 U12585 ( .A1(n9743), .A2(n10053), .ZN(n9758) );
  NAND2_X1 U12586 ( .A1(n14552), .A2(n10756), .ZN(n9759) );
  INV_X1 U12587 ( .A(n14824), .ZN(n10049) );
  AND2_X1 U12588 ( .A1(n10194), .A2(n9741), .ZN(n9760) );
  BUF_X1 U12589 ( .A(n9671), .Z(n12192) );
  NOR2_X1 U12590 ( .A1(n13556), .A2(n13555), .ZN(n9761) );
  AND2_X1 U12591 ( .A1(n14223), .A2(n11011), .ZN(n13285) );
  INV_X1 U12592 ( .A(n10333), .ZN(n13122) );
  INV_X1 U12593 ( .A(n13500), .ZN(n9834) );
  NAND2_X1 U12594 ( .A1(n13542), .A2(n13541), .ZN(n13550) );
  NAND2_X1 U12595 ( .A1(n10095), .A2(n9745), .ZN(n13628) );
  OR2_X1 U12596 ( .A1(n13285), .A2(n10086), .ZN(n13353) );
  AND2_X1 U12597 ( .A1(n12060), .A2(n12037), .ZN(n9762) );
  NOR2_X1 U12598 ( .A1(n13088), .A2(n13636), .ZN(n13635) );
  OR2_X1 U12599 ( .A1(n17978), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9763) );
  AND2_X1 U12600 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9764) );
  AND2_X1 U12601 ( .A1(n13111), .A2(n10990), .ZN(n9765) );
  AND2_X1 U12602 ( .A1(n13455), .A2(n13456), .ZN(n13453) );
  NAND2_X1 U12603 ( .A1(n13561), .A2(n13560), .ZN(n13619) );
  OR2_X1 U12604 ( .A1(n15841), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9766) );
  NAND2_X1 U12605 ( .A1(n13985), .A2(n13986), .ZN(n9801) );
  AND2_X1 U12606 ( .A1(n10125), .A2(n10206), .ZN(n9767) );
  INV_X1 U12607 ( .A(n14453), .ZN(n10125) );
  AND2_X1 U12608 ( .A1(n9961), .A2(n9963), .ZN(n9768) );
  NAND2_X1 U12609 ( .A1(n10180), .A2(n9762), .ZN(n9769) );
  NAND2_X1 U12610 ( .A1(n16004), .A2(n13373), .ZN(n20167) );
  INV_X1 U12611 ( .A(n20167), .ZN(n20343) );
  NOR2_X1 U12612 ( .A1(n13443), .A2(n10001), .ZN(n9770) );
  AND2_X1 U12613 ( .A1(n10990), .A2(n10085), .ZN(n9771) );
  AND2_X1 U12614 ( .A1(n11289), .A2(n10115), .ZN(n9772) );
  AND2_X1 U12615 ( .A1(n9704), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9773) );
  AND2_X1 U12616 ( .A1(n9763), .A2(n9990), .ZN(n9774) );
  AND2_X1 U12617 ( .A1(n9710), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9775) );
  AND2_X1 U12618 ( .A1(n10125), .A2(n10124), .ZN(n9776) );
  INV_X1 U12619 ( .A(n14836), .ZN(n10182) );
  NAND2_X1 U12620 ( .A1(n12462), .A2(n11625), .ZN(n13012) );
  AND2_X1 U12621 ( .A1(n17739), .A2(n9966), .ZN(n9777) );
  INV_X1 U12622 ( .A(n15386), .ZN(n9819) );
  NAND2_X1 U12623 ( .A1(n11245), .A2(n11244), .ZN(n9778) );
  AND2_X1 U12624 ( .A1(n15247), .A2(n9710), .ZN(n13071) );
  AND2_X1 U12625 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13491) );
  INV_X1 U12626 ( .A(n16773), .ZN(n9977) );
  NAND3_X1 U12627 ( .A1(n9984), .A2(n9715), .A3(n18032), .ZN(n18030) );
  AND2_X1 U12628 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9779) );
  AND2_X1 U12629 ( .A1(n12119), .A2(n12118), .ZN(n9780) );
  NOR2_X1 U12630 ( .A1(n9711), .A2(n11196), .ZN(n9781) );
  INV_X1 U12631 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U12632 ( .A1(n11318), .A2(n11317), .ZN(n9782) );
  INV_X1 U12633 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10117) );
  AND4_X1 U12634 ( .A1(n12407), .A2(n15135), .A3(n15138), .A4(n15127), .ZN(
        n9783) );
  OR2_X1 U12635 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U12636 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9785) );
  AND2_X1 U12637 ( .A1(n12405), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9786) );
  AND2_X1 U12638 ( .A1(n10170), .A2(n15755), .ZN(n9787) );
  INV_X1 U12639 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9991) );
  INV_X1 U12640 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9990) );
  INV_X1 U12641 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10035) );
  INV_X1 U12642 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10108) );
  OR2_X1 U12643 ( .A1(n11318), .A2(n11317), .ZN(n9788) );
  INV_X1 U12644 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9982) );
  OR2_X2 U12645 ( .A1(n12321), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20351) );
  OAI21_X2 U12646 ( .B1(n16544), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16036), 
        .ZN(n19964) );
  OAI22_X2 U12647 ( .A1(n21120), .A2(n13763), .B1(n19484), .B2(n13764), .ZN(
        n20842) );
  NOR3_X2 U12648 ( .A1(n18927), .A2(n18679), .A3(n18540), .ZN(n18510) );
  INV_X1 U12649 ( .A(n20850), .ZN(n9789) );
  INV_X1 U12650 ( .A(n9789), .ZN(n9790) );
  INV_X1 U12651 ( .A(n20830), .ZN(n9791) );
  INV_X1 U12652 ( .A(n9791), .ZN(n9792) );
  INV_X1 U12653 ( .A(n20836), .ZN(n9793) );
  INV_X1 U12654 ( .A(n9793), .ZN(n9794) );
  NOR3_X2 U12655 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18927), .A3(
        n18630), .ZN(n18601) );
  OAI22_X2 U12656 ( .A1(n19497), .A2(n13764), .B1(n21079), .B2(n13763), .ZN(
        n20858) );
  NAND2_X1 U12657 ( .A1(n13542), .A2(n9706), .ZN(n13640) );
  NOR2_X2 U12658 ( .A1(n9801), .A2(n10129), .ZN(n14306) );
  AND2_X2 U12659 ( .A1(n9802), .A2(n14333), .ZN(n10309) );
  AND2_X2 U12660 ( .A1(n10447), .A2(n9802), .ZN(n14359) );
  NAND3_X1 U12661 ( .A1(n10122), .A2(n9732), .A3(n9926), .ZN(n9803) );
  NAND2_X1 U12662 ( .A1(n9804), .A2(n10866), .ZN(n9926) );
  NAND2_X2 U12663 ( .A1(n9805), .A2(n10396), .ZN(n10122) );
  NOR2_X2 U12664 ( .A1(n15415), .A2(n14392), .ZN(n14414) );
  NAND3_X1 U12665 ( .A1(n9815), .A2(n9813), .A3(n9776), .ZN(n9806) );
  NAND2_X2 U12666 ( .A1(n10408), .A2(n10392), .ZN(n10396) );
  NAND2_X2 U12667 ( .A1(n9807), .A2(n10383), .ZN(n10408) );
  NAND2_X1 U12668 ( .A1(n10404), .A2(n10412), .ZN(n9807) );
  AND2_X2 U12669 ( .A1(n9809), .A2(n9808), .ZN(n15396) );
  NAND2_X1 U12670 ( .A1(n9815), .A2(n9813), .ZN(n15401) );
  NAND2_X1 U12671 ( .A1(n14434), .A2(n10206), .ZN(n9810) );
  INV_X1 U12672 ( .A(n9815), .ZN(n9811) );
  NAND2_X1 U12673 ( .A1(n9813), .A2(n10124), .ZN(n9812) );
  NAND2_X1 U12674 ( .A1(n15407), .A2(n10207), .ZN(n14434) );
  NAND2_X1 U12675 ( .A1(n15407), .A2(n9814), .ZN(n9813) );
  INV_X1 U12676 ( .A(n9816), .ZN(n9815) );
  NAND2_X1 U12677 ( .A1(n9820), .A2(n9819), .ZN(n15451) );
  OAI21_X2 U12678 ( .B1(n15423), .B2(n10126), .A(n9822), .ZN(n15415) );
  XNOR2_X2 U12679 ( .A(n14369), .B(n14391), .ZN(n15423) );
  INV_X1 U12680 ( .A(n13640), .ZN(n13642) );
  NAND3_X1 U12681 ( .A1(n9828), .A2(n10830), .A3(n9826), .ZN(n10829) );
  NAND2_X1 U12682 ( .A1(n9827), .A2(n13080), .ZN(n9826) );
  NAND2_X1 U12683 ( .A1(n9830), .A2(n10828), .ZN(n9827) );
  NAND3_X1 U12684 ( .A1(n10824), .A2(n9829), .A3(n10825), .ZN(n9828) );
  INV_X1 U12685 ( .A(n9830), .ZN(n9829) );
  INV_X2 U12686 ( .A(n10960), .ZN(n10499) );
  NAND2_X2 U12687 ( .A1(n10281), .A2(n9831), .ZN(n10960) );
  NAND2_X1 U12688 ( .A1(n9832), .A2(n10275), .ZN(n9831) );
  NAND3_X1 U12689 ( .A1(n10272), .A2(n10274), .A3(n9730), .ZN(n9832) );
  NAND2_X1 U12690 ( .A1(n13502), .A2(n9833), .ZN(n10858) );
  NAND2_X1 U12691 ( .A1(n13488), .A2(n14487), .ZN(n13221) );
  NOR2_X2 U12692 ( .A1(n15897), .A2(n15891), .ZN(n15877) );
  NAND2_X2 U12693 ( .A1(n15812), .A2(n15814), .ZN(n19434) );
  NAND3_X1 U12694 ( .A1(n10580), .A2(n10579), .A3(n10997), .ZN(n10626) );
  NAND3_X1 U12695 ( .A1(n11187), .A2(n9957), .A3(n10536), .ZN(n9847) );
  NOR2_X1 U12696 ( .A1(n9853), .A2(n9849), .ZN(n9848) );
  NOR2_X1 U12697 ( .A1(n9850), .A2(n9854), .ZN(n19599) );
  INV_X1 U12698 ( .A(n9853), .ZN(n9851) );
  NAND3_X1 U12699 ( .A1(n10122), .A2(n9639), .A3(n19321), .ZN(n9853) );
  INV_X1 U12700 ( .A(n10000), .ZN(n9854) );
  NAND2_X1 U12701 ( .A1(n10596), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n9856) );
  NAND2_X1 U12702 ( .A1(n9862), .A2(n12644), .ZN(n12645) );
  NOR2_X2 U12703 ( .A1(n17977), .A2(n12658), .ZN(n17917) );
  OR2_X2 U12704 ( .A1(n12672), .A2(n17978), .ZN(n16022) );
  INV_X1 U12705 ( .A(n9867), .ZN(n17586) );
  NAND2_X1 U12706 ( .A1(n9867), .A2(n17593), .ZN(n12637) );
  NOR2_X1 U12707 ( .A1(n12824), .A2(n9867), .ZN(n12822) );
  OR2_X2 U12708 ( .A1(n17754), .A2(n18107), .ZN(n9996) );
  NAND2_X1 U12709 ( .A1(n14013), .A2(n14024), .ZN(n14023) );
  NAND2_X1 U12710 ( .A1(n14013), .A2(n9872), .ZN(n9871) );
  NAND2_X1 U12711 ( .A1(n11620), .A2(n11636), .ZN(n9881) );
  NAND2_X1 U12712 ( .A1(n9879), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11662) );
  NAND3_X1 U12713 ( .A1(n12449), .A2(n9880), .A3(n11637), .ZN(n9879) );
  NOR2_X1 U12714 ( .A1(n9881), .A2(n11626), .ZN(n9880) );
  NAND2_X1 U12715 ( .A1(n12449), .A2(n11620), .ZN(n13011) );
  NOR2_X2 U12716 ( .A1(n14828), .A2(n9769), .ZN(n14765) );
  NAND3_X1 U12717 ( .A1(n11359), .A2(n10041), .A3(
        P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n9886) );
  NAND4_X1 U12718 ( .A1(n10041), .A2(n11347), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n9885) );
  OAI21_X2 U12719 ( .B1(n11662), .B2(n11347), .A(n11639), .ZN(n9888) );
  NAND2_X1 U12720 ( .A1(n12278), .A2(n11624), .ZN(n11527) );
  INV_X1 U12721 ( .A(n11621), .ZN(n9889) );
  OAI21_X1 U12722 ( .B1(n15085), .B2(n20167), .A(n14252), .ZN(P1_U2970) );
  NAND2_X1 U12723 ( .A1(n9893), .A2(n14247), .ZN(n9892) );
  INV_X1 U12724 ( .A(n9894), .ZN(n9893) );
  NAND2_X1 U12725 ( .A1(n12494), .A2(n15087), .ZN(n9896) );
  NAND2_X1 U12726 ( .A1(n12494), .A2(n9753), .ZN(n9894) );
  NAND2_X1 U12727 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  NAND2_X1 U12728 ( .A1(n10147), .A2(n9746), .ZN(n9897) );
  NAND2_X1 U12729 ( .A1(n20618), .A2(n20865), .ZN(n9898) );
  NAND3_X1 U12730 ( .A1(n9903), .A2(n12405), .A3(n9901), .ZN(n12406) );
  NAND3_X1 U12731 ( .A1(n9903), .A2(n9786), .A3(n9901), .ZN(n9905) );
  NAND2_X1 U12732 ( .A1(n9904), .A2(n10154), .ZN(n15154) );
  NAND2_X1 U12733 ( .A1(n9906), .A2(n10157), .ZN(n9904) );
  AND2_X1 U12734 ( .A1(n10156), .A2(n14991), .ZN(n9906) );
  NAND2_X1 U12735 ( .A1(n11867), .A2(n11866), .ZN(n11890) );
  NAND2_X2 U12736 ( .A1(n11867), .A2(n9907), .ZN(n12324) );
  NAND2_X1 U12737 ( .A1(n10151), .A2(n10150), .ZN(n9910) );
  NAND4_X1 U12738 ( .A1(n10476), .A2(n9914), .A3(n9912), .A4(n10475), .ZN(
        n10514) );
  NAND4_X1 U12739 ( .A1(n10465), .A2(n10466), .A3(n10467), .A4(n10464), .ZN(
        n9913) );
  NAND2_X1 U12740 ( .A1(n9919), .A2(n9920), .ZN(n10578) );
  NAND2_X1 U12741 ( .A1(n10548), .A2(n9922), .ZN(n9919) );
  NAND3_X1 U12742 ( .A1(n10000), .A2(n10426), .A3(n10122), .ZN(n10415) );
  AND2_X2 U12743 ( .A1(n9926), .A2(n10121), .ZN(n10000) );
  AND2_X2 U12744 ( .A1(n10411), .A2(n9927), .ZN(n10590) );
  NAND2_X1 U12745 ( .A1(n15578), .A2(n9931), .ZN(n9933) );
  INV_X1 U12746 ( .A(n9933), .ZN(n15565) );
  NAND2_X1 U12747 ( .A1(n15578), .A2(n9929), .ZN(n12849) );
  INV_X1 U12748 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9930) );
  INV_X1 U12749 ( .A(n15598), .ZN(n11206) );
  NAND2_X1 U12750 ( .A1(n9937), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12840) );
  NOR2_X2 U12751 ( .A1(n12532), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12602) );
  NAND3_X1 U12752 ( .A1(n18159), .A2(n9944), .A3(n18141), .ZN(n9943) );
  AND2_X1 U12753 ( .A1(n9946), .A2(n10368), .ZN(n10369) );
  NAND2_X1 U12754 ( .A1(n10936), .A2(n9946), .ZN(n10943) );
  NAND2_X1 U12755 ( .A1(n10357), .A2(n10356), .ZN(n9946) );
  NAND2_X1 U12756 ( .A1(n9948), .A2(n14487), .ZN(n9947) );
  NAND4_X1 U12757 ( .A1(n9949), .A2(n10438), .A3(n10439), .A4(n10440), .ZN(
        n9948) );
  AND4_X1 U12758 ( .A1(n10423), .A2(n10421), .A3(n10420), .A4(n10422), .ZN(
        n9949) );
  INV_X2 U12759 ( .A(n10321), .ZN(n10837) );
  NAND2_X2 U12760 ( .A1(n10257), .A2(n10256), .ZN(n10321) );
  NAND2_X1 U12761 ( .A1(n10689), .A2(n11180), .ZN(n9957) );
  NAND2_X2 U12762 ( .A1(n9956), .A2(n10688), .ZN(n11187) );
  INV_X1 U12763 ( .A(n10689), .ZN(n9956) );
  AOI21_X2 U12764 ( .B1(n15701), .B2(n16519), .A(n9958), .ZN(n15702) );
  OR2_X2 U12765 ( .A1(n10068), .A2(n10070), .ZN(n10067) );
  NAND3_X1 U12766 ( .A1(n16770), .A2(n16769), .A3(n9960), .ZN(P3_U2641) );
  INV_X1 U12767 ( .A(n9965), .ZN(n16875) );
  INV_X1 U12768 ( .A(n9964), .ZN(n16857) );
  NOR2_X1 U12769 ( .A1(n16785), .A2(n17710), .ZN(n16784) );
  NAND2_X1 U12770 ( .A1(n16785), .A2(n9976), .ZN(n9972) );
  NAND3_X1 U12771 ( .A1(n9981), .A2(n18013), .A3(n9726), .ZN(n17867) );
  NAND2_X1 U12772 ( .A1(n18040), .A2(n18354), .ZN(n9984) );
  NAND2_X1 U12773 ( .A1(n17876), .A2(n9986), .ZN(n9985) );
  NAND2_X2 U12774 ( .A1(n17993), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17992) );
  AND2_X1 U12775 ( .A1(n9722), .A2(n17992), .ZN(n12658) );
  INV_X1 U12776 ( .A(n9992), .ZN(n16588) );
  NOR2_X1 U12777 ( .A1(n12669), .A2(n9993), .ZN(n9988) );
  INV_X1 U12778 ( .A(n13619), .ZN(n10005) );
  NAND2_X1 U12779 ( .A1(n10005), .A2(n10006), .ZN(n13088) );
  OR2_X1 U12780 ( .A1(n15699), .A2(n16527), .ZN(n10012) );
  XNOR2_X2 U12781 ( .A(n14560), .B(n14559), .ZN(n15699) );
  INV_X1 U12782 ( .A(n10013), .ZN(n15410) );
  INV_X1 U12783 ( .A(n15426), .ZN(n10018) );
  NOR2_X4 U12784 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10041) );
  AOI21_X2 U12785 ( .B1(n14999), .B2(n12401), .A(n12400), .ZN(n16124) );
  NAND3_X1 U12786 ( .A1(n10027), .A2(n11613), .A3(n13900), .ZN(n12460) );
  NAND2_X1 U12787 ( .A1(n11809), .A2(n10028), .ZN(n11865) );
  INV_X1 U12788 ( .A(n11865), .ZN(n11867) );
  NOR2_X1 U12789 ( .A1(n15019), .A2(n15017), .ZN(n10029) );
  NAND2_X2 U12790 ( .A1(n12324), .A2(n12326), .ZN(n12396) );
  NAND3_X1 U12791 ( .A1(n12371), .A2(n12324), .A3(n12383), .ZN(n12380) );
  NAND2_X1 U12792 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10037) );
  NAND3_X1 U12793 ( .A1(n10038), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U12794 ( .A1(n15247), .A2(n9775), .ZN(n13072) );
  AND2_X2 U12795 ( .A1(n13656), .A2(n10041), .ZN(n11562) );
  NAND2_X1 U12796 ( .A1(n14610), .A2(n10043), .ZN(n10042) );
  NOR2_X1 U12797 ( .A1(n13774), .A2(n9716), .ZN(n13700) );
  NAND3_X1 U12798 ( .A1(n14824), .A2(n14768), .A3(n10048), .ZN(n10047) );
  NAND2_X1 U12799 ( .A1(n10050), .A2(n16305), .ZN(n14781) );
  AND2_X1 U12800 ( .A1(n15647), .A2(n15648), .ZN(n15651) );
  AND2_X2 U12801 ( .A1(n10960), .A2(n19854), .ZN(n11032) );
  NAND2_X1 U12802 ( .A1(n13111), .A2(n10084), .ZN(n13848) );
  NAND2_X1 U12803 ( .A1(n15520), .A2(n10097), .ZN(n15323) );
  NOR3_X1 U12804 ( .A1(n15483), .A2(n10100), .A3(n15307), .ZN(n12858) );
  INV_X1 U12805 ( .A(n12859), .ZN(n10102) );
  INV_X1 U12806 ( .A(n10103), .ZN(n15482) );
  OR2_X2 U12807 ( .A1(n15564), .A2(n19449), .ZN(n10104) );
  NAND2_X1 U12808 ( .A1(n10700), .A2(n10699), .ZN(n10704) );
  AND2_X2 U12809 ( .A1(n10724), .A2(n10111), .ZN(n10770) );
  NAND2_X1 U12810 ( .A1(n11288), .A2(n9772), .ZN(n11314) );
  NAND2_X1 U12811 ( .A1(n11288), .A2(n11289), .ZN(n11298) );
  NAND2_X1 U12812 ( .A1(n10396), .A2(n10395), .ZN(n10867) );
  INV_X1 U12813 ( .A(n10395), .ZN(n10119) );
  INV_X1 U12814 ( .A(n15403), .ZN(n10124) );
  AND2_X2 U12815 ( .A1(n13803), .A2(n10426), .ZN(n10427) );
  NAND2_X1 U12816 ( .A1(n11313), .A2(n11312), .ZN(n12851) );
  AND2_X2 U12817 ( .A1(n11358), .A2(n13656), .ZN(n11559) );
  NAND2_X2 U12818 ( .A1(n10149), .A2(n9733), .ZN(n16145) );
  NAND2_X1 U12819 ( .A1(n16166), .A2(n16165), .ZN(n16164) );
  INV_X1 U12820 ( .A(n16165), .ZN(n10150) );
  NAND2_X1 U12821 ( .A1(n15035), .A2(n9784), .ZN(n10159) );
  NAND2_X1 U12822 ( .A1(n14160), .A2(n10166), .ZN(n15681) );
  NAND2_X1 U12823 ( .A1(n10162), .A2(n10160), .ZN(n15685) );
  NAND2_X1 U12824 ( .A1(n14233), .A2(n11192), .ZN(n10161) );
  NAND2_X1 U12825 ( .A1(n10167), .A2(n9737), .ZN(n10169) );
  NAND2_X2 U12826 ( .A1(n10945), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10899) );
  AND2_X2 U12827 ( .A1(n15565), .A2(n10173), .ZN(n15542) );
  INV_X1 U12828 ( .A(n11723), .ZN(n10174) );
  NAND2_X1 U12829 ( .A1(n10174), .A2(n11774), .ZN(n10175) );
  NAND2_X1 U12830 ( .A1(n10175), .A2(n10176), .ZN(n11746) );
  NAND2_X1 U12831 ( .A1(n11723), .A2(n11722), .ZN(n11773) );
  NAND2_X1 U12832 ( .A1(n10183), .A2(n10181), .ZN(n14828) );
  AND2_X2 U12834 ( .A1(n13326), .A2(n13900), .ZN(n13895) );
  INV_X1 U12835 ( .A(n10190), .ZN(n14683) );
  NAND2_X1 U12836 ( .A1(n14629), .A2(n9760), .ZN(n12448) );
  XNOR2_X1 U12837 ( .A(n14544), .B(n14543), .ZN(n14593) );
  NAND2_X1 U12838 ( .A1(n10328), .A2(n10537), .ZN(n10844) );
  XNOR2_X1 U12839 ( .A(n14530), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15068) );
  NOR2_X1 U12840 ( .A1(n10499), .A2(n19097), .ZN(n10341) );
  INV_X1 U12841 ( .A(n10387), .ZN(n10903) );
  AND2_X1 U12842 ( .A1(n15685), .A2(n15684), .ZN(n16497) );
  NAND2_X1 U12843 ( .A1(n10286), .A2(n10275), .ZN(n10292) );
  AOI22_X1 U12844 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U12845 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10265) );
  XOR2_X1 U12846 ( .A(n14536), .B(n14535), .Z(n14844) );
  AND2_X1 U12847 ( .A1(n10246), .A2(n10275), .ZN(n10247) );
  AOI22_X1 U12848 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10246) );
  INV_X1 U12849 ( .A(n12530), .ZN(n12531) );
  NAND2_X1 U12850 ( .A1(n13688), .A2(n20431), .ZN(n20764) );
  INV_X1 U12851 ( .A(n20431), .ZN(n15191) );
  OR2_X1 U12852 ( .A1(n13688), .A2(n20431), .ZN(n20653) );
  OAI21_X1 U12853 ( .B1(n14285), .B2(n15054), .A(n12529), .ZN(n12530) );
  AOI22_X1 U12854 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n14500), .ZN(n10262) );
  NAND2_X1 U12855 ( .A1(n10427), .A2(n9639), .ZN(n19963) );
  NAND2_X1 U12856 ( .A1(n12899), .A2(n13895), .ZN(n12967) );
  NAND2_X1 U12857 ( .A1(n11560), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11603) );
  AOI21_X1 U12858 ( .B1(n14253), .B2(n20344), .A(n12323), .ZN(n12414) );
  INV_X1 U12859 ( .A(n14904), .ZN(n16119) );
  AND2_X2 U12860 ( .A1(n12873), .A2(n13373), .ZN(n20270) );
  AND2_X2 U12861 ( .A1(n20167), .A2(n12317), .ZN(n20338) );
  AND2_X1 U12862 ( .A1(n11201), .A2(n20139), .ZN(n16519) );
  NOR2_X1 U12863 ( .A1(n20683), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10195) );
  AND2_X1 U12864 ( .A1(n10332), .A2(n10837), .ZN(n10196) );
  OR2_X1 U12865 ( .A1(n12396), .A2(n16272), .ZN(n10197) );
  AND2_X1 U12866 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10199) );
  AND2_X2 U12867 ( .A1(n10410), .A2(n15374), .ZN(n10588) );
  OR2_X1 U12868 ( .A1(n15273), .A2(n19302), .ZN(n10201) );
  OR2_X1 U12869 ( .A1(n11619), .A2(n13900), .ZN(n10202) );
  OR2_X1 U12870 ( .A1(n15692), .A2(n16526), .ZN(n10203) );
  NAND2_X1 U12871 ( .A1(n11831), .A2(n11830), .ZN(n13698) );
  INV_X1 U12872 ( .A(n11777), .ZN(n11899) );
  INV_X1 U12873 ( .A(n11899), .ZN(n12524) );
  INV_X1 U12874 ( .A(n18069), .ZN(n18080) );
  NOR2_X2 U12875 ( .A1(n16733), .A2(n16713), .ZN(n18069) );
  INV_X2 U12876 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20865) );
  INV_X1 U12877 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14528) );
  AND2_X1 U12878 ( .A1(n11281), .A2(n11272), .ZN(n10204) );
  INV_X1 U12879 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11318) );
  AND2_X1 U12880 ( .A1(n10287), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10205) );
  AND2_X1 U12881 ( .A1(n14431), .A2(n14449), .ZN(n10206) );
  INV_X1 U12882 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14247) );
  NOR2_X1 U12883 ( .A1(n14589), .A2(n14588), .ZN(n10208) );
  INV_X1 U12884 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U12885 ( .A1(n18024), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18023) );
  AND4_X1 U12886 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n10209) );
  INV_X1 U12887 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12653) );
  INV_X1 U12888 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13651) );
  INV_X1 U12889 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14543) );
  AND2_X1 U12890 ( .A1(n13644), .A2(n13641), .ZN(n10210) );
  INV_X1 U12891 ( .A(n15437), .ZN(n15444) );
  INV_X1 U12892 ( .A(n10997), .ZN(n11156) );
  AND4_X1 U12893 ( .A1(n10587), .A2(n10586), .A3(n10585), .A4(n10584), .ZN(
        n10211) );
  INV_X1 U12894 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20109) );
  NOR2_X1 U12895 ( .A1(n18937), .A2(n18022), .ZN(n17780) );
  AND3_X1 U12896 ( .A1(n12847), .A2(n12846), .A3(n12845), .ZN(n10212) );
  AND2_X1 U12897 ( .A1(n17437), .A2(n17564), .ZN(n17435) );
  AND4_X1 U12898 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10213) );
  INV_X1 U12899 ( .A(n11530), .ZN(n11561) );
  INV_X1 U12900 ( .A(n11559), .ZN(n11576) );
  AND2_X1 U12901 ( .A1(n11532), .A2(n11531), .ZN(n10216) );
  AND2_X1 U12902 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10217) );
  INV_X1 U12903 ( .A(n11539), .ZN(n11552) );
  AND2_X1 U12904 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10218) );
  INV_X1 U12905 ( .A(n11550), .ZN(n11731) );
  OR2_X1 U12906 ( .A1(n12198), .A2(n11601), .ZN(n10219) );
  AND2_X1 U12907 ( .A1(n13023), .A2(n9654), .ZN(n12462) );
  INV_X1 U12908 ( .A(n11634), .ZN(n13028) );
  INV_X1 U12909 ( .A(n12280), .ZN(n12298) );
  OR3_X1 U12910 ( .A1(n12298), .A2(n12297), .A3(n12453), .ZN(n12299) );
  OR2_X1 U12911 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12290), .ZN(
        n12266) );
  NAND2_X1 U12912 ( .A1(n11528), .A2(n11629), .ZN(n13021) );
  AND2_X1 U12913 ( .A1(n11633), .A2(n11649), .ZN(n11637) );
  AOI22_X1 U12914 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11456) );
  OR2_X1 U12915 ( .A1(n10899), .A2(n10345), .ZN(n10346) );
  AND2_X1 U12916 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20125), .ZN(
        n10539) );
  INV_X1 U12917 ( .A(n10570), .ZN(n10574) );
  OR2_X1 U12918 ( .A1(n11857), .A2(n11856), .ZN(n12373) );
  INV_X1 U12919 ( .A(n12206), .ZN(n11523) );
  INV_X1 U12920 ( .A(n12161), .ZN(n11522) );
  INV_X1 U12921 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11511) );
  INV_X1 U12922 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U12923 ( .A1(n15587), .A2(n11309), .ZN(n11310) );
  AND2_X1 U12924 ( .A1(n10844), .A2(n19470), .ZN(n10318) );
  INV_X1 U12925 ( .A(n12639), .ZN(n12640) );
  OR2_X1 U12926 ( .A1(n12275), .A2(n12281), .ZN(n12277) );
  AND2_X1 U12927 ( .A1(n13698), .A2(n13773), .ZN(n11841) );
  INV_X1 U12928 ( .A(n12227), .ZN(n11524) );
  NAND2_X1 U12929 ( .A1(n11522), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12184) );
  INV_X1 U12930 ( .A(n14830), .ZN(n12037) );
  INV_X1 U12931 ( .A(n13998), .ZN(n11921) );
  OR2_X1 U12932 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20386), .ZN(
        n12304) );
  INV_X1 U12933 ( .A(n12854), .ZN(n11321) );
  OR2_X1 U12934 ( .A1(n11279), .A2(n11278), .ZN(n11283) );
  AOI22_X1 U12935 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10284) );
  AND2_X1 U12936 ( .A1(n19470), .A2(n10939), .ZN(n10349) );
  AND2_X1 U12937 ( .A1(n14611), .A2(n12962), .ZN(n12882) );
  OR2_X1 U12938 ( .A1(n14596), .A2(n12461), .ZN(n12464) );
  NOR2_X1 U12939 ( .A1(n12246), .A2(n14646), .ZN(n12256) );
  OR2_X1 U12940 ( .A1(n12215), .A2(n14686), .ZN(n12227) );
  INV_X1 U12941 ( .A(n15247), .ZN(n15248) );
  INV_X1 U12942 ( .A(n14413), .ZN(n14410) );
  AND4_X1 U12943 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  NOR2_X1 U12944 ( .A1(n10852), .A2(n10334), .ZN(n10317) );
  OAI21_X1 U12945 ( .B1(n10370), .B2(n10369), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10371) );
  NAND2_X1 U12946 ( .A1(n11190), .A2(n11189), .ZN(n11194) );
  INV_X1 U12948 ( .A(n13581), .ZN(n13567) );
  NAND2_X1 U12949 ( .A1(n17955), .A2(n18212), .ZN(n12659) );
  AND2_X1 U12950 ( .A1(n18423), .A2(n12783), .ZN(n12781) );
  AND2_X1 U12951 ( .A1(n11993), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11998) );
  INV_X1 U12952 ( .A(n13775), .ZN(n12889) );
  NAND2_X1 U12953 ( .A1(n12922), .A2(n14611), .ZN(n12932) );
  OR2_X1 U12954 ( .A1(n12441), .A2(n12440), .ZN(n13891) );
  NOR2_X1 U12955 ( .A1(n11570), .A2(n10199), .ZN(n11571) );
  NAND2_X1 U12956 ( .A1(n9654), .A2(n13900), .ZN(n11643) );
  NOR2_X1 U12957 ( .A1(n13891), .A2(n13890), .ZN(n13892) );
  NAND2_X1 U12958 ( .A1(n12256), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12439) );
  OR2_X1 U12959 ( .A1(n12236), .A2(n12235), .ZN(n12246) );
  AND2_X1 U12960 ( .A1(n11521), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12139) );
  NOR2_X1 U12961 ( .A1(n12039), .A2(n16057), .ZN(n12062) );
  NOR2_X1 U12962 ( .A1(n16198), .A2(n16241), .ZN(n16206) );
  AND2_X1 U12963 ( .A1(n16286), .A2(n16287), .ZN(n12903) );
  NAND2_X1 U12964 ( .A1(n13895), .A2(n12962), .ZN(n12952) );
  NAND2_X1 U12965 ( .A1(n13372), .A2(n13371), .ZN(n15993) );
  INV_X1 U12966 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12290) );
  NOR2_X1 U12967 ( .A1(n9689), .A2(n13711), .ZN(n20800) );
  NAND2_X1 U12968 ( .A1(n10794), .A2(n10793), .ZN(n10830) );
  AND2_X1 U12969 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13393) );
  INV_X1 U12970 ( .A(n10358), .ZN(n13080) );
  INV_X1 U12971 ( .A(n11151), .ZN(n13592) );
  INV_X1 U12972 ( .A(n10582), .ZN(n19720) );
  INV_X1 U12973 ( .A(n18432), .ZN(n14072) );
  NOR2_X1 U12974 ( .A1(n16730), .A2(n18885), .ZN(n15939) );
  NOR2_X1 U12975 ( .A1(n18448), .A2(n18427), .ZN(n12806) );
  AOI211_X1 U12976 ( .C1(n12790), .C2(n12803), .A(n12789), .B(n15940), .ZN(
        n12795) );
  NAND4_X1 U12977 ( .A1(n12806), .A2(n18436), .A3(n12781), .A4(n17600), .ZN(
        n12776) );
  OR2_X1 U12978 ( .A1(n14640), .A2(n14276), .ZN(n14615) );
  AND2_X1 U12979 ( .A1(n11998), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12018) );
  INV_X1 U12980 ( .A(n20203), .ZN(n14788) );
  INV_X1 U12981 ( .A(n14538), .ZN(n13907) );
  AND3_X1 U12982 ( .A1(n12930), .A2(n12929), .A3(n12928), .ZN(n14824) );
  AND2_X1 U12983 ( .A1(n14979), .A2(n13889), .ZN(n12162) );
  AOI21_X1 U12984 ( .B1(n12362), .B2(n12052), .A(n11864), .ZN(n13814) );
  XNOR2_X1 U12985 ( .A(n13892), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14538) );
  NAND2_X1 U12986 ( .A1(n12139), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12161) );
  OR2_X1 U12987 ( .A1(n16146), .A2(n16232), .ZN(n16138) );
  OR2_X1 U12988 ( .A1(n13056), .A2(n13658), .ZN(n20369) );
  NAND2_X1 U12989 ( .A1(n11791), .A2(n11790), .ZN(n20506) );
  INV_X1 U12990 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20686) );
  NOR2_X1 U12991 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20677) );
  NOR2_X1 U12992 ( .A1(n15217), .A2(n20560), .ZN(n20688) );
  INV_X1 U12993 ( .A(n20758), .ZN(n15238) );
  NAND3_X1 U12994 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20865), .A3(n13720), 
        .ZN(n13765) );
  OR2_X2 U12995 ( .A1(n10704), .A2(n14552), .ZN(n14554) );
  AND3_X1 U12996 ( .A1(n10996), .A2(n10995), .A3(n10994), .ZN(n13783) );
  INV_X1 U12997 ( .A(n13635), .ZN(n13821) );
  INV_X1 U12998 ( .A(n15667), .ZN(n10750) );
  INV_X1 U12999 ( .A(n19420), .ZN(n16466) );
  INV_X1 U13000 ( .A(n10809), .ZN(n11200) );
  NOR2_X1 U13001 ( .A1(n10934), .A2(n10933), .ZN(n13583) );
  OR2_X1 U13002 ( .A1(n19096), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19178) );
  AND2_X1 U13003 ( .A1(n20103), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19687) );
  AND2_X1 U13004 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19812) );
  INV_X1 U13005 ( .A(n19493), .ZN(n19496) );
  INV_X1 U13006 ( .A(n10843), .ZN(n13613) );
  AOI21_X1 U13007 ( .B1(n12686), .B2(n12685), .A(n12684), .ZN(n12801) );
  OR3_X1 U13008 ( .A1(n18996), .A2(n18997), .A3(n16854), .ZN(n16845) );
  NOR2_X1 U13009 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16890), .ZN(n16872) );
  NOR2_X1 U13010 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17057), .ZN(n17041) );
  NOR2_X1 U13011 ( .A1(n17403), .A2(n17413), .ZN(n17402) );
  AOI211_X1 U13012 ( .C1(n17394), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n12772), .B(n12771), .ZN(n12773) );
  INV_X1 U13013 ( .A(n12562), .ZN(n12572) );
  INV_X1 U13014 ( .A(n18217), .ZN(n17886) );
  AND2_X1 U13015 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17914) );
  NAND2_X1 U13016 ( .A1(n16021), .A2(n12670), .ZN(n12677) );
  NAND2_X1 U13017 ( .A1(n12646), .A2(n17569), .ZN(n12623) );
  INV_X1 U13018 ( .A(n12667), .ZN(n12668) );
  NOR2_X1 U13019 ( .A1(n17964), .A2(n17960), .ZN(n17935) );
  NOR2_X2 U13020 ( .A1(n18248), .A2(n18864), .ZN(n18345) );
  OR2_X1 U13021 ( .A1(n19053), .A2(n18934), .ZN(n18414) );
  INV_X1 U13022 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18679) );
  OR2_X1 U13023 ( .A1(n18453), .A2(n18654), .ZN(n18444) );
  AND2_X1 U13024 ( .A1(n12476), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14848)
         );
  NOR2_X1 U13025 ( .A1(n14706), .A2(n14273), .ZN(n14679) );
  AND2_X1 U13026 ( .A1(n20203), .A2(n14263), .ZN(n14718) );
  NOR2_X1 U13027 ( .A1(n14772), .A2(n16226), .ZN(n16044) );
  NOR2_X1 U13028 ( .A1(n16100), .A2(n14269), .ZN(n16089) );
  NOR2_X2 U13029 ( .A1(n13908), .A2(n14538), .ZN(n20210) );
  INV_X1 U13030 ( .A(n16102), .ZN(n20250) );
  INV_X1 U13031 ( .A(n13403), .ZN(n20314) );
  NAND2_X1 U13032 ( .A1(n11884), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11894) );
  INV_X1 U13033 ( .A(n20349), .ZN(n16152) );
  OR2_X1 U13034 ( .A1(n13056), .A2(n13055), .ZN(n20352) );
  INV_X1 U13035 ( .A(n16239), .ZN(n16198) );
  OR2_X1 U13036 ( .A1(n15134), .A2(n13046), .ZN(n16239) );
  NAND2_X1 U13037 ( .A1(n13010), .A2(n13373), .ZN(n13056) );
  OR2_X1 U13038 ( .A1(n15183), .A2(n15170), .ZN(n20379) );
  NOR2_X1 U13039 ( .A1(n13056), .A2(n13676), .ZN(n15183) );
  OAI22_X1 U13040 ( .A1(n13927), .A2(n13926), .B1(n20508), .B2(n20621), .ZN(
        n20402) );
  NOR2_X2 U13041 ( .A1(n20485), .A2(n20616), .ZN(n20427) );
  OAI21_X1 U13042 ( .B1(n20439), .B2(n20438), .A(n20437), .ZN(n20471) );
  INV_X1 U13043 ( .A(n20484), .ZN(n20502) );
  NOR2_X2 U13044 ( .A1(n20485), .A2(n20586), .ZN(n20529) );
  OR2_X1 U13045 ( .A1(n13688), .A2(n15191), .ZN(n20616) );
  OAI211_X1 U13046 ( .C1(n20580), .C2(n20689), .A(n20769), .B(n20565), .ZN(
        n20582) );
  NOR2_X2 U13047 ( .A1(n20587), .A2(n20764), .ZN(n20612) );
  INV_X1 U13048 ( .A(n20693), .ZN(n20722) );
  AND2_X1 U13049 ( .A1(n20680), .A2(n20679), .ZN(n20751) );
  OAI211_X1 U13050 ( .C1(n20757), .C2(n20689), .A(n20769), .B(n15221), .ZN(
        n20760) );
  AND2_X1 U13051 ( .A1(n13651), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16015) );
  INV_X1 U13052 ( .A(n20911), .ZN(n20923) );
  INV_X1 U13053 ( .A(n20909), .ZN(n20924) );
  AND2_X1 U13054 ( .A1(n13579), .A2(n16538), .ZN(n13119) );
  NAND2_X1 U13055 ( .A1(n15275), .A2(n15274), .ZN(n15276) );
  OR2_X1 U13056 ( .A1(n19098), .A2(n13079), .ZN(n19262) );
  AND2_X1 U13057 ( .A1(n19098), .A2(n13612), .ZN(n19305) );
  NAND2_X1 U13058 ( .A1(n13272), .A2(n16538), .ZN(n13273) );
  NAND2_X1 U13059 ( .A1(n21164), .A2(n13282), .ZN(n20121) );
  INV_X1 U13060 ( .A(n15522), .ZN(n16364) );
  OAI21_X1 U13061 ( .B1(n12990), .B2(n12989), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13201) );
  INV_X1 U13062 ( .A(n13219), .ZN(n13168) );
  INV_X1 U13063 ( .A(n13171), .ZN(n13204) );
  INV_X1 U13064 ( .A(n19423), .ZN(n16449) );
  AOI21_X1 U13065 ( .B1(n16338), .B2(n19440), .A(n12864), .ZN(n12865) );
  AND2_X1 U13066 ( .A1(n11201), .A2(n10930), .ZN(n19440) );
  AND2_X1 U13067 ( .A1(n11201), .A2(n11153), .ZN(n19436) );
  AND2_X1 U13068 ( .A1(n13398), .A2(n13321), .ZN(n20111) );
  OAI21_X1 U13069 ( .B1(n19464), .B2(n19463), .A(n19462), .ZN(n19502) );
  AND2_X1 U13070 ( .A1(n19755), .A2(n19693), .ZN(n19554) );
  INV_X1 U13071 ( .A(n19572), .ZN(n19588) );
  INV_X1 U13072 ( .A(n19607), .ZN(n19619) );
  AND2_X1 U13073 ( .A1(n19693), .A2(n19894), .ZN(n19682) );
  OAI21_X1 U13074 ( .B1(n19719), .B2(n19854), .A(n19692), .ZN(n19709) );
  AND2_X1 U13075 ( .A1(n20103), .A2(n19713), .ZN(n19693) );
  INV_X1 U13076 ( .A(n19773), .ZN(n19776) );
  NOR2_X1 U13077 ( .A1(n20111), .A2(n20099), .ZN(n19822) );
  INV_X1 U13078 ( .A(n19989), .ZN(n19865) );
  INV_X1 U13079 ( .A(n19958), .ZN(n19949) );
  XNOR2_X1 U13080 ( .A(n16733), .B(n17600), .ZN(n19077) );
  NOR2_X1 U13081 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16866), .ZN(n16852) );
  NOR2_X1 U13082 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16909), .ZN(n16893) );
  NOR2_X1 U13083 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16934), .ZN(n16918) );
  OR2_X1 U13084 ( .A1(n16955), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n16956) );
  NOR2_X1 U13085 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16994), .ZN(n16993) );
  NOR2_X1 U13086 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17031), .ZN(n17010) );
  NOR2_X1 U13087 ( .A1(n19067), .A2(n18416), .ZN(n16737) );
  NOR2_X2 U13088 ( .A1(n19028), .A2(n17115), .ZN(n17121) );
  AND2_X1 U13089 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17236), .ZN(n17223) );
  AND2_X1 U13090 ( .A1(n18448), .A2(n17252), .ZN(n17236) );
  NAND2_X1 U13091 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17416), .ZN(n17413) );
  INV_X1 U13092 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17423) );
  NAND2_X1 U13093 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17467), .ZN(n17462) );
  NOR2_X1 U13094 ( .A1(n17564), .A2(n17481), .ZN(n17477) );
  NOR3_X1 U13095 ( .A1(n17564), .A2(n17517), .A3(n17644), .ZN(n17509) );
  INV_X1 U13096 ( .A(n17491), .ZN(n17515) );
  NOR2_X1 U13097 ( .A1(n17563), .A2(n17523), .ZN(n17559) );
  OAI21_X1 U13098 ( .B1(n16040), .B2(n16039), .A(n19069), .ZN(n17563) );
  NOR2_X1 U13099 ( .A1(n18022), .A2(n17907), .ZN(n18012) );
  INV_X1 U13100 ( .A(n17903), .ZN(n18274) );
  NOR2_X1 U13101 ( .A1(n15962), .A2(n15941), .ZN(n15969) );
  INV_X1 U13102 ( .A(n18312), .ZN(n18299) );
  NOR2_X1 U13103 ( .A1(n16729), .A2(n18382), .ZN(n18359) );
  NAND2_X1 U13104 ( .A1(n18926), .A2(n18414), .ZN(n18453) );
  INV_X1 U13105 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19086) );
  INV_X1 U13106 ( .A(n14848), .ZN(n13718) );
  OR2_X1 U13107 ( .A1(n13328), .A2(n9686), .ZN(n13296) );
  OR3_X1 U13108 ( .A1(n14748), .A2(n20989), .A3(n14717), .ZN(n14706) );
  INV_X1 U13109 ( .A(n20210), .ZN(n16093) );
  OR2_X1 U13110 ( .A1(n16115), .A2(n12482), .ZN(n16122) );
  INV_X1 U13111 ( .A(n16115), .ZN(n14903) );
  INV_X1 U13112 ( .A(n20274), .ZN(n20303) );
  NOR2_X1 U13113 ( .A1(n13296), .A2(n13295), .ZN(n13402) );
  OR2_X1 U13114 ( .A1(n13056), .A2(n13015), .ZN(n16278) );
  OR2_X1 U13115 ( .A1(n20485), .A2(n20653), .ZN(n20469) );
  AOI22_X1 U13116 ( .A1(n20435), .A2(n20438), .B1(n20685), .B2(n10195), .ZN(
        n20474) );
  OR2_X1 U13117 ( .A1(n20587), .A2(n20616), .ZN(n20557) );
  AOI22_X1 U13118 ( .A1(n20564), .A2(n20561), .B1(n20560), .B2(n10195), .ZN(
        n20585) );
  OR2_X1 U13119 ( .A1(n20587), .A2(n20586), .ZN(n20622) );
  NAND2_X1 U13120 ( .A1(n20680), .A2(n20617), .ZN(n20675) );
  AOI22_X1 U13121 ( .A1(n20692), .A2(n20687), .B1(n20685), .B2(n20684), .ZN(
        n20726) );
  NAND2_X1 U13122 ( .A1(n20680), .A2(n15212), .ZN(n20763) );
  INV_X1 U13123 ( .A(n20759), .ZN(n15242) );
  INV_X1 U13124 ( .A(n13717), .ZN(n13772) );
  OR2_X1 U13125 ( .A1(n20807), .A2(n20764), .ZN(n20846) );
  OR2_X1 U13126 ( .A1(n20807), .A2(n20586), .ZN(n20863) );
  INV_X1 U13127 ( .A(n20934), .ZN(n20868) );
  INV_X1 U13128 ( .A(n20916), .ZN(n20962) );
  AND2_X1 U13129 ( .A1(n13287), .A2(n13119), .ZN(n19098) );
  INV_X1 U13130 ( .A(n19317), .ZN(n19302) );
  INV_X1 U13131 ( .A(n19305), .ZN(n19315) );
  INV_X1 U13132 ( .A(n13273), .ZN(n15442) );
  INV_X1 U13133 ( .A(n13273), .ZN(n15440) );
  INV_X1 U13134 ( .A(n19379), .ZN(n19349) );
  OR2_X1 U13135 ( .A1(n19379), .A2(n13291), .ZN(n19356) );
  AND2_X1 U13136 ( .A1(n15522), .A2(n13990), .ZN(n19386) );
  NAND2_X1 U13137 ( .A1(n19388), .A2(n13224), .ZN(n13387) );
  INV_X1 U13138 ( .A(n19388), .ZN(n19419) );
  NAND2_X1 U13139 ( .A1(n13127), .A2(n10458), .ZN(n13219) );
  INV_X1 U13140 ( .A(n11344), .ZN(n11345) );
  INV_X1 U13141 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16418) );
  INV_X1 U13142 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16438) );
  XNOR2_X1 U13143 ( .A(n10789), .B(n10204), .ZN(n15630) );
  NAND2_X1 U13144 ( .A1(n11201), .A2(n20138), .ZN(n16524) );
  INV_X1 U13145 ( .A(n16519), .ZN(n19449) );
  NAND2_X1 U13146 ( .A1(n19755), .A2(n19656), .ZN(n19530) );
  AND2_X1 U13147 ( .A1(n19562), .A2(n19561), .ZN(n19572) );
  INV_X1 U13148 ( .A(n19583), .ZN(n19591) );
  NAND2_X1 U13149 ( .A1(n19656), .A2(n19894), .ZN(n19638) );
  INV_X1 U13150 ( .A(n19682), .ZN(n19655) );
  NAND2_X1 U13151 ( .A1(n19920), .A2(n19656), .ZN(n19712) );
  NAND2_X1 U13152 ( .A1(n19693), .A2(n19920), .ZN(n19743) );
  NAND2_X1 U13153 ( .A1(n19921), .A2(n19822), .ZN(n19835) );
  AND2_X1 U13154 ( .A1(n19818), .A2(n19817), .ZN(n19848) );
  NAND2_X1 U13155 ( .A1(n19921), .A2(n19894), .ZN(n19919) );
  INV_X1 U13156 ( .A(n20021), .ZN(n19959) );
  NAND2_X1 U13157 ( .A1(n19921), .A2(n19920), .ZN(n20001) );
  AND2_X1 U13158 ( .A1(n13615), .A2(n13614), .ZN(n16540) );
  INV_X1 U13159 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20043) );
  NOR2_X1 U13160 ( .A1(n18855), .A2(n17638), .ZN(n19089) );
  INV_X1 U13161 ( .A(n12808), .ZN(n16713) );
  INV_X1 U13162 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18020) );
  INV_X1 U13163 ( .A(n18448), .ZN(n17564) );
  NOR2_X1 U13164 ( .A1(n17239), .A2(n17238), .ZN(n17252) );
  INV_X1 U13165 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17415) );
  OR2_X1 U13166 ( .A1(n17530), .A2(n17558), .ZN(n17548) );
  NOR2_X2 U13167 ( .A1(n12549), .A2(n12548), .ZN(n17565) );
  NOR2_X1 U13168 ( .A1(n12560), .A2(n12559), .ZN(n17573) );
  INV_X1 U13169 ( .A(n17594), .ZN(n17587) );
  NOR2_X1 U13170 ( .A1(n19071), .A2(n17618), .ZN(n17615) );
  INV_X1 U13171 ( .A(n17618), .ZN(n17637) );
  NAND2_X1 U13172 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18012), .ZN(n17911) );
  INV_X1 U13173 ( .A(n17973), .ZN(n17991) );
  NAND2_X1 U13174 ( .A1(n12808), .A2(n16733), .ZN(n18079) );
  INV_X1 U13175 ( .A(n18396), .ZN(n18374) );
  INV_X1 U13176 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18906) );
  INV_X1 U13177 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18908) );
  INV_X1 U13178 ( .A(n19069), .ZN(n18924) );
  INV_X1 U13179 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19028) );
  INV_X1 U13180 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18952) );
  OAI21_X1 U13181 ( .B1(n15630), .B2(n19449), .A(n11204), .ZN(P2_U3025) );
  AOI22_X1 U13182 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10226) );
  AND2_X4 U13183 ( .A1(n13491), .A2(n10222), .ZN(n14503) );
  AOI22_X1 U13184 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10225) );
  INV_X2 U13185 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10222) );
  AND3_X4 U13186 ( .A1(n10222), .A2(n10221), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14504) );
  AOI22_X1 U13187 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10224) );
  AND2_X4 U13188 ( .A1(n13489), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10451) );
  AOI22_X1 U13189 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10223) );
  NAND4_X1 U13190 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10232) );
  AOI22_X1 U13191 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U13192 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U13193 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U13194 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10227) );
  NAND4_X1 U13195 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10231) );
  MUX2_X2 U13196 ( .A(n10232), .B(n10231), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10332) );
  INV_X1 U13197 ( .A(n10332), .ZN(n19499) );
  AOI22_X1 U13198 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13199 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13200 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U13201 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10233) );
  NAND4_X1 U13202 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10237) );
  NAND2_X1 U13203 ( .A1(n10237), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10244) );
  AOI22_X1 U13204 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13205 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13206 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13207 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10238) );
  NAND4_X1 U13208 ( .A1(n10241), .A2(n10240), .A3(n10239), .A4(n10238), .ZN(
        n10242) );
  NAND2_X1 U13209 ( .A1(n10242), .A2(n10275), .ZN(n10243) );
  AOI22_X1 U13210 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U13211 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10248) );
  NAND4_X1 U13212 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10257) );
  AOI22_X1 U13213 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13214 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10251) );
  AND2_X1 U13215 ( .A1(n10251), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10254) );
  AOI22_X1 U13216 ( .A1(n9644), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13217 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10252) );
  NAND4_X1 U13218 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10256) );
  AOI22_X1 U13219 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13220 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13221 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10259) );
  NAND4_X1 U13222 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10263) );
  NAND2_X1 U13223 ( .A1(n10263), .A2(n10275), .ZN(n10270) );
  AOI22_X1 U13224 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13225 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10266) );
  NAND4_X1 U13226 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  NAND2_X1 U13227 ( .A1(n10268), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10269) );
  NAND4_X1 U13228 ( .A1(n19499), .A2(n9653), .A3(n10321), .A4(n10328), .ZN(
        n10355) );
  INV_X1 U13229 ( .A(n10355), .ZN(n10343) );
  AOI22_X1 U13230 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U13231 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13232 ( .A1(n9644), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13233 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13234 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13235 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13236 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13237 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10276) );
  NAND4_X1 U13238 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10280) );
  AOI22_X1 U13239 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13240 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13241 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13242 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13243 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13244 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13245 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10288) );
  NAND4_X1 U13246 ( .A1(n10205), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10291) );
  NAND2_X1 U13247 ( .A1(n10499), .A2(n19470), .ZN(n10852) );
  AOI22_X1 U13248 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13249 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13250 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U13251 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13252 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13253 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13254 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13255 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10297) );
  NAND4_X1 U13256 ( .A1(n10300), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n10301) );
  AOI22_X1 U13257 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13258 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13259 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13260 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10304) );
  NAND4_X1 U13261 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10308) );
  AOI22_X1 U13262 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14504), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13263 ( .A1(n10309), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13264 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13265 ( .A1(n9644), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10310) );
  NAND4_X1 U13266 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10314) );
  INV_X4 U13267 ( .A(n10325), .ZN(n20152) );
  NAND2_X1 U13268 ( .A1(n19474), .A2(n20152), .ZN(n10334) );
  NAND2_X1 U13269 ( .A1(n10343), .A2(n10317), .ZN(n13289) );
  MUX2_X1 U13270 ( .A(n10328), .B(n10332), .S(n10837), .Z(n10319) );
  NAND3_X1 U13271 ( .A1(n10320), .A2(n10319), .A3(n10318), .ZN(n10323) );
  INV_X1 U13272 ( .A(n19470), .ZN(n10857) );
  AND2_X1 U13273 ( .A1(n19474), .A2(n10857), .ZN(n10322) );
  NAND2_X1 U13274 ( .A1(n10321), .A2(n10332), .ZN(n10330) );
  NAND2_X1 U13275 ( .A1(n10322), .A2(n10350), .ZN(n10833) );
  NAND3_X1 U13276 ( .A1(n10323), .A2(n10833), .A3(n20152), .ZN(n10352) );
  NAND2_X1 U13277 ( .A1(n10857), .A2(n11330), .ZN(n10324) );
  AND3_X2 U13278 ( .A1(n13289), .A2(n10352), .A3(n10324), .ZN(n10944) );
  NAND2_X1 U13279 ( .A1(n10499), .A2(n20152), .ZN(n10326) );
  NAND2_X2 U13280 ( .A1(n10960), .A2(n10325), .ZN(n10358) );
  NAND2_X1 U13282 ( .A1(n10342), .A2(n10321), .ZN(n10327) );
  NAND2_X1 U13283 ( .A1(n13122), .A2(n10327), .ZN(n10942) );
  NAND2_X2 U13284 ( .A1(n10944), .A2(n10329), .ZN(n10361) );
  INV_X1 U13285 ( .A(n10330), .ZN(n10331) );
  NAND3_X2 U13286 ( .A1(n10846), .A2(n10349), .A3(n10331), .ZN(n10843) );
  NAND2_X1 U13287 ( .A1(n10340), .A2(n10499), .ZN(n10339) );
  INV_X1 U13288 ( .A(n13291), .ZN(n10965) );
  NAND2_X1 U13289 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  INV_X1 U13290 ( .A(n10342), .ZN(n10839) );
  NAND2_X1 U13291 ( .A1(n11151), .A2(n10839), .ZN(n10928) );
  NAND2_X4 U13292 ( .A1(n10341), .A2(n10340), .ZN(n14517) );
  INV_X1 U13293 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U13294 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10347) );
  NOR2_X1 U13295 ( .A1(n10342), .A2(n10358), .ZN(n10344) );
  AND2_X2 U13296 ( .A1(n10344), .A2(n10343), .ZN(n10945) );
  INV_X1 U13297 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10345) );
  OAI211_X1 U13298 ( .C1(n14517), .C2(n13256), .A(n10347), .B(n10346), .ZN(
        n10348) );
  NAND2_X1 U13299 ( .A1(n10350), .A2(n10349), .ZN(n10809) );
  NAND3_X1 U13300 ( .A1(n14487), .A2(n10809), .A3(n19470), .ZN(n10351) );
  NAND2_X1 U13301 ( .A1(n10351), .A2(n10843), .ZN(n11150) );
  INV_X1 U13302 ( .A(n10935), .ZN(n10368) );
  NAND3_X1 U13303 ( .A1(n10844), .A2(n10321), .A3(n10354), .ZN(n10849) );
  NAND3_X1 U13304 ( .A1(n10849), .A2(n10835), .A3(n10332), .ZN(n10937) );
  NAND2_X1 U13305 ( .A1(n10937), .A2(n10939), .ZN(n10357) );
  NAND2_X1 U13306 ( .A1(n10355), .A2(n19474), .ZN(n10356) );
  OAI21_X2 U13307 ( .B1(n10370), .B2(n10359), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10384) );
  INV_X1 U13308 ( .A(n10384), .ZN(n10360) );
  NAND2_X1 U13309 ( .A1(n10360), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10363) );
  NAND2_X2 U13310 ( .A1(n10361), .A2(n11149), .ZN(n10927) );
  NOR2_X1 U13311 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16539) );
  INV_X1 U13312 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10375) );
  INV_X1 U13313 ( .A(n16539), .ZN(n10366) );
  NAND2_X1 U13314 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U13315 ( .A1(n10366), .A2(n10365), .ZN(n10367) );
  AOI21_X1 U13316 ( .B1(n10400), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10367), .ZN(
        n10372) );
  INV_X1 U13317 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19115) );
  NOR2_X1 U13319 ( .A1(n10342), .A2(n19097), .ZN(n10377) );
  INV_X1 U13320 ( .A(n10380), .ZN(n10382) );
  NAND2_X1 U13321 ( .A1(n10382), .A2(n10381), .ZN(n10383) );
  AOI21_X1 U13322 ( .B1(n19097), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U13323 ( .A1(n10903), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10391) );
  AOI22_X1 U13324 ( .A1(n10400), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10389) );
  NAND2_X1 U13325 ( .A1(n14562), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10388) );
  NAND2_X1 U13326 ( .A1(n13302), .A2(n10393), .ZN(n10392) );
  INV_X1 U13327 ( .A(n13302), .ZN(n10394) );
  NAND2_X1 U13328 ( .A1(n10394), .A2(n13304), .ZN(n10395) );
  NAND2_X1 U13329 ( .A1(n16539), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10397) );
  INV_X1 U13330 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13804) );
  NAND2_X1 U13331 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U13332 ( .A1(n10400), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10401) );
  OAI211_X1 U13333 ( .C1(n14517), .C2(n13804), .A(n10402), .B(n10401), .ZN(
        n10403) );
  NOR2_X1 U13335 ( .A1(n10404), .A2(n19321), .ZN(n10417) );
  AOI22_X1 U13336 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19885), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10423) );
  XNOR2_X2 U13337 ( .A(n10412), .B(n10414), .ZN(n13277) );
  NAND2_X1 U13338 ( .A1(n10590), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10422) );
  NOR2_X2 U13339 ( .A1(n13803), .A2(n10413), .ZN(n10589) );
  NOR2_X1 U13340 ( .A1(n10414), .A2(n19321), .ZN(n10426) );
  AOI22_X1 U13341 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10589), .B1(
        n19566), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10421) );
  AND2_X2 U13342 ( .A1(n13399), .A2(n10418), .ZN(n19631) );
  AND2_X1 U13343 ( .A1(n9639), .A2(n10426), .ZN(n10419) );
  AND2_X2 U13344 ( .A1(n10419), .A2(n13399), .ZN(n10591) );
  AOI22_X1 U13345 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19631), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U13346 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10596), .B1(
        n19855), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10440) );
  INV_X1 U13347 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10425) );
  NAND2_X1 U13348 ( .A1(n15374), .A2(n13277), .ZN(n10433) );
  INV_X1 U13349 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10424) );
  OAI22_X1 U13350 ( .A1(n10425), .A2(n19454), .B1(n19789), .B2(n10424), .ZN(
        n10430) );
  INV_X1 U13351 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n19832) );
  INV_X1 U13352 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10428) );
  OAI22_X1 U13353 ( .A1(n19832), .A2(n19815), .B1(n19963), .B2(n10428), .ZN(
        n10429) );
  NOR2_X1 U13354 ( .A1(n10430), .A2(n10429), .ZN(n10439) );
  INV_X1 U13355 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10436) );
  INV_X1 U13356 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10435) );
  AOI21_X1 U13357 ( .B1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n19599), .A(
        n10437), .ZN(n10438) );
  INV_X4 U13358 ( .A(n10499), .ZN(n14487) );
  AND2_X2 U13359 ( .A1(n9646), .A2(n10275), .ZN(n10653) );
  AOI22_X1 U13360 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13361 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10445) );
  AND2_X2 U13362 ( .A1(n14499), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10658) );
  AOI22_X1 U13363 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10444) );
  AND2_X2 U13364 ( .A1(n9681), .A2(n10275), .ZN(n14353) );
  AOI22_X1 U13365 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10443) );
  NAND4_X1 U13366 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10457) );
  AND2_X2 U13367 ( .A1(n10441), .A2(n10275), .ZN(n11015) );
  AOI22_X1 U13368 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U13369 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14334) );
  INV_X1 U13370 ( .A(n14334), .ZN(n10447) );
  NAND3_X1 U13371 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10799) );
  INV_X1 U13372 ( .A(n10799), .ZN(n10448) );
  AOI22_X1 U13373 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n14358), .ZN(n10450) );
  AND2_X1 U13374 ( .A1(n14504), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13375 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10449) );
  AND2_X1 U13376 ( .A1(n10450), .A2(n10449), .ZN(n10454) );
  AOI22_X1 U13378 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10453) );
  INV_X1 U13379 ( .A(n10451), .ZN(n13570) );
  NAND2_X1 U13380 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10452) );
  NAND4_X1 U13381 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10456) );
  INV_X1 U13382 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10463) );
  INV_X1 U13383 ( .A(n19631), .ZN(n19624) );
  INV_X1 U13384 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10460) );
  OR2_X2 U13385 ( .A1(n19624), .A2(n10460), .ZN(n10461) );
  OAI211_X1 U13386 ( .C1(n10581), .C2(n10463), .A(n10462), .B(n10461), .ZN(
        n10468) );
  NAND2_X1 U13387 ( .A1(n10591), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13388 ( .A1(n19885), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10467) );
  NAND2_X1 U13389 ( .A1(n10588), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10466) );
  INV_X1 U13390 ( .A(n19963), .ZN(n10583) );
  NAND2_X1 U13391 ( .A1(n10583), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10465) );
  INV_X1 U13392 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10470) );
  INV_X1 U13393 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10469) );
  OAI22_X1 U13394 ( .A1(n10470), .A2(n10582), .B1(n19789), .B2(n10469), .ZN(
        n10474) );
  INV_X1 U13395 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10472) );
  INV_X1 U13396 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10471) );
  OAI22_X1 U13397 ( .A1(n10472), .A2(n19454), .B1(n19815), .B2(n10471), .ZN(
        n10473) );
  NOR2_X1 U13398 ( .A1(n10474), .A2(n10473), .ZN(n10476) );
  AOI22_X1 U13399 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19855), .B1(
        n10590), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13400 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n14358), .ZN(n10480) );
  AOI22_X1 U13401 ( .A1(n11033), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13402 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14352), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13403 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n10659), .ZN(n10477) );
  NAND4_X1 U13404 ( .A1(n10480), .A2(n10479), .A3(n10478), .A4(n10477), .ZN(
        n10486) );
  AOI22_X1 U13405 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13406 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n14359), .ZN(n10483) );
  AOI22_X1 U13407 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U13408 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10658), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10481) );
  NAND4_X1 U13409 ( .A1(n10484), .A2(n10483), .A3(n10482), .A4(n10481), .ZN(
        n10485) );
  AOI22_X1 U13410 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13411 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U13412 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10488) );
  NAND2_X1 U13413 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10487) );
  AND3_X1 U13414 ( .A1(n10489), .A2(n10488), .A3(n10487), .ZN(n10491) );
  AOI22_X1 U13415 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10490) );
  NAND3_X1 U13416 ( .A1(n10492), .A2(n10491), .A3(n10490), .ZN(n10498) );
  AOI22_X1 U13417 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13418 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10495) );
  INV_X1 U13419 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n19977) );
  AOI22_X1 U13420 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13421 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10493) );
  NAND4_X1 U13422 ( .A1(n10496), .A2(n10495), .A3(n10494), .A4(n10493), .ZN(
        n10497) );
  NAND2_X1 U13423 ( .A1(n10499), .A2(n13242), .ZN(n10500) );
  OR2_X1 U13424 ( .A1(n11159), .A2(n10500), .ZN(n11163) );
  AOI22_X1 U13425 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13426 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n14358), .ZN(n10503) );
  NAND2_X1 U13427 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13428 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10501) );
  AND3_X1 U13429 ( .A1(n10503), .A2(n10502), .A3(n10501), .ZN(n10505) );
  AOI22_X1 U13430 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10504) );
  NAND3_X1 U13431 ( .A1(n10506), .A2(n10505), .A3(n10504), .ZN(n10513) );
  AOI22_X1 U13432 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13433 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13434 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14351), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13435 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10508) );
  NAND4_X1 U13436 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10512) );
  NAND2_X1 U13437 ( .A1(n11163), .A2(n11162), .ZN(n11161) );
  AND2_X2 U13438 ( .A1(n10514), .A2(n11161), .ZN(n10579) );
  NAND2_X1 U13439 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10519) );
  NAND2_X1 U13440 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10518) );
  NAND2_X1 U13441 ( .A1(n11033), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10517) );
  NAND2_X1 U13442 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10516) );
  NAND2_X1 U13443 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10523) );
  NAND2_X1 U13444 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U13445 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13446 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10520) );
  AOI22_X1 U13447 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n14358), .ZN(n10527) );
  NAND2_X1 U13448 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10526) );
  INV_X1 U13449 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19847) );
  NAND2_X1 U13450 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10525) );
  AND3_X1 U13451 ( .A1(n10527), .A2(n10526), .A3(n10525), .ZN(n10533) );
  NAND2_X1 U13452 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10531) );
  NAND2_X1 U13453 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13454 ( .A1(n14353), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10529) );
  NAND2_X1 U13455 ( .A1(n10644), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10528) );
  NAND4_X1 U13456 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n11010) );
  INV_X1 U13457 ( .A(n11010), .ZN(n10536) );
  NAND2_X1 U13458 ( .A1(n13798), .A2(n10536), .ZN(n10548) );
  INV_X1 U13459 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U13460 ( .A1(n10345), .A2(n13274), .ZN(n10538) );
  MUX2_X1 U13461 ( .A(n10538), .B(n11159), .S(n11295), .Z(n10552) );
  MUX2_X1 U13462 ( .A(n20125), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10817) );
  INV_X1 U13463 ( .A(n10795), .ZN(n10540) );
  NAND2_X1 U13464 ( .A1(n14333), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10544) );
  OAI21_X1 U13465 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14333), .A(
        n10544), .ZN(n10541) );
  XNOR2_X1 U13466 ( .A(n10543), .B(n10541), .ZN(n10815) );
  NAND2_X1 U13467 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20116), .ZN(
        n10542) );
  NAND2_X1 U13468 ( .A1(n10543), .A2(n10542), .ZN(n10545) );
  MUX2_X1 U13469 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20109), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10571) );
  XNOR2_X1 U13470 ( .A(n10570), .B(n10571), .ZN(n10826) );
  INV_X1 U13471 ( .A(n10826), .ZN(n10825) );
  MUX2_X1 U13472 ( .A(n10993), .B(n10825), .S(n10358), .Z(n10806) );
  INV_X1 U13473 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13864) );
  MUX2_X1 U13474 ( .A(n10806), .B(n13864), .S(n14552), .Z(n10546) );
  OAI21_X1 U13475 ( .B1(n10547), .B2(n10546), .A(n10618), .ZN(n13863) );
  XNOR2_X1 U13476 ( .A(n10549), .B(n10552), .ZN(n10556) );
  XNOR2_X1 U13477 ( .A(n10556), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13100) );
  AND2_X1 U13478 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10550) );
  NAND2_X1 U13479 ( .A1(n14552), .A2(n10550), .ZN(n10551) );
  NAND2_X1 U13480 ( .A1(n10552), .A2(n10551), .ZN(n19301) );
  INV_X1 U13481 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19441) );
  INV_X1 U13482 ( .A(n13242), .ZN(n13241) );
  OAI21_X1 U13483 ( .B1(n20135), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10795), .ZN(n10812) );
  MUX2_X1 U13484 ( .A(n13241), .B(n10812), .S(n10358), .Z(n10804) );
  INV_X1 U13485 ( .A(n10804), .ZN(n10553) );
  MUX2_X1 U13486 ( .A(n10553), .B(P2_EBX_REG_0__SCAN_IN), .S(n14552), .Z(
        n19318) );
  NAND2_X1 U13487 ( .A1(n19318), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13254) );
  OAI21_X1 U13488 ( .B1(n19301), .B2(n19441), .A(n13254), .ZN(n10555) );
  NAND2_X1 U13489 ( .A1(n19301), .A2(n19441), .ZN(n10554) );
  AND2_X1 U13490 ( .A1(n10555), .A2(n10554), .ZN(n13099) );
  NAND2_X1 U13491 ( .A1(n13100), .A2(n13099), .ZN(n13098) );
  INV_X1 U13492 ( .A(n10556), .ZN(n15368) );
  NAND2_X1 U13493 ( .A1(n15368), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10557) );
  NAND2_X1 U13494 ( .A1(n13098), .A2(n10557), .ZN(n13800) );
  AOI22_X1 U13495 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13496 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n14358), .ZN(n10560) );
  NAND2_X1 U13497 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10559) );
  NAND2_X1 U13498 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10558) );
  AND3_X1 U13499 ( .A1(n10560), .A2(n10559), .A3(n10558), .ZN(n10562) );
  AOI22_X1 U13500 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n10659), .ZN(n10561) );
  NAND3_X1 U13501 ( .A1(n10563), .A2(n10562), .A3(n10561), .ZN(n10569) );
  AOI22_X1 U13502 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11033), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13503 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13504 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14351), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13505 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14353), .B1(
        n14352), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10564) );
  NAND4_X1 U13506 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10568) );
  INV_X1 U13508 ( .A(n10571), .ZN(n10573) );
  NOR2_X1 U13509 ( .A1(n10275), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10572) );
  NOR2_X1 U13510 ( .A1(n16037), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10575) );
  AND2_X1 U13511 ( .A1(n10790), .A2(n10575), .ZN(n10827) );
  MUX2_X1 U13512 ( .A(n11156), .B(n10827), .S(n10358), .Z(n10805) );
  MUX2_X1 U13513 ( .A(P2_EBX_REG_4__SCAN_IN), .B(n10805), .S(n11295), .Z(
        n10617) );
  XNOR2_X1 U13514 ( .A(n10618), .B(n10617), .ZN(n19283) );
  XNOR2_X1 U13515 ( .A(n19283), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13870) );
  INV_X1 U13516 ( .A(n19283), .ZN(n10576) );
  NAND2_X1 U13517 ( .A1(n10576), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10577) );
  NAND2_X1 U13518 ( .A1(n10578), .A2(n10577), .ZN(n16441) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19461), .B1(
        n19783), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13520 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19532), .B1(
        n19720), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10586) );
  INV_X1 U13521 ( .A(n19815), .ZN(n10677) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n10677), .B1(
        n10583), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13523 ( .A1(n19599), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10584) );
  AOI22_X1 U13524 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19885), .B1(
        n10588), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13525 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10589), .B1(
        n19566), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U13526 ( .A1(n10590), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10593) );
  AOI22_X1 U13527 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19631), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10592) );
  INV_X1 U13528 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10599) );
  INV_X1 U13529 ( .A(n19855), .ZN(n10598) );
  INV_X1 U13530 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10597) );
  OAI22_X1 U13531 ( .A1(n10599), .A2(n19659), .B1(n10598), .B2(n10597), .ZN(
        n10600) );
  INV_X1 U13532 ( .A(n10600), .ZN(n10601) );
  NAND3_X1 U13533 ( .A1(n10211), .A2(n10213), .A3(n10601), .ZN(n10616) );
  AOI22_X1 U13534 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13535 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13536 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13537 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10602) );
  NAND4_X1 U13538 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n10613) );
  AOI22_X1 U13539 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13540 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13541 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10606) );
  AND2_X1 U13542 ( .A1(n10607), .A2(n10606), .ZN(n10610) );
  AOI22_X1 U13543 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13544 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10608) );
  NAND4_X1 U13545 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10612) );
  INV_X1 U13546 ( .A(n11001), .ZN(n10614) );
  NAND2_X1 U13547 ( .A1(n10614), .A2(n10458), .ZN(n10615) );
  NAND2_X1 U13548 ( .A1(n11175), .A2(n10536), .ZN(n10623) );
  INV_X1 U13549 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10619) );
  MUX2_X1 U13550 ( .A(n10619), .B(n11001), .S(n11295), .Z(n10620) );
  NOR2_X1 U13551 ( .A1(n10621), .A2(n10620), .ZN(n10622) );
  OR2_X1 U13552 ( .A1(n10693), .A2(n10622), .ZN(n13853) );
  NAND2_X1 U13553 ( .A1(n10623), .A2(n13853), .ZN(n10624) );
  INV_X1 U13554 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16506) );
  XNOR2_X1 U13555 ( .A(n10624), .B(n16506), .ZN(n16442) );
  NAND2_X1 U13556 ( .A1(n10624), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10625) );
  INV_X1 U13557 ( .A(n11015), .ZN(n10631) );
  INV_X1 U13558 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10630) );
  INV_X1 U13559 ( .A(n11033), .ZN(n10629) );
  INV_X1 U13560 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10628) );
  OAI22_X1 U13561 ( .A1(n10631), .A2(n10630), .B1(n10629), .B2(n10628), .ZN(
        n10638) );
  INV_X1 U13562 ( .A(n10507), .ZN(n10636) );
  INV_X1 U13563 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10635) );
  INV_X1 U13564 ( .A(n10632), .ZN(n10634) );
  INV_X1 U13565 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10633) );
  OAI22_X1 U13566 ( .A1(n10636), .A2(n10635), .B1(n10634), .B2(n10633), .ZN(
        n10637) );
  OR2_X1 U13567 ( .A1(n10638), .A2(n10637), .ZN(n10652) );
  INV_X1 U13568 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10643) );
  INV_X1 U13569 ( .A(n10639), .ZN(n10642) );
  INV_X1 U13570 ( .A(n14353), .ZN(n10641) );
  INV_X1 U13571 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10640) );
  OAI22_X1 U13572 ( .A1(n10643), .A2(n10642), .B1(n10641), .B2(n10640), .ZN(
        n10650) );
  INV_X1 U13573 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10648) );
  INV_X1 U13574 ( .A(n14351), .ZN(n10647) );
  INV_X1 U13575 ( .A(n10644), .ZN(n10646) );
  INV_X1 U13576 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10645) );
  OAI22_X1 U13577 ( .A1(n10648), .A2(n10647), .B1(n10646), .B2(n10645), .ZN(
        n10649) );
  OR2_X1 U13578 ( .A1(n10650), .A2(n10649), .ZN(n10651) );
  NOR2_X1 U13579 ( .A1(n10652), .A2(n10651), .ZN(n10672) );
  INV_X1 U13580 ( .A(n10653), .ZN(n10657) );
  INV_X1 U13581 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10683) );
  INV_X1 U13582 ( .A(n10654), .ZN(n10656) );
  INV_X1 U13583 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10655) );
  OAI22_X1 U13584 ( .A1(n10657), .A2(n10683), .B1(n10656), .B2(n10655), .ZN(
        n10665) );
  INV_X1 U13585 ( .A(n10658), .ZN(n10663) );
  INV_X1 U13586 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10662) );
  INV_X1 U13587 ( .A(n10659), .ZN(n10661) );
  INV_X1 U13588 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10660) );
  OAI22_X1 U13589 ( .A1(n10663), .A2(n10662), .B1(n10661), .B2(n10660), .ZN(
        n10664) );
  OR2_X1 U13590 ( .A1(n10665), .A2(n10664), .ZN(n10670) );
  AOI22_X1 U13591 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n14358), .ZN(n10668) );
  NAND2_X1 U13592 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10667) );
  NAND2_X1 U13593 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10666) );
  NAND3_X1 U13594 ( .A1(n10668), .A2(n10667), .A3(n10666), .ZN(n10669) );
  NOR2_X1 U13595 ( .A1(n10670), .A2(n10669), .ZN(n10671) );
  INV_X1 U13596 ( .A(n10690), .ZN(n11005) );
  AOI22_X1 U13597 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19461), .B1(
        n19783), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13598 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19532), .B1(
        n19720), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13599 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10588), .B1(
        n10583), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13600 ( .A1(n19599), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10673) );
  NAND4_X1 U13601 ( .A1(n10676), .A2(n10675), .A3(n10674), .A4(n10673), .ZN(
        n10686) );
  AOI22_X1 U13602 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19885), .B1(
        n10677), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13603 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19631), .B1(
        n10589), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10680) );
  NAND2_X1 U13604 ( .A1(n19855), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10679) );
  AOI22_X1 U13605 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19566), .B1(
        n10591), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10678) );
  NAND4_X1 U13606 ( .A1(n10681), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        n10685) );
  INV_X1 U13607 ( .A(n10590), .ZN(n19922) );
  INV_X1 U13608 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10682) );
  OAI22_X1 U13609 ( .A1(n10683), .A2(n19659), .B1(n19922), .B2(n10682), .ZN(
        n10684) );
  MUX2_X1 U13610 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n10690), .S(n11295), .Z(
        n10691) );
  INV_X1 U13611 ( .A(n10691), .ZN(n10692) );
  AND2_X2 U13612 ( .A1(n10693), .A2(n10692), .ZN(n10700) );
  NOR2_X1 U13613 ( .A1(n10693), .A2(n10692), .ZN(n10694) );
  OR2_X1 U13614 ( .A1(n10700), .A2(n10694), .ZN(n19274) );
  INV_X1 U13615 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14218) );
  NAND2_X1 U13616 ( .A1(n10695), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10696) );
  INV_X1 U13617 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10698) );
  MUX2_X1 U13618 ( .A(n10698), .B(n11010), .S(n11295), .Z(n10699) );
  XNOR2_X1 U13619 ( .A(n10700), .B(n10110), .ZN(n19260) );
  INV_X1 U13620 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10701) );
  NOR2_X1 U13621 ( .A1(n11295), .A2(n10701), .ZN(n10703) );
  INV_X1 U13622 ( .A(n10703), .ZN(n10702) );
  XNOR2_X1 U13623 ( .A(n10704), .B(n10702), .ZN(n19245) );
  AND2_X1 U13624 ( .A1(n19245), .A2(n11189), .ZN(n15675) );
  INV_X1 U13625 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U13626 ( .A1(n14552), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10705) );
  OAI21_X1 U13627 ( .B1(n9748), .B2(n10705), .A(n14554), .ZN(n10706) );
  OR2_X1 U13628 ( .A1(n10714), .A2(n10706), .ZN(n19236) );
  INV_X1 U13629 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15867) );
  OAI21_X1 U13630 ( .B1(n19236), .B2(n10536), .A(n15867), .ZN(n15872) );
  NAND2_X1 U13631 ( .A1(n19245), .A2(n14550), .ZN(n10707) );
  INV_X1 U13632 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U13633 ( .A1(n10707), .A2(n11188), .ZN(n15676) );
  INV_X1 U13634 ( .A(n19260), .ZN(n10708) );
  INV_X1 U13635 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11192) );
  NAND2_X1 U13636 ( .A1(n10708), .A2(n11192), .ZN(n15674) );
  AND2_X1 U13637 ( .A1(n15676), .A2(n15674), .ZN(n15868) );
  NAND2_X1 U13638 ( .A1(n14552), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10709) );
  XNOR2_X1 U13639 ( .A(n10710), .B(n10709), .ZN(n15362) );
  NAND2_X1 U13640 ( .A1(n15362), .A2(n14550), .ZN(n10711) );
  INV_X1 U13641 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15891) );
  NAND2_X1 U13642 ( .A1(n10711), .A2(n15891), .ZN(n15886) );
  AND3_X1 U13643 ( .A1(n15872), .A2(n15868), .A3(n15886), .ZN(n10712) );
  NAND2_X1 U13644 ( .A1(n14552), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10713) );
  OR2_X1 U13645 ( .A1(n10714), .A2(n10713), .ZN(n10716) );
  INV_X1 U13646 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13630) );
  INV_X1 U13647 ( .A(n10724), .ZN(n10715) );
  NAND2_X1 U13648 ( .A1(n10716), .A2(n10715), .ZN(n10721) );
  INV_X1 U13649 ( .A(n10721), .ZN(n13086) );
  AOI21_X1 U13650 ( .B1(n13086), .B2(n14550), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16408) );
  INV_X1 U13651 ( .A(n19236), .ZN(n10718) );
  AND2_X1 U13652 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U13653 ( .A1(n10718), .A2(n10717), .ZN(n15871) );
  AND2_X1 U13654 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10719) );
  NAND2_X1 U13655 ( .A1(n15362), .A2(n10719), .ZN(n15885) );
  NAND2_X1 U13656 ( .A1(n15871), .A2(n15885), .ZN(n16406) );
  NAND2_X1 U13657 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10720) );
  NOR2_X1 U13658 ( .A1(n10721), .A2(n10720), .ZN(n16407) );
  NOR2_X1 U13659 ( .A1(n16406), .A2(n16407), .ZN(n10722) );
  NAND2_X1 U13660 ( .A1(n14552), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10723) );
  NAND3_X1 U13661 ( .A1(n14552), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n10725), 
        .ZN(n10726) );
  NAND2_X1 U13662 ( .A1(n10733), .A2(n10726), .ZN(n19225) );
  NAND2_X1 U13663 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10727) );
  NOR2_X1 U13664 ( .A1(n19225), .A2(n10727), .ZN(n15855) );
  OR2_X1 U13665 ( .A1(n19225), .A2(n10536), .ZN(n10728) );
  INV_X1 U13666 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16387) );
  NAND2_X1 U13667 ( .A1(n10728), .A2(n16387), .ZN(n11267) );
  INV_X1 U13668 ( .A(n11267), .ZN(n15856) );
  INV_X1 U13669 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10729) );
  NOR2_X1 U13670 ( .A1(n11295), .A2(n10729), .ZN(n10732) );
  INV_X1 U13671 ( .A(n10732), .ZN(n10730) );
  XNOR2_X1 U13672 ( .A(n10733), .B(n10730), .ZN(n19216) );
  NAND2_X1 U13673 ( .A1(n19216), .A2(n14550), .ZN(n10731) );
  INV_X1 U13674 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16468) );
  NAND2_X1 U13675 ( .A1(n10731), .A2(n16468), .ZN(n16390) );
  NAND2_X1 U13676 ( .A1(n10743), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10734) );
  MUX2_X1 U13677 ( .A(n10734), .B(n10743), .S(n11295), .Z(n10736) );
  INV_X1 U13678 ( .A(n10743), .ZN(n10735) );
  INV_X1 U13679 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U13680 ( .A1(n10735), .A2(n13841), .ZN(n10741) );
  NAND2_X1 U13681 ( .A1(n10736), .A2(n10741), .ZN(n19204) );
  INV_X1 U13682 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15842) );
  OAI21_X1 U13683 ( .B1(n19204), .B2(n10536), .A(n15842), .ZN(n15834) );
  INV_X1 U13684 ( .A(n19204), .ZN(n10738) );
  AND2_X1 U13685 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13686 ( .A1(n10738), .A2(n10737), .ZN(n16371) );
  INV_X1 U13687 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10739) );
  NOR2_X1 U13688 ( .A1(n11295), .A2(n10739), .ZN(n10740) );
  NAND2_X1 U13689 ( .A1(n10741), .A2(n10740), .ZN(n10744) );
  NOR2_X1 U13690 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n10742) );
  NAND2_X1 U13691 ( .A1(n10744), .A2(n9713), .ZN(n15356) );
  NAND2_X1 U13692 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10745) );
  OR2_X1 U13693 ( .A1(n15356), .A2(n10745), .ZN(n16373) );
  OR2_X1 U13694 ( .A1(n15356), .A2(n10536), .ZN(n10746) );
  INV_X1 U13695 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16455) );
  NAND2_X1 U13696 ( .A1(n10746), .A2(n16455), .ZN(n16374) );
  INV_X1 U13697 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10755) );
  NOR2_X1 U13698 ( .A1(n11295), .A2(n10755), .ZN(n10747) );
  INV_X1 U13699 ( .A(n14554), .ZN(n11296) );
  AOI21_X1 U13700 ( .B1(n9713), .B2(n10747), .A(n11296), .ZN(n10748) );
  NAND2_X1 U13701 ( .A1(n19191), .A2(n14550), .ZN(n10749) );
  INV_X1 U13702 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15818) );
  XNOR2_X1 U13703 ( .A(n10749), .B(n15818), .ZN(n15667) );
  AND2_X1 U13704 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U13705 ( .A1(n19191), .A2(n10751), .ZN(n11276) );
  NAND2_X1 U13706 ( .A1(n15668), .A2(n11276), .ZN(n15659) );
  INV_X1 U13707 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10752) );
  NOR2_X1 U13708 ( .A1(n11295), .A2(n10752), .ZN(n10753) );
  NAND2_X1 U13709 ( .A1(n10754), .A2(n10753), .ZN(n10757) );
  NAND2_X1 U13710 ( .A1(n10755), .A2(n10752), .ZN(n10756) );
  INV_X1 U13711 ( .A(n10770), .ZN(n10762) );
  NAND2_X1 U13712 ( .A1(n10757), .A2(n10762), .ZN(n10759) );
  INV_X1 U13713 ( .A(n10759), .ZN(n19183) );
  AND2_X1 U13714 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10758) );
  NAND2_X1 U13715 ( .A1(n19183), .A2(n10758), .ZN(n15657) );
  INV_X1 U13716 ( .A(n15657), .ZN(n10760) );
  INV_X1 U13717 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11196) );
  OAI21_X1 U13718 ( .B1(n10759), .B2(n10536), .A(n11196), .ZN(n15658) );
  OAI21_X2 U13719 ( .B1(n15659), .B2(n10760), .A(n15658), .ZN(n15647) );
  NAND2_X1 U13720 ( .A1(n14552), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10761) );
  MUX2_X1 U13721 ( .A(n14552), .B(n10761), .S(n10762), .Z(n10763) );
  NAND2_X1 U13722 ( .A1(n10763), .A2(n10767), .ZN(n19165) );
  NAND2_X1 U13723 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10764) );
  INV_X1 U13724 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10765) );
  NOR2_X1 U13725 ( .A1(n11295), .A2(n10765), .ZN(n10766) );
  NAND2_X1 U13726 ( .A1(n10767), .A2(n10766), .ZN(n10771) );
  INV_X1 U13727 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19164) );
  NAND2_X1 U13728 ( .A1(n19164), .A2(n10765), .ZN(n10768) );
  NAND2_X1 U13729 ( .A1(n14552), .A2(n10768), .ZN(n10769) );
  AND2_X2 U13730 ( .A1(n10770), .A2(n10769), .ZN(n10782) );
  INV_X1 U13731 ( .A(n10782), .ZN(n10776) );
  NAND2_X1 U13732 ( .A1(n10771), .A2(n10776), .ZN(n19156) );
  NOR2_X1 U13733 ( .A1(n19156), .A2(n10536), .ZN(n10773) );
  NAND2_X1 U13734 ( .A1(n10773), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15637) );
  OR2_X1 U13735 ( .A1(n19165), .A2(n10536), .ZN(n10772) );
  INV_X1 U13736 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15802) );
  INV_X1 U13737 ( .A(n15638), .ZN(n15650) );
  OR2_X1 U13738 ( .A1(n10773), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15636) );
  NAND2_X1 U13739 ( .A1(n15650), .A2(n15636), .ZN(n10774) );
  NAND2_X1 U13740 ( .A1(n14552), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10775) );
  XNOR2_X1 U13741 ( .A(n10776), .B(n10775), .ZN(n19142) );
  NAND2_X1 U13742 ( .A1(n19142), .A2(n14550), .ZN(n10778) );
  INV_X1 U13743 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U13744 ( .A1(n10778), .A2(n10777), .ZN(n10780) );
  AND2_X1 U13745 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10779) );
  NAND2_X1 U13746 ( .A1(n19142), .A2(n10779), .ZN(n11280) );
  INV_X1 U13747 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13748 ( .A1(n10782), .A2(n10781), .ZN(n10785) );
  INV_X1 U13749 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10783) );
  NOR2_X1 U13750 ( .A1(n11295), .A2(n10783), .ZN(n10784) );
  AOI21_X1 U13751 ( .B1(n10785), .B2(n10784), .A(n11296), .ZN(n10786) );
  OR2_X2 U13752 ( .A1(n10785), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11286) );
  AND2_X1 U13753 ( .A1(n10786), .A2(n11286), .ZN(n19129) );
  NAND2_X1 U13754 ( .A1(n19129), .A2(n14550), .ZN(n10788) );
  INV_X1 U13755 ( .A(n10788), .ZN(n10787) );
  NAND2_X1 U13756 ( .A1(n10787), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11281) );
  INV_X1 U13757 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U13758 ( .A1(n10788), .A2(n11231), .ZN(n11272) );
  NOR3_X1 U13759 ( .A1(n10827), .A2(n10815), .A3(n10826), .ZN(n10796) );
  INV_X1 U13760 ( .A(n10796), .ZN(n10798) );
  INV_X1 U13761 ( .A(n10790), .ZN(n10792) );
  AND2_X1 U13762 ( .A1(n16037), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10791) );
  INV_X1 U13763 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15955) );
  NAND2_X1 U13764 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15955), .ZN(
        n10793) );
  XNOR2_X1 U13765 ( .A(n10817), .B(n10795), .ZN(n10813) );
  NAND2_X1 U13766 ( .A1(n10813), .A2(n10796), .ZN(n10797) );
  OAI21_X1 U13767 ( .B1(n10812), .B2(n10798), .A(n13579), .ZN(n10801) );
  INV_X1 U13768 ( .A(n14359), .ZN(n10800) );
  AND2_X1 U13769 ( .A1(n15955), .A2(n10799), .ZN(n13586) );
  AOI21_X1 U13770 ( .B1(n10800), .B2(n13586), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n20128) );
  MUX2_X1 U13771 ( .A(n10801), .B(n20128), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20140) );
  INV_X1 U13772 ( .A(n10817), .ZN(n10803) );
  OAI21_X1 U13773 ( .B1(n10804), .B2(n10803), .A(n10802), .ZN(n10807) );
  INV_X1 U13774 ( .A(n10805), .ZN(n10824) );
  NAND3_X1 U13775 ( .A1(n10807), .A2(n10824), .A3(n10806), .ZN(n10808) );
  NAND2_X1 U13776 ( .A1(n10808), .A2(n10830), .ZN(n20137) );
  NAND2_X1 U13777 ( .A1(n10458), .A2(n11330), .ZN(n10847) );
  OAI22_X1 U13778 ( .A1(n20140), .A2(n10458), .B1(n20137), .B2(n10847), .ZN(
        n10810) );
  INV_X1 U13779 ( .A(n11332), .ZN(n10860) );
  NAND2_X1 U13780 ( .A1(n11330), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13223) );
  NAND2_X1 U13781 ( .A1(n13223), .A2(n14487), .ZN(n10811) );
  MUX2_X1 U13782 ( .A(n10358), .B(n10811), .S(n10815), .Z(n10823) );
  INV_X1 U13783 ( .A(n10812), .ZN(n10818) );
  OAI21_X1 U13784 ( .B1(n14487), .B2(n10818), .A(n10813), .ZN(n10814) );
  OAI21_X1 U13785 ( .B1(n10815), .B2(n14487), .A(n10814), .ZN(n10816) );
  NAND2_X1 U13786 ( .A1(n10816), .A2(n20152), .ZN(n10821) );
  NAND2_X1 U13787 ( .A1(n10818), .A2(n10817), .ZN(n10819) );
  NAND2_X1 U13788 ( .A1(n13080), .A2(n10819), .ZN(n10820) );
  NAND2_X1 U13789 ( .A1(n10821), .A2(n10820), .ZN(n10822) );
  NOR2_X1 U13790 ( .A1(n10827), .A2(n10826), .ZN(n10828) );
  MUX2_X1 U13791 ( .A(n10829), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19097), .Z(n10832) );
  AOI21_X1 U13792 ( .B1(n10832), .B2(n20152), .A(n10321), .ZN(n10856) );
  INV_X1 U13793 ( .A(n10833), .ZN(n10834) );
  NAND2_X1 U13794 ( .A1(n10834), .A2(n20152), .ZN(n13587) );
  NAND2_X1 U13795 ( .A1(n10835), .A2(n19470), .ZN(n10836) );
  NAND2_X1 U13796 ( .A1(n13587), .A2(n10836), .ZN(n10842) );
  NAND2_X1 U13797 ( .A1(n10837), .A2(n10458), .ZN(n10931) );
  NAND2_X1 U13798 ( .A1(n10931), .A2(n20152), .ZN(n10838) );
  NAND2_X1 U13799 ( .A1(n10838), .A2(n10332), .ZN(n10840) );
  AOI21_X1 U13800 ( .B1(n10840), .B2(n19470), .A(n10839), .ZN(n10841) );
  NAND2_X1 U13801 ( .A1(n10842), .A2(n10841), .ZN(n10934) );
  NAND2_X1 U13802 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20150) );
  INV_X1 U13803 ( .A(n20150), .ZN(n20029) );
  NAND2_X1 U13804 ( .A1(n20043), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20160) );
  INV_X2 U13805 ( .A(n20160), .ZN(n20159) );
  NAND2_X2 U13806 ( .A1(n20159), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20086) );
  NOR2_X1 U13807 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20040) );
  INV_X1 U13808 ( .A(n20040), .ZN(n20030) );
  NAND3_X1 U13809 ( .A1(n20043), .A2(n20086), .A3(n20030), .ZN(n20035) );
  NOR2_X1 U13810 ( .A1(n20029), .A2(n20035), .ZN(n13500) );
  NAND3_X1 U13811 ( .A1(n13613), .A2(n13579), .A3(n13500), .ZN(n10850) );
  INV_X1 U13812 ( .A(n10844), .ZN(n10845) );
  OAI21_X1 U13813 ( .B1(n10846), .B2(n10845), .A(n10332), .ZN(n10848) );
  INV_X1 U13814 ( .A(n10847), .ZN(n13082) );
  NAND2_X1 U13815 ( .A1(n10848), .A2(n13082), .ZN(n10938) );
  NAND3_X1 U13816 ( .A1(n10850), .A2(n10849), .A3(n10938), .ZN(n10851) );
  NOR2_X1 U13817 ( .A1(n10934), .A2(n10851), .ZN(n13504) );
  NAND2_X1 U13818 ( .A1(n10843), .A2(n14487), .ZN(n10853) );
  NAND4_X1 U13819 ( .A1(n10853), .A2(n13579), .A3(n10852), .A4(n20150), .ZN(
        n10854) );
  NAND2_X1 U13820 ( .A1(n13504), .A2(n10854), .ZN(n10855) );
  AOI21_X1 U13821 ( .B1(n13221), .B2(n10856), .A(n10855), .ZN(n10859) );
  NAND3_X1 U13822 ( .A1(n10860), .A2(n10859), .A3(n10858), .ZN(n10861) );
  NAND2_X1 U13823 ( .A1(n16035), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13077) );
  AND2_X1 U13824 ( .A1(n11200), .A2(n13080), .ZN(n20139) );
  NAND2_X1 U13825 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10865) );
  AOI22_X1 U13826 ( .A1(n14561), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10863) );
  NAND2_X1 U13827 ( .A1(n14562), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10862) );
  AND2_X1 U13828 ( .A1(n10863), .A2(n10862), .ZN(n10864) );
  NAND2_X1 U13829 ( .A1(n10865), .A2(n10864), .ZN(n13545) );
  NAND2_X1 U13830 ( .A1(n10867), .A2(n10866), .ZN(n10872) );
  INV_X1 U13831 ( .A(n10868), .ZN(n10870) );
  NAND2_X1 U13832 ( .A1(n10870), .A2(n10869), .ZN(n10871) );
  NAND2_X1 U13833 ( .A1(n10872), .A2(n10871), .ZN(n13443) );
  INV_X1 U13834 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11000) );
  NAND2_X1 U13835 ( .A1(n14561), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U13836 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10873) );
  OAI211_X1 U13837 ( .C1(n14517), .C2(n11000), .A(n10874), .B(n10873), .ZN(
        n10875) );
  AOI21_X1 U13838 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10875), .ZN(n13444) );
  INV_X1 U13839 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13852) );
  NAND2_X1 U13840 ( .A1(n14561), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U13841 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10877) );
  OAI211_X1 U13842 ( .C1(n14517), .C2(n13852), .A(n10878), .B(n10877), .ZN(
        n10879) );
  AOI21_X1 U13843 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10879), .ZN(n13448) );
  INV_X1 U13844 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U13845 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10881) );
  AOI22_X1 U13846 ( .A1(n14561), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10880) );
  OAI211_X1 U13847 ( .C1(n14517), .C2(n11007), .A(n10881), .B(n10880), .ZN(
        n13531) );
  INV_X1 U13848 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U13849 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10883) );
  AOI22_X1 U13850 ( .A1(n14561), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10882) );
  OAI211_X1 U13851 ( .C1(n14517), .C2(n11012), .A(n10883), .B(n10882), .ZN(
        n13560) );
  INV_X1 U13852 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11030) );
  NAND2_X1 U13853 ( .A1(n14561), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U13854 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10884) );
  OAI211_X1 U13855 ( .C1(n14517), .C2(n11030), .A(n10885), .B(n10884), .ZN(
        n10886) );
  AOI21_X1 U13856 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10886), .ZN(n13620) );
  INV_X1 U13857 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U13858 ( .A1(n14561), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U13859 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10887) );
  OAI211_X1 U13860 ( .C1(n14517), .C2(n11063), .A(n10888), .B(n10887), .ZN(
        n10889) );
  AOI21_X1 U13861 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10889), .ZN(n13553) );
  INV_X1 U13862 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16488) );
  AOI22_X1 U13863 ( .A1(n14561), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10891) );
  NAND2_X1 U13864 ( .A1(n14562), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10890) );
  OAI211_X1 U13865 ( .C1(n10387), .C2(n16488), .A(n10891), .B(n10890), .ZN(
        n13089) );
  INV_X1 U13866 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U13867 ( .A1(n14561), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13868 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10892) );
  OAI211_X1 U13869 ( .C1(n14517), .C2(n11094), .A(n10893), .B(n10892), .ZN(
        n10894) );
  AOI21_X1 U13870 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10894), .ZN(n13636) );
  INV_X1 U13871 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13872 ( .A1(n10400), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U13873 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10895) );
  OAI211_X1 U13874 ( .C1(n14517), .C2(n11095), .A(n10896), .B(n10895), .ZN(
        n10897) );
  AOI21_X1 U13875 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10897), .ZN(n13820) );
  NAND2_X1 U13876 ( .A1(n13635), .A2(n10898), .ZN(n13837) );
  INV_X1 U13877 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n15845) );
  NAND2_X1 U13878 ( .A1(n14561), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10901) );
  NAND2_X1 U13879 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10900) );
  OAI211_X1 U13880 ( .C1(n14517), .C2(n15845), .A(n10901), .B(n10900), .ZN(
        n10902) );
  AOI21_X1 U13881 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10902), .ZN(n13838) );
  INV_X1 U13882 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U13883 ( .A1(n14561), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10905) );
  NAND2_X1 U13884 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10904) );
  OAI211_X1 U13885 ( .C1(n14517), .C2(n11140), .A(n10905), .B(n10904), .ZN(
        n10906) );
  AOI21_X1 U13886 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10906), .ZN(n13963) );
  INV_X1 U13887 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20062) );
  NAND2_X1 U13888 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10909) );
  AOI22_X1 U13889 ( .A1(n10400), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10908) );
  OAI211_X1 U13890 ( .C1(n14517), .C2(n20062), .A(n10909), .B(n10908), .ZN(
        n14003) );
  INV_X1 U13891 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U13892 ( .A1(n14561), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U13893 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10910) );
  OAI211_X1 U13894 ( .C1(n14517), .C2(n10912), .A(n10911), .B(n10910), .ZN(
        n10913) );
  AOI21_X1 U13895 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10913), .ZN(n14067) );
  INV_X1 U13896 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20065) );
  NAND2_X1 U13897 ( .A1(n14561), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U13898 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10914) );
  OAI211_X1 U13899 ( .C1(n14517), .C2(n20065), .A(n10915), .B(n10914), .ZN(
        n10916) );
  AOI21_X1 U13900 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10916), .ZN(n14185) );
  INV_X1 U13901 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15791) );
  AOI22_X1 U13902 ( .A1(n10400), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10918) );
  NAND2_X1 U13903 ( .A1(n14562), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10917) );
  OAI211_X1 U13904 ( .C1(n10387), .C2(n15791), .A(n10918), .B(n10917), .ZN(
        n14189) );
  INV_X1 U13905 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20068) );
  NAND2_X1 U13906 ( .A1(n14561), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U13907 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10919) );
  OAI211_X1 U13908 ( .C1(n14517), .C2(n20068), .A(n10920), .B(n10919), .ZN(
        n10921) );
  AOI21_X1 U13909 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10921), .ZN(n15446) );
  OR2_X2 U13910 ( .A1(n14188), .A2(n15446), .ZN(n15448) );
  INV_X1 U13911 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20070) );
  NAND2_X1 U13912 ( .A1(n14561), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U13913 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10922) );
  OAI211_X1 U13914 ( .C1(n14517), .C2(n20070), .A(n10923), .B(n10922), .ZN(
        n10924) );
  AOI21_X1 U13915 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10924), .ZN(n10925) );
  AND2_X1 U13916 ( .A1(n15448), .A2(n10925), .ZN(n10926) );
  NOR2_X1 U13917 ( .A1(n15427), .A2(n10926), .ZN(n19128) );
  NAND2_X1 U13918 ( .A1(n10927), .A2(n10458), .ZN(n10929) );
  NAND2_X1 U13919 ( .A1(n10929), .A2(n10928), .ZN(n10930) );
  INV_X1 U13920 ( .A(n10931), .ZN(n10932) );
  NAND2_X1 U13921 ( .A1(n10938), .A2(n10932), .ZN(n10933) );
  NOR2_X1 U13922 ( .A1(n10935), .A2(n10342), .ZN(n10936) );
  NAND2_X1 U13923 ( .A1(n10937), .A2(n14487), .ZN(n13591) );
  NAND2_X1 U13924 ( .A1(n13591), .A2(n10938), .ZN(n10940) );
  NAND2_X1 U13925 ( .A1(n10940), .A2(n10939), .ZN(n10941) );
  AND4_X1 U13926 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n13597) );
  INV_X1 U13927 ( .A(n10945), .ZN(n13494) );
  NAND2_X1 U13928 ( .A1(n13597), .A2(n13494), .ZN(n10946) );
  NAND2_X1 U13929 ( .A1(n11201), .A2(n10946), .ZN(n15812) );
  NAND3_X1 U13930 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10957) );
  NOR2_X1 U13931 ( .A1(n14218), .A2(n10957), .ZN(n14215) );
  INV_X1 U13932 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13103) );
  NAND2_X1 U13933 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19433) );
  NAND2_X1 U13934 ( .A1(n13103), .A2(n19433), .ZN(n13104) );
  NAND4_X1 U13935 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n14215), .A4(n13104), .ZN(
        n10947) );
  NAND2_X1 U13936 ( .A1(n19434), .A2(n10947), .ZN(n10951) );
  NOR2_X1 U13937 ( .A1(n13103), .A2(n19433), .ZN(n13105) );
  OR2_X1 U13938 ( .A1(n15812), .A2(n13105), .ZN(n10949) );
  INV_X1 U13939 ( .A(n11201), .ZN(n10948) );
  NOR2_X2 U13940 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20107) );
  NAND2_X1 U13941 ( .A1(n20107), .A2(n16035), .ZN(n19096) );
  NAND2_X1 U13942 ( .A1(n10948), .A2(n19178), .ZN(n19442) );
  NAND2_X1 U13943 ( .A1(n10949), .A2(n19442), .ZN(n13875) );
  INV_X1 U13944 ( .A(n13875), .ZN(n10950) );
  AND2_X1 U13945 ( .A1(n10951), .A2(n10950), .ZN(n15892) );
  NOR2_X1 U13946 ( .A1(n15867), .A2(n16488), .ZN(n16479) );
  NAND3_X1 U13947 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16479), .ZN(n15846) );
  INV_X1 U13948 ( .A(n15846), .ZN(n10952) );
  NAND2_X1 U13949 ( .A1(n10952), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11195) );
  OAI21_X1 U13950 ( .B1(n11195), .B2(n15891), .A(n19434), .ZN(n10953) );
  NAND2_X1 U13951 ( .A1(n15892), .A2(n10953), .ZN(n16460) );
  AND3_X1 U13952 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10958) );
  NAND2_X1 U13953 ( .A1(n10958), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10954) );
  AND2_X1 U13954 ( .A1(n19434), .A2(n10954), .ZN(n10955) );
  OR2_X1 U13955 ( .A1(n16460), .A2(n10955), .ZN(n15807) );
  NAND2_X1 U13956 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15782) );
  AND2_X1 U13957 ( .A1(n19434), .A2(n15782), .ZN(n10956) );
  NOR2_X1 U13958 ( .A1(n15807), .A2(n10956), .ZN(n11233) );
  OAI211_X1 U13959 ( .C1(n13877), .C2(n13105), .A(n13104), .B(n19434), .ZN(
        n16523) );
  NAND3_X1 U13960 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n16491), .ZN(n15897) );
  INV_X1 U13961 ( .A(n10958), .ZN(n10959) );
  INV_X1 U13962 ( .A(n15782), .ZN(n11197) );
  NOR2_X1 U13963 ( .A1(n19178), .A2(n20070), .ZN(n15624) );
  AOI21_X1 U13964 ( .B1(n11237), .B2(n11231), .A(n15624), .ZN(n11155) );
  NAND2_X1 U13965 ( .A1(n11251), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10962) );
  NOR2_X1 U13966 ( .A1(n10332), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10984) );
  INV_X1 U13967 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U13968 ( .A1(n14577), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10961) );
  AND2_X1 U13969 ( .A1(n10962), .A2(n10961), .ZN(n11242) );
  AND2_X2 U13970 ( .A1(n10963), .A2(n11295), .ZN(n11137) );
  NAND2_X1 U13971 ( .A1(n11137), .A2(n13242), .ZN(n10967) );
  AND2_X1 U13972 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10964) );
  NOR2_X1 U13973 ( .A1(n10984), .A2(n10964), .ZN(n10966) );
  NAND2_X1 U13974 ( .A1(n10965), .A2(n11032), .ZN(n10982) );
  NAND3_X1 U13975 ( .A1(n10967), .A2(n10966), .A3(n10982), .ZN(n13782) );
  INV_X1 U13976 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U13977 ( .A1(n14487), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10968) );
  OAI211_X1 U13978 ( .C1(n10332), .C2(n13182), .A(n10968), .B(n19854), .ZN(
        n10969) );
  INV_X1 U13979 ( .A(n10969), .ZN(n10971) );
  NAND2_X1 U13980 ( .A1(n10971), .A2(n10970), .ZN(n13781) );
  NAND2_X1 U13981 ( .A1(n13782), .A2(n13781), .ZN(n13780) );
  OR2_X1 U13982 ( .A1(n14579), .A2(n13256), .ZN(n10973) );
  AOI22_X1 U13983 ( .A1(n10984), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10972) );
  INV_X1 U13984 ( .A(n10979), .ZN(n10974) );
  XNOR2_X1 U13985 ( .A(n13780), .B(n10974), .ZN(n13779) );
  INV_X1 U13986 ( .A(n11137), .ZN(n10975) );
  OR2_X1 U13987 ( .A1(n11159), .A2(n10975), .ZN(n10978) );
  NAND2_X1 U13988 ( .A1(n13291), .A2(n10332), .ZN(n10976) );
  MUX2_X1 U13989 ( .A(n10976), .B(n20125), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10977) );
  AND2_X1 U13990 ( .A1(n10978), .A2(n10977), .ZN(n13778) );
  NAND2_X1 U13991 ( .A1(n13779), .A2(n13778), .ZN(n13777) );
  NAND2_X1 U13992 ( .A1(n10979), .A2(n13780), .ZN(n10980) );
  NAND2_X1 U13993 ( .A1(n13777), .A2(n10980), .ZN(n10988) );
  NAND2_X1 U13994 ( .A1(n11137), .A2(n10981), .ZN(n10983) );
  OAI211_X1 U13995 ( .C1(n19854), .C2(n20116), .A(n10983), .B(n10982), .ZN(
        n10987) );
  XNOR2_X1 U13996 ( .A(n10988), .B(n10987), .ZN(n13110) );
  INV_X1 U13997 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n15371) );
  OR2_X1 U13998 ( .A1(n14579), .A2(n15371), .ZN(n10986) );
  AOI22_X1 U13999 ( .A1(n14577), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10985) );
  AND2_X1 U14000 ( .A1(n10986), .A2(n10985), .ZN(n13109) );
  INV_X1 U14001 ( .A(n10987), .ZN(n10989) );
  NAND2_X1 U14002 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  OR2_X1 U14003 ( .A1(n14579), .A2(n13804), .ZN(n10996) );
  AOI22_X1 U14004 ( .A1(n11032), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n10992) );
  NAND2_X1 U14005 ( .A1(n14577), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10991) );
  AND2_X1 U14006 ( .A1(n10992), .A2(n10991), .ZN(n10995) );
  NAND2_X1 U14007 ( .A1(n11137), .A2(n10993), .ZN(n10994) );
  AOI22_X1 U14008 ( .A1(n14577), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10999) );
  NAND2_X1 U14009 ( .A1(n11137), .A2(n10997), .ZN(n10998) );
  OAI211_X1 U14010 ( .C1(n14579), .C2(n11000), .A(n10999), .B(n10998), .ZN(
        n13785) );
  INV_X1 U14011 ( .A(n13848), .ZN(n11004) );
  AOI22_X1 U14012 ( .A1(n14577), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11003) );
  NAND2_X1 U14013 ( .A1(n11137), .A2(n11001), .ZN(n11002) );
  OAI211_X1 U14014 ( .C1(n14579), .C2(n13852), .A(n11003), .B(n11002), .ZN(
        n13845) );
  NAND2_X1 U14015 ( .A1(n11004), .A2(n13845), .ZN(n13846) );
  NAND2_X1 U14016 ( .A1(n11137), .A2(n11005), .ZN(n11006) );
  OR2_X1 U14017 ( .A1(n14579), .A2(n11007), .ZN(n11009) );
  AOI22_X1 U14018 ( .A1(n14577), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U14019 ( .A1(n11009), .A2(n11008), .ZN(n14220) );
  NAND2_X1 U14020 ( .A1(n14221), .A2(n14220), .ZN(n14223) );
  NAND2_X1 U14021 ( .A1(n11137), .A2(n11010), .ZN(n11011) );
  OR2_X1 U14022 ( .A1(n14579), .A2(n11012), .ZN(n11014) );
  AOI22_X1 U14023 ( .A1(n14577), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14024 ( .A1(n14577), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14025 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14026 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14027 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14028 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11016) );
  NAND4_X1 U14029 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11027) );
  AOI22_X1 U14030 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U14031 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11020) );
  AND2_X1 U14032 ( .A1(n11021), .A2(n11020), .ZN(n11025) );
  AOI22_X1 U14033 ( .A1(n10632), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U14034 ( .A1(n11033), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U14035 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11022) );
  NAND4_X1 U14036 ( .A1(n11025), .A2(n11024), .A3(n11023), .A4(n11022), .ZN(
        n11026) );
  NAND2_X1 U14037 ( .A1(n11137), .A2(n13623), .ZN(n11028) );
  OAI211_X1 U14038 ( .C1(n14579), .C2(n11030), .A(n11029), .B(n11028), .ZN(
        n13352) );
  INV_X1 U14039 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11031) );
  OR2_X1 U14040 ( .A1(n14579), .A2(n11031), .ZN(n11048) );
  AOI22_X1 U14041 ( .A1(n14577), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11032), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U14042 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14043 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14045 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11034) );
  NAND4_X1 U14046 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n11045) );
  AOI22_X1 U14047 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U14048 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14358), .ZN(n11039) );
  NAND2_X1 U14049 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11038) );
  AND2_X1 U14050 ( .A1(n11039), .A2(n11038), .ZN(n11042) );
  AOI22_X1 U14051 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11041) );
  NAND2_X1 U14052 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11040) );
  NAND4_X1 U14053 ( .A1(n11043), .A2(n11042), .A3(n11041), .A4(n11040), .ZN(
        n11044) );
  NAND2_X1 U14054 ( .A1(n11137), .A2(n13543), .ZN(n11046) );
  AOI22_X1 U14055 ( .A1(n14577), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U14056 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14057 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14358), .ZN(n11050) );
  NAND2_X1 U14058 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11049) );
  AND2_X1 U14059 ( .A1(n11050), .A2(n11049), .ZN(n11053) );
  AOI22_X1 U14060 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U14061 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11051) );
  NAND4_X1 U14062 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(
        n11060) );
  AOI22_X1 U14063 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14064 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14065 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U14066 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14353), .B1(
        n14352), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11055) );
  NAND4_X1 U14067 ( .A1(n11058), .A2(n11057), .A3(n11056), .A4(n11055), .ZN(
        n11059) );
  NAND2_X1 U14068 ( .A1(n11137), .A2(n13551), .ZN(n11061) );
  OAI211_X1 U14069 ( .C1(n14579), .C2(n11063), .A(n11062), .B(n11061), .ZN(
        n13430) );
  NAND2_X1 U14070 ( .A1(n13429), .A2(n13430), .ZN(n13083) );
  INV_X1 U14071 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11064) );
  OR2_X1 U14072 ( .A1(n14579), .A2(n11064), .ZN(n11079) );
  AOI22_X1 U14073 ( .A1(n14577), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14074 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14075 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14076 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14077 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11065) );
  NAND4_X1 U14078 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(
        n11076) );
  AOI22_X1 U14079 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14080 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14358), .ZN(n11070) );
  NAND2_X1 U14081 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11069) );
  AND2_X1 U14082 ( .A1(n11070), .A2(n11069), .ZN(n11073) );
  AOI22_X1 U14083 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11072) );
  NAND2_X1 U14084 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11071) );
  NAND4_X1 U14085 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11075) );
  NAND2_X1 U14086 ( .A1(n11137), .A2(n13641), .ZN(n11077) );
  AOI22_X1 U14087 ( .A1(n14577), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14088 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11015), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14089 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14090 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U14091 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11080) );
  NAND4_X1 U14092 ( .A1(n11083), .A2(n11082), .A3(n11081), .A4(n11080), .ZN(
        n11091) );
  AOI22_X1 U14093 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10632), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14094 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14358), .ZN(n11085) );
  NAND2_X1 U14095 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11084) );
  AND2_X1 U14096 ( .A1(n11085), .A2(n11084), .ZN(n11088) );
  AOI22_X1 U14097 ( .A1(n10654), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U14098 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11086) );
  NAND4_X1 U14099 ( .A1(n11089), .A2(n11088), .A3(n11087), .A4(n11086), .ZN(
        n11090) );
  NAND2_X1 U14100 ( .A1(n11137), .A2(n13644), .ZN(n11092) );
  OAI211_X1 U14101 ( .C1(n14579), .C2(n11094), .A(n11093), .B(n11092), .ZN(
        n13627) );
  OR2_X1 U14102 ( .A1(n14579), .A2(n11095), .ZN(n11110) );
  AOI22_X1 U14103 ( .A1(n14577), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14104 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14105 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14106 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14107 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11096) );
  NAND4_X1 U14108 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11107) );
  AOI22_X1 U14109 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14110 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U14111 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11100) );
  AND2_X1 U14112 ( .A1(n11101), .A2(n11100), .ZN(n11104) );
  AOI22_X1 U14113 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U14114 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11102) );
  NAND4_X1 U14115 ( .A1(n11105), .A2(n11104), .A3(n11103), .A4(n11102), .ZN(
        n11106) );
  OR2_X1 U14116 ( .A1(n11107), .A2(n11106), .ZN(n13833) );
  NAND2_X1 U14117 ( .A1(n11137), .A2(n13833), .ZN(n11108) );
  AOI22_X1 U14118 ( .A1(n14577), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11124) );
  AOI22_X1 U14119 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14120 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14121 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14122 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11111) );
  NAND4_X1 U14123 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n11122) );
  AOI22_X1 U14124 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14125 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14358), .ZN(n11116) );
  NAND2_X1 U14126 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11115) );
  AND2_X1 U14127 ( .A1(n11116), .A2(n11115), .ZN(n11119) );
  AOI22_X1 U14128 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U14129 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11117) );
  NAND4_X1 U14130 ( .A1(n11120), .A2(n11119), .A3(n11118), .A4(n11117), .ZN(
        n11121) );
  OR2_X1 U14131 ( .A1(n11122), .A2(n11121), .ZN(n13834) );
  NAND2_X1 U14132 ( .A1(n11137), .A2(n13834), .ZN(n11123) );
  OAI211_X1 U14133 ( .C1(n14579), .C2(n15845), .A(n11124), .B(n11123), .ZN(
        n15844) );
  AOI22_X1 U14134 ( .A1(n14577), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14135 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14136 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14137 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n14351), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14138 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11125) );
  NAND4_X1 U14139 ( .A1(n11128), .A2(n11127), .A3(n11126), .A4(n11125), .ZN(
        n11136) );
  AOI22_X1 U14140 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11134) );
  AOI22_X1 U14141 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n14358), .ZN(n11130) );
  NAND2_X1 U14142 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11129) );
  AND2_X1 U14143 ( .A1(n11130), .A2(n11129), .ZN(n11133) );
  AOI22_X1 U14144 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U14145 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11131) );
  NAND4_X1 U14146 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(
        n11135) );
  NAND2_X1 U14147 ( .A1(n11137), .A2(n13961), .ZN(n11138) );
  OAI211_X1 U14148 ( .C1(n14579), .C2(n11140), .A(n11139), .B(n11138), .ZN(
        n15349) );
  AOI22_X1 U14149 ( .A1(n14577), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11141) );
  OAI21_X1 U14150 ( .B1(n14579), .B2(n20062), .A(n11141), .ZN(n13988) );
  NAND2_X1 U14151 ( .A1(n11251), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14152 ( .A1(n14577), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11142) );
  AND2_X1 U14153 ( .A1(n11143), .A2(n11142), .ZN(n14059) );
  NAND2_X1 U14154 ( .A1(n11251), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14155 ( .A1(n14577), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11144) );
  INV_X1 U14156 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14157 ( .A1(n14577), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11146) );
  OAI21_X1 U14158 ( .B1(n14579), .B2(n11147), .A(n11146), .ZN(n15518) );
  AOI22_X1 U14159 ( .A1(n14577), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11148) );
  OAI21_X1 U14160 ( .B1(n14579), .B2(n20068), .A(n11148), .ZN(n15509) );
  XOR2_X1 U14161 ( .A(n11242), .B(n11243), .Z(n19133) );
  NAND2_X1 U14162 ( .A1(n13587), .A2(n11149), .ZN(n13287) );
  NAND2_X1 U14163 ( .A1(n13287), .A2(n14487), .ZN(n11152) );
  NAND2_X1 U14164 ( .A1(n11151), .A2(n11150), .ZN(n13581) );
  NAND2_X1 U14165 ( .A1(n11152), .A2(n13581), .ZN(n11153) );
  NAND2_X1 U14166 ( .A1(n19133), .A2(n19436), .ZN(n11154) );
  OAI211_X1 U14167 ( .C1(n11233), .C2(n11231), .A(n11155), .B(n11154), .ZN(
        n11203) );
  INV_X1 U14168 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16507) );
  NAND2_X1 U14169 ( .A1(n13872), .A2(n16507), .ZN(n11170) );
  OR3_X1 U14170 ( .A1(n11159), .A2(n13242), .A3(n10375), .ZN(n11160) );
  NOR2_X1 U14171 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13242), .ZN(
        n11158) );
  XOR2_X1 U14172 ( .A(n11159), .B(n11158), .Z(n13258) );
  NAND2_X1 U14173 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13258), .ZN(
        n13257) );
  NAND2_X1 U14174 ( .A1(n11160), .A2(n13257), .ZN(n11164) );
  XOR2_X1 U14175 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11164), .Z(
        n13107) );
  OAI21_X1 U14176 ( .B1(n11163), .B2(n11162), .A(n11161), .ZN(n13106) );
  NAND2_X1 U14177 ( .A1(n13107), .A2(n13106), .ZN(n11166) );
  NAND2_X1 U14178 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11164), .ZN(
        n11165) );
  NAND2_X1 U14179 ( .A1(n11166), .A2(n11165), .ZN(n11167) );
  INV_X1 U14180 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16522) );
  XNOR2_X1 U14181 ( .A(n11167), .B(n16522), .ZN(n13799) );
  NAND2_X1 U14182 ( .A1(n13798), .A2(n13799), .ZN(n11169) );
  NAND2_X1 U14183 ( .A1(n11167), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11168) );
  NAND2_X1 U14184 ( .A1(n11170), .A2(n13874), .ZN(n11173) );
  INV_X1 U14185 ( .A(n13872), .ZN(n11171) );
  NAND2_X1 U14186 ( .A1(n11171), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11172) );
  NAND2_X2 U14187 ( .A1(n11173), .A2(n11172), .ZN(n16444) );
  INV_X1 U14188 ( .A(n11175), .ZN(n11174) );
  NAND2_X2 U14189 ( .A1(n16444), .A2(n16445), .ZN(n16443) );
  INV_X1 U14190 ( .A(n11184), .ZN(n11177) );
  INV_X1 U14191 ( .A(n11183), .ZN(n11176) );
  NAND2_X1 U14192 ( .A1(n11177), .A2(n11176), .ZN(n11178) );
  NAND2_X1 U14193 ( .A1(n11178), .A2(n16443), .ZN(n11179) );
  OAI21_X1 U14194 ( .B1(n16443), .B2(n11184), .A(n11179), .ZN(n11182) );
  NAND2_X1 U14195 ( .A1(n11183), .A2(n11180), .ZN(n11181) );
  NAND2_X1 U14196 ( .A1(n16443), .A2(n11176), .ZN(n11185) );
  NAND2_X1 U14197 ( .A1(n11185), .A2(n11177), .ZN(n11186) );
  XNOR2_X1 U14198 ( .A(n11187), .B(n10536), .ZN(n14233) );
  OAI21_X1 U14199 ( .B1(n11187), .B2(n10536), .A(n11188), .ZN(n11191) );
  INV_X1 U14200 ( .A(n11187), .ZN(n11190) );
  NAND2_X1 U14201 ( .A1(n11191), .A2(n11194), .ZN(n15682) );
  INV_X1 U14202 ( .A(n15682), .ZN(n11193) );
  INV_X1 U14203 ( .A(n11199), .ZN(n11198) );
  INV_X1 U14204 ( .A(n11205), .ZN(n15605) );
  OAI21_X1 U14205 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n11198), .A(
        n15605), .ZN(n15626) );
  AND2_X1 U14206 ( .A1(n11200), .A2(n13082), .ZN(n20138) );
  NOR2_X1 U14207 ( .A1(n15626), .A2(n16524), .ZN(n11202) );
  AOI211_X1 U14208 ( .C1(n19128), .C2(n19440), .A(n11203), .B(n11202), .ZN(
        n11204) );
  INV_X1 U14209 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14582) );
  AND2_X1 U14210 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15755) );
  INV_X1 U14211 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15745) );
  INV_X1 U14212 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15732) );
  NAND2_X1 U14213 ( .A1(n11333), .A2(n19438), .ZN(n11329) );
  INV_X1 U14214 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n16328) );
  NAND2_X1 U14215 ( .A1(n14561), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14216 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11207) );
  OAI211_X1 U14217 ( .C1(n14517), .C2(n16328), .A(n11208), .B(n11207), .ZN(
        n11209) );
  AOI21_X1 U14218 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11209), .ZN(n11230) );
  INV_X1 U14219 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20072) );
  NAND2_X1 U14220 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11212) );
  AOI22_X1 U14221 ( .A1(n14561), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11211) );
  OAI211_X1 U14222 ( .C1(n14517), .C2(n20072), .A(n11212), .B(n11211), .ZN(
        n15426) );
  INV_X1 U14223 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20074) );
  NAND2_X1 U14224 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11214) );
  AOI22_X1 U14225 ( .A1(n10400), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11213) );
  OAI211_X1 U14226 ( .C1(n14517), .C2(n20074), .A(n11214), .B(n11213), .ZN(
        n15340) );
  INV_X1 U14227 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20076) );
  NAND2_X1 U14228 ( .A1(n14561), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U14229 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11215) );
  OAI211_X1 U14230 ( .C1(n14517), .C2(n20076), .A(n11216), .B(n11215), .ZN(
        n11217) );
  AOI21_X1 U14231 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11217), .ZN(n15322) );
  INV_X1 U14232 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n11220) );
  NAND2_X1 U14233 ( .A1(n14561), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U14234 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11218) );
  OAI211_X1 U14235 ( .C1(n14517), .C2(n11220), .A(n11219), .B(n11218), .ZN(
        n11221) );
  AOI21_X1 U14236 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11221), .ZN(n15409) );
  INV_X1 U14237 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20079) );
  NAND2_X1 U14238 ( .A1(n14561), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U14239 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11222) );
  OAI211_X1 U14240 ( .C1(n14517), .C2(n20079), .A(n11223), .B(n11222), .ZN(
        n11224) );
  AOI21_X1 U14241 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11224), .ZN(n15310) );
  NOR2_X2 U14242 ( .A1(n15412), .A2(n15310), .ZN(n15311) );
  INV_X1 U14243 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20082) );
  NAND2_X1 U14244 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11226) );
  AOI22_X1 U14245 ( .A1(n14561), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11225) );
  OAI211_X1 U14246 ( .C1(n14517), .C2(n20082), .A(n11226), .B(n11225), .ZN(
        n15289) );
  NAND2_X1 U14247 ( .A1(n15311), .A2(n15289), .ZN(n15291) );
  INV_X1 U14248 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20083) );
  NAND2_X1 U14249 ( .A1(n14561), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U14250 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11227) );
  OAI211_X1 U14251 ( .C1(n14517), .C2(n20083), .A(n11228), .B(n11227), .ZN(
        n11229) );
  AOI21_X1 U14252 ( .B1(n11210), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11229), .ZN(n12856) );
  NOR2_X4 U14253 ( .A1(n9712), .A2(n11230), .ZN(n14560) );
  AOI21_X1 U14254 ( .B1(n11230), .B2(n9712), .A(n14560), .ZN(n15385) );
  NAND2_X1 U14255 ( .A1(n19434), .A2(n11231), .ZN(n11232) );
  NAND2_X1 U14256 ( .A1(n11233), .A2(n11232), .ZN(n15772) );
  INV_X1 U14257 ( .A(n15755), .ZN(n11238) );
  AND2_X1 U14258 ( .A1(n19434), .A2(n11238), .ZN(n11234) );
  OR2_X1 U14259 ( .A1(n15772), .A2(n11234), .ZN(n15742) );
  AND2_X1 U14260 ( .A1(n19434), .A2(n15745), .ZN(n11235) );
  NOR2_X1 U14261 ( .A1(n15742), .A2(n11235), .ZN(n15733) );
  NAND2_X1 U14262 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U14263 ( .A1(n19434), .A2(n11239), .ZN(n11236) );
  AND2_X1 U14264 ( .A1(n15733), .A2(n11236), .ZN(n15710) );
  INV_X1 U14265 ( .A(n11239), .ZN(n15720) );
  NAND2_X1 U14266 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14581) );
  NAND2_X1 U14267 ( .A1(n15705), .A2(n14581), .ZN(n11240) );
  AND2_X1 U14268 ( .A1(n15710), .A2(n11240), .ZN(n12863) );
  NOR2_X1 U14269 ( .A1(n12863), .A2(n14582), .ZN(n11263) );
  AOI22_X1 U14270 ( .A1(n14577), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11241) );
  OAI21_X1 U14271 ( .B1(n14579), .B2(n16328), .A(n11241), .ZN(n11256) );
  INV_X1 U14272 ( .A(n11256), .ZN(n11259) );
  NAND2_X1 U14273 ( .A1(n11251), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14274 ( .A1(n14577), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14275 ( .A1(n14577), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11246) );
  OAI21_X1 U14276 ( .B1(n14579), .B2(n20074), .A(n11246), .ZN(n15335) );
  NAND2_X1 U14277 ( .A1(n11251), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14278 ( .A1(n14577), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11247) );
  AND2_X1 U14279 ( .A1(n11248), .A2(n11247), .ZN(n15324) );
  NAND2_X1 U14280 ( .A1(n11251), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14281 ( .A1(n14577), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11249) );
  AND2_X1 U14282 ( .A1(n11250), .A2(n11249), .ZN(n15484) );
  NAND2_X1 U14283 ( .A1(n11251), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14284 ( .A1(n14577), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11252) );
  AND2_X1 U14285 ( .A1(n11253), .A2(n11252), .ZN(n15307) );
  AOI22_X1 U14286 ( .A1(n14577), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11254) );
  OAI21_X1 U14287 ( .B1(n14579), .B2(n20082), .A(n11254), .ZN(n15292) );
  AOI22_X1 U14288 ( .A1(n14577), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11255) );
  OAI21_X1 U14289 ( .B1(n14579), .B2(n20083), .A(n11255), .ZN(n12859) );
  INV_X1 U14290 ( .A(n11257), .ZN(n11258) );
  AOI21_X1 U14291 ( .B1(n11259), .B2(n11258), .A(n14576), .ZN(n16335) );
  INV_X1 U14292 ( .A(n16335), .ZN(n15458) );
  INV_X2 U14293 ( .A(n19178), .ZN(n19420) );
  NAND2_X1 U14294 ( .A1(n19420), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11338) );
  INV_X1 U14295 ( .A(n14581), .ZN(n11260) );
  NAND3_X1 U14296 ( .A1(n15705), .A2(n14582), .A3(n11260), .ZN(n11261) );
  OAI211_X1 U14297 ( .C1(n15458), .C2(n16526), .A(n11338), .B(n11261), .ZN(
        n11262) );
  AOI211_X1 U14298 ( .C1(n15385), .C2(n19440), .A(n11263), .B(n11262), .ZN(
        n11327) );
  INV_X1 U14299 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15979) );
  NOR2_X1 U14300 ( .A1(n11295), .A2(n15979), .ZN(n11287) );
  AOI21_X4 U14301 ( .B1(n11286), .B2(n14554), .A(n11287), .ZN(n11288) );
  NAND2_X1 U14302 ( .A1(n14552), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11289) );
  INV_X1 U14303 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11302) );
  INV_X1 U14304 ( .A(n11303), .ZN(n11265) );
  NAND2_X1 U14305 ( .A1(n14552), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11264) );
  INV_X1 U14306 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n16343) );
  NOR2_X1 U14307 ( .A1(n11295), .A2(n16343), .ZN(n11320) );
  NAND2_X1 U14308 ( .A1(n14552), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14547) );
  XNOR2_X1 U14309 ( .A(n14548), .B(n14547), .ZN(n11266) );
  INV_X1 U14310 ( .A(n11266), .ZN(n16330) );
  NAND3_X1 U14311 ( .A1(n16330), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14550), .ZN(n15543) );
  OAI21_X1 U14312 ( .B1(n11266), .B2(n10536), .A(n14582), .ZN(n14545) );
  NAND2_X1 U14313 ( .A1(n15543), .A2(n14545), .ZN(n11324) );
  NAND2_X1 U14314 ( .A1(n10536), .A2(n15782), .ZN(n11268) );
  AND4_X1 U14315 ( .A1(n16374), .A2(n16390), .A3(n11268), .A4(n11267), .ZN(
        n11270) );
  NAND2_X1 U14316 ( .A1(n19156), .A2(n15791), .ZN(n11269) );
  AND4_X1 U14317 ( .A1(n11270), .A2(n15658), .A3(n15834), .A4(n11269), .ZN(
        n11271) );
  OAI211_X1 U14318 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n19142), .A(
        n11272), .B(n11271), .ZN(n11273) );
  INV_X1 U14319 ( .A(n11273), .ZN(n11275) );
  NAND4_X1 U14320 ( .A1(n15637), .A2(n16391), .A3(n11276), .A4(n15657), .ZN(
        n11279) );
  NAND2_X1 U14321 ( .A1(n15648), .A2(n11277), .ZN(n11278) );
  NAND2_X1 U14322 ( .A1(n11281), .A2(n11280), .ZN(n11282) );
  NOR2_X1 U14323 ( .A1(n11283), .A2(n11282), .ZN(n11284) );
  AOI21_X1 U14324 ( .B1(n11287), .B2(n11286), .A(n11288), .ZN(n15978) );
  AOI21_X1 U14325 ( .B1(n15978), .B2(n14550), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15617) );
  NAND3_X1 U14326 ( .A1(n15978), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14550), .ZN(n15615) );
  INV_X1 U14327 ( .A(n11288), .ZN(n11291) );
  INV_X1 U14328 ( .A(n11289), .ZN(n11290) );
  NAND2_X1 U14329 ( .A1(n11291), .A2(n11290), .ZN(n11292) );
  NAND2_X1 U14330 ( .A1(n11298), .A2(n11292), .ZN(n15346) );
  OR2_X1 U14331 ( .A1(n15346), .A2(n10536), .ZN(n11293) );
  XNOR2_X1 U14332 ( .A(n11293), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15607) );
  INV_X1 U14333 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15757) );
  NOR3_X1 U14334 ( .A1(n15346), .A2(n10536), .A3(n15757), .ZN(n11294) );
  NOR2_X1 U14335 ( .A1(n11295), .A2(n10117), .ZN(n11297) );
  AOI21_X1 U14336 ( .B1(n11298), .B2(n11297), .A(n11296), .ZN(n11299) );
  NAND2_X1 U14337 ( .A1(n11299), .A2(n11305), .ZN(n15331) );
  INV_X1 U14338 ( .A(n15595), .ZN(n11300) );
  OR3_X1 U14339 ( .A1(n11308), .A2(n11302), .A3(n11295), .ZN(n11304) );
  NAND3_X1 U14340 ( .A1(n11305), .A2(P2_EBX_REG_25__SCAN_IN), .A3(n14552), 
        .ZN(n11306) );
  NAND2_X1 U14341 ( .A1(n11306), .A2(n14554), .ZN(n11307) );
  NAND2_X1 U14342 ( .A1(n15595), .A2(n15745), .ZN(n11309) );
  NOR2_X2 U14343 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  NAND3_X1 U14344 ( .A1(n14552), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n11314), 
        .ZN(n11315) );
  AND2_X1 U14345 ( .A1(n11319), .A2(n11315), .ZN(n15294) );
  NAND2_X1 U14346 ( .A1(n15294), .A2(n14550), .ZN(n12853) );
  AOI21_X1 U14347 ( .B1(n11320), .B2(n11319), .A(n14548), .ZN(n16342) );
  NAND2_X1 U14348 ( .A1(n16342), .A2(n14550), .ZN(n12854) );
  NAND2_X1 U14349 ( .A1(n14550), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11322) );
  NOR2_X1 U14350 ( .A1(n16350), .A2(n11322), .ZN(n15586) );
  AOI21_X1 U14351 ( .B1(n11323), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15586), .ZN(n12850) );
  XOR2_X1 U14352 ( .A(n11324), .B(n14546), .Z(n11343) );
  NAND2_X1 U14353 ( .A1(n11329), .A2(n11328), .ZN(P2_U3017) );
  AND2_X1 U14354 ( .A1(n11330), .A2(n16538), .ZN(n11331) );
  INV_X1 U14355 ( .A(n13124), .ZN(n11334) );
  NAND2_X1 U14356 ( .A1(n11334), .A2(n10458), .ZN(n19423) );
  NAND2_X1 U14357 ( .A1(n11333), .A2(n16449), .ZN(n11346) );
  NAND2_X1 U14358 ( .A1(n11334), .A2(n14487), .ZN(n19424) );
  NAND2_X1 U14359 ( .A1(n16035), .A2(n19854), .ZN(n20100) );
  INV_X1 U14360 ( .A(n20100), .ZN(n15911) );
  OR2_X1 U14361 ( .A1(n20107), .A2(n15911), .ZN(n20126) );
  NAND2_X1 U14362 ( .A1(n20126), .A2(n19097), .ZN(n11335) );
  AND2_X1 U14363 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20117) );
  INV_X1 U14364 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11340) );
  NAND2_X1 U14365 ( .A1(n19097), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13307) );
  INV_X1 U14366 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20098) );
  NAND2_X1 U14367 ( .A1(n20098), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U14368 ( .A1(n13307), .A2(n11336), .ZN(n13245) );
  INV_X1 U14369 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16399) );
  NAND2_X1 U14370 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n15259), .ZN(
        n15258) );
  INV_X1 U14371 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16381) );
  INV_X1 U14372 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15661) );
  INV_X1 U14373 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15642) );
  NAND2_X1 U14374 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n15264), .ZN(
        n15263) );
  INV_X1 U14375 ( .A(n15263), .ZN(n11337) );
  INV_X1 U14376 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16349) );
  AOI21_X1 U14377 ( .B1(n11340), .B2(n15244), .A(n13071), .ZN(n16326) );
  NAND2_X1 U14378 ( .A1(n16440), .A2(n16326), .ZN(n11339) );
  OAI211_X1 U14379 ( .C1(n16453), .C2(n11340), .A(n11339), .B(n11338), .ZN(
        n11341) );
  AOI21_X1 U14380 ( .B1(n15385), .B2(n19428), .A(n11341), .ZN(n11342) );
  OAI21_X1 U14381 ( .B1(n11343), .B2(n19424), .A(n11342), .ZN(n11344) );
  NAND2_X1 U14382 ( .A1(n11346), .A2(n11345), .ZN(P2_U2985) );
  INV_X1 U14383 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11357) );
  NAND2_X4 U14384 ( .A1(n13660), .A2(n11350), .ZN(n11703) );
  INV_X1 U14385 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11349) );
  INV_X1 U14386 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11347) );
  OAI22_X1 U14387 ( .A1(n11349), .A2(n11348), .B1(n11731), .B2(n11511), .ZN(
        n11352) );
  AND2_X2 U14388 ( .A1(n13669), .A2(n11360), .ZN(n11539) );
  INV_X1 U14389 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11981) );
  INV_X1 U14390 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13942) );
  OAI22_X1 U14391 ( .A1(n11552), .A2(n11981), .B1(n11569), .B2(n13942), .ZN(
        n11351) );
  AOI211_X1 U14392 ( .C1(n12124), .C2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n11352), .B(n11351), .ZN(n11356) );
  INV_X1 U14393 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14394 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n9685), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11355) );
  OAI211_X1 U14395 ( .C1(n11357), .C2(n11703), .A(n11356), .B(n11355), .ZN(
        n11366) );
  INV_X2 U14396 ( .A(n11576), .ZN(n12146) );
  AOI22_X1 U14397 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14398 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12511), .B1(
        n12145), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14399 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n9687), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11362) );
  AND2_X2 U14400 ( .A1(n13669), .A2(n13656), .ZN(n11530) );
  INV_X2 U14401 ( .A(n11561), .ZN(n12415) );
  AOI22_X1 U14402 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11361) );
  NAND4_X1 U14403 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11365) );
  NOR2_X1 U14404 ( .A1(n11366), .A2(n11365), .ZN(n12251) );
  INV_X1 U14405 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11372) );
  INV_X1 U14406 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11537) );
  INV_X1 U14407 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13938) );
  OAI22_X1 U14408 ( .A1(n11731), .A2(n11537), .B1(n11569), .B2(n13938), .ZN(
        n11369) );
  INV_X1 U14409 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12110) );
  INV_X1 U14410 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11367) );
  OAI22_X1 U14411 ( .A1(n9674), .A2(n12110), .B1(n12503), .B2(n11367), .ZN(
        n11368) );
  AOI211_X1 U14412 ( .C1(n12124), .C2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11369), .B(n11368), .ZN(n11371) );
  AOI22_X1 U14413 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11370) );
  OAI211_X1 U14414 ( .C1(n11703), .C2(n11372), .A(n11371), .B(n11370), .ZN(
        n11378) );
  AOI22_X1 U14415 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14416 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11375) );
  INV_X2 U14417 ( .A(n11552), .ZN(n12510) );
  AOI22_X1 U14418 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14419 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14420 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  NOR2_X1 U14421 ( .A1(n11378), .A2(n11377), .ZN(n12230) );
  INV_X1 U14422 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11384) );
  INV_X1 U14423 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13934) );
  INV_X1 U14424 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11379) );
  OAI22_X1 U14425 ( .A1(n11348), .A2(n13934), .B1(n11569), .B2(n11379), .ZN(
        n11381) );
  INV_X1 U14426 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12046) );
  INV_X1 U14427 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12502) );
  OAI22_X1 U14428 ( .A1(n9674), .A2(n12046), .B1(n9684), .B2(n12502), .ZN(
        n11380) );
  AOI211_X1 U14429 ( .C1(n12124), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11381), .B(n11380), .ZN(n11383) );
  AOI22_X1 U14430 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9685), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11382) );
  OAI211_X1 U14431 ( .C1(n11690), .C2(n11384), .A(n11383), .B(n11382), .ZN(
        n11390) );
  AOI22_X1 U14432 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14433 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14434 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11386) );
  AOI22_X1 U14435 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11385) );
  NAND4_X1 U14436 ( .A1(n11388), .A2(n11387), .A3(n11386), .A4(n11385), .ZN(
        n11389) );
  NOR2_X1 U14437 ( .A1(n11390), .A2(n11389), .ZN(n12209) );
  INV_X1 U14438 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11397) );
  INV_X1 U14439 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11391) );
  OAI22_X1 U14440 ( .A1(n11348), .A2(n11391), .B1(n11731), .B2(n11587), .ZN(
        n11394) );
  INV_X1 U14441 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11392) );
  INV_X1 U14442 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20391) );
  OAI22_X1 U14443 ( .A1(n11576), .A2(n11392), .B1(n11569), .B2(n20391), .ZN(
        n11393) );
  AOI211_X1 U14444 ( .C1(n12124), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n11394), .B(n11393), .ZN(n11396) );
  AOI22_X1 U14445 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9685), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11395) );
  OAI211_X1 U14446 ( .C1(n11703), .C2(n11397), .A(n11396), .B(n11395), .ZN(
        n11403) );
  AOI22_X1 U14447 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14448 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14449 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14450 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14451 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11402) );
  NOR2_X1 U14452 ( .A1(n11403), .A2(n11402), .ZN(n12210) );
  NOR2_X1 U14453 ( .A1(n12209), .A2(n12210), .ZN(n12221) );
  INV_X1 U14454 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11406) );
  NAND2_X1 U14455 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11405) );
  NAND2_X1 U14456 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11404) );
  OAI211_X1 U14457 ( .C1(n11703), .C2(n11406), .A(n11405), .B(n11404), .ZN(
        n11407) );
  INV_X1 U14458 ( .A(n11407), .ZN(n11411) );
  AOI22_X1 U14459 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11410) );
  INV_X1 U14460 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20395) );
  AOI22_X1 U14461 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11409) );
  NAND2_X1 U14462 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11408) );
  NAND4_X1 U14463 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11417) );
  AOI22_X1 U14464 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14465 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14466 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14467 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11412) );
  NAND4_X1 U14468 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11416) );
  OR2_X1 U14469 ( .A1(n11417), .A2(n11416), .ZN(n12219) );
  NAND2_X1 U14470 ( .A1(n12221), .A2(n12219), .ZN(n12231) );
  NOR2_X1 U14471 ( .A1(n12230), .A2(n12231), .ZN(n12243) );
  INV_X1 U14472 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11420) );
  NAND2_X1 U14473 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11419) );
  NAND2_X1 U14474 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11418) );
  OAI211_X1 U14475 ( .C1(n11703), .C2(n11420), .A(n11419), .B(n11418), .ZN(
        n11421) );
  INV_X1 U14476 ( .A(n11421), .ZN(n11425) );
  AOI22_X1 U14477 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14478 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U14479 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11422) );
  NAND4_X1 U14480 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11431) );
  AOI22_X1 U14481 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14482 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14483 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14484 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11426) );
  NAND4_X1 U14485 ( .A1(n11429), .A2(n11428), .A3(n11427), .A4(n11426), .ZN(
        n11430) );
  OR2_X1 U14486 ( .A1(n11431), .A2(n11430), .ZN(n12241) );
  NAND2_X1 U14487 ( .A1(n12243), .A2(n12241), .ZN(n12250) );
  NOR2_X1 U14488 ( .A1(n12251), .A2(n12250), .ZN(n12432) );
  INV_X1 U14489 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11434) );
  NAND2_X1 U14490 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11433) );
  NAND2_X1 U14491 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11432) );
  OAI211_X1 U14492 ( .C1(n11690), .C2(n11434), .A(n11433), .B(n11432), .ZN(
        n11435) );
  INV_X1 U14493 ( .A(n11435), .ZN(n11439) );
  AOI22_X1 U14494 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11438) );
  INV_X1 U14495 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20399) );
  AOI22_X1 U14496 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11437) );
  NAND2_X1 U14497 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11436) );
  NAND4_X1 U14498 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(
        n11445) );
  AOI22_X1 U14499 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14500 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14501 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14502 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11440) );
  NAND4_X1 U14503 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11444) );
  OR2_X1 U14504 ( .A1(n11445), .A2(n11444), .ZN(n12431) );
  XNOR2_X1 U14505 ( .A(n12432), .B(n12431), .ZN(n11519) );
  INV_X1 U14506 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U14507 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11447) );
  NAND2_X1 U14508 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11446) );
  OAI211_X1 U14509 ( .C1(n11703), .C2(n11448), .A(n11447), .B(n11446), .ZN(
        n11449) );
  INV_X1 U14510 ( .A(n11449), .ZN(n11453) );
  NAND2_X1 U14511 ( .A1(n11553), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11450) );
  AOI22_X1 U14512 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14513 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n9673), .ZN(n11454) );
  NAND2_X1 U14514 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11463) );
  NAND2_X1 U14515 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U14516 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11461) );
  NAND2_X1 U14517 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11460) );
  NAND4_X1 U14518 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11466) );
  INV_X1 U14519 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11464) );
  NOR2_X1 U14520 ( .A1(n12198), .A2(n11464), .ZN(n11465) );
  NAND2_X1 U14521 ( .A1(n9683), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11469) );
  NAND2_X1 U14522 ( .A1(n9677), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11468) );
  NAND2_X1 U14523 ( .A1(n11562), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11467) );
  NAND3_X1 U14524 ( .A1(n11469), .A2(n11468), .A3(n11467), .ZN(n11470) );
  NAND2_X1 U14525 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11474) );
  NAND2_X1 U14526 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11473) );
  NAND2_X1 U14527 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11472) );
  NAND2_X1 U14528 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11471) );
  INV_X1 U14529 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U14530 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11475) );
  OAI21_X1 U14531 ( .B1(n11703), .B2(n11476), .A(n11475), .ZN(n11478) );
  INV_X1 U14532 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11485) );
  NAND2_X1 U14533 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11484) );
  NAND2_X1 U14534 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11483) );
  OAI211_X1 U14535 ( .C1(n11703), .C2(n11485), .A(n11484), .B(n11483), .ZN(
        n11486) );
  INV_X1 U14536 ( .A(n11486), .ZN(n11490) );
  AOI22_X1 U14537 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14538 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U14539 ( .A1(n11553), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11487) );
  AOI22_X1 U14540 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9683), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14541 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11559), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14542 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11560), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14543 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11562), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U14544 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14545 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U14546 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11498) );
  NAND2_X1 U14547 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11497) );
  NAND4_X1 U14548 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11503) );
  NAND2_X1 U14549 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11505) );
  NAND2_X1 U14550 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11504) );
  NAND2_X1 U14551 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U14552 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14553 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14554 ( .A1(n11562), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11506) );
  NAND2_X1 U14555 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11510) );
  NAND3_X1 U14556 ( .A1(n11627), .A2(n11567), .A3(n11682), .ZN(n11614) );
  NOR2_X2 U14557 ( .A1(n11567), .A2(n11760), .ZN(n11777) );
  NAND2_X1 U14558 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11516) );
  NAND2_X1 U14559 ( .A1(n12434), .A2(n11516), .ZN(n11517) );
  AOI21_X1 U14560 ( .B1(n12524), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11517), .ZN(
        n11518) );
  OAI21_X1 U14561 ( .B1(n11519), .B2(n12437), .A(n11518), .ZN(n11526) );
  INV_X1 U14562 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14710) );
  INV_X1 U14563 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14686) );
  INV_X1 U14564 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12235) );
  INV_X1 U14565 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14646) );
  XNOR2_X1 U14566 ( .A(n12439), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12320) );
  NAND2_X1 U14567 ( .A1(n12320), .A2(n12523), .ZN(n11525) );
  NAND2_X1 U14568 ( .A1(n11526), .A2(n11525), .ZN(n12445) );
  NAND2_X1 U14569 ( .A1(n11627), .A2(n13013), .ZN(n11528) );
  AND2_X2 U14570 ( .A1(n11527), .A2(n11567), .ZN(n11629) );
  AOI22_X1 U14571 ( .A1(n9691), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14572 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11562), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14573 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11560), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14574 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11559), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14575 ( .A1(n9692), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11536) );
  OAI211_X1 U14576 ( .C1(n11703), .C2(n11537), .A(n11536), .B(n11535), .ZN(
        n11538) );
  INV_X1 U14577 ( .A(n11538), .ZN(n11543) );
  AOI22_X1 U14578 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14579 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U14580 ( .A1(n11553), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11540) );
  INV_X1 U14581 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U14582 ( .A1(n11596), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14583 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11546) );
  OAI211_X1 U14584 ( .C1(n11703), .C2(n11548), .A(n11547), .B(n11546), .ZN(
        n11549) );
  INV_X1 U14585 ( .A(n11549), .ZN(n11557) );
  AOI22_X1 U14586 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14587 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11555) );
  NAND2_X1 U14588 ( .A1(n11553), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11554) );
  AOI22_X1 U14589 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11559), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14590 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11560), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14591 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9683), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14592 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11562), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14593 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11574) );
  NAND2_X1 U14594 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U14595 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11572) );
  NAND2_X1 U14596 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11580) );
  NAND2_X1 U14597 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11579) );
  NAND2_X1 U14598 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11578) );
  NAND2_X1 U14599 ( .A1(n11562), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11577) );
  NAND2_X1 U14600 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11584) );
  NAND2_X1 U14601 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11583) );
  NAND2_X1 U14602 ( .A1(n11560), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11582) );
  NAND2_X1 U14603 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11581) );
  NAND2_X1 U14604 ( .A1(n9692), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11586) );
  NAND2_X1 U14605 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11585) );
  OAI211_X1 U14606 ( .C1(n11703), .C2(n11587), .A(n11586), .B(n11585), .ZN(
        n11588) );
  INV_X1 U14607 ( .A(n11588), .ZN(n11589) );
  NAND4_X4 U14608 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n13900) );
  NAND2_X1 U14609 ( .A1(n11539), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11595) );
  NAND2_X1 U14610 ( .A1(n11530), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11594) );
  NAND2_X1 U14611 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11593) );
  INV_X1 U14612 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U14613 ( .A1(n9692), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U14614 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11597) );
  OAI211_X1 U14615 ( .C1(n11703), .C2(n11599), .A(n11598), .B(n11597), .ZN(
        n11600) );
  INV_X1 U14616 ( .A(n11600), .ZN(n11602) );
  NAND2_X1 U14617 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14618 ( .A1(n11559), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14619 ( .A1(n11545), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U14620 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11610) );
  NAND2_X1 U14621 ( .A1(n11558), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14622 ( .A1(n9671), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14623 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11607) );
  NAND4_X4 U14624 ( .A1(n9714), .A2(n9637), .A3(n11612), .A4(n11611), .ZN(
        n13326) );
  NAND2_X1 U14625 ( .A1(n11615), .A2(n11624), .ZN(n11616) );
  INV_X1 U14626 ( .A(n11619), .ZN(n13018) );
  XNOR2_X1 U14627 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12993) );
  NAND2_X1 U14628 ( .A1(n11624), .A2(n11567), .ZN(n12997) );
  NOR2_X1 U14629 ( .A1(n12997), .A2(n13357), .ZN(n11625) );
  INV_X1 U14630 ( .A(n11628), .ZN(n11641) );
  NAND3_X1 U14631 ( .A1(n11641), .A2(n11629), .A3(n13013), .ZN(n13004) );
  NAND2_X1 U14632 ( .A1(n13004), .A2(n15194), .ZN(n11650) );
  INV_X1 U14633 ( .A(n13023), .ZN(n11645) );
  NAND2_X1 U14634 ( .A1(n12927), .A2(n12457), .ZN(n13017) );
  NAND2_X1 U14635 ( .A1(n11635), .A2(n13326), .ZN(n20955) );
  NAND2_X1 U14636 ( .A1(n13900), .A2(n13749), .ZN(n11631) );
  NAND2_X1 U14637 ( .A1(n11634), .A2(n11635), .ZN(n11636) );
  NAND2_X1 U14638 ( .A1(n20937), .A2(n20865), .ZN(n12321) );
  NAND2_X1 U14639 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11660) );
  OAI21_X1 U14640 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11660), .ZN(n20683) );
  OR2_X1 U14641 ( .A1(n16015), .A2(n20686), .ZN(n11655) );
  OAI21_X1 U14642 ( .B1(n12321), .B2(n20683), .A(n11655), .ZN(n11638) );
  INV_X1 U14643 ( .A(n11638), .ZN(n11639) );
  MUX2_X1 U14644 ( .A(n12321), .B(n16015), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11640) );
  OAI21_X2 U14645 ( .B1(n11662), .B2(n11353), .A(n11640), .ZN(n11687) );
  INV_X1 U14646 ( .A(n12874), .ZN(n12899) );
  AOI21_X1 U14647 ( .B1(n11641), .B2(n11630), .A(n12899), .ZN(n11642) );
  OR2_X1 U14648 ( .A1(n13900), .A2(n13326), .ZN(n14603) );
  MUX2_X1 U14649 ( .A(n11634), .B(n11642), .S(n14603), .Z(n11652) );
  NAND2_X1 U14650 ( .A1(n20937), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20165) );
  INV_X1 U14651 ( .A(n20165), .ZN(n11644) );
  AND2_X1 U14652 ( .A1(n20955), .A2(n11644), .ZN(n11646) );
  OR2_X1 U14653 ( .A1(n11645), .A2(n11624), .ZN(n13030) );
  OAI211_X1 U14654 ( .C1(n11629), .C2(n11643), .A(n11646), .B(n13030), .ZN(
        n11647) );
  INV_X1 U14655 ( .A(n11647), .ZN(n11648) );
  OAI211_X1 U14656 ( .C1(n11650), .C2(n9654), .A(n11649), .B(n11648), .ZN(
        n11651) );
  INV_X1 U14657 ( .A(n11686), .ZN(n11653) );
  NAND2_X1 U14658 ( .A1(n11687), .A2(n11653), .ZN(n11748) );
  INV_X1 U14659 ( .A(n11748), .ZN(n11654) );
  INV_X1 U14660 ( .A(n11655), .ZN(n11657) );
  INV_X1 U14661 ( .A(n11660), .ZN(n11659) );
  NAND2_X1 U14662 ( .A1(n11659), .A2(n12290), .ZN(n20728) );
  NAND2_X1 U14663 ( .A1(n11660), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11661) );
  INV_X1 U14664 ( .A(n16015), .ZN(n11663) );
  NAND2_X1 U14665 ( .A1(n11663), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11664) );
  INV_X1 U14666 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11670) );
  NAND2_X1 U14667 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11669) );
  NAND2_X1 U14668 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11668) );
  OAI211_X1 U14669 ( .C1(n11690), .C2(n11670), .A(n11669), .B(n11668), .ZN(
        n11671) );
  INV_X1 U14670 ( .A(n11671), .ZN(n11675) );
  AOI22_X1 U14671 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14672 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11673) );
  NAND2_X1 U14673 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11672) );
  NAND4_X1 U14674 ( .A1(n11675), .A2(n11674), .A3(n11673), .A4(n11672), .ZN(
        n11681) );
  AOI22_X1 U14675 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14676 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14677 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14678 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11676) );
  NAND4_X1 U14679 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11680) );
  NOR2_X1 U14680 ( .A1(n11681), .A2(n11680), .ZN(n12331) );
  OAI22_X1 U14681 ( .A1(n13657), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12331), 
        .B2(n11793), .ZN(n11685) );
  OAI22_X1 U14682 ( .A1(n12301), .A2(n13938), .B1(n11792), .B2(n12331), .ZN(
        n11683) );
  INV_X1 U14683 ( .A(n11683), .ZN(n11684) );
  XNOR2_X1 U14684 ( .A(n11685), .B(n11684), .ZN(n11757) );
  INV_X1 U14685 ( .A(n11757), .ZN(n11756) );
  INV_X1 U14686 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U14687 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11689) );
  NAND2_X1 U14688 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11688) );
  OAI211_X1 U14689 ( .C1(n11690), .C2(n12501), .A(n11689), .B(n11688), .ZN(
        n11691) );
  INV_X1 U14690 ( .A(n11691), .ZN(n11696) );
  INV_X1 U14691 ( .A(n11731), .ZN(n11692) );
  AOI22_X1 U14692 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14693 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U14694 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11693) );
  NAND4_X1 U14695 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11702) );
  AOI22_X1 U14696 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14697 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14698 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14699 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11697) );
  NAND4_X1 U14700 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11701) );
  INV_X1 U14701 ( .A(n12389), .ZN(n11720) );
  INV_X1 U14702 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11706) );
  NAND2_X1 U14703 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U14704 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11704) );
  OAI211_X1 U14705 ( .C1(n11690), .C2(n11706), .A(n11705), .B(n11704), .ZN(
        n11707) );
  INV_X1 U14706 ( .A(n11707), .ZN(n11712) );
  INV_X1 U14707 ( .A(n11731), .ZN(n11708) );
  AOI22_X1 U14708 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14709 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U14710 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11709) );
  NAND4_X1 U14711 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11719) );
  AOI22_X1 U14712 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14713 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14714 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14715 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11714) );
  NAND4_X1 U14716 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11718) );
  XNOR2_X1 U14717 ( .A(n11720), .B(n12342), .ZN(n11721) );
  NAND2_X1 U14718 ( .A1(n11721), .A2(n12325), .ZN(n11722) );
  AOI21_X1 U14719 ( .B1(n13013), .B2(n12389), .A(n20865), .ZN(n11725) );
  NAND2_X1 U14720 ( .A1(n11635), .A2(n12342), .ZN(n11724) );
  NAND2_X1 U14721 ( .A1(n12325), .A2(n12389), .ZN(n11726) );
  INV_X1 U14722 ( .A(n11792), .ZN(n11742) );
  INV_X1 U14723 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U14724 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11728) );
  NAND2_X1 U14725 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11727) );
  OAI211_X1 U14726 ( .C1(n11690), .C2(n11729), .A(n11728), .B(n11727), .ZN(
        n11730) );
  INV_X1 U14727 ( .A(n11730), .ZN(n11735) );
  AOI22_X1 U14728 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14729 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U14730 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11732) );
  NAND4_X1 U14731 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11741) );
  AOI22_X1 U14732 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14733 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14734 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14735 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11736) );
  NAND4_X1 U14736 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n11740) );
  NAND2_X1 U14737 ( .A1(n11742), .A2(n12341), .ZN(n11744) );
  OR2_X1 U14738 ( .A1(n12301), .A2(n20395), .ZN(n11743) );
  OAI211_X1 U14739 ( .C1(n11793), .C2(n12389), .A(n11744), .B(n11743), .ZN(
        n11745) );
  NAND2_X1 U14740 ( .A1(n11746), .A2(n11745), .ZN(n11747) );
  NAND2_X1 U14741 ( .A1(n11754), .A2(n11747), .ZN(n11768) );
  NAND2_X1 U14742 ( .A1(n11749), .A2(n11748), .ZN(n13712) );
  NAND2_X1 U14743 ( .A1(n11750), .A2(n13712), .ZN(n13702) );
  NAND2_X1 U14744 ( .A1(n11751), .A2(n20865), .ZN(n11753) );
  NAND2_X1 U14745 ( .A1(n12325), .A2(n12341), .ZN(n11752) );
  OAI21_X1 U14746 ( .B1(n11768), .B2(n12339), .A(n11754), .ZN(n11755) );
  INV_X1 U14747 ( .A(n11755), .ZN(n11758) );
  NAND2_X1 U14748 ( .A1(n11756), .A2(n11755), .ZN(n11759) );
  NAND2_X1 U14749 ( .A1(n11758), .A2(n11757), .ZN(n11832) );
  NAND2_X1 U14750 ( .A1(n12330), .A2(n12052), .ZN(n11761) );
  NOR2_X1 U14751 ( .A1(n12997), .A2(n11760), .ZN(n11776) );
  NAND2_X1 U14752 ( .A1(n11776), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11767) );
  INV_X1 U14753 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11764) );
  OAI21_X1 U14754 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11762), .ZN(n20348) );
  NAND2_X1 U14755 ( .A1(n13889), .A2(n20348), .ZN(n11763) );
  OAI21_X1 U14756 ( .B1(n11764), .B2(n12097), .A(n11763), .ZN(n11765) );
  AOI21_X1 U14757 ( .B1(n12524), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11765), .ZN(
        n11766) );
  AND2_X1 U14758 ( .A1(n11767), .A2(n11766), .ZN(n11782) );
  XNOR2_X1 U14759 ( .A(n11768), .B(n12339), .ZN(n13688) );
  NAND2_X1 U14760 ( .A1(n13688), .A2(n12052), .ZN(n11772) );
  NAND2_X1 U14761 ( .A1(n11776), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11770) );
  AOI22_X1 U14762 ( .A1(n12524), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11760), .ZN(n11769) );
  AND2_X1 U14763 ( .A1(n11770), .A2(n11769), .ZN(n11771) );
  NAND2_X1 U14764 ( .A1(n11772), .A2(n11771), .ZN(n13455) );
  AOI21_X1 U14765 ( .B1(n20431), .B2(n9669), .A(n11760), .ZN(n13427) );
  INV_X1 U14766 ( .A(n11776), .ZN(n11838) );
  NAND2_X1 U14767 ( .A1(n11777), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11779) );
  NAND2_X1 U14768 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11778) );
  OAI211_X1 U14769 ( .C1(n11838), .C2(n11353), .A(n11779), .B(n11778), .ZN(
        n11780) );
  AOI21_X1 U14770 ( .B1(n11775), .B2(n12052), .A(n11780), .ZN(n13428) );
  MUX2_X1 U14771 ( .A(n13427), .B(n12523), .S(n13428), .Z(n13456) );
  NAND2_X1 U14772 ( .A1(n13755), .A2(n13453), .ZN(n11785) );
  INV_X1 U14773 ( .A(n11782), .ZN(n11783) );
  NAND2_X1 U14774 ( .A1(n11781), .A2(n11783), .ZN(n11784) );
  INV_X1 U14775 ( .A(n11832), .ZN(n11809) );
  NAND3_X1 U14776 ( .A1(n20727), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20590) );
  INV_X1 U14777 ( .A(n20590), .ZN(n20595) );
  NAND2_X1 U14778 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20595), .ZN(
        n20588) );
  NAND2_X1 U14779 ( .A1(n20727), .A2(n20588), .ZN(n11788) );
  NOR3_X1 U14780 ( .A1(n20727), .A2(n12290), .A3(n20686), .ZN(n20811) );
  NAND2_X1 U14781 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20811), .ZN(
        n20798) );
  NAND2_X1 U14782 ( .A1(n11788), .A2(n20798), .ZN(n15214) );
  OAI22_X1 U14783 ( .A1(n12321), .A2(n15214), .B1(n16015), .B2(n20727), .ZN(
        n11789) );
  INV_X1 U14784 ( .A(n11789), .ZN(n11790) );
  INV_X1 U14785 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U14786 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U14787 ( .A1(n12192), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11794) );
  OAI211_X1 U14788 ( .C1(n11690), .C2(n11796), .A(n11795), .B(n11794), .ZN(
        n11797) );
  INV_X1 U14789 ( .A(n11797), .ZN(n11801) );
  AOI22_X1 U14790 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U14791 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U14792 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11798) );
  NAND4_X1 U14793 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11807) );
  AOI22_X1 U14794 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U14795 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9685), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U14796 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14797 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11802) );
  NAND4_X1 U14798 ( .A1(n11805), .A2(n11804), .A3(n11803), .A4(n11802), .ZN(
        n11806) );
  AOI22_X1 U14799 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12307), .B1(
        n12280), .B2(n12355), .ZN(n11808) );
  INV_X1 U14800 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11812) );
  NAND2_X1 U14801 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11811) );
  NAND2_X1 U14802 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11810) );
  OAI211_X1 U14803 ( .C1(n11690), .C2(n11812), .A(n11811), .B(n11810), .ZN(
        n11813) );
  INV_X1 U14804 ( .A(n11813), .ZN(n11817) );
  AOI22_X1 U14805 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9690), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14806 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12510), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11815) );
  NAND2_X1 U14807 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11814) );
  NAND4_X1 U14808 ( .A1(n11817), .A2(n11816), .A3(n11815), .A4(n11814), .ZN(
        n11823) );
  AOI22_X1 U14809 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14810 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14811 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14812 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11818) );
  NAND4_X1 U14813 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11822) );
  NAND2_X1 U14814 ( .A1(n12280), .A2(n12364), .ZN(n11825) );
  OR2_X1 U14815 ( .A1(n12301), .A2(n13942), .ZN(n11824) );
  NAND2_X1 U14816 ( .A1(n11825), .A2(n11824), .ZN(n11843) );
  NAND2_X1 U14817 ( .A1(n12354), .A2(n12052), .ZN(n11831) );
  INV_X1 U14818 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U14819 ( .A1(n12524), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11827) );
  INV_X1 U14820 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21022) );
  OAI21_X1 U14821 ( .B1(n21022), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11760), .ZN(n11826) );
  OAI211_X1 U14822 ( .C1(n11838), .C2(n13652), .A(n11827), .B(n11826), .ZN(
        n11829) );
  AOI21_X1 U14823 ( .B1(n20235), .B2(n11834), .A(n11861), .ZN(n20230) );
  NAND2_X1 U14824 ( .A1(n20230), .A2(n12523), .ZN(n11828) );
  NAND2_X1 U14825 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  INV_X1 U14826 ( .A(n13691), .ZN(n13692) );
  NAND2_X1 U14827 ( .A1(n11832), .A2(n13692), .ZN(n11833) );
  INV_X1 U14828 ( .A(n12052), .ZN(n11997) );
  OAI21_X1 U14829 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11835), .A(
        n11834), .ZN(n20337) );
  AOI22_X1 U14830 ( .A1(n12523), .A2(n20337), .B1(n14531), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U14831 ( .A1(n12524), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11836) );
  OAI211_X1 U14832 ( .C1(n11838), .C2(n11350), .A(n11837), .B(n11836), .ZN(
        n11839) );
  INV_X1 U14833 ( .A(n11839), .ZN(n11840) );
  INV_X1 U14834 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11846) );
  NAND2_X1 U14835 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11845) );
  NAND2_X1 U14836 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11844) );
  OAI211_X1 U14837 ( .C1(n11690), .C2(n11846), .A(n11845), .B(n11844), .ZN(
        n11847) );
  INV_X1 U14838 ( .A(n11847), .ZN(n11851) );
  AOI22_X1 U14839 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14840 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U14841 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11848) );
  NAND4_X1 U14842 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(
        n11857) );
  AOI22_X1 U14843 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14844 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14845 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14846 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11852) );
  NAND4_X1 U14847 ( .A1(n11855), .A2(n11854), .A3(n11853), .A4(n11852), .ZN(
        n11856) );
  NAND2_X1 U14848 ( .A1(n12280), .A2(n12373), .ZN(n11859) );
  OR2_X1 U14849 ( .A1(n12301), .A2(n20399), .ZN(n11858) );
  NAND2_X1 U14850 ( .A1(n11859), .A2(n11858), .ZN(n11866) );
  XNOR2_X1 U14851 ( .A(n11865), .B(n11866), .ZN(n12362) );
  INV_X1 U14852 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11863) );
  OAI21_X1 U14853 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11861), .A(
        n11860), .ZN(n20226) );
  AOI22_X1 U14854 ( .A1(n12523), .A2(n20226), .B1(n14531), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11862) );
  OAI21_X1 U14855 ( .B1(n11899), .B2(n11863), .A(n11862), .ZN(n11864) );
  INV_X1 U14856 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U14857 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U14858 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11869) );
  OAI211_X1 U14859 ( .C1(n11690), .C2(n12417), .A(n11870), .B(n11869), .ZN(
        n11871) );
  INV_X1 U14860 ( .A(n11871), .ZN(n11875) );
  AOI22_X1 U14861 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14862 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11873) );
  NAND2_X1 U14863 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11872) );
  NAND4_X1 U14864 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11881) );
  AOI22_X1 U14865 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9687), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14866 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14867 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14868 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U14869 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11880) );
  NAND2_X1 U14870 ( .A1(n12280), .A2(n12377), .ZN(n11883) );
  INV_X1 U14871 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20405) );
  OR2_X1 U14872 ( .A1(n12301), .A2(n20405), .ZN(n11882) );
  INV_X1 U14873 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11886) );
  OAI21_X1 U14874 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11884), .A(
        n11894), .ZN(n20207) );
  NAND2_X1 U14875 ( .A1(n20207), .A2(n12523), .ZN(n11885) );
  OAI21_X1 U14876 ( .B1(n11886), .B2(n12097), .A(n11885), .ZN(n11887) );
  AOI21_X1 U14877 ( .B1(n12524), .B2(P1_EAX_REG_6__SCAN_IN), .A(n11887), .ZN(
        n11888) );
  NAND2_X1 U14878 ( .A1(n12280), .A2(n12389), .ZN(n11892) );
  OAI21_X1 U14879 ( .B1(n13934), .B2(n12301), .A(n11892), .ZN(n11893) );
  NAND2_X1 U14880 ( .A1(n12384), .A2(n12052), .ZN(n11902) );
  INV_X1 U14881 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11898) );
  INV_X1 U14882 ( .A(n11894), .ZN(n11896) );
  INV_X1 U14883 ( .A(n11917), .ZN(n11895) );
  OAI21_X1 U14884 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11896), .A(
        n11895), .ZN(n20195) );
  AOI22_X1 U14885 ( .A1(n13889), .A2(n20195), .B1(n14531), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11897) );
  OAI21_X1 U14886 ( .B1(n11899), .B2(n11898), .A(n11897), .ZN(n11900) );
  AOI22_X1 U14887 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14888 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14889 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14890 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11903) );
  NAND4_X1 U14891 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11916) );
  INV_X1 U14892 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11909) );
  NAND2_X1 U14893 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11908) );
  NAND2_X1 U14894 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11907) );
  OAI211_X1 U14895 ( .C1(n11690), .C2(n11909), .A(n11908), .B(n11907), .ZN(
        n11910) );
  INV_X1 U14896 ( .A(n11910), .ZN(n11914) );
  AOI22_X1 U14897 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14898 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U14899 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11911) );
  NAND4_X1 U14900 ( .A1(n11914), .A2(n11913), .A3(n11912), .A4(n11911), .ZN(
        n11915) );
  OAI21_X1 U14901 ( .B1(n11916), .B2(n11915), .A(n12052), .ZN(n11920) );
  XOR2_X1 U14902 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11917), .Z(n20185) );
  INV_X1 U14903 ( .A(n20185), .ZN(n14041) );
  AOI22_X1 U14904 ( .A1(n14531), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13889), .B2(n14041), .ZN(n11919) );
  NAND2_X1 U14905 ( .A1(n11777), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U14906 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14907 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U14908 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U14909 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11922) );
  NAND4_X1 U14910 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11935) );
  INV_X1 U14911 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U14912 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U14913 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11926) );
  OAI211_X1 U14914 ( .C1(n11690), .C2(n11928), .A(n11927), .B(n11926), .ZN(
        n11929) );
  INV_X1 U14915 ( .A(n11929), .ZN(n11933) );
  AOI22_X1 U14916 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14917 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11931) );
  NAND2_X1 U14918 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11930) );
  NAND4_X1 U14919 ( .A1(n11933), .A2(n11932), .A3(n11931), .A4(n11930), .ZN(
        n11934) );
  OAI21_X1 U14920 ( .B1(n11935), .B2(n11934), .A(n12052), .ZN(n11940) );
  INV_X1 U14921 ( .A(n11936), .ZN(n11937) );
  XNOR2_X1 U14922 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11937), .ZN(
        n15049) );
  AOI22_X1 U14923 ( .A1(n13889), .A2(n15049), .B1(n14531), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U14924 ( .A1(n11777), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11938) );
  XOR2_X1 U14925 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n11941), .Z(
        n16153) );
  INV_X1 U14926 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11944) );
  NAND2_X1 U14927 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11943) );
  NAND2_X1 U14928 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11942) );
  OAI211_X1 U14929 ( .C1(n11690), .C2(n11944), .A(n11943), .B(n11942), .ZN(
        n11945) );
  INV_X1 U14930 ( .A(n11945), .ZN(n11949) );
  AOI22_X1 U14931 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14932 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11947) );
  NAND2_X1 U14933 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11946) );
  NAND4_X1 U14934 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n11955) );
  AOI22_X1 U14935 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U14936 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14937 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U14938 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11950) );
  NAND4_X1 U14939 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n11954) );
  OR2_X1 U14940 ( .A1(n11955), .A2(n11954), .ZN(n11956) );
  AOI22_X1 U14941 ( .A1(n12052), .A2(n11956), .B1(n14531), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U14942 ( .A1(n11777), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11957) );
  OAI211_X1 U14943 ( .C1(n16153), .C2(n12434), .A(n11958), .B(n11957), .ZN(
        n14024) );
  XNOR2_X1 U14944 ( .A(n11959), .B(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15041) );
  NOR2_X1 U14945 ( .A1(n12097), .A2(n15038), .ZN(n11960) );
  AOI21_X1 U14946 ( .B1(n12524), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11960), .ZN(
        n11961) );
  OAI21_X1 U14947 ( .B1(n15041), .B2(n12434), .A(n11961), .ZN(n11977) );
  INV_X1 U14948 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U14949 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U14950 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11962) );
  OAI211_X1 U14951 ( .C1(n11690), .C2(n11964), .A(n11963), .B(n11962), .ZN(
        n11965) );
  INV_X1 U14952 ( .A(n11965), .ZN(n11969) );
  AOI22_X1 U14953 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U14954 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U14955 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11966) );
  NAND4_X1 U14956 ( .A1(n11969), .A2(n11968), .A3(n11967), .A4(n11966), .ZN(
        n11975) );
  AOI22_X1 U14957 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12145), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U14958 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9685), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U14959 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U14960 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11970) );
  NAND4_X1 U14961 ( .A1(n11973), .A2(n11972), .A3(n11971), .A4(n11970), .ZN(
        n11974) );
  OR2_X1 U14962 ( .A1(n11975), .A2(n11974), .ZN(n11976) );
  AND2_X1 U14963 ( .A1(n12052), .A2(n11976), .ZN(n14778) );
  INV_X1 U14964 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U14965 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11980) );
  NAND2_X1 U14966 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11979) );
  OAI211_X1 U14967 ( .C1(n11690), .C2(n11981), .A(n11980), .B(n11979), .ZN(
        n11982) );
  INV_X1 U14968 ( .A(n11982), .ZN(n11986) );
  AOI22_X1 U14969 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n9690), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U14970 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12510), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U14971 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11983) );
  NAND4_X1 U14972 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n11983), .ZN(
        n11992) );
  AOI22_X1 U14973 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U14974 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12511), .B1(
        n12145), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U14975 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U14976 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n9687), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U14977 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11991) );
  NOR2_X1 U14978 ( .A1(n11992), .A2(n11991), .ZN(n11996) );
  XNOR2_X1 U14979 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11993), .ZN(
        n16092) );
  AOI22_X1 U14980 ( .A1(n13889), .A2(n16092), .B1(n14531), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11995) );
  NAND2_X1 U14981 ( .A1(n11777), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11994) );
  OAI211_X1 U14982 ( .C1(n11997), .C2(n11996), .A(n11995), .B(n11994), .ZN(
        n14836) );
  XOR2_X1 U14983 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11998), .Z(
        n16083) );
  INV_X1 U14984 ( .A(n16083), .ZN(n15022) );
  AOI22_X1 U14985 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U14986 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12415), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U14987 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U14988 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U14989 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12012) );
  INV_X1 U14990 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12005) );
  NAND2_X1 U14991 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12004) );
  NAND2_X1 U14992 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12003) );
  OAI211_X1 U14993 ( .C1(n11690), .C2(n12005), .A(n12004), .B(n12003), .ZN(
        n12006) );
  INV_X1 U14994 ( .A(n12006), .ZN(n12010) );
  AOI22_X1 U14995 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U14996 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U14997 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12007) );
  NAND4_X1 U14998 ( .A1(n12010), .A2(n12009), .A3(n12008), .A4(n12007), .ZN(
        n12011) );
  OAI21_X1 U14999 ( .B1(n12012), .B2(n12011), .A(n12052), .ZN(n12015) );
  NAND2_X1 U15000 ( .A1(n11777), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U15001 ( .A1(n14531), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12013) );
  NAND3_X1 U15002 ( .A1(n12015), .A2(n12014), .A3(n12013), .ZN(n12016) );
  AOI21_X1 U15003 ( .B1(n15022), .B2(n12523), .A(n12016), .ZN(n14894) );
  INV_X1 U15004 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12017) );
  XNOR2_X1 U15005 ( .A(n12018), .B(n12017), .ZN(n16066) );
  INV_X1 U15006 ( .A(n16066), .ZN(n15014) );
  AOI22_X1 U15007 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15008 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15009 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15010 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U15011 ( .A1(n12022), .A2(n12021), .A3(n12020), .A4(n12019), .ZN(
        n12032) );
  INV_X1 U15012 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12025) );
  NAND2_X1 U15013 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12024) );
  NAND2_X1 U15014 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12023) );
  OAI211_X1 U15015 ( .C1(n11690), .C2(n12025), .A(n12024), .B(n12023), .ZN(
        n12026) );
  INV_X1 U15016 ( .A(n12026), .ZN(n12030) );
  AOI22_X1 U15017 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15018 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12028) );
  NAND2_X1 U15019 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12027) );
  NAND4_X1 U15020 ( .A1(n12030), .A2(n12029), .A3(n12028), .A4(n12027), .ZN(
        n12031) );
  OAI21_X1 U15021 ( .B1(n12032), .B2(n12031), .A(n12052), .ZN(n12035) );
  NAND2_X1 U15022 ( .A1(n11777), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U15023 ( .A1(n14531), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12033) );
  NAND3_X1 U15024 ( .A1(n12035), .A2(n12034), .A3(n12033), .ZN(n12036) );
  AOI21_X1 U15025 ( .B1(n15014), .B2(n12523), .A(n12036), .ZN(n14830) );
  XOR2_X1 U15026 ( .A(n16057), .B(n12039), .Z(n16141) );
  INV_X1 U15027 ( .A(n16141), .ZN(n12059) );
  AOI22_X1 U15028 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15029 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15030 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15031 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12040) );
  NAND4_X1 U15032 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(
        n12054) );
  NAND2_X1 U15033 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12045) );
  NAND2_X1 U15034 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12044) );
  OAI211_X1 U15035 ( .C1(n11690), .C2(n12046), .A(n12045), .B(n12044), .ZN(
        n12047) );
  INV_X1 U15036 ( .A(n12047), .ZN(n12051) );
  AOI22_X1 U15037 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15038 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U15039 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12048) );
  NAND4_X1 U15040 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12053) );
  OAI21_X1 U15041 ( .B1(n12054), .B2(n12053), .A(n12052), .ZN(n12057) );
  NAND2_X1 U15042 ( .A1(n11777), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U15043 ( .A1(n14531), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12055) );
  NAND3_X1 U15044 ( .A1(n12057), .A2(n12056), .A3(n12055), .ZN(n12058) );
  AOI21_X1 U15045 ( .B1(n12059), .B2(n12523), .A(n12058), .ZN(n14823) );
  INV_X1 U15046 ( .A(n14823), .ZN(n12060) );
  INV_X1 U15047 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12061) );
  XNOR2_X1 U15048 ( .A(n12062), .B(n12061), .ZN(n15002) );
  NAND2_X1 U15049 ( .A1(n15002), .A2(n12523), .ZN(n12081) );
  INV_X1 U15050 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12065) );
  NAND2_X1 U15051 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U15052 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12063) );
  OAI211_X1 U15053 ( .C1(n11703), .C2(n12065), .A(n12064), .B(n12063), .ZN(
        n12066) );
  INV_X1 U15054 ( .A(n12066), .ZN(n12070) );
  AOI22_X1 U15055 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15056 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12068) );
  NAND2_X1 U15057 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12067) );
  NAND4_X1 U15058 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12076) );
  AOI22_X1 U15059 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15060 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15061 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15062 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12071) );
  NAND4_X1 U15063 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n12071), .ZN(
        n12075) );
  NOR2_X1 U15064 ( .A1(n12076), .A2(n12075), .ZN(n12079) );
  AOI21_X1 U15065 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n12061), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12077) );
  AOI21_X1 U15066 ( .B1(n12524), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12077), .ZN(
        n12078) );
  OAI21_X1 U15067 ( .B1(n12437), .B2(n12079), .A(n12078), .ZN(n12080) );
  NAND2_X1 U15068 ( .A1(n12081), .A2(n12080), .ZN(n14767) );
  INV_X1 U15069 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12084) );
  NAND2_X1 U15070 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12083) );
  NAND2_X1 U15071 ( .A1(n11491), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12082) );
  OAI211_X1 U15072 ( .C1(n11690), .C2(n12084), .A(n12083), .B(n12082), .ZN(
        n12085) );
  INV_X1 U15073 ( .A(n12085), .ZN(n12089) );
  AOI22_X1 U15074 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15075 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12087) );
  NAND2_X1 U15076 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12086) );
  NAND4_X1 U15077 ( .A1(n12089), .A2(n12088), .A3(n12087), .A4(n12086), .ZN(
        n12095) );
  AOI22_X1 U15078 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15079 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15080 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9671), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15081 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12090) );
  NAND4_X1 U15082 ( .A1(n12093), .A2(n12092), .A3(n12091), .A4(n12090), .ZN(
        n12094) );
  NOR2_X1 U15083 ( .A1(n12095), .A2(n12094), .ZN(n12100) );
  INV_X1 U15084 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16045) );
  XOR2_X1 U15085 ( .A(n16045), .B(n12096), .Z(n16130) );
  OAI22_X1 U15086 ( .A1(n16130), .A2(n12434), .B1(n12097), .B2(n16045), .ZN(
        n12098) );
  AOI21_X1 U15087 ( .B1(n12524), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12098), .ZN(
        n12099) );
  OAI21_X1 U15088 ( .B1(n12437), .B2(n12100), .A(n12099), .ZN(n16047) );
  NAND2_X1 U15089 ( .A1(n12437), .A2(n12434), .ZN(n12203) );
  AOI22_X1 U15090 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9687), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15091 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15092 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15093 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15094 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12113) );
  AOI22_X1 U15095 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15096 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12107) );
  AOI21_X1 U15097 ( .B1(n12510), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n12523), .ZN(n12106) );
  NAND2_X1 U15098 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12105) );
  NAND4_X1 U15099 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        n12112) );
  INV_X1 U15100 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12109) );
  OAI22_X1 U15101 ( .A1(n11690), .A2(n12110), .B1(n12198), .B2(n12109), .ZN(
        n12111) );
  OR3_X1 U15102 ( .A1(n12113), .A2(n12112), .A3(n12111), .ZN(n12114) );
  NAND2_X1 U15103 ( .A1(n12203), .A2(n12114), .ZN(n12116) );
  AOI22_X1 U15104 ( .A1(n11777), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11760), .ZN(n12115) );
  NAND2_X1 U15105 ( .A1(n12116), .A2(n12115), .ZN(n12119) );
  XNOR2_X1 U15106 ( .A(n12117), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14995) );
  NAND2_X1 U15107 ( .A1(n14995), .A2(n12523), .ZN(n12118) );
  INV_X1 U15108 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12122) );
  NAND2_X1 U15109 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U15110 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12120) );
  OAI211_X1 U15111 ( .C1(n11690), .C2(n12122), .A(n12121), .B(n12120), .ZN(
        n12123) );
  INV_X1 U15112 ( .A(n12123), .ZN(n12128) );
  AOI22_X1 U15113 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15114 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12126) );
  NAND2_X1 U15115 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12125) );
  NAND4_X1 U15116 ( .A1(n12128), .A2(n12127), .A3(n12126), .A4(n12125), .ZN(
        n12134) );
  AOI22_X1 U15117 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15118 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15119 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15120 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12129) );
  NAND4_X1 U15121 ( .A1(n12132), .A2(n12131), .A3(n12130), .A4(n12129), .ZN(
        n12133) );
  NOR2_X1 U15122 ( .A1(n12134), .A2(n12133), .ZN(n12138) );
  OAI21_X1 U15123 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n21022), .A(
        n11760), .ZN(n12135) );
  INV_X1 U15124 ( .A(n12135), .ZN(n12136) );
  AOI21_X1 U15125 ( .B1(n12524), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12136), .ZN(
        n12137) );
  OAI21_X1 U15126 ( .B1(n12437), .B2(n12138), .A(n12137), .ZN(n12144) );
  INV_X1 U15127 ( .A(n12139), .ZN(n12141) );
  INV_X1 U15128 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U15129 ( .A1(n12141), .A2(n12140), .ZN(n12142) );
  AND2_X1 U15130 ( .A1(n12161), .A2(n12142), .ZN(n14984) );
  NAND2_X1 U15131 ( .A1(n14984), .A2(n12523), .ZN(n12143) );
  NAND2_X1 U15132 ( .A1(n12144), .A2(n12143), .ZN(n14734) );
  AOI22_X1 U15133 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12145), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15134 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15135 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9685), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15136 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15137 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12159) );
  AOI22_X1 U15138 ( .A1(n12173), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15139 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11491), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12153) );
  AOI21_X1 U15140 ( .B1(n12510), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12523), .ZN(n12152) );
  NAND2_X1 U15141 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12151) );
  NAND4_X1 U15142 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12158) );
  INV_X1 U15143 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12156) );
  INV_X1 U15144 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12155) );
  OAI22_X1 U15145 ( .A1(n12156), .A2(n11690), .B1(n12198), .B2(n12155), .ZN(
        n12157) );
  OR3_X1 U15146 ( .A1(n12159), .A2(n12158), .A3(n12157), .ZN(n12160) );
  NAND2_X1 U15147 ( .A1(n12203), .A2(n12160), .ZN(n12164) );
  AOI22_X1 U15148 ( .A1(n11777), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11760), .ZN(n12163) );
  XNOR2_X1 U15149 ( .A(n12161), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14979) );
  INV_X1 U15150 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12167) );
  NAND2_X1 U15151 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15152 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12165) );
  OAI211_X1 U15153 ( .C1(n11703), .C2(n12167), .A(n12166), .B(n12165), .ZN(
        n12168) );
  INV_X1 U15154 ( .A(n12168), .ZN(n12172) );
  AOI22_X1 U15155 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15156 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12170) );
  NAND2_X1 U15157 ( .A1(n12124), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12169) );
  NAND4_X1 U15158 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12179) );
  AOI22_X1 U15159 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12415), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15160 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15161 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15162 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12174) );
  NAND4_X1 U15163 ( .A1(n12177), .A2(n12176), .A3(n12175), .A4(n12174), .ZN(
        n12178) );
  NOR2_X1 U15164 ( .A1(n12179), .A2(n12178), .ZN(n12183) );
  NAND2_X1 U15165 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12180) );
  NAND2_X1 U15166 ( .A1(n12434), .A2(n12180), .ZN(n12181) );
  AOI21_X1 U15167 ( .B1(n12524), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12181), .ZN(
        n12182) );
  OAI21_X1 U15168 ( .B1(n12437), .B2(n12183), .A(n12182), .ZN(n12187) );
  NAND2_X1 U15169 ( .A1(n12184), .A2(n14710), .ZN(n12185) );
  AND2_X1 U15170 ( .A1(n12206), .A2(n12185), .ZN(n14709) );
  NAND2_X1 U15171 ( .A1(n14709), .A2(n12523), .ZN(n12186) );
  AOI22_X1 U15172 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15173 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12190) );
  AOI21_X1 U15174 ( .B1(n11708), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n12523), .ZN(n12189) );
  NAND2_X1 U15175 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12188) );
  NAND4_X1 U15176 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12201) );
  AOI22_X1 U15177 ( .A1(n12415), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9685), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15178 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15179 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12173), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15180 ( .A1(n12145), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12193) );
  NAND4_X1 U15181 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12200) );
  INV_X1 U15182 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12418) );
  INV_X1 U15183 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12197) );
  OAI22_X1 U15184 ( .A1(n11690), .A2(n12418), .B1(n12198), .B2(n12197), .ZN(
        n12199) );
  OR3_X1 U15185 ( .A1(n12201), .A2(n12200), .A3(n12199), .ZN(n12202) );
  NAND2_X1 U15186 ( .A1(n12203), .A2(n12202), .ZN(n12205) );
  AOI22_X1 U15187 ( .A1(n11777), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11760), .ZN(n12204) );
  NAND2_X1 U15188 ( .A1(n12205), .A2(n12204), .ZN(n12208) );
  XNOR2_X1 U15189 ( .A(n12206), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14952) );
  NAND2_X1 U15190 ( .A1(n14952), .A2(n12523), .ZN(n12207) );
  NAND2_X1 U15191 ( .A1(n12208), .A2(n12207), .ZN(n14696) );
  XNOR2_X1 U15192 ( .A(n12210), .B(n12209), .ZN(n12214) );
  NAND2_X1 U15193 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12211) );
  NAND2_X1 U15194 ( .A1(n12434), .A2(n12211), .ZN(n12212) );
  AOI21_X1 U15195 ( .B1(n12524), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12212), .ZN(
        n12213) );
  OAI21_X1 U15196 ( .B1(n12214), .B2(n12437), .A(n12213), .ZN(n12218) );
  NAND2_X1 U15197 ( .A1(n12215), .A2(n14686), .ZN(n12216) );
  AND2_X1 U15198 ( .A1(n12227), .A2(n12216), .ZN(n14685) );
  NAND2_X1 U15199 ( .A1(n14685), .A2(n12523), .ZN(n12217) );
  NAND2_X1 U15200 ( .A1(n12218), .A2(n12217), .ZN(n14684) );
  INV_X1 U15201 ( .A(n12219), .ZN(n12220) );
  XNOR2_X1 U15202 ( .A(n12221), .B(n12220), .ZN(n12222) );
  INV_X1 U15203 ( .A(n12437), .ZN(n12520) );
  NAND2_X1 U15204 ( .A1(n12222), .A2(n12520), .ZN(n12226) );
  NAND2_X1 U15205 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12223) );
  NAND2_X1 U15206 ( .A1(n12434), .A2(n12223), .ZN(n12224) );
  AOI21_X1 U15207 ( .B1(n12524), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12224), .ZN(
        n12225) );
  NAND2_X1 U15208 ( .A1(n12226), .A2(n12225), .ZN(n12229) );
  XNOR2_X1 U15209 ( .A(n12227), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14937) );
  NAND2_X1 U15210 ( .A1(n14937), .A2(n12523), .ZN(n12228) );
  NAND2_X1 U15211 ( .A1(n12229), .A2(n12228), .ZN(n14673) );
  XNOR2_X1 U15212 ( .A(n12231), .B(n12230), .ZN(n12234) );
  AOI21_X1 U15213 ( .B1(n12235), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12232) );
  AOI21_X1 U15214 ( .B1(n12524), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12232), .ZN(
        n12233) );
  OAI21_X1 U15215 ( .B1(n12234), .B2(n12437), .A(n12233), .ZN(n12239) );
  NAND2_X1 U15216 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  NAND2_X1 U15217 ( .A1(n12246), .A2(n12237), .ZN(n14929) );
  NAND2_X1 U15218 ( .A1(n12239), .A2(n12238), .ZN(n14660) );
  INV_X1 U15219 ( .A(n12241), .ZN(n12242) );
  XNOR2_X1 U15220 ( .A(n12243), .B(n12242), .ZN(n12244) );
  NAND2_X1 U15221 ( .A1(n12244), .A2(n12520), .ZN(n12249) );
  AOI21_X1 U15222 ( .B1(n14646), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12245) );
  AOI21_X1 U15223 ( .B1(n11777), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12245), .ZN(
        n12248) );
  XNOR2_X1 U15224 ( .A(n12246), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14913) );
  XNOR2_X1 U15225 ( .A(n12251), .B(n12250), .ZN(n12255) );
  NAND2_X1 U15226 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12252) );
  NAND2_X1 U15227 ( .A1(n12434), .A2(n12252), .ZN(n12253) );
  AOI21_X1 U15228 ( .B1(n12524), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12253), .ZN(
        n12254) );
  OAI21_X1 U15229 ( .B1(n12255), .B2(n12437), .A(n12254), .ZN(n12260) );
  INV_X1 U15230 ( .A(n12256), .ZN(n12257) );
  INV_X1 U15231 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14632) );
  NAND2_X1 U15232 ( .A1(n12257), .A2(n14632), .ZN(n12258) );
  NAND2_X1 U15233 ( .A1(n12439), .A2(n12258), .ZN(n14909) );
  INV_X1 U15234 ( .A(n12448), .ZN(n12261) );
  AOI21_X1 U15235 ( .B1(n12445), .B2(n14630), .A(n12261), .ZN(n14253) );
  NOR2_X1 U15236 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13651), .ZN(n20952) );
  AND2_X1 U15237 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20952), .ZN(n12262) );
  NAND2_X1 U15238 ( .A1(n15194), .A2(n11635), .ZN(n12263) );
  NAND2_X1 U15239 ( .A1(n10027), .A2(n12263), .ZN(n13005) );
  OR2_X1 U15240 ( .A1(n13005), .A2(n11619), .ZN(n14595) );
  NAND2_X1 U15241 ( .A1(n13326), .A2(n13357), .ZN(n12338) );
  NAND2_X1 U15242 ( .A1(n20686), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12265) );
  NAND2_X1 U15243 ( .A1(n11347), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12264) );
  NAND2_X1 U15244 ( .A1(n12265), .A2(n12264), .ZN(n12275) );
  NAND2_X1 U15245 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20647), .ZN(
        n12281) );
  NAND2_X1 U15246 ( .A1(n12277), .A2(n12265), .ZN(n12292) );
  NAND2_X1 U15247 ( .A1(n12292), .A2(n12266), .ZN(n12268) );
  NAND2_X1 U15248 ( .A1(n12290), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12267) );
  NAND2_X1 U15249 ( .A1(n12268), .A2(n12267), .ZN(n12274) );
  XNOR2_X1 U15250 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U15251 ( .A1(n12274), .A2(n12273), .ZN(n12270) );
  NAND2_X1 U15252 ( .A1(n20727), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U15253 ( .A1(n12270), .A2(n12269), .ZN(n12305) );
  NOR2_X1 U15254 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13652), .ZN(
        n12271) );
  NAND2_X1 U15255 ( .A1(n12303), .A2(n12450), .ZN(n12316) );
  NAND2_X1 U15256 ( .A1(n12450), .A2(n12280), .ZN(n12314) );
  XNOR2_X1 U15257 ( .A(n12274), .B(n12273), .ZN(n12452) );
  NAND2_X1 U15258 ( .A1(n12275), .A2(n12281), .ZN(n12276) );
  NAND2_X1 U15259 ( .A1(n12277), .A2(n12276), .ZN(n12451) );
  AOI22_X1 U15260 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12278), .B1(n12280), 
        .B2(n13326), .ZN(n12289) );
  INV_X1 U15261 ( .A(n12289), .ZN(n12279) );
  NOR2_X1 U15262 ( .A1(n12451), .A2(n12279), .ZN(n12287) );
  OAI21_X1 U15263 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20647), .A(
        n12281), .ZN(n12283) );
  NOR2_X1 U15264 ( .A1(n12298), .A2(n12283), .ZN(n12286) );
  NAND2_X1 U15265 ( .A1(n12278), .A2(n13900), .ZN(n12282) );
  NAND2_X1 U15266 ( .A1(n12282), .A2(n9654), .ZN(n12297) );
  INV_X1 U15267 ( .A(n12283), .ZN(n12284) );
  OAI211_X1 U15268 ( .C1(n11635), .C2(n11619), .A(n12297), .B(n12284), .ZN(
        n12285) );
  OAI21_X1 U15269 ( .B1(n12303), .B2(n12286), .A(n12285), .ZN(n12288) );
  NAND2_X1 U15270 ( .A1(n12287), .A2(n12288), .ZN(n12296) );
  NAND2_X1 U15271 ( .A1(n12289), .A2(n13326), .ZN(n12309) );
  OAI211_X1 U15272 ( .C1(n12289), .C2(n12288), .A(n12451), .B(n12309), .ZN(
        n12295) );
  MUX2_X1 U15273 ( .A(n12290), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12291) );
  XNOR2_X1 U15274 ( .A(n12292), .B(n12291), .ZN(n12453) );
  NAND2_X1 U15275 ( .A1(n12307), .A2(n12453), .ZN(n12293) );
  OAI211_X1 U15276 ( .C1(n12298), .C2(n12453), .A(n12293), .B(n12297), .ZN(
        n12294) );
  NAND3_X1 U15277 ( .A1(n12296), .A2(n12295), .A3(n12294), .ZN(n12300) );
  AOI22_X1 U15278 ( .A1(n12301), .A2(n12452), .B1(n12300), .B2(n12299), .ZN(
        n12302) );
  AOI21_X1 U15279 ( .B1(n12303), .B2(n12452), .A(n12302), .ZN(n12311) );
  NOR2_X1 U15280 ( .A1(n12305), .A2(n12304), .ZN(n12454) );
  INV_X1 U15281 ( .A(n12454), .ZN(n12306) );
  NOR2_X1 U15282 ( .A1(n12307), .A2(n12306), .ZN(n12310) );
  NAND2_X1 U15283 ( .A1(n12307), .A2(n12454), .ZN(n12308) );
  OAI22_X1 U15284 ( .A1(n12311), .A2(n12310), .B1(n12309), .B2(n12308), .ZN(
        n12312) );
  AOI21_X1 U15285 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20865), .A(
        n12312), .ZN(n12313) );
  NAND2_X1 U15286 ( .A1(n12314), .A2(n12313), .ZN(n12315) );
  NAND2_X1 U15287 ( .A1(n20802), .A2(n12321), .ZN(n20950) );
  NAND2_X1 U15288 ( .A1(n20950), .A2(n20865), .ZN(n12317) );
  NAND2_X1 U15289 ( .A1(n20865), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U15290 ( .A1(n21022), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12318) );
  AND2_X1 U15291 ( .A1(n12319), .A2(n12318), .ZN(n13517) );
  INV_X1 U15292 ( .A(n12320), .ZN(n14622) );
  INV_X1 U15293 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21134) );
  NOR2_X1 U15294 ( .A1(n20351), .A2(n21134), .ZN(n15091) );
  AOI21_X1 U15295 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15091), .ZN(n12322) );
  OAI21_X1 U15296 ( .B1(n20349), .B2(n14622), .A(n12322), .ZN(n12323) );
  INV_X1 U15297 ( .A(n12338), .ZN(n12383) );
  AND3_X1 U15298 ( .A1(n12383), .A2(n12325), .A3(n12389), .ZN(n12326) );
  NAND2_X1 U15299 ( .A1(n12341), .A2(n12342), .ZN(n12340) );
  NAND2_X1 U15300 ( .A1(n12340), .A2(n12331), .ZN(n12356) );
  INV_X1 U15301 ( .A(n12355), .ZN(n12327) );
  XNOR2_X1 U15302 ( .A(n12356), .B(n12327), .ZN(n12328) );
  INV_X1 U15303 ( .A(n11643), .ZN(n12390) );
  NAND2_X1 U15304 ( .A1(n12328), .A2(n12390), .ZN(n12329) );
  INV_X1 U15305 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20364) );
  XNOR2_X1 U15306 ( .A(n12352), .B(n20364), .ZN(n20332) );
  XNOR2_X1 U15307 ( .A(n12340), .B(n12331), .ZN(n12333) );
  NAND2_X1 U15308 ( .A1(n11635), .A2(n11630), .ZN(n12335) );
  INV_X1 U15309 ( .A(n12335), .ZN(n12332) );
  AOI21_X1 U15310 ( .B1(n12333), .B2(n12390), .A(n12332), .ZN(n12334) );
  OAI21_X1 U15311 ( .B1(n11643), .B2(n12342), .A(n12335), .ZN(n12336) );
  INV_X1 U15312 ( .A(n12336), .ZN(n12337) );
  OAI21_X1 U15313 ( .B1(n20431), .B2(n12338), .A(n12337), .ZN(n13513) );
  NAND2_X1 U15314 ( .A1(n13513), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13512) );
  OAI21_X1 U15315 ( .B1(n12342), .B2(n12341), .A(n12340), .ZN(n12343) );
  INV_X1 U15316 ( .A(n12457), .ZN(n12866) );
  OAI211_X1 U15317 ( .C1(n12343), .C2(n11643), .A(n12866), .B(n13357), .ZN(
        n12344) );
  INV_X1 U15318 ( .A(n12344), .ZN(n12345) );
  NAND2_X1 U15319 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  XNOR2_X1 U15320 ( .A(n13512), .B(n12347), .ZN(n13828) );
  NAND2_X1 U15321 ( .A1(n13828), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15166) );
  INV_X1 U15322 ( .A(n12347), .ZN(n12348) );
  OR2_X1 U15323 ( .A1(n13512), .A2(n12348), .ZN(n12349) );
  NAND2_X1 U15324 ( .A1(n15166), .A2(n12349), .ZN(n12350) );
  INV_X1 U15325 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20380) );
  XNOR2_X1 U15326 ( .A(n12350), .B(n20380), .ZN(n20341) );
  NAND2_X1 U15327 ( .A1(n20340), .A2(n20341), .ZN(n20339) );
  NAND2_X1 U15328 ( .A1(n12350), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12351) );
  NAND2_X1 U15329 ( .A1(n20339), .A2(n12351), .ZN(n20331) );
  NAND2_X1 U15330 ( .A1(n20332), .A2(n20331), .ZN(n20330) );
  NAND2_X1 U15331 ( .A1(n12352), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12353) );
  NAND2_X1 U15332 ( .A1(n20330), .A2(n12353), .ZN(n13955) );
  NAND2_X1 U15333 ( .A1(n12354), .A2(n12383), .ZN(n12359) );
  NAND2_X1 U15334 ( .A1(n12356), .A2(n12355), .ZN(n12363) );
  XNOR2_X1 U15335 ( .A(n12363), .B(n12364), .ZN(n12357) );
  NAND2_X1 U15336 ( .A1(n12357), .A2(n12390), .ZN(n12358) );
  NAND2_X1 U15337 ( .A1(n12359), .A2(n12358), .ZN(n12360) );
  INV_X1 U15338 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20359) );
  XNOR2_X1 U15339 ( .A(n12360), .B(n20359), .ZN(n13954) );
  NAND2_X1 U15340 ( .A1(n13955), .A2(n13954), .ZN(n13953) );
  NAND2_X1 U15341 ( .A1(n12360), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12361) );
  NAND2_X1 U15342 ( .A1(n13953), .A2(n12361), .ZN(n16173) );
  NAND2_X1 U15343 ( .A1(n12362), .A2(n12383), .ZN(n12368) );
  INV_X1 U15344 ( .A(n12363), .ZN(n12365) );
  NAND2_X1 U15345 ( .A1(n12365), .A2(n12364), .ZN(n12372) );
  XNOR2_X1 U15346 ( .A(n12372), .B(n12373), .ZN(n12366) );
  NAND2_X1 U15347 ( .A1(n12366), .A2(n12390), .ZN(n12367) );
  NAND2_X1 U15348 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  INV_X1 U15349 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16309) );
  XNOR2_X1 U15350 ( .A(n12369), .B(n16309), .ZN(n16172) );
  NAND2_X1 U15351 ( .A1(n16173), .A2(n16172), .ZN(n16171) );
  NAND2_X1 U15352 ( .A1(n12369), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12370) );
  INV_X1 U15353 ( .A(n12372), .ZN(n12374) );
  NAND2_X1 U15354 ( .A1(n12374), .A2(n12373), .ZN(n12376) );
  INV_X1 U15355 ( .A(n12376), .ZN(n12378) );
  INV_X1 U15356 ( .A(n12377), .ZN(n12375) );
  OR2_X1 U15357 ( .A1(n12376), .A2(n12375), .ZN(n12392) );
  OAI211_X1 U15358 ( .C1(n12378), .C2(n12377), .A(n12392), .B(n12390), .ZN(
        n12379) );
  NAND2_X1 U15359 ( .A1(n12380), .A2(n12379), .ZN(n12381) );
  INV_X1 U15360 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14033) );
  XNOR2_X1 U15361 ( .A(n12381), .B(n14033), .ZN(n16165) );
  NAND2_X1 U15362 ( .A1(n12381), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12382) );
  NAND2_X1 U15363 ( .A1(n12384), .A2(n12383), .ZN(n12387) );
  XNOR2_X1 U15364 ( .A(n12392), .B(n12389), .ZN(n12385) );
  NAND2_X1 U15365 ( .A1(n12385), .A2(n12390), .ZN(n12386) );
  NAND2_X1 U15366 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  AND2_X1 U15367 ( .A1(n12388), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16157) );
  NAND2_X1 U15368 ( .A1(n12390), .A2(n12389), .ZN(n12391) );
  OR2_X1 U15369 ( .A1(n12392), .A2(n12391), .ZN(n12393) );
  NAND2_X1 U15370 ( .A1(n16146), .A2(n12393), .ZN(n12394) );
  NAND2_X1 U15371 ( .A1(n12394), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14027) );
  INV_X1 U15372 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16272) );
  NAND2_X1 U15373 ( .A1(n16146), .A2(n16272), .ZN(n12395) );
  NAND2_X2 U15374 ( .A1(n16145), .A2(n12395), .ZN(n14998) );
  INV_X2 U15375 ( .A(n12396), .ZN(n14933) );
  INV_X1 U15376 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16241) );
  INV_X1 U15377 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12403) );
  INV_X1 U15378 ( .A(n15009), .ZN(n12398) );
  INV_X1 U15379 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12923) );
  NAND2_X1 U15380 ( .A1(n16146), .A2(n12923), .ZN(n12397) );
  NAND2_X1 U15381 ( .A1(n12398), .A2(n12397), .ZN(n14999) );
  OR2_X1 U15382 ( .A1(n16146), .A2(n12923), .ZN(n12399) );
  INV_X1 U15383 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16232) );
  XNOR2_X1 U15384 ( .A(n15046), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15001) );
  NAND2_X1 U15385 ( .A1(n16146), .A2(n16232), .ZN(n16137) );
  NAND2_X1 U15386 ( .A1(n15001), .A2(n16137), .ZN(n12400) );
  NOR2_X1 U15387 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15388 ( .A1(n15026), .A2(n15028), .ZN(n15018) );
  NOR2_X1 U15389 ( .A1(n16125), .A2(n15018), .ZN(n12404) );
  XNOR2_X1 U15390 ( .A(n15046), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14991) );
  NAND2_X1 U15391 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15125) );
  INV_X1 U15392 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U15393 ( .A1(n15125), .A2(n15127), .ZN(n12405) );
  INV_X1 U15394 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12407) );
  INV_X1 U15395 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15135) );
  INV_X1 U15396 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15138) );
  NAND2_X1 U15397 ( .A1(n12491), .A2(n15035), .ZN(n14924) );
  AND3_X1 U15398 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15060) );
  NAND2_X1 U15399 ( .A1(n14924), .A2(n12488), .ZN(n12410) );
  INV_X1 U15400 ( .A(n12410), .ZN(n12408) );
  NOR2_X1 U15401 ( .A1(n12408), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12411) );
  INV_X1 U15402 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16183) );
  INV_X1 U15403 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14925) );
  INV_X1 U15404 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14926) );
  NAND3_X1 U15405 ( .A1(n16183), .A2(n14925), .A3(n14926), .ZN(n12492) );
  NOR2_X1 U15406 ( .A1(n12492), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12409) );
  OAI22_X1 U15407 ( .A1(n12410), .A2(n12409), .B1(n15035), .B2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14905) );
  AOI211_X1 U15408 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15035), .A(
        n12411), .B(n14905), .ZN(n12412) );
  XNOR2_X1 U15409 ( .A(n12412), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15096) );
  OR2_X1 U15410 ( .A1(n15096), .A2(n20167), .ZN(n12413) );
  NAND2_X1 U15411 ( .A1(n12414), .A2(n12413), .ZN(P1_U2971) );
  INV_X1 U15412 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12424) );
  INV_X1 U15413 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12416) );
  OAI22_X1 U15414 ( .A1(n11561), .A2(n12417), .B1(n12503), .B2(n12416), .ZN(
        n12421) );
  INV_X1 U15415 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12419) );
  OAI22_X1 U15416 ( .A1(n9688), .A2(n12419), .B1(n9674), .B2(n12418), .ZN(
        n12420) );
  AOI211_X1 U15417 ( .C1(n12124), .C2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n12421), .B(n12420), .ZN(n12423) );
  AOI22_X1 U15418 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12422) );
  OAI211_X1 U15419 ( .C1(n11703), .C2(n12424), .A(n12423), .B(n12422), .ZN(
        n12430) );
  AOI22_X1 U15420 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U15421 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15422 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15423 ( .A1(n12510), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12192), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12425) );
  NAND4_X1 U15424 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12429) );
  NOR2_X1 U15425 ( .A1(n12430), .A2(n12429), .ZN(n12500) );
  NAND2_X1 U15426 ( .A1(n12432), .A2(n12431), .ZN(n12499) );
  XNOR2_X1 U15427 ( .A(n12500), .B(n12499), .ZN(n12438) );
  NAND2_X1 U15428 ( .A1(n11760), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12433) );
  NAND2_X1 U15429 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  AOI21_X1 U15430 ( .B1(n12524), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12435), .ZN(
        n12436) );
  OAI21_X1 U15431 ( .B1(n12438), .B2(n12437), .A(n12436), .ZN(n12444) );
  INV_X1 U15432 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14621) );
  INV_X1 U15433 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12440) );
  NAND2_X1 U15434 ( .A1(n12441), .A2(n12440), .ZN(n12442) );
  AND2_X1 U15435 ( .A1(n13891), .A2(n12442), .ZN(n14287) );
  NAND2_X1 U15436 ( .A1(n14287), .A2(n12523), .ZN(n12443) );
  NAND2_X1 U15437 ( .A1(n12444), .A2(n12443), .ZN(n12447) );
  NOR2_X1 U15438 ( .A1(n12447), .A2(n12445), .ZN(n12446) );
  NAND2_X1 U15439 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20953) );
  INV_X1 U15440 ( .A(n20953), .ZN(n20948) );
  INV_X1 U15441 ( .A(n12450), .ZN(n12456) );
  OR4_X1 U15442 ( .A1(n12454), .A2(n12453), .A3(n12452), .A4(n12451), .ZN(
        n12455) );
  NAND2_X1 U15443 ( .A1(n12456), .A2(n12455), .ZN(n14600) );
  NOR2_X1 U15444 ( .A1(n20948), .A2(n14600), .ZN(n12996) );
  INV_X1 U15445 ( .A(n12996), .ZN(n12459) );
  INV_X1 U15446 ( .A(n15194), .ZN(n13663) );
  NOR2_X1 U15447 ( .A1(n12457), .A2(n14603), .ZN(n12458) );
  NAND2_X1 U15448 ( .A1(n13663), .A2(n12458), .ZN(n14594) );
  OAI22_X1 U15449 ( .A1(n12449), .A2(n12459), .B1(n14596), .B2(n14594), .ZN(
        n13370) );
  NAND2_X1 U15450 ( .A1(n13326), .A2(n20953), .ZN(n12461) );
  INV_X1 U15451 ( .A(n12462), .ZN(n12463) );
  INV_X1 U15452 ( .A(n11567), .ZN(n14843) );
  NAND4_X1 U15453 ( .A1(n12278), .A2(n13013), .A3(n14843), .A4(n11624), .ZN(
        n12868) );
  OAI22_X1 U15454 ( .A1(n9686), .A2(n12464), .B1(n12463), .B2(n12868), .ZN(
        n12465) );
  NOR2_X1 U15455 ( .A1(n11628), .A2(n14843), .ZN(n13511) );
  OR2_X2 U15456 ( .A1(n16115), .A2(n13511), .ZN(n14904) );
  NOR4_X1 U15457 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12470) );
  NOR4_X1 U15458 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12469) );
  NOR4_X1 U15459 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12468) );
  NOR4_X1 U15460 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12467) );
  AND4_X1 U15461 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        n12475) );
  NOR4_X1 U15462 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12473) );
  NOR4_X1 U15463 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12472) );
  NOR4_X1 U15464 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12471) );
  INV_X1 U15465 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20886) );
  AND4_X1 U15466 ( .A1(n12473), .A2(n12472), .A3(n12471), .A4(n20886), .ZN(
        n12474) );
  NAND2_X1 U15467 ( .A1(n12475), .A2(n12474), .ZN(n12476) );
  NOR3_X1 U15468 ( .A1(n16115), .A2(n14848), .A3(n12997), .ZN(n12477) );
  AOI22_X1 U15469 ( .A1(n16118), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16115), .ZN(n12478) );
  INV_X1 U15470 ( .A(n12478), .ZN(n12485) );
  NOR3_X1 U15471 ( .A1(n16115), .A2(n14843), .A3(n13357), .ZN(n12479) );
  INV_X1 U15472 ( .A(DATAI_13_), .ZN(n21091) );
  NAND2_X1 U15473 ( .A1(n14848), .A2(BUF1_REG_13__SCAN_IN), .ZN(n12480) );
  OAI21_X1 U15474 ( .B1(n14260), .B2(n21091), .A(n12480), .ZN(n20311) );
  INV_X1 U15475 ( .A(n12997), .ZN(n12481) );
  NAND2_X1 U15476 ( .A1(n12481), .A2(n14848), .ZN(n12482) );
  AOI22_X1 U15477 ( .A1(n16117), .A2(n20311), .B1(BUF1_REG_29__SCAN_IN), .B2(
        n14885), .ZN(n12483) );
  INV_X1 U15478 ( .A(n12483), .ZN(n12484) );
  NOR2_X1 U15479 ( .A1(n12485), .A2(n12484), .ZN(n12486) );
  OAI21_X1 U15480 ( .B1(n14293), .B2(n14904), .A(n12486), .ZN(P1_U2875) );
  OR2_X1 U15481 ( .A1(n16146), .A2(n12492), .ZN(n12487) );
  NAND2_X1 U15482 ( .A1(n12488), .A2(n12487), .ZN(n12489) );
  INV_X1 U15483 ( .A(n13016), .ZN(n12490) );
  INV_X1 U15484 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15061) );
  NAND2_X1 U15485 ( .A1(n12490), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12992) );
  OAI21_X1 U15486 ( .B1(n12491), .B2(n12492), .A(n15035), .ZN(n12493) );
  NOR2_X1 U15487 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15088) );
  INV_X1 U15488 ( .A(n14529), .ZN(n12497) );
  AND2_X1 U15489 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15087) );
  NAND2_X1 U15490 ( .A1(n12396), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12495) );
  INV_X1 U15491 ( .A(n14527), .ZN(n12496) );
  NOR2_X1 U15492 ( .A1(n12500), .A2(n12499), .ZN(n12519) );
  INV_X1 U15493 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12509) );
  OAI22_X1 U15494 ( .A1(n11561), .A2(n12501), .B1(n11569), .B2(n13934), .ZN(
        n12506) );
  INV_X1 U15495 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12504) );
  OAI22_X1 U15496 ( .A1(n11576), .A2(n12504), .B1(n12503), .B2(n12502), .ZN(
        n12505) );
  AOI211_X1 U15497 ( .C1(n12124), .C2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12506), .B(n12505), .ZN(n12508) );
  AOI22_X1 U15498 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11491), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12507) );
  OAI211_X1 U15499 ( .C1(n11690), .C2(n12509), .A(n12508), .B(n12507), .ZN(
        n12517) );
  AOI22_X1 U15500 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12510), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15501 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15502 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11545), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15503 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12512) );
  NAND4_X1 U15504 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12516) );
  NOR2_X1 U15505 ( .A1(n12517), .A2(n12516), .ZN(n12518) );
  XNOR2_X1 U15506 ( .A(n12519), .B(n12518), .ZN(n12521) );
  NAND2_X1 U15507 ( .A1(n12521), .A2(n12520), .ZN(n12526) );
  INV_X1 U15508 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13890) );
  NOR2_X1 U15509 ( .A1(n13890), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12522) );
  AOI211_X1 U15510 ( .C1(n12524), .C2(P1_EAX_REG_30__SCAN_IN), .A(n12523), .B(
        n12522), .ZN(n12525) );
  XNOR2_X1 U15511 ( .A(n13891), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14278) );
  AOI22_X1 U15512 ( .A1(n12526), .A2(n12525), .B1(n13889), .B2(n14278), .ZN(
        n14532) );
  XNOR2_X2 U15513 ( .A(n12527), .B(n14532), .ZN(n14285) );
  INV_X1 U15514 ( .A(n20344), .ZN(n15054) );
  INV_X1 U15515 ( .A(n20338), .ZN(n15039) );
  INV_X2 U15516 ( .A(n20351), .ZN(n20377) );
  NAND2_X1 U15517 ( .A1(n20377), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15070) );
  OAI21_X1 U15518 ( .B1(n15039), .B2(n13890), .A(n15070), .ZN(n12528) );
  OAI21_X1 U15519 ( .B1(n15077), .B2(n20167), .A(n12531), .ZN(P1_U2969) );
  BUF_X4 U15520 ( .A(n12582), .Z(n17365) );
  AOI22_X1 U15521 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12538) );
  NAND2_X1 U15522 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18875), .ZN(
        n18877) );
  AOI22_X1 U15523 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15524 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12536) );
  INV_X4 U15525 ( .A(n17150), .ZN(n17386) );
  AND2_X2 U15526 ( .A1(n12534), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17387) );
  AOI22_X1 U15527 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12535) );
  NAND4_X1 U15528 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12549) );
  NOR2_X2 U15529 ( .A1(n12539), .A2(n18884), .ZN(n12574) );
  BUF_X2 U15530 ( .A(n12574), .Z(n17394) );
  AOI22_X1 U15531 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12574), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12547) );
  NOR2_X2 U15532 ( .A1(n12543), .A2(n12540), .ZN(n12585) );
  INV_X4 U15533 ( .A(n12541), .ZN(n17384) );
  AOI22_X1 U15534 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12546) );
  NOR3_X4 U15535 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n12540), .ZN(n12581) );
  NOR2_X2 U15536 ( .A1(n18888), .A2(n12543), .ZN(n12584) );
  AOI22_X1 U15537 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12545) );
  NOR2_X2 U15538 ( .A1(n18884), .A2(n12543), .ZN(n12563) );
  AOI22_X1 U15539 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12544) );
  NAND4_X1 U15540 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12544), .ZN(
        n12548) );
  AOI22_X1 U15541 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15542 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15543 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15544 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12551) );
  NAND4_X1 U15545 ( .A1(n12554), .A2(n12553), .A3(n12552), .A4(n12551), .ZN(
        n12560) );
  AOI22_X1 U15546 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15547 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15548 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15549 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12555) );
  NAND4_X1 U15550 ( .A1(n12558), .A2(n12557), .A3(n12556), .A4(n12555), .ZN(
        n12559) );
  INV_X1 U15551 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14133) );
  AOI22_X1 U15552 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12573), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12561) );
  OAI21_X1 U15553 ( .B1(n14110), .B2(n14133), .A(n12561), .ZN(n12562) );
  AOI22_X1 U15554 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12583), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15555 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15556 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15557 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15558 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12575), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15559 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12582), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15560 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12550), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17387), .ZN(n12580) );
  INV_X1 U15561 ( .A(n12573), .ZN(n17197) );
  AOI22_X1 U15562 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17367), .B1(
        n17369), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15563 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15564 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12575), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12577) );
  NAND4_X1 U15565 ( .A1(n12580), .A2(n12579), .A3(n12578), .A4(n12577), .ZN(
        n12591) );
  AOI22_X1 U15566 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12563), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15567 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12582), .ZN(n12588) );
  AOI22_X1 U15568 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12583), .ZN(n12587) );
  AOI22_X1 U15569 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12584), .B1(
        n12585), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12586) );
  NAND4_X1 U15570 ( .A1(n12589), .A2(n12588), .A3(n12587), .A4(n12586), .ZN(
        n12590) );
  OR2_X2 U15571 ( .A1(n12591), .A2(n12590), .ZN(n17593) );
  AOI22_X1 U15572 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15573 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15574 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15575 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12592) );
  NAND4_X1 U15576 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12601) );
  AOI22_X1 U15577 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12582), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15578 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15579 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15580 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12596) );
  NAND4_X1 U15581 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12600) );
  AOI22_X1 U15582 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12612) );
  BUF_X2 U15583 ( .A(n12563), .Z(n17374) );
  AOI22_X1 U15584 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12611) );
  INV_X1 U15585 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U15586 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12603) );
  OAI21_X1 U15587 ( .B1(n14110), .B2(n17424), .A(n12603), .ZN(n12609) );
  AOI22_X1 U15588 ( .A1(n12584), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12582), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15589 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15590 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15591 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12604) );
  NAND4_X1 U15592 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n12608) );
  AOI211_X1 U15593 ( .C1(n17350), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n12609), .B(n12608), .ZN(n12610) );
  NAND3_X1 U15594 ( .A1(n12612), .A2(n12611), .A3(n12610), .ZN(n17577) );
  NAND2_X1 U15595 ( .A1(n12638), .A2(n17577), .ZN(n12642) );
  NOR2_X1 U15596 ( .A1(n17573), .A2(n12642), .ZN(n12646) );
  AOI22_X1 U15597 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15598 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15599 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12613) );
  OAI21_X1 U15600 ( .B1(n14110), .B2(n17415), .A(n12613), .ZN(n12619) );
  AOI22_X1 U15601 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15602 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15603 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15604 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12614) );
  NAND4_X1 U15605 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n12618) );
  AOI211_X1 U15606 ( .C1(n17350), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n12619), .B(n12618), .ZN(n12620) );
  NAND3_X1 U15607 ( .A1(n12622), .A2(n12621), .A3(n12620), .ZN(n17569) );
  NOR2_X4 U15608 ( .A1(n17565), .A2(n12623), .ZN(n17955) );
  NAND2_X1 U15609 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18083) );
  INV_X1 U15610 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18107) );
  INV_X1 U15611 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12657) );
  INV_X1 U15612 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12656) );
  INV_X1 U15613 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18354) );
  INV_X1 U15614 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18380) );
  NAND2_X1 U15615 ( .A1(n12816), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12634) );
  AOI22_X1 U15616 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15617 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U15618 ( .A1(n12576), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15619 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12624) );
  NAND4_X1 U15620 ( .A1(n12627), .A2(n12626), .A3(n12625), .A4(n12624), .ZN(
        n12633) );
  AOI22_X1 U15621 ( .A1(n12583), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15622 ( .A1(n12581), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12582), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15623 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15624 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12628) );
  NAND4_X1 U15625 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12632) );
  INV_X1 U15626 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18385) );
  NAND2_X1 U15627 ( .A1(n18067), .A2(n18075), .ZN(n18066) );
  NAND2_X1 U15628 ( .A1(n12634), .A2(n18066), .ZN(n18056) );
  NAND2_X1 U15629 ( .A1(n18057), .A2(n18056), .ZN(n18055) );
  OR2_X1 U15630 ( .A1(n18380), .A2(n12635), .ZN(n12636) );
  XOR2_X1 U15631 ( .A(n17581), .B(n12637), .Z(n18041) );
  NAND2_X1 U15632 ( .A1(n18042), .A2(n18041), .ZN(n18040) );
  NAND2_X1 U15633 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12640), .ZN(
        n12641) );
  XOR2_X1 U15634 ( .A(n17573), .B(n12642), .Z(n12644) );
  INV_X1 U15635 ( .A(n12644), .ZN(n12643) );
  XOR2_X1 U15636 ( .A(n17569), .B(n12646), .Z(n12647) );
  XOR2_X1 U15637 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12647), .Z(
        n18009) );
  NAND2_X1 U15638 ( .A1(n18008), .A2(n18009), .ZN(n18007) );
  NAND2_X1 U15639 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12647), .ZN(
        n12648) );
  NAND2_X1 U15640 ( .A1(n12649), .A2(n12651), .ZN(n12652) );
  INV_X1 U15641 ( .A(n12649), .ZN(n12650) );
  XNOR2_X1 U15642 ( .A(n12651), .B(n12650), .ZN(n17993) );
  INV_X1 U15643 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12655) );
  NAND2_X1 U15644 ( .A1(n17935), .A2(n12655), .ZN(n17922) );
  INV_X1 U15645 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18269) );
  INV_X1 U15646 ( .A(n12664), .ZN(n12662) );
  NOR2_X1 U15647 ( .A1(n12654), .A2(n12653), .ZN(n18281) );
  NAND2_X1 U15648 ( .A1(n18281), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18263) );
  INV_X1 U15649 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18229) );
  NOR3_X1 U15650 ( .A1(n18263), .A2(n18229), .A3(n12656), .ZN(n17877) );
  NAND2_X1 U15651 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17877), .ZN(
        n18218) );
  NOR2_X1 U15652 ( .A1(n18218), .A2(n12657), .ZN(n17863) );
  NAND2_X1 U15653 ( .A1(n17863), .A2(n17917), .ZN(n12663) );
  NAND2_X1 U15654 ( .A1(n12663), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12660) );
  INV_X1 U15655 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18212) );
  NAND2_X1 U15656 ( .A1(n12660), .A2(n12659), .ZN(n12661) );
  NOR2_X2 U15657 ( .A1(n12662), .A2(n12661), .ZN(n17857) );
  INV_X1 U15658 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17861) );
  NAND2_X1 U15659 ( .A1(n17857), .A2(n17861), .ZN(n17856) );
  NAND2_X2 U15660 ( .A1(n17856), .A2(n17978), .ZN(n17824) );
  NAND2_X1 U15661 ( .A1(n12664), .A2(n12663), .ZN(n17864) );
  NOR2_X1 U15662 ( .A1(n18212), .A2(n17861), .ZN(n18184) );
  INV_X1 U15663 ( .A(n18184), .ZN(n17847) );
  INV_X1 U15664 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18182) );
  INV_X1 U15665 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18148) );
  NOR2_X1 U15666 ( .A1(n18182), .A2(n18148), .ZN(n18160) );
  NAND3_X1 U15667 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18160), .ZN(n17790) );
  NOR2_X1 U15668 ( .A1(n17847), .A2(n17790), .ZN(n18146) );
  INV_X1 U15669 ( .A(n18146), .ZN(n18150) );
  INV_X1 U15670 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18151) );
  NOR2_X1 U15671 ( .A1(n18150), .A2(n18151), .ZN(n18105) );
  INV_X1 U15672 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18139) );
  NOR2_X1 U15673 ( .A1(n18135), .A2(n18139), .ZN(n17764) );
  NOR2_X1 U15674 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17955), .ZN(
        n17840) );
  NAND2_X1 U15675 ( .A1(n17840), .A2(n18182), .ZN(n12665) );
  NOR2_X1 U15676 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12665), .ZN(
        n17812) );
  INV_X1 U15677 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18149) );
  NAND2_X1 U15678 ( .A1(n17812), .A2(n18149), .ZN(n17789) );
  NOR3_X1 U15679 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17789), .ZN(n12666) );
  NAND2_X1 U15680 ( .A1(n18184), .A2(n17864), .ZN(n17809) );
  OR2_X1 U15681 ( .A1(n17955), .A2(n17765), .ZN(n17753) );
  NOR2_X1 U15682 ( .A1(n17754), .A2(n17978), .ZN(n12669) );
  NAND2_X1 U15683 ( .A1(n16588), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17726) );
  INV_X1 U15684 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16587) );
  AOI22_X1 U15685 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17955), .B1(
        n17978), .B2(n16587), .ZN(n17721) );
  AOI21_X2 U15686 ( .B1(n16592), .B2(n9718), .A(n17721), .ZN(n15971) );
  INV_X1 U15687 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16563) );
  NAND2_X1 U15688 ( .A1(n15971), .A2(n16563), .ZN(n15970) );
  NAND2_X2 U15689 ( .A1(n15970), .A2(n17978), .ZN(n16021) );
  INV_X1 U15690 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19037) );
  NAND3_X1 U15691 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16578) );
  AOI21_X1 U15692 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n19037), .A(
        n12672), .ZN(n12670) );
  NOR2_X1 U15693 ( .A1(n19037), .A2(n17978), .ZN(n12674) );
  AOI22_X1 U15694 ( .A1(n19037), .A2(n17978), .B1(n12674), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12671) );
  INV_X1 U15695 ( .A(n12671), .ZN(n12676) );
  NOR2_X1 U15696 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17955), .ZN(
        n12673) );
  AOI22_X1 U15697 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18679), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19048), .ZN(n12797) );
  OAI22_X1 U15698 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18908), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12682), .ZN(n12687) );
  NOR2_X1 U15699 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18908), .ZN(
        n12683) );
  NAND2_X1 U15700 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12682), .ZN(
        n12688) );
  AOI22_X1 U15701 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12687), .B1(
        n12683), .B2(n12688), .ZN(n12692) );
  AOI21_X1 U15702 ( .B1(n12679), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12796), .ZN(n12800) );
  AND2_X1 U15703 ( .A1(n12797), .A2(n12800), .ZN(n12691) );
  OAI21_X1 U15704 ( .B1(n12686), .B2(n12685), .A(n12692), .ZN(n12684) );
  AOI21_X1 U15705 ( .B1(n12688), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n12687), .ZN(n12689) );
  AOI21_X1 U15706 ( .B1(n18908), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n12689), .ZN(n12690) );
  INV_X1 U15707 ( .A(n12690), .ZN(n12798) );
  AOI22_X1 U15708 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15709 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U15710 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U15711 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12693) );
  NAND4_X1 U15712 ( .A1(n12696), .A2(n12695), .A3(n12694), .A4(n12693), .ZN(
        n12704) );
  AOI22_X1 U15713 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17395), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15714 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15715 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12700) );
  INV_X2 U15716 ( .A(n14122), .ZN(n17349) );
  AOI22_X1 U15717 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12699) );
  NAND4_X1 U15718 ( .A1(n12702), .A2(n12701), .A3(n12700), .A4(n12699), .ZN(
        n12703) );
  AOI22_X1 U15719 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15720 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15721 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15722 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12705) );
  NAND4_X1 U15723 ( .A1(n12708), .A2(n12707), .A3(n12706), .A4(n12705), .ZN(
        n12714) );
  AOI22_X1 U15724 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15725 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17395), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15726 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15727 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12709) );
  NAND4_X1 U15728 ( .A1(n12712), .A2(n12711), .A3(n12710), .A4(n12709), .ZN(
        n12713) );
  AOI22_X1 U15729 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15730 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15731 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15732 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12715) );
  NAND4_X1 U15733 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        n12725) );
  AOI22_X1 U15734 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15735 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15736 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15737 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12720) );
  NAND4_X1 U15738 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12724) );
  AOI22_X1 U15739 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15740 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15741 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15742 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12726) );
  NAND4_X1 U15743 ( .A1(n12729), .A2(n12728), .A3(n12727), .A4(n12726), .ZN(
        n12735) );
  AOI22_X1 U15744 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15745 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15746 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15747 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12730) );
  NAND4_X1 U15748 ( .A1(n12733), .A2(n12732), .A3(n12731), .A4(n12730), .ZN(
        n12734) );
  AOI22_X1 U15749 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U15750 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U15751 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U15752 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12736) );
  NAND4_X1 U15753 ( .A1(n12739), .A2(n12738), .A3(n12737), .A4(n12736), .ZN(
        n12745) );
  AOI22_X1 U15754 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U15755 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15756 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15757 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12740) );
  NAND4_X1 U15758 ( .A1(n12743), .A2(n12742), .A3(n12741), .A4(n12740), .ZN(
        n12744) );
  AOI22_X1 U15759 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15760 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15761 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12746) );
  OAI21_X1 U15762 ( .B1(n14122), .B2(n14133), .A(n12746), .ZN(n12752) );
  AOI22_X1 U15763 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15764 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15765 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U15766 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12747) );
  NAND4_X1 U15767 ( .A1(n12750), .A2(n12749), .A3(n12748), .A4(n12747), .ZN(
        n12751) );
  AOI211_X1 U15768 ( .C1(n17384), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n12752), .B(n12751), .ZN(n12753) );
  NAND3_X1 U15769 ( .A1(n12755), .A2(n12754), .A3(n12753), .ZN(n12802) );
  AOI22_X1 U15770 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15771 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17350), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15772 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U15773 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12756) );
  NAND4_X1 U15774 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n12765) );
  AOI22_X1 U15775 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15776 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U15777 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U15778 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12760) );
  NAND4_X1 U15779 ( .A1(n12763), .A2(n12762), .A3(n12761), .A4(n12760), .ZN(
        n12764) );
  AOI22_X1 U15780 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U15781 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15782 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12766) );
  OAI21_X1 U15783 ( .B1(n14122), .B2(n17415), .A(n12766), .ZN(n12772) );
  AOI22_X1 U15784 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U15785 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U15786 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U15787 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12767) );
  NAND4_X1 U15788 ( .A1(n12770), .A2(n12769), .A3(n12768), .A4(n12767), .ZN(
        n12771) );
  NOR2_X1 U15789 ( .A1(n18432), .A2(n17444), .ZN(n18870) );
  NAND3_X1 U15790 ( .A1(n12806), .A2(n15961), .A3(n18870), .ZN(n14074) );
  INV_X1 U15791 ( .A(n18427), .ZN(n12787) );
  NOR2_X1 U15792 ( .A1(n12787), .A2(n12802), .ZN(n18869) );
  INV_X1 U15793 ( .A(n17444), .ZN(n18441) );
  NAND2_X1 U15794 ( .A1(n18869), .A2(n12804), .ZN(n14073) );
  NOR2_X1 U15795 ( .A1(n12777), .A2(n14073), .ZN(n12778) );
  INV_X1 U15796 ( .A(n12802), .ZN(n18423) );
  NOR2_X1 U15797 ( .A1(n14072), .A2(n17444), .ZN(n12783) );
  NOR4_X2 U15798 ( .A1(n12787), .A2(n14072), .A3(n12790), .A4(n12777), .ZN(
        n12791) );
  AND2_X1 U15799 ( .A1(n12802), .A2(n12791), .ZN(n15943) );
  NOR2_X4 U15800 ( .A1(n17640), .A2(n15943), .ZN(n16712) );
  NOR2_X4 U15801 ( .A1(n19077), .A2(n16712), .ZN(n16731) );
  AOI211_X2 U15802 ( .C1(n19074), .C2(n12778), .A(n16730), .B(n16731), .ZN(
        n18879) );
  NAND2_X1 U15803 ( .A1(n18416), .A2(n16733), .ZN(n12779) );
  NAND2_X1 U15804 ( .A1(n18423), .A2(n12779), .ZN(n12803) );
  NOR2_X1 U15805 ( .A1(n18416), .A2(n16733), .ZN(n12780) );
  NOR2_X1 U15806 ( .A1(n17444), .A2(n18436), .ZN(n12807) );
  INV_X1 U15807 ( .A(n12807), .ZN(n18893) );
  NAND2_X1 U15808 ( .A1(n17564), .A2(n18893), .ZN(n16041) );
  NAND2_X1 U15809 ( .A1(n12780), .A2(n16041), .ZN(n15942) );
  AOI221_X1 U15810 ( .B1(n15961), .B2(n15942), .C1(n12781), .C2(n15942), .A(
        n18427), .ZN(n12789) );
  INV_X1 U15811 ( .A(n12790), .ZN(n12784) );
  OAI21_X1 U15812 ( .B1(n12802), .B2(n17600), .A(n18893), .ZN(n12782) );
  OAI21_X1 U15813 ( .B1(n12784), .B2(n12783), .A(n12782), .ZN(n12786) );
  OAI21_X1 U15814 ( .B1(n18448), .B2(n12784), .A(n14072), .ZN(n12785) );
  OAI211_X1 U15815 ( .C1(n12788), .C2(n12787), .A(n12786), .B(n12785), .ZN(
        n15940) );
  NAND2_X1 U15816 ( .A1(n12791), .A2(n12795), .ZN(n18865) );
  NAND2_X1 U15817 ( .A1(n18879), .A2(n18865), .ZN(n18897) );
  INV_X1 U15818 ( .A(n12806), .ZN(n12793) );
  INV_X1 U15819 ( .A(n16731), .ZN(n12792) );
  NAND3_X1 U15820 ( .A1(n12793), .A2(n16733), .A3(n12792), .ZN(n12794) );
  NAND2_X1 U15821 ( .A1(n12795), .A2(n12794), .ZN(n18868) );
  AOI21_X2 U15822 ( .B1(n18869), .B2(n18879), .A(n18868), .ZN(n18894) );
  XOR2_X1 U15823 ( .A(n12797), .B(n12796), .Z(n12799) );
  AOI21_X1 U15824 ( .B1(n12801), .B2(n12800), .A(n16710), .ZN(n18857) );
  NOR2_X1 U15825 ( .A1(n19074), .A2(n12802), .ZN(n15958) );
  NAND2_X1 U15826 ( .A1(n15958), .A2(n17444), .ZN(n15962) );
  NOR2_X1 U15827 ( .A1(n12804), .A2(n12803), .ZN(n12805) );
  OAI211_X1 U15828 ( .C1(n18432), .C2(n12807), .A(n12806), .B(n12805), .ZN(
        n15941) );
  NAND2_X1 U15829 ( .A1(n19049), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18929) );
  NOR2_X2 U15830 ( .A1(n18861), .A2(n18924), .ZN(n12808) );
  NAND2_X1 U15831 ( .A1(n16582), .A2(n17973), .ZN(n12848) );
  NAND2_X1 U15832 ( .A1(n19049), .A2(n19028), .ZN(n19032) );
  NAND2_X1 U15833 ( .A1(n19086), .A2(n19028), .ZN(n16707) );
  AND2_X1 U15834 ( .A1(n19032), .A2(n16707), .ZN(n19068) );
  INV_X1 U15835 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19073) );
  NOR2_X1 U15836 ( .A1(n19049), .A2(n19073), .ZN(n17907) );
  INV_X1 U15837 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16760) );
  INV_X1 U15838 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18070) );
  NAND2_X1 U15839 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17979) );
  NAND4_X1 U15840 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17938), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17906) );
  NAND2_X1 U15841 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17868) );
  NAND2_X1 U15842 ( .A1(n17851), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17829) );
  NAND2_X1 U15843 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17830) );
  NAND2_X1 U15844 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17796) );
  NAND2_X1 U15845 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17758) );
  NAND2_X1 U15846 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17712) );
  NAND2_X1 U15847 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16567), .ZN(
        n12809) );
  INV_X1 U15848 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19014) );
  NOR3_X1 U15849 ( .A1(n19032), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n16729) );
  NOR2_X1 U15850 ( .A1(n19014), .A2(n9655), .ZN(n16580) );
  INV_X1 U15851 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18926) );
  NAND2_X1 U15852 ( .A1(n18926), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18937) );
  NOR2_X1 U15853 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19028), .ZN(
        n19053) );
  NOR2_X1 U15854 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19078) );
  AOI21_X1 U15855 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19078), .ZN(n18934) );
  NAND3_X1 U15856 ( .A1(n19086), .A2(n19028), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18654) );
  INV_X2 U15857 ( .A(n18444), .ZN(n18798) );
  OR2_X1 U15858 ( .A1(n12810), .A2(n17910), .ZN(n16550) );
  XNOR2_X1 U15859 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12812) );
  INV_X1 U15860 ( .A(n17780), .ZN(n17817) );
  NOR2_X1 U15861 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17817), .ZN(
        n16569) );
  NAND2_X1 U15862 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9777), .ZN(
        n16568) );
  INV_X1 U15863 ( .A(n16568), .ZN(n16738) );
  NAND2_X1 U15864 ( .A1(n18798), .A2(n12810), .ZN(n12811) );
  OAI211_X1 U15865 ( .C1(n16738), .C2(n18937), .A(n9676), .B(n12811), .ZN(
        n16570) );
  NOR2_X1 U15866 ( .A1(n16569), .A2(n16570), .ZN(n16549) );
  OAI22_X1 U15867 ( .A1(n16550), .A2(n12812), .B1(n16549), .B2(n16760), .ZN(
        n12813) );
  AOI211_X1 U15868 ( .C1(n17927), .C2(n17083), .A(n16580), .B(n12813), .ZN(
        n12847) );
  NAND2_X1 U15869 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18103) );
  INV_X1 U15870 ( .A(n18103), .ZN(n18106) );
  NAND3_X1 U15871 ( .A1(n18106), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16552) );
  NOR2_X1 U15872 ( .A1(n18135), .A2(n16552), .ZN(n18081) );
  NAND2_X1 U15873 ( .A1(n17904), .A2(n17863), .ZN(n18217) );
  NAND2_X1 U15874 ( .A1(n18081), .A2(n17886), .ZN(n18090) );
  NOR2_X1 U15875 ( .A1(n16578), .A2(n18090), .ZN(n16561) );
  NAND2_X1 U15876 ( .A1(n16561), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12814) );
  XOR2_X1 U15877 ( .A(n12814), .B(n19037), .Z(n16583) );
  INV_X1 U15878 ( .A(n17565), .ZN(n16594) );
  NOR2_X2 U15879 ( .A1(n16594), .A2(n18079), .ZN(n17945) );
  NAND2_X1 U15880 ( .A1(n16583), .A2(n17945), .ZN(n12846) );
  INV_X1 U15881 ( .A(n18218), .ZN(n17896) );
  NOR2_X1 U15882 ( .A1(n12822), .A2(n17581), .ZN(n12821) );
  NAND2_X1 U15883 ( .A1(n12821), .A2(n17577), .ZN(n12819) );
  NOR2_X1 U15884 ( .A1(n17573), .A2(n12819), .ZN(n12818) );
  NAND2_X1 U15885 ( .A1(n12818), .A2(n17569), .ZN(n12817) );
  NOR2_X1 U15886 ( .A1(n17565), .A2(n12817), .ZN(n12841) );
  XOR2_X1 U15887 ( .A(n12817), .B(n17565), .Z(n18000) );
  XOR2_X1 U15888 ( .A(n12818), .B(n17569), .Z(n12834) );
  XOR2_X1 U15889 ( .A(n12819), .B(n17573), .Z(n12820) );
  NAND2_X1 U15890 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12820), .ZN(
        n12833) );
  XOR2_X1 U15891 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12820), .Z(
        n18019) );
  XOR2_X1 U15892 ( .A(n12821), .B(n17577), .Z(n12831) );
  XOR2_X1 U15893 ( .A(n17581), .B(n12822), .Z(n12823) );
  NAND2_X1 U15894 ( .A1(n12823), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12829) );
  XOR2_X1 U15895 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12823), .Z(
        n18046) );
  OR2_X1 U15896 ( .A1(n18380), .A2(n12825), .ZN(n12828) );
  INV_X1 U15897 ( .A(n12815), .ZN(n16042) );
  AOI21_X1 U15898 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17593), .A(
        n16042), .ZN(n12827) );
  NOR2_X1 U15899 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17593), .ZN(
        n12826) );
  AOI221_X1 U15900 ( .B1(n16042), .B2(n17593), .C1(n12827), .C2(n18385), .A(
        n12826), .ZN(n18059) );
  NAND2_X1 U15901 ( .A1(n18060), .A2(n18059), .ZN(n18058) );
  NAND2_X1 U15902 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  NAND2_X1 U15903 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18034), .ZN(
        n18033) );
  NAND2_X1 U15904 ( .A1(n12832), .A2(n18033), .ZN(n18018) );
  NAND2_X1 U15905 ( .A1(n18019), .A2(n18018), .ZN(n18017) );
  NAND2_X1 U15906 ( .A1(n12833), .A2(n18017), .ZN(n12835) );
  NAND2_X1 U15907 ( .A1(n12834), .A2(n12835), .ZN(n12836) );
  XOR2_X1 U15908 ( .A(n12835), .B(n12834), .Z(n18006) );
  NAND2_X1 U15909 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18006), .ZN(
        n18005) );
  INV_X1 U15910 ( .A(n12840), .ZN(n12837) );
  NAND2_X1 U15911 ( .A1(n12841), .A2(n12837), .ZN(n12842) );
  NAND2_X1 U15912 ( .A1(n18000), .A2(n17999), .ZN(n12839) );
  NAND2_X1 U15913 ( .A1(n12841), .A2(n12840), .ZN(n12838) );
  OAI211_X1 U15914 ( .C1(n12841), .C2(n12840), .A(n12839), .B(n12838), .ZN(
        n17985) );
  NAND2_X1 U15915 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17985), .ZN(
        n17984) );
  NAND2_X1 U15916 ( .A1(n17885), .A2(n18081), .ZN(n18087) );
  NAND2_X1 U15917 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16558), .ZN(
        n12843) );
  XNOR2_X1 U15918 ( .A(n19037), .B(n12843), .ZN(n16586) );
  INV_X1 U15919 ( .A(n16586), .ZN(n12844) );
  NAND2_X1 U15920 ( .A1(n12844), .A2(n18069), .ZN(n12845) );
  NAND2_X1 U15921 ( .A1(n12848), .A2(n10212), .ZN(P3_U2799) );
  NAND2_X1 U15922 ( .A1(n12851), .A2(n12850), .ZN(n12852) );
  XNOR2_X1 U15923 ( .A(n12854), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12855) );
  NAND2_X1 U15924 ( .A1(n15291), .A2(n12856), .ZN(n12857) );
  AOI21_X1 U15925 ( .B1(n15705), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12862) );
  NOR2_X1 U15926 ( .A1(n12858), .A2(n12859), .ZN(n12860) );
  OR2_X1 U15927 ( .A1(n11257), .A2(n12860), .ZN(n15464) );
  INV_X1 U15928 ( .A(n15464), .ZN(n16337) );
  NOR2_X1 U15929 ( .A1(n16466), .A2(n20083), .ZN(n15557) );
  AOI21_X1 U15930 ( .B1(n16337), .B2(n19436), .A(n15557), .ZN(n12861) );
  OAI21_X1 U15931 ( .B1(n12863), .B2(n12862), .A(n12861), .ZN(n12864) );
  NAND2_X1 U15932 ( .A1(n12866), .A2(n13895), .ZN(n12867) );
  OR2_X1 U15933 ( .A1(n15194), .A2(n12867), .ZN(n13658) );
  INV_X1 U15934 ( .A(n13658), .ZN(n14598) );
  NAND2_X1 U15935 ( .A1(n14596), .A2(n14598), .ZN(n12872) );
  INV_X1 U15936 ( .A(n12868), .ZN(n12870) );
  NAND4_X1 U15937 ( .A1(n12870), .A2(n11622), .A3(n12869), .A4(n13895), .ZN(
        n12871) );
  NAND2_X1 U15938 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  INV_X1 U15939 ( .A(n14842), .ZN(n12977) );
  NAND2_X1 U15940 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12876) );
  INV_X1 U15941 ( .A(n12886), .ZN(n12922) );
  MUX2_X1 U15943 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12875) );
  NAND3_X1 U15944 ( .A1(n12876), .A2(n12932), .A3(n12875), .ZN(n12880) );
  NAND2_X1 U15945 ( .A1(n12953), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12879) );
  INV_X1 U15946 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12877) );
  NAND2_X1 U15947 ( .A1(n12962), .A2(n12877), .ZN(n12878) );
  NAND2_X1 U15948 ( .A1(n12879), .A2(n12878), .ZN(n13425) );
  INV_X1 U15949 ( .A(n12880), .ZN(n12881) );
  MUX2_X1 U15950 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12885) );
  NAND2_X1 U15951 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12883) );
  AND2_X1 U15952 ( .A1(n12932), .A2(n12883), .ZN(n12884) );
  NAND2_X1 U15953 ( .A1(n12885), .A2(n12884), .ZN(n13792) );
  NAND2_X1 U15954 ( .A1(n13793), .A2(n13792), .ZN(n13795) );
  INV_X1 U15955 ( .A(n13795), .ZN(n12890) );
  NAND2_X1 U15956 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12887) );
  OAI211_X1 U15957 ( .C1(n14611), .C2(P1_EBX_REG_3__SCAN_IN), .A(n12953), .B(
        n12887), .ZN(n12888) );
  OAI21_X1 U15958 ( .B1(n12952), .B2(P1_EBX_REG_3__SCAN_IN), .A(n12888), .ZN(
        n13775) );
  MUX2_X1 U15959 ( .A(n12946), .B(n12922), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12892) );
  INV_X1 U15960 ( .A(n12882), .ZN(n12924) );
  OAI21_X1 U15961 ( .B1(n12924), .B2(n20359), .A(n12932), .ZN(n12891) );
  INV_X1 U15962 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20269) );
  NAND2_X1 U15963 ( .A1(n12961), .A2(n20269), .ZN(n12895) );
  NAND2_X1 U15964 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12893) );
  OAI211_X1 U15965 ( .C1(n14611), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12953), .B(
        n12893), .ZN(n12894) );
  MUX2_X1 U15966 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12898) );
  NAND2_X1 U15967 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12896) );
  AND2_X1 U15968 ( .A1(n12932), .A2(n12896), .ZN(n12897) );
  NAND2_X1 U15969 ( .A1(n12898), .A2(n12897), .ZN(n16286) );
  INV_X1 U15970 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20263) );
  NAND2_X1 U15971 ( .A1(n12961), .A2(n20263), .ZN(n12902) );
  NAND2_X1 U15972 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12900) );
  OAI211_X1 U15973 ( .C1(n14611), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12953), .B(
        n12900), .ZN(n12901) );
  MUX2_X1 U15974 ( .A(n12946), .B(n12922), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12905) );
  INV_X1 U15975 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14034) );
  OAI21_X1 U15976 ( .B1(n12924), .B2(n14034), .A(n12932), .ZN(n12904) );
  NOR2_X1 U15977 ( .A1(n12905), .A2(n12904), .ZN(n14009) );
  NAND2_X1 U15978 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12906) );
  OAI211_X1 U15979 ( .C1(n14611), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12953), .B(
        n12906), .ZN(n12907) );
  OAI21_X1 U15980 ( .B1(n12952), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12907), .ZN(
        n14015) );
  INV_X1 U15981 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n16103) );
  NAND2_X1 U15982 ( .A1(n12946), .A2(n16103), .ZN(n12912) );
  INV_X1 U15983 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12908) );
  NAND2_X1 U15984 ( .A1(n12953), .A2(n12908), .ZN(n12910) );
  NAND2_X1 U15985 ( .A1(n13895), .A2(n16103), .ZN(n12909) );
  NAND3_X1 U15986 ( .A1(n12910), .A2(n12962), .A3(n12909), .ZN(n12911) );
  NAND2_X1 U15987 ( .A1(n12912), .A2(n12911), .ZN(n14210) );
  NAND2_X1 U15988 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12913) );
  OAI211_X1 U15989 ( .C1(n14611), .C2(P1_EBX_REG_11__SCAN_IN), .A(n12953), .B(
        n12913), .ZN(n12914) );
  OAI21_X1 U15990 ( .B1(n12952), .B2(P1_EBX_REG_11__SCAN_IN), .A(n12914), .ZN(
        n14782) );
  MUX2_X1 U15991 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12917) );
  NAND2_X1 U15992 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12915) );
  AND2_X1 U15993 ( .A1(n12932), .A2(n12915), .ZN(n12916) );
  NAND2_X1 U15994 ( .A1(n12917), .A2(n12916), .ZN(n16076) );
  INV_X1 U15995 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n16114) );
  NAND2_X1 U15996 ( .A1(n12961), .A2(n16114), .ZN(n12920) );
  NAND2_X1 U15997 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12918) );
  OAI211_X1 U15998 ( .C1(n14611), .C2(P1_EBX_REG_13__SCAN_IN), .A(n12953), .B(
        n12918), .ZN(n12919) );
  NAND2_X1 U15999 ( .A1(n16076), .A2(n16077), .ZN(n12921) );
  MUX2_X1 U16000 ( .A(n12946), .B(n12922), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12926) );
  OAI21_X1 U16001 ( .B1(n12924), .B2(n12923), .A(n12932), .ZN(n12925) );
  NOR2_X1 U16002 ( .A1(n12926), .A2(n12925), .ZN(n14833) );
  OR2_X1 U16003 ( .A1(n12927), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12930) );
  INV_X1 U16004 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14827) );
  NAND2_X1 U16005 ( .A1(n12961), .A2(n14827), .ZN(n12929) );
  NAND2_X1 U16006 ( .A1(n12899), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n12928) );
  MUX2_X1 U16007 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12934) );
  NAND2_X1 U16008 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12931) );
  AND2_X1 U16009 ( .A1(n12932), .A2(n12931), .ZN(n12933) );
  NAND2_X1 U16010 ( .A1(n12934), .A2(n12933), .ZN(n14768) );
  NAND2_X1 U16011 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12935) );
  OAI211_X1 U16012 ( .C1(n14611), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12953), .B(
        n12935), .ZN(n12936) );
  OAI21_X1 U16013 ( .B1(n12952), .B2(P1_EBX_REG_17__SCAN_IN), .A(n12936), .ZN(
        n16049) );
  MUX2_X1 U16014 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12938) );
  NAND2_X1 U16015 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12937) );
  NOR2_X2 U16016 ( .A1(n9693), .A2(n14751), .ZN(n14752) );
  INV_X1 U16017 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U16018 ( .A1(n12961), .A2(n14818), .ZN(n12941) );
  NAND2_X1 U16019 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12939) );
  OAI211_X1 U16020 ( .C1(n14611), .C2(P1_EBX_REG_19__SCAN_IN), .A(n12953), .B(
        n12939), .ZN(n12940) );
  AND2_X2 U16021 ( .A1(n14752), .A2(n14735), .ZN(n14737) );
  MUX2_X1 U16022 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12943) );
  NAND2_X1 U16023 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12942) );
  NAND2_X1 U16024 ( .A1(n12943), .A2(n12942), .ZN(n14724) );
  INV_X1 U16025 ( .A(n12899), .ZN(n12962) );
  NAND2_X1 U16026 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12944) );
  OAI211_X1 U16027 ( .C1(n14611), .C2(P1_EBX_REG_21__SCAN_IN), .A(n12953), .B(
        n12944), .ZN(n12945) );
  OAI21_X1 U16028 ( .B1(n12952), .B2(P1_EBX_REG_21__SCAN_IN), .A(n12945), .ZN(
        n14712) );
  INV_X1 U16029 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U16030 ( .A1(n12946), .A2(n14812), .ZN(n12949) );
  INV_X1 U16031 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U16032 ( .A1(n12953), .A2(n16189), .ZN(n12947) );
  OAI211_X1 U16033 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n14611), .A(n12947), .B(
        n12962), .ZN(n12948) );
  AND2_X1 U16034 ( .A1(n12949), .A2(n12948), .ZN(n14697) );
  NAND2_X1 U16035 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12950) );
  OAI211_X1 U16036 ( .C1(n14611), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12953), .B(
        n12950), .ZN(n12951) );
  OAI21_X1 U16037 ( .B1(n12952), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12951), .ZN(
        n14688) );
  MUX2_X1 U16038 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12955) );
  NAND2_X1 U16039 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12954) );
  NAND2_X1 U16040 ( .A1(n12955), .A2(n12954), .ZN(n14674) );
  INV_X1 U16041 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U16042 ( .A1(n12961), .A2(n14808), .ZN(n12958) );
  NAND2_X1 U16043 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12956) );
  OAI211_X1 U16044 ( .C1(n14611), .C2(P1_EBX_REG_25__SCAN_IN), .A(n12953), .B(
        n12956), .ZN(n12957) );
  AND2_X1 U16045 ( .A1(n12958), .A2(n12957), .ZN(n14663) );
  MUX2_X1 U16046 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12960) );
  NAND2_X1 U16047 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12959) );
  NAND2_X1 U16048 ( .A1(n12960), .A2(n12959), .ZN(n14633) );
  INV_X1 U16049 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14805) );
  NAND2_X1 U16050 ( .A1(n12961), .A2(n14805), .ZN(n12965) );
  NAND2_X1 U16051 ( .A1(n12962), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12963) );
  OAI211_X1 U16052 ( .C1(n14611), .C2(P1_EBX_REG_27__SCAN_IN), .A(n12953), .B(
        n12963), .ZN(n12964) );
  AND2_X1 U16053 ( .A1(n12965), .A2(n12964), .ZN(n14635) );
  AND2_X1 U16054 ( .A1(n14633), .A2(n14635), .ZN(n12966) );
  MUX2_X1 U16055 ( .A(n12967), .B(n12953), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12969) );
  NAND2_X1 U16056 ( .A1(n12882), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12968) );
  AND2_X1 U16057 ( .A1(n12969), .A2(n12968), .ZN(n14254) );
  OR2_X1 U16058 ( .A1(n12927), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12970) );
  OR2_X1 U16059 ( .A1(n14611), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U16060 ( .A1(n12970), .A2(n12971), .ZN(n14257) );
  MUX2_X1 U16061 ( .A(n14257), .B(n12971), .S(n12899), .Z(n12972) );
  NOR2_X2 U16062 ( .A1(n14256), .A2(n12972), .ZN(n14610) );
  INV_X1 U16063 ( .A(n14610), .ZN(n12974) );
  NAND2_X1 U16064 ( .A1(n14256), .A2(n12972), .ZN(n12973) );
  NAND2_X1 U16065 ( .A1(n12974), .A2(n12973), .ZN(n15081) );
  INV_X1 U16066 ( .A(n15081), .ZN(n12976) );
  INV_X1 U16067 ( .A(n20265), .ZN(n12975) );
  NOR2_X1 U16068 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12979) );
  NOR4_X1 U16069 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12978) );
  NAND4_X1 U16070 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12979), .A4(n12978), .ZN(n12991) );
  NOR2_X1 U16071 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12991), .ZN(n16692)
         );
  INV_X1 U16072 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21068) );
  NOR3_X1 U16073 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21068), .ZN(n12981) );
  NOR4_X1 U16074 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12980)
         );
  NAND4_X1 U16075 ( .A1(n14260), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12981), .A4(
        n12980), .ZN(U214) );
  NOR4_X1 U16076 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12985) );
  NOR4_X1 U16077 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12984) );
  NOR4_X1 U16078 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12983) );
  NOR4_X1 U16079 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12982) );
  NAND4_X1 U16080 ( .A1(n12985), .A2(n12984), .A3(n12983), .A4(n12982), .ZN(
        n12990) );
  NOR4_X1 U16081 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12988) );
  NOR4_X1 U16082 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12987) );
  NOR4_X1 U16083 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12986) );
  INV_X1 U16084 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20049) );
  NAND4_X1 U16085 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n20049), .ZN(
        n12989) );
  NOR2_X1 U16086 ( .A1(n19451), .A2(n12991), .ZN(n16605) );
  NAND2_X1 U16087 ( .A1(n16605), .A2(U214), .ZN(U212) );
  INV_X1 U16088 ( .A(n12993), .ZN(n12995) );
  INV_X1 U16089 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12994) );
  NAND2_X1 U16090 ( .A1(n12995), .A2(n12994), .ZN(n16029) );
  INV_X1 U16091 ( .A(n16029), .ZN(n20954) );
  OAI21_X1 U16092 ( .B1(n9654), .B2(n20954), .A(n12996), .ZN(n13001) );
  OR2_X1 U16093 ( .A1(n13326), .A2(n20954), .ZN(n13899) );
  NAND2_X1 U16094 ( .A1(n13899), .A2(n20953), .ZN(n12998) );
  OAI211_X1 U16095 ( .C1(n11621), .C2(n12998), .A(n13900), .B(n12997), .ZN(
        n12999) );
  INV_X1 U16096 ( .A(n14596), .ZN(n14604) );
  NAND2_X1 U16097 ( .A1(n12999), .A2(n14604), .ZN(n13000) );
  MUX2_X1 U16098 ( .A(n13001), .B(n13000), .S(n12869), .Z(n13009) );
  INV_X1 U16099 ( .A(n13002), .ZN(n13007) );
  AOI21_X1 U16100 ( .B1(n11628), .B2(n13326), .A(n11635), .ZN(n13003) );
  AND2_X1 U16101 ( .A1(n13004), .A2(n13003), .ZN(n13020) );
  OR2_X1 U16102 ( .A1(n13005), .A2(n13020), .ZN(n13006) );
  NAND2_X1 U16103 ( .A1(n13007), .A2(n13006), .ZN(n13368) );
  NAND3_X1 U16104 ( .A1(n14596), .A2(n13663), .A3(n13326), .ZN(n13008) );
  NAND3_X1 U16105 ( .A1(n13009), .A2(n13368), .A3(n13008), .ZN(n13010) );
  OAI211_X1 U16106 ( .C1(n13013), .C2(n13012), .A(n14595), .B(n14594), .ZN(
        n13014) );
  NOR2_X1 U16107 ( .A1(n13011), .A2(n13014), .ZN(n13015) );
  NAND2_X1 U16108 ( .A1(n13016), .A2(n15061), .ZN(n14914) );
  AND3_X1 U16109 ( .A1(n12992), .A2(n20375), .A3(n14914), .ZN(n13062) );
  INV_X1 U16110 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16207) );
  NAND2_X1 U16111 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16217) );
  NOR3_X1 U16112 ( .A1(n12923), .A2(n16207), .A3(n16217), .ZN(n15148) );
  NAND2_X1 U16113 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15148), .ZN(
        n13034) );
  INV_X1 U16114 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16296) );
  NOR2_X1 U16115 ( .A1(n14034), .A2(n16296), .ZN(n16271) );
  NAND2_X1 U16116 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16271), .ZN(
        n16266) );
  OR3_X1 U16117 ( .A1(n12908), .A2(n16272), .A3(n16266), .ZN(n15159) );
  NOR2_X1 U16118 ( .A1(n20359), .A2(n20364), .ZN(n20354) );
  AND2_X1 U16119 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20354), .ZN(
        n14032) );
  INV_X1 U16120 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20368) );
  INV_X1 U16121 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20367) );
  OAI21_X1 U16122 ( .B1(n20368), .B2(n20367), .A(n20380), .ZN(n14031) );
  NAND2_X1 U16123 ( .A1(n14032), .A2(n14031), .ZN(n16265) );
  NOR2_X1 U16124 ( .A1(n15159), .A2(n16265), .ZN(n16246) );
  NAND3_X1 U16125 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16246), .ZN(n13045) );
  OR2_X1 U16126 ( .A1(n16241), .A2(n13045), .ZN(n15147) );
  NOR2_X1 U16127 ( .A1(n13034), .A2(n15147), .ZN(n13036) );
  OAI21_X1 U16128 ( .B1(n13018), .B2(n20955), .A(n13017), .ZN(n13019) );
  NOR2_X1 U16129 ( .A1(n13020), .A2(n13019), .ZN(n13027) );
  NAND2_X1 U16130 ( .A1(n13021), .A2(n12899), .ZN(n13025) );
  OAI21_X1 U16131 ( .B1(n12869), .B2(n11624), .A(n11567), .ZN(n13022) );
  OAI21_X1 U16132 ( .B1(n13023), .B2(n13022), .A(n13326), .ZN(n13024) );
  AND2_X1 U16133 ( .A1(n13025), .A2(n13024), .ZN(n13026) );
  OAI211_X1 U16134 ( .C1(n13028), .C2(n14603), .A(n13027), .B(n13026), .ZN(
        n13360) );
  MUX2_X1 U16135 ( .A(n13029), .B(n12869), .S(n13900), .Z(n13031) );
  NAND2_X1 U16136 ( .A1(n13031), .A2(n13030), .ZN(n13032) );
  NOR2_X1 U16137 ( .A1(n13360), .A2(n13032), .ZN(n13033) );
  NAND2_X1 U16138 ( .A1(n20351), .A2(n13056), .ZN(n15171) );
  INV_X1 U16139 ( .A(n15171), .ZN(n15182) );
  AOI21_X1 U16140 ( .B1(n15170), .B2(n20368), .A(n15182), .ZN(n16268) );
  NAND3_X1 U16141 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14032), .ZN(n16267) );
  OR2_X1 U16142 ( .A1(n16267), .A2(n15159), .ZN(n16249) );
  NAND2_X1 U16143 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15161) );
  NOR2_X1 U16144 ( .A1(n16249), .A2(n15161), .ZN(n15145) );
  INV_X1 U16145 ( .A(n15145), .ZN(n13044) );
  INV_X1 U16146 ( .A(n13034), .ZN(n13047) );
  NAND2_X1 U16147 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n13047), .ZN(
        n16197) );
  NAND2_X1 U16148 ( .A1(n13002), .A2(n13326), .ZN(n13676) );
  OAI21_X1 U16149 ( .B1(n13044), .B2(n16197), .A(n20379), .ZN(n13035) );
  OAI211_X1 U16150 ( .C1(n13036), .C2(n20369), .A(n16268), .B(n13035), .ZN(
        n16199) );
  INV_X1 U16151 ( .A(n20369), .ZN(n15169) );
  NAND2_X1 U16152 ( .A1(n16269), .A2(n16268), .ZN(n13037) );
  OAI21_X1 U16153 ( .B1(n16199), .B2(n15125), .A(n13037), .ZN(n16190) );
  NOR2_X1 U16154 ( .A1(n15127), .A2(n16189), .ZN(n16196) );
  INV_X1 U16155 ( .A(n16196), .ZN(n13038) );
  NAND2_X1 U16156 ( .A1(n15175), .A2(n13038), .ZN(n13039) );
  NAND2_X1 U16157 ( .A1(n16190), .A2(n13039), .ZN(n16182) );
  NOR2_X1 U16158 ( .A1(n20369), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13040) );
  NAND2_X1 U16159 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13050) );
  NAND2_X1 U16160 ( .A1(n13050), .A2(n20379), .ZN(n13041) );
  OAI21_X1 U16161 ( .B1(n20369), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n13041), .ZN(n13042) );
  NOR2_X1 U16162 ( .A1(n15055), .A2(n13042), .ZN(n15110) );
  INV_X1 U16163 ( .A(n15125), .ZN(n13049) );
  NAND2_X1 U16164 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15170), .ZN(
        n13043) );
  OAI22_X1 U16165 ( .A1(n20369), .A2(n13045), .B1(n13044), .B2(n13043), .ZN(
        n15134) );
  AND2_X1 U16166 ( .A1(n15183), .A2(n15145), .ZN(n13046) );
  NAND2_X1 U16167 ( .A1(n13049), .A2(n13048), .ZN(n15116) );
  INV_X1 U16168 ( .A(n13050), .ZN(n13051) );
  NAND2_X1 U16169 ( .A1(n14926), .A2(n13051), .ZN(n13052) );
  NOR2_X1 U16170 ( .A1(n15116), .A2(n13052), .ZN(n15107) );
  INV_X1 U16171 ( .A(n15107), .ZN(n13053) );
  AOI21_X1 U16172 ( .B1(n15110), .B2(n13053), .A(n15061), .ZN(n13061) );
  XNOR2_X1 U16173 ( .A(n14665), .B(n14633), .ZN(n14806) );
  OAI22_X1 U16174 ( .A1(n9686), .A2(n13326), .B1(n11682), .B2(n13012), .ZN(
        n13054) );
  INV_X1 U16175 ( .A(n13054), .ZN(n13055) );
  INV_X1 U16176 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n13057) );
  NOR2_X1 U16177 ( .A1(n20351), .A2(n13057), .ZN(n14915) );
  INV_X1 U16178 ( .A(n14915), .ZN(n13059) );
  INV_X1 U16179 ( .A(n15116), .ZN(n16184) );
  NAND3_X1 U16180 ( .A1(n16184), .A2(n15060), .A3(n15061), .ZN(n13058) );
  OAI211_X1 U16181 ( .C1(n14806), .C2(n20352), .A(n13059), .B(n13058), .ZN(
        n13060) );
  OR3_X1 U16182 ( .A1(n13062), .A2(n13061), .A3(n13060), .ZN(P1_U3005) );
  AOI21_X1 U16183 ( .B1(n16418), .B2(n13069), .A(n15257), .ZN(n16405) );
  AOI21_X1 U16184 ( .B1(n16430), .B2(n13068), .A(n13070), .ZN(n16424) );
  AOI21_X1 U16185 ( .B1(n16438), .B2(n13067), .A(n13063), .ZN(n19258) );
  AOI21_X1 U16186 ( .B1(n16454), .B2(n13065), .A(n9695), .ZN(n16439) );
  AOI21_X1 U16187 ( .B1(n13807), .B2(n13064), .A(n13066), .ZN(n13860) );
  OAI22_X1 U16188 ( .A1(n19097), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19330) );
  INV_X1 U16189 ( .A(n19330), .ZN(n15909) );
  AOI22_X1 U16190 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19441), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19097), .ZN(n15908) );
  NOR2_X1 U16191 ( .A1(n15909), .A2(n15908), .ZN(n15907) );
  OAI21_X1 U16192 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13064), .ZN(n15376) );
  NAND2_X1 U16193 ( .A1(n15907), .A2(n15376), .ZN(n13858) );
  NOR2_X1 U16194 ( .A1(n13860), .A2(n13858), .ZN(n19287) );
  OAI21_X1 U16195 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13066), .A(
        n13065), .ZN(n19431) );
  NAND2_X1 U16196 ( .A1(n19287), .A2(n19431), .ZN(n13842) );
  NOR2_X1 U16197 ( .A1(n16439), .A2(n13842), .ZN(n19270) );
  OAI21_X1 U16198 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9695), .A(
        n13067), .ZN(n19271) );
  NAND2_X1 U16199 ( .A1(n19270), .A2(n19271), .ZN(n19256) );
  NOR2_X1 U16200 ( .A1(n19258), .A2(n19256), .ZN(n19248) );
  OAI21_X1 U16201 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13063), .A(
        n13068), .ZN(n19249) );
  NAND2_X1 U16202 ( .A1(n19248), .A2(n19249), .ZN(n15359) );
  NOR2_X1 U16203 ( .A1(n16424), .A2(n15359), .ZN(n19238) );
  OAI21_X1 U16204 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13070), .A(
        n13069), .ZN(n19239) );
  NAND2_X1 U16205 ( .A1(n19238), .A2(n19239), .ZN(n13073) );
  NAND4_X1 U16206 ( .A1(n19884), .A2(n19097), .A3(n20098), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19289) );
  INV_X1 U16207 ( .A(n19289), .ZN(n19306) );
  NAND2_X1 U16208 ( .A1(n19257), .A2(n19306), .ZN(n19329) );
  AOI211_X1 U16209 ( .C1(n16405), .C2(n13073), .A(n19227), .B(n19329), .ZN(
        n13097) );
  AND2_X1 U16210 ( .A1(n10340), .A2(n13119), .ZN(n13127) );
  NAND2_X1 U16211 ( .A1(n20150), .A2(n20098), .ZN(n13091) );
  INV_X1 U16212 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15384) );
  NAND2_X1 U16213 ( .A1(n13091), .A2(n15384), .ZN(n13074) );
  AOI22_X1 U16214 ( .A1(n14487), .A2(n13074), .B1(n13500), .B2(n20098), .ZN(
        n13075) );
  AND2_X2 U16215 ( .A1(n13127), .A2(n13075), .ZN(n19311) );
  INV_X1 U16216 ( .A(n19311), .ZN(n19180) );
  NOR2_X1 U16217 ( .A1(n19854), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19686) );
  INV_X1 U16218 ( .A(n19686), .ZN(n13076) );
  NOR2_X1 U16219 ( .A1(n13077), .A2(n13076), .ZN(n16533) );
  NAND2_X1 U16220 ( .A1(n16466), .A2(n19289), .ZN(n13078) );
  OR2_X1 U16221 ( .A1(n16533), .A2(n13078), .ZN(n13079) );
  NAND2_X1 U16222 ( .A1(n19262), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19297) );
  OAI22_X1 U16223 ( .A1(n13630), .A2(n19180), .B1(n16418), .B2(n19297), .ZN(
        n13096) );
  AND2_X1 U16224 ( .A1(n19098), .A2(n13080), .ZN(n13090) );
  AND2_X1 U16225 ( .A1(n13091), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13081) );
  AND3_X1 U16226 ( .A1(n13082), .A2(n20098), .A3(n13500), .ZN(n13612) );
  AOI21_X1 U16227 ( .B1(n13085), .B2(n13083), .A(n13084), .ZN(n19345) );
  AOI22_X1 U16228 ( .A1(n13086), .A2(n19317), .B1(n19305), .B2(n19345), .ZN(
        n13087) );
  OAI211_X1 U16229 ( .C1(n11064), .C2(n19262), .A(n13087), .B(n19178), .ZN(
        n13095) );
  OAI21_X1 U16230 ( .B1(n13556), .B2(n13089), .A(n13637), .ZN(n16411) );
  INV_X1 U16231 ( .A(n13090), .ZN(n13092) );
  INV_X1 U16232 ( .A(n16405), .ZN(n13093) );
  NOR2_X1 U16233 ( .A1(n19257), .A2(n19289), .ZN(n19322) );
  INV_X1 U16234 ( .A(n19322), .ZN(n19310) );
  OAI22_X1 U16235 ( .A1(n16411), .A2(n19320), .B1(n13093), .B2(n19310), .ZN(
        n13094) );
  OR4_X1 U16236 ( .A1(n13097), .A2(n13096), .A3(n13095), .A4(n13094), .ZN(
        P2_U2844) );
  OAI21_X1 U16237 ( .B1(n13100), .B2(n13099), .A(n13098), .ZN(n13101) );
  INV_X1 U16238 ( .A(n13101), .ZN(n13252) );
  AOI22_X1 U16239 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19420), .B1(n16519), 
        .B2(n13252), .ZN(n13102) );
  OAI21_X1 U16240 ( .B1(n13103), .B2(n19442), .A(n13102), .ZN(n13118) );
  NOR2_X1 U16241 ( .A1(n16527), .A2(n15374), .ZN(n13117) );
  INV_X1 U16242 ( .A(n13104), .ZN(n13876) );
  NOR2_X1 U16243 ( .A1(n13105), .A2(n13876), .ZN(n13114) );
  INV_X1 U16244 ( .A(n13114), .ZN(n13108) );
  XNOR2_X1 U16245 ( .A(n13107), .B(n13106), .ZN(n13248) );
  OAI22_X1 U16246 ( .A1(n13108), .A2(n15812), .B1(n16524), .B2(n13248), .ZN(
        n13116) );
  OR2_X1 U16247 ( .A1(n13110), .A2(n13109), .ZN(n13112) );
  NAND2_X1 U16248 ( .A1(n13112), .A2(n13111), .ZN(n20110) );
  INV_X1 U16249 ( .A(n20110), .ZN(n13113) );
  OAI22_X1 U16250 ( .A1(n13114), .A2(n15814), .B1(n16526), .B2(n13113), .ZN(
        n13115) );
  OR4_X1 U16251 ( .A1(n13118), .A2(n13117), .A3(n13116), .A4(n13115), .ZN(
        P2_U3044) );
  INV_X1 U16252 ( .A(n13119), .ZN(n13120) );
  NOR2_X1 U16253 ( .A1(n13587), .A2(n13120), .ZN(n19327) );
  INV_X1 U16254 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13121) );
  INV_X1 U16255 ( .A(n13127), .ZN(n13126) );
  OAI211_X1 U16256 ( .C1(n19327), .C2(n13121), .A(n19096), .B(n13126), .ZN(
        P2_U2814) );
  INV_X1 U16257 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13125) );
  INV_X1 U16258 ( .A(n13287), .ZN(n13580) );
  NOR2_X1 U16259 ( .A1(n13122), .A2(n20029), .ZN(n13286) );
  INV_X1 U16260 ( .A(n13579), .ZN(n13123) );
  NOR4_X1 U16261 ( .A1(n13580), .A2(n13286), .A3(n13500), .A4(n13123), .ZN(
        n13585) );
  NOR2_X1 U16262 ( .A1(n13585), .A2(n13508), .ZN(n20143) );
  OAI21_X1 U16263 ( .B1(n13125), .B2(n20143), .A(n13124), .ZN(P2_U2819) );
  OAI21_X2 U16264 ( .B1(n13126), .B2(n20029), .A(n13219), .ZN(n13177) );
  INV_X1 U16265 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13129) );
  NAND3_X1 U16266 ( .A1(n13127), .A2(n14487), .A3(n20150), .ZN(n13171) );
  AOI22_X1 U16267 ( .A1(n19453), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19451), .ZN(n19486) );
  NOR2_X1 U16268 ( .A1(n13171), .A2(n19486), .ZN(n13147) );
  AOI21_X1 U16269 ( .B1(n13168), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13147), .ZN(
        n13128) );
  OAI21_X1 U16270 ( .B1(n13177), .B2(n13129), .A(n13128), .ZN(P2_U2957) );
  INV_X1 U16271 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13131) );
  INV_X1 U16272 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16653) );
  INV_X1 U16273 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18431) );
  OAI22_X1 U16274 ( .A1(n19451), .A2(n16653), .B1(n18431), .B2(n19453), .ZN(
        n13788) );
  INV_X1 U16275 ( .A(n13788), .ZN(n19480) );
  NOR2_X1 U16276 ( .A1(n13171), .A2(n19480), .ZN(n13141) );
  AOI21_X1 U16277 ( .B1(n13168), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13141), .ZN(
        n13130) );
  OAI21_X1 U16278 ( .B1(n13177), .B2(n13131), .A(n13130), .ZN(P2_U2956) );
  INV_X1 U16279 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13133) );
  AOI22_X1 U16280 ( .A1(n19453), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19451), .ZN(n19475) );
  NOR2_X1 U16281 ( .A1(n13171), .A2(n19475), .ZN(n13134) );
  AOI21_X1 U16282 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n13168), .A(n13134), .ZN(
        n13132) );
  OAI21_X1 U16283 ( .B1(n13177), .B2(n13133), .A(n13132), .ZN(P2_U2970) );
  INV_X1 U16284 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13136) );
  AOI21_X1 U16285 ( .B1(n13168), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13134), .ZN(
        n13135) );
  OAI21_X1 U16286 ( .B1(n13177), .B2(n13136), .A(n13135), .ZN(P2_U2955) );
  INV_X1 U16287 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13138) );
  AOI22_X1 U16288 ( .A1(n19453), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19451), .ZN(n19467) );
  NOR2_X1 U16289 ( .A1(n13171), .A2(n19467), .ZN(n13150) );
  AOI21_X1 U16290 ( .B1(n13168), .B2(P2_EAX_REG_1__SCAN_IN), .A(n13150), .ZN(
        n13137) );
  OAI21_X1 U16291 ( .B1(n13177), .B2(n13138), .A(n13137), .ZN(P2_U2968) );
  INV_X1 U16292 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13140) );
  AOI22_X1 U16293 ( .A1(n19453), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19451), .ZN(n19471) );
  NOR2_X1 U16294 ( .A1(n13171), .A2(n19471), .ZN(n13144) );
  AOI21_X1 U16295 ( .B1(n13168), .B2(P2_EAX_REG_2__SCAN_IN), .A(n13144), .ZN(
        n13139) );
  OAI21_X1 U16296 ( .B1(n13177), .B2(n13140), .A(n13139), .ZN(P2_U2969) );
  INV_X1 U16297 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13143) );
  AOI21_X1 U16298 ( .B1(n13168), .B2(P2_EAX_REG_4__SCAN_IN), .A(n13141), .ZN(
        n13142) );
  OAI21_X1 U16299 ( .B1(n13177), .B2(n13143), .A(n13142), .ZN(P2_U2971) );
  INV_X1 U16300 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13146) );
  AOI21_X1 U16301 ( .B1(n13168), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13144), .ZN(
        n13145) );
  OAI21_X1 U16302 ( .B1(n13177), .B2(n13146), .A(n13145), .ZN(P2_U2954) );
  INV_X1 U16303 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13149) );
  AOI21_X1 U16304 ( .B1(n13168), .B2(P2_EAX_REG_5__SCAN_IN), .A(n13147), .ZN(
        n13148) );
  OAI21_X1 U16305 ( .B1(n13177), .B2(n13149), .A(n13148), .ZN(P2_U2972) );
  INV_X1 U16306 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13152) );
  AOI21_X1 U16307 ( .B1(n13168), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13150), .ZN(
        n13151) );
  OAI21_X1 U16308 ( .B1(n13177), .B2(n13152), .A(n13151), .ZN(P2_U2953) );
  INV_X1 U16309 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n13155) );
  AOI22_X1 U16310 ( .A1(n19453), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19451), .ZN(n15460) );
  INV_X1 U16311 ( .A(n15460), .ZN(n13153) );
  NAND2_X1 U16312 ( .A1(n13204), .A2(n13153), .ZN(n13208) );
  NAND2_X1 U16313 ( .A1(n13168), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n13154) );
  OAI211_X1 U16314 ( .C1(n13177), .C2(n13155), .A(n13208), .B(n13154), .ZN(
        P2_U2979) );
  INV_X1 U16315 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n13159) );
  INV_X1 U16316 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16643) );
  NOR2_X1 U16317 ( .A1(n19451), .A2(n16643), .ZN(n13156) );
  AOI21_X1 U16318 ( .B1(n13201), .B2(BUF2_REG_10__SCAN_IN), .A(n13156), .ZN(
        n15477) );
  INV_X1 U16319 ( .A(n15477), .ZN(n13157) );
  NAND2_X1 U16320 ( .A1(n13204), .A2(n13157), .ZN(n13189) );
  NAND2_X1 U16321 ( .A1(n13168), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n13158) );
  OAI211_X1 U16322 ( .C1(n13177), .C2(n13159), .A(n13189), .B(n13158), .ZN(
        P2_U2977) );
  INV_X1 U16323 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13164) );
  NAND2_X1 U16324 ( .A1(n19451), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13162) );
  INV_X1 U16325 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13160) );
  OR2_X1 U16326 ( .A1(n19451), .A2(n13160), .ZN(n13161) );
  NAND2_X1 U16327 ( .A1(n13162), .A2(n13161), .ZN(n15499) );
  NAND2_X1 U16328 ( .A1(n13204), .A2(n15499), .ZN(n13210) );
  NAND2_X1 U16329 ( .A1(n13168), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n13163) );
  OAI211_X1 U16330 ( .C1(n13177), .C2(n13164), .A(n13210), .B(n13163), .ZN(
        P2_U2974) );
  INV_X1 U16331 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n13170) );
  INV_X1 U16332 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13165) );
  OR2_X1 U16333 ( .A1(n19451), .A2(n13165), .ZN(n13167) );
  NAND2_X1 U16334 ( .A1(n13201), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13166) );
  NAND2_X1 U16335 ( .A1(n13167), .A2(n13166), .ZN(n15495) );
  NAND2_X1 U16336 ( .A1(n13204), .A2(n15495), .ZN(n13195) );
  NAND2_X1 U16337 ( .A1(n13168), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n13169) );
  OAI211_X1 U16338 ( .C1(n13177), .C2(n13170), .A(n13195), .B(n13169), .ZN(
        P2_U2975) );
  INV_X1 U16339 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13172) );
  AOI22_X1 U16340 ( .A1(n19453), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19451), .ZN(n19340) );
  INV_X1 U16341 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19336) );
  OAI222_X1 U16342 ( .A1(n13172), .A2(n13177), .B1(n13171), .B2(n19340), .C1(
        n19336), .C2(n13219), .ZN(P2_U2982) );
  INV_X1 U16343 ( .A(n14600), .ZN(n13173) );
  AND2_X1 U16344 ( .A1(n13002), .A2(n13173), .ZN(n14607) );
  NAND2_X1 U16345 ( .A1(n14607), .A2(n13373), .ZN(n13264) );
  INV_X1 U16346 ( .A(n13264), .ZN(n13176) );
  INV_X1 U16347 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13175) );
  INV_X1 U16348 ( .A(n13373), .ZN(n20162) );
  AND2_X1 U16349 ( .A1(n20810), .A2(n13651), .ZN(n13263) );
  INV_X1 U16350 ( .A(n13263), .ZN(n13174) );
  OAI211_X1 U16351 ( .C1(n13176), .C2(n13175), .A(n13296), .B(n13174), .ZN(
        P1_U2801) );
  INV_X1 U16352 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19391) );
  INV_X1 U16353 ( .A(n13177), .ZN(n13216) );
  NAND2_X1 U16354 ( .A1(n13216), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13180) );
  INV_X1 U16355 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16636) );
  OR2_X1 U16356 ( .A1(n19451), .A2(n16636), .ZN(n13179) );
  NAND2_X1 U16357 ( .A1(n19451), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13178) );
  NAND2_X1 U16358 ( .A1(n13179), .A2(n13178), .ZN(n19341) );
  NAND2_X1 U16359 ( .A1(n13204), .A2(n19341), .ZN(n13217) );
  OAI211_X1 U16360 ( .C1(n19391), .C2(n13219), .A(n13180), .B(n13217), .ZN(
        P2_U2981) );
  NAND2_X1 U16361 ( .A1(n13216), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U16362 ( .A1(n19453), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19451), .ZN(n19459) );
  INV_X1 U16363 ( .A(n19459), .ZN(n13991) );
  NAND2_X1 U16364 ( .A1(n13204), .A2(n13991), .ZN(n13197) );
  OAI211_X1 U16365 ( .C1(n13219), .C2(n13182), .A(n13181), .B(n13197), .ZN(
        P2_U2967) );
  INV_X1 U16366 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n13188) );
  NAND2_X1 U16367 ( .A1(n13216), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13187) );
  INV_X1 U16368 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13183) );
  OR2_X1 U16369 ( .A1(n19451), .A2(n13183), .ZN(n13185) );
  NAND2_X1 U16370 ( .A1(n19451), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13184) );
  AND2_X1 U16371 ( .A1(n13185), .A2(n13184), .ZN(n19347) );
  INV_X1 U16372 ( .A(n19347), .ZN(n13186) );
  NAND2_X1 U16373 ( .A1(n13204), .A2(n13186), .ZN(n13212) );
  OAI211_X1 U16374 ( .C1(n13219), .C2(n13188), .A(n13187), .B(n13212), .ZN(
        P2_U2978) );
  INV_X1 U16375 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15476) );
  NAND2_X1 U16376 ( .A1(n13216), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13190) );
  OAI211_X1 U16377 ( .C1(n13219), .C2(n15476), .A(n13190), .B(n13189), .ZN(
        P2_U2962) );
  INV_X1 U16378 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19400) );
  NAND2_X1 U16379 ( .A1(n13216), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13193) );
  INV_X1 U16380 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16645) );
  OR2_X1 U16381 ( .A1(n19451), .A2(n16645), .ZN(n13192) );
  NAND2_X1 U16382 ( .A1(n13201), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13191) );
  NAND2_X1 U16383 ( .A1(n13192), .A2(n13191), .ZN(n15487) );
  NAND2_X1 U16384 ( .A1(n13204), .A2(n15487), .ZN(n13206) );
  OAI211_X1 U16385 ( .C1(n19400), .C2(n13219), .A(n13193), .B(n13206), .ZN(
        P2_U2976) );
  INV_X1 U16386 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19348) );
  NAND2_X1 U16387 ( .A1(n13216), .A2(P2_LWORD_REG_6__SCAN_IN), .ZN(n13194) );
  OAI22_X1 U16388 ( .A1(n19451), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19453), .ZN(n19489) );
  INV_X1 U16389 ( .A(n19489), .ZN(n16363) );
  NAND2_X1 U16390 ( .A1(n13204), .A2(n16363), .ZN(n13199) );
  OAI211_X1 U16391 ( .C1(n13219), .C2(n19348), .A(n13194), .B(n13199), .ZN(
        P2_U2973) );
  INV_X1 U16392 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15492) );
  NAND2_X1 U16393 ( .A1(n13216), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13196) );
  OAI211_X1 U16394 ( .C1(n13219), .C2(n15492), .A(n13196), .B(n13195), .ZN(
        P2_U2960) );
  INV_X1 U16395 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U16396 ( .A1(n13216), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13198) );
  OAI211_X1 U16397 ( .C1(n13219), .C2(n13381), .A(n13198), .B(n13197), .ZN(
        P2_U2952) );
  INV_X1 U16398 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13235) );
  NAND2_X1 U16399 ( .A1(n13216), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13200) );
  OAI211_X1 U16400 ( .C1(n13219), .C2(n13235), .A(n13200), .B(n13199), .ZN(
        P2_U2958) );
  INV_X1 U16401 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19393) );
  NAND2_X1 U16402 ( .A1(n13216), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13205) );
  INV_X1 U16403 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16638) );
  OR2_X1 U16404 ( .A1(n19451), .A2(n16638), .ZN(n13203) );
  NAND2_X1 U16405 ( .A1(n13201), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U16406 ( .A1(n13203), .A2(n13202), .ZN(n15452) );
  NAND2_X1 U16407 ( .A1(n13204), .A2(n15452), .ZN(n13214) );
  OAI211_X1 U16408 ( .C1(n19393), .C2(n13219), .A(n13205), .B(n13214), .ZN(
        P2_U2980) );
  INV_X1 U16409 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13226) );
  NAND2_X1 U16410 ( .A1(n13216), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13207) );
  OAI211_X1 U16411 ( .C1(n13226), .C2(n13219), .A(n13207), .B(n13206), .ZN(
        P2_U2961) );
  INV_X1 U16412 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13230) );
  NAND2_X1 U16413 ( .A1(n13216), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13209) );
  OAI211_X1 U16414 ( .C1(n13219), .C2(n13230), .A(n13209), .B(n13208), .ZN(
        P2_U2964) );
  INV_X1 U16415 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13232) );
  NAND2_X1 U16416 ( .A1(n13216), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13211) );
  OAI211_X1 U16417 ( .C1(n13219), .C2(n13232), .A(n13211), .B(n13210), .ZN(
        P2_U2959) );
  INV_X1 U16418 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13239) );
  NAND2_X1 U16419 ( .A1(n13216), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13213) );
  OAI211_X1 U16420 ( .C1(n13219), .C2(n13239), .A(n13213), .B(n13212), .ZN(
        P2_U2963) );
  INV_X1 U16421 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13228) );
  NAND2_X1 U16422 ( .A1(n13216), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13215) );
  OAI211_X1 U16423 ( .C1(n13228), .C2(n13219), .A(n13215), .B(n13214), .ZN(
        P2_U2965) );
  INV_X1 U16424 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U16425 ( .A1(n13216), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13218) );
  OAI211_X1 U16426 ( .C1(n13388), .C2(n13219), .A(n13218), .B(n13217), .ZN(
        P2_U2966) );
  OR2_X1 U16427 ( .A1(n13587), .A2(n13508), .ZN(n13220) );
  OAI21_X1 U16428 ( .B1(n13221), .B2(n13220), .A(n13219), .ZN(n13222) );
  INV_X1 U16429 ( .A(n20035), .ZN(n20151) );
  INV_X1 U16430 ( .A(n13223), .ZN(n13224) );
  NAND2_X1 U16431 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20127) );
  NOR2_X1 U16432 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20127), .ZN(n19417) );
  AOI22_X1 U16433 ( .A1(n20146), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13225) );
  OAI21_X1 U16434 ( .B1(n13226), .B2(n13387), .A(n13225), .ZN(P2_U2926) );
  AOI22_X1 U16435 ( .A1(n20146), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13227) );
  OAI21_X1 U16436 ( .B1(n13228), .B2(n13387), .A(n13227), .ZN(P2_U2922) );
  AOI22_X1 U16437 ( .A1(n20146), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13229) );
  OAI21_X1 U16438 ( .B1(n13230), .B2(n13387), .A(n13229), .ZN(P2_U2923) );
  AOI22_X1 U16439 ( .A1(n20146), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U16440 ( .B1(n13232), .B2(n13387), .A(n13231), .ZN(P2_U2928) );
  INV_X1 U16441 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15521) );
  AOI22_X1 U16442 ( .A1(n20146), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U16443 ( .B1(n15521), .B2(n13387), .A(n13233), .ZN(P2_U2932) );
  AOI22_X1 U16444 ( .A1(n20146), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13234) );
  OAI21_X1 U16445 ( .B1(n13235), .B2(n13387), .A(n13234), .ZN(P2_U2929) );
  AOI22_X1 U16446 ( .A1(n20146), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13236) );
  OAI21_X1 U16447 ( .B1(n15492), .B2(n13387), .A(n13236), .ZN(P2_U2927) );
  INV_X1 U16448 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U16449 ( .A1(n20146), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13237) );
  OAI21_X1 U16450 ( .B1(n15511), .B2(n13387), .A(n13237), .ZN(P2_U2931) );
  AOI22_X1 U16451 ( .A1(n20146), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U16452 ( .B1(n13239), .B2(n13387), .A(n13238), .ZN(P2_U2924) );
  INV_X1 U16453 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U16454 ( .A1(n20146), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19387), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13240) );
  OAI21_X1 U16455 ( .B1(n15504), .B2(n13387), .A(n13240), .ZN(P2_U2930) );
  OAI21_X1 U16456 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19318), .A(
        n13254), .ZN(n16532) );
  INV_X1 U16457 ( .A(n16532), .ZN(n13244) );
  AOI22_X1 U16458 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13242), .B1(
        n13241), .B2(n10375), .ZN(n16525) );
  OR2_X1 U16459 ( .A1(n19178), .A2(n19115), .ZN(n16530) );
  OAI21_X1 U16460 ( .B1(n19423), .B2(n16525), .A(n16530), .ZN(n13243) );
  AOI21_X1 U16461 ( .B1(n16450), .B2(n13244), .A(n13243), .ZN(n13247) );
  OAI21_X1 U16462 ( .B1(n19421), .B2(n13245), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13246) );
  OAI211_X1 U16463 ( .C1(n15688), .C2(n19321), .A(n13247), .B(n13246), .ZN(
        P2_U3014) );
  OAI22_X1 U16464 ( .A1(n19423), .A2(n13248), .B1(n15371), .B2(n19178), .ZN(
        n13249) );
  AOI21_X1 U16465 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19421), .A(
        n13249), .ZN(n13250) );
  OAI21_X1 U16466 ( .B1(n15376), .B2(n19432), .A(n13250), .ZN(n13251) );
  AOI21_X1 U16467 ( .B1(n16450), .B2(n13252), .A(n13251), .ZN(n13253) );
  OAI21_X1 U16468 ( .B1(n15374), .B2(n15688), .A(n13253), .ZN(P2_U3012) );
  INV_X1 U16469 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13261) );
  XNOR2_X1 U16470 ( .A(n19301), .B(n19441), .ZN(n13255) );
  XNOR2_X1 U16471 ( .A(n13255), .B(n13254), .ZN(n19450) );
  OR2_X1 U16472 ( .A1(n19178), .A2(n13256), .ZN(n19447) );
  OAI21_X1 U16473 ( .B1(n19424), .B2(n19450), .A(n19447), .ZN(n13260) );
  OAI21_X1 U16474 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13258), .A(
        n13257), .ZN(n19435) );
  OAI22_X1 U16475 ( .A1(n19423), .A2(n19435), .B1(n16453), .B2(n13261), .ZN(
        n13259) );
  AOI211_X1 U16476 ( .C1(n16440), .C2(n13261), .A(n13260), .B(n13259), .ZN(
        n13262) );
  OAI21_X1 U16477 ( .B1(n13277), .B2(n15688), .A(n13262), .ZN(P2_U3013) );
  NOR2_X1 U16478 ( .A1(n13263), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13266)
         );
  INV_X1 U16479 ( .A(n14603), .ZN(n14605) );
  OAI21_X1 U16480 ( .B1(n12899), .B2(n14605), .A(n20949), .ZN(n13265) );
  OAI21_X1 U16481 ( .B1(n13266), .B2(n20949), .A(n13265), .ZN(P1_U3487) );
  NAND2_X1 U16482 ( .A1(n13434), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U16483 ( .A1(n13391), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20107), .B2(n20135), .ZN(n13268) );
  NAND2_X1 U16484 ( .A1(n14487), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13270) );
  AND4_X1 U16485 ( .A1(n13269), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13270), 
        .A4(n19854), .ZN(n13271) );
  INV_X1 U16486 ( .A(n13488), .ZN(n13584) );
  NAND2_X1 U16487 ( .A1(n13584), .A2(n13567), .ZN(n13503) );
  NAND2_X1 U16488 ( .A1(n13503), .A2(n13494), .ZN(n13272) );
  INV_X1 U16489 ( .A(n15442), .ZN(n13322) );
  MUX2_X1 U16490 ( .A(n19321), .B(n13274), .S(n13322), .Z(n13275) );
  OAI21_X1 U16491 ( .B1(n20130), .B2(n15450), .A(n13275), .ZN(P2_U2887) );
  NAND2_X1 U16492 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20125), .ZN(
        n19745) );
  NAND2_X1 U16493 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20135), .ZN(
        n19782) );
  NAND2_X1 U16494 ( .A1(n19745), .A2(n19782), .ZN(n19593) );
  AND2_X1 U16495 ( .A1(n20107), .A2(n19593), .ZN(n19531) );
  AOI21_X1 U16496 ( .B1(n13391), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19531), .ZN(n13276) );
  NOR2_X1 U16497 ( .A1(n13434), .A2(n19097), .ZN(n13278) );
  XNOR2_X1 U16498 ( .A(n13314), .B(n13313), .ZN(n13280) );
  NAND2_X1 U16501 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  MUX2_X1 U16502 ( .A(n13277), .B(n10345), .S(n13322), .Z(n13283) );
  OAI21_X1 U16503 ( .B1(n20099), .B2(n15450), .A(n13283), .ZN(P2_U2886) );
  XNOR2_X1 U16504 ( .A(n13285), .B(n13284), .ZN(n19264) );
  AND3_X1 U16505 ( .A1(n13287), .A2(n13579), .A3(n13286), .ZN(n13288) );
  AOI21_X1 U16506 ( .B1(n13488), .B2(n13583), .A(n13288), .ZN(n13505) );
  NAND2_X1 U16507 ( .A1(n13505), .A2(n13289), .ZN(n13290) );
  OR2_X1 U16508 ( .A1(n19379), .A2(n10332), .ZN(n15538) );
  INV_X1 U16509 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19404) );
  INV_X1 U16510 ( .A(n13292), .ZN(n13293) );
  NAND2_X1 U16511 ( .A1(n13434), .A2(n10332), .ZN(n13294) );
  INV_X1 U16512 ( .A(n15499), .ZN(n19501) );
  OAI222_X1 U16513 ( .A1(n19264), .A2(n19351), .B1(n19349), .B2(n19404), .C1(
        n19386), .C2(n19501), .ZN(P2_U2912) );
  AND2_X1 U16514 ( .A1(n11643), .A2(n20948), .ZN(n13295) );
  NAND2_X1 U16515 ( .A1(n13402), .A2(n9654), .ZN(n13458) );
  INV_X1 U16516 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14890) );
  NAND2_X1 U16517 ( .A1(n13402), .A2(n13326), .ZN(n13403) );
  INV_X1 U16518 ( .A(DATAI_15_), .ZN(n13298) );
  INV_X1 U16519 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13297) );
  MUX2_X1 U16520 ( .A(n13298), .B(n13297), .S(n14260), .Z(n14889) );
  INV_X1 U16521 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20273) );
  OAI222_X1 U16522 ( .A1(n13458), .A2(n14890), .B1(n13403), .B2(n14889), .C1(
        n13402), .C2(n20273), .ZN(P1_U2967) );
  NAND2_X1 U16523 ( .A1(n19812), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19456) );
  OAI21_X1 U16524 ( .B1(n19812), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n19456), .ZN(n19594) );
  NOR2_X1 U16525 ( .A1(n19594), .A2(n19969), .ZN(n13299) );
  AOI21_X1 U16526 ( .B1(n13391), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13299), .ZN(n13306) );
  INV_X1 U16527 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13300) );
  AND2_X1 U16528 ( .A1(n13306), .A2(n13394), .ZN(n13301) );
  NAND2_X1 U16529 ( .A1(n13302), .A2(n13301), .ZN(n13311) );
  INV_X1 U16530 ( .A(n13301), .ZN(n13303) );
  OAI22_X1 U16531 ( .A1(n13311), .A2(n13304), .B1(n13303), .B2(n13302), .ZN(
        n13305) );
  NAND2_X1 U16532 ( .A1(n13312), .A2(n13305), .ZN(n13310) );
  INV_X1 U16533 ( .A(n13306), .ZN(n13395) );
  INV_X1 U16534 ( .A(n13307), .ZN(n13389) );
  OAI21_X1 U16535 ( .B1(n13395), .B2(n13389), .A(n13394), .ZN(n13308) );
  OAI21_X1 U16536 ( .B1(n13394), .B2(n13395), .A(n13308), .ZN(n13309) );
  OAI211_X1 U16537 ( .C1(n13312), .C2(n13311), .A(n13310), .B(n13309), .ZN(
        n13319) );
  INV_X1 U16538 ( .A(n13319), .ZN(n13315) );
  OR2_X1 U16539 ( .A1(n13314), .A2(n13313), .ZN(n13318) );
  NAND2_X1 U16540 ( .A1(n21164), .A2(n13318), .ZN(n13320) );
  NAND2_X1 U16541 ( .A1(n13320), .A2(n13319), .ZN(n13321) );
  INV_X1 U16542 ( .A(n20111), .ZN(n13325) );
  INV_X1 U16543 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13323) );
  MUX2_X1 U16544 ( .A(n15374), .B(n13323), .S(n13322), .Z(n13324) );
  OAI21_X1 U16545 ( .B1(n13325), .B2(n15450), .A(n13324), .ZN(P2_U2885) );
  INV_X1 U16546 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13332) );
  OR2_X1 U16547 ( .A1(n13326), .A2(n16029), .ZN(n13327) );
  OR2_X1 U16548 ( .A1(n9686), .A2(n13327), .ZN(n16011) );
  OAI21_X1 U16549 ( .B1(n13676), .B2(n16029), .A(n16011), .ZN(n13330) );
  INV_X1 U16550 ( .A(n13328), .ZN(n13329) );
  NAND2_X1 U16551 ( .A1(n20274), .A2(n13900), .ZN(n13529) );
  NAND2_X1 U16552 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16318) );
  INV_X1 U16553 ( .A(n16318), .ZN(n15188) );
  NAND2_X1 U16554 ( .A1(n20865), .A2(n15188), .ZN(n20272) );
  INV_X2 U16555 ( .A(n20272), .ZN(n20301) );
  NOR2_X4 U16556 ( .A1(n20274), .A2(n20301), .ZN(n16031) );
  AOI22_X1 U16557 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13331) );
  OAI21_X1 U16558 ( .B1(n13332), .B2(n13529), .A(n13331), .ZN(P1_U2914) );
  INV_X1 U16559 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13334) );
  AOI22_X1 U16560 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16561 ( .B1(n13334), .B2(n13529), .A(n13333), .ZN(P1_U2911) );
  INV_X1 U16562 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13336) );
  AOI22_X1 U16563 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13335) );
  OAI21_X1 U16564 ( .B1(n13336), .B2(n13529), .A(n13335), .ZN(P1_U2907) );
  INV_X1 U16565 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U16566 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13337) );
  OAI21_X1 U16567 ( .B1(n13338), .B2(n13529), .A(n13337), .ZN(P1_U2915) );
  INV_X1 U16568 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13340) );
  AOI22_X1 U16569 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13339) );
  OAI21_X1 U16570 ( .B1(n13340), .B2(n13529), .A(n13339), .ZN(P1_U2916) );
  INV_X1 U16571 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U16572 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13341) );
  OAI21_X1 U16573 ( .B1(n13342), .B2(n13529), .A(n13341), .ZN(P1_U2909) );
  INV_X1 U16574 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U16575 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13343) );
  OAI21_X1 U16576 ( .B1(n13344), .B2(n13529), .A(n13343), .ZN(P1_U2920) );
  INV_X1 U16577 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U16578 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13345) );
  OAI21_X1 U16579 ( .B1(n13346), .B2(n13529), .A(n13345), .ZN(P1_U2908) );
  INV_X1 U16580 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U16581 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13347) );
  OAI21_X1 U16582 ( .B1(n13348), .B2(n13529), .A(n13347), .ZN(P1_U2913) );
  INV_X1 U16583 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U16584 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13349) );
  OAI21_X1 U16585 ( .B1(n13350), .B2(n13529), .A(n13349), .ZN(P1_U2912) );
  OR2_X1 U16586 ( .A1(n13352), .A2(n13351), .ZN(n13354) );
  NAND2_X1 U16587 ( .A1(n13354), .A2(n13353), .ZN(n19255) );
  INV_X1 U16588 ( .A(n15495), .ZN(n13355) );
  INV_X1 U16589 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19402) );
  OAI222_X1 U16590 ( .A1(n19255), .A2(n19351), .B1(n13355), .B2(n19386), .C1(
        n19402), .C2(n19349), .ZN(P2_U2911) );
  INV_X1 U16591 ( .A(n13356), .ZN(n13358) );
  NAND2_X1 U16592 ( .A1(n13358), .A2(n13357), .ZN(n13359) );
  NOR2_X1 U16593 ( .A1(n13360), .A2(n13359), .ZN(n13361) );
  AND2_X1 U16594 ( .A1(n12449), .A2(n13361), .ZN(n13679) );
  INV_X1 U16595 ( .A(n13679), .ZN(n15197) );
  NOR2_X1 U16596 ( .A1(n15194), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13362) );
  AOI21_X1 U16597 ( .B1(n11775), .B2(n15197), .A(n13362), .ZN(n15992) );
  INV_X1 U16598 ( .A(n15992), .ZN(n13364) );
  INV_X1 U16599 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20689) );
  OAI22_X1 U16600 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13651), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15199), .ZN(n13363) );
  AOI21_X1 U16601 ( .B1(n13364), .B2(n20937), .A(n13363), .ZN(n13379) );
  AOI21_X1 U16602 ( .B1(n13676), .B2(n11621), .A(n16029), .ZN(n13366) );
  OAI21_X1 U16603 ( .B1(n13366), .B2(n13365), .A(n20953), .ZN(n13367) );
  MUX2_X1 U16604 ( .A(n13658), .B(n13367), .S(n14604), .Z(n13372) );
  OAI21_X1 U16605 ( .B1(n20955), .B2(n13749), .A(n13368), .ZN(n13369) );
  NOR2_X1 U16606 ( .A1(n13370), .A2(n13369), .ZN(n13371) );
  NAND2_X1 U16607 ( .A1(n15993), .A2(n13373), .ZN(n13376) );
  NAND2_X1 U16608 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15188), .ZN(n16322) );
  INV_X1 U16609 ( .A(n16322), .ZN(n13374) );
  NAND2_X1 U16610 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13374), .ZN(n13375) );
  NAND2_X1 U16611 ( .A1(n13376), .A2(n13375), .ZN(n16314) );
  AND2_X1 U16612 ( .A1(n20865), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13377) );
  OR2_X1 U16613 ( .A1(n16314), .A2(n13377), .ZN(n16317) );
  INV_X1 U16614 ( .A(n16317), .ZN(n20940) );
  INV_X1 U16615 ( .A(n13676), .ZN(n15990) );
  AOI21_X1 U16616 ( .B1(n15990), .B2(n20937), .A(n20940), .ZN(n13378) );
  OAI22_X1 U16617 ( .A1(n13379), .A2(n20940), .B1(n13378), .B2(n11353), .ZN(
        P1_U3474) );
  AOI22_X1 U16618 ( .A1(n19417), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13380) );
  OAI21_X1 U16619 ( .B1(n13381), .B2(n13387), .A(n13380), .ZN(P2_U2935) );
  INV_X1 U16620 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U16621 ( .A1(n20146), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13382) );
  OAI21_X1 U16622 ( .B1(n14062), .B2(n13387), .A(n13382), .ZN(P2_U2934) );
  INV_X1 U16623 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13384) );
  AOI22_X1 U16624 ( .A1(n20146), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13383) );
  OAI21_X1 U16625 ( .B1(n13384), .B2(n13387), .A(n13383), .ZN(P2_U2933) );
  AOI22_X1 U16626 ( .A1(n20146), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13385) );
  OAI21_X1 U16627 ( .B1(n15476), .B2(n13387), .A(n13385), .ZN(P2_U2925) );
  AOI22_X1 U16628 ( .A1(n20146), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n19416), .ZN(n13386) );
  OAI21_X1 U16629 ( .B1(n13388), .B2(n13387), .A(n13386), .ZN(P2_U2921) );
  NOR2_X1 U16630 ( .A1(n20116), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19625) );
  INV_X1 U16631 ( .A(n19719), .ZN(n19716) );
  NAND2_X1 U16632 ( .A1(n19456), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13390) );
  AOI21_X1 U16633 ( .B1(n19716), .B2(n13390), .A(n19969), .ZN(n19849) );
  AOI21_X1 U16634 ( .B1(n13391), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19849), .ZN(n13392) );
  NAND2_X1 U16635 ( .A1(n13438), .A2(n13393), .ZN(n13437) );
  INV_X1 U16636 ( .A(n13394), .ZN(n13396) );
  NAND2_X1 U16637 ( .A1(n13396), .A2(n13395), .ZN(n13397) );
  NOR2_X1 U16638 ( .A1(n16512), .A2(n13322), .ZN(n13400) );
  AOI21_X1 U16639 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n13273), .A(n13400), .ZN(
        n13401) );
  OAI21_X1 U16640 ( .B1(n20103), .B2(n15450), .A(n13401), .ZN(P2_U2884) );
  INV_X2 U16641 ( .A(n13402), .ZN(n20326) );
  AOI22_X1 U16642 ( .A1(n20327), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13406) );
  INV_X1 U16643 ( .A(DATAI_4_), .ZN(n13405) );
  NAND2_X1 U16644 ( .A1(n14848), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13404) );
  OAI21_X1 U16645 ( .B1(n14848), .B2(n13405), .A(n13404), .ZN(n14874) );
  NAND2_X1 U16646 ( .A1(n20314), .A2(n14874), .ZN(n13462) );
  NAND2_X1 U16647 ( .A1(n13406), .A2(n13462), .ZN(P1_U2956) );
  AOI22_X1 U16648 ( .A1(n20327), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13409) );
  INV_X1 U16649 ( .A(DATAI_5_), .ZN(n13408) );
  NAND2_X1 U16650 ( .A1(n14260), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13407) );
  OAI21_X1 U16651 ( .B1(n14848), .B2(n13408), .A(n13407), .ZN(n14871) );
  NAND2_X1 U16652 ( .A1(n20314), .A2(n14871), .ZN(n13472) );
  NAND2_X1 U16653 ( .A1(n13409), .A2(n13472), .ZN(P1_U2957) );
  AOI22_X1 U16654 ( .A1(n20327), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13412) );
  INV_X1 U16655 ( .A(DATAI_3_), .ZN(n13411) );
  NAND2_X1 U16656 ( .A1(n14848), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13410) );
  OAI21_X1 U16657 ( .B1(n14260), .B2(n13411), .A(n13410), .ZN(n14877) );
  NAND2_X1 U16658 ( .A1(n20314), .A2(n14877), .ZN(n13464) );
  NAND2_X1 U16659 ( .A1(n13412), .A2(n13464), .ZN(P1_U2955) );
  AOI22_X1 U16660 ( .A1(n20327), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13415) );
  INV_X1 U16661 ( .A(DATAI_7_), .ZN(n13414) );
  NAND2_X1 U16662 ( .A1(n14848), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13413) );
  OAI21_X1 U16663 ( .B1(n14260), .B2(n13414), .A(n13413), .ZN(n14863) );
  NAND2_X1 U16664 ( .A1(n20314), .A2(n14863), .ZN(n13482) );
  NAND2_X1 U16665 ( .A1(n13415), .A2(n13482), .ZN(P1_U2959) );
  AOI22_X1 U16666 ( .A1(n20327), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13418) );
  INV_X1 U16667 ( .A(DATAI_6_), .ZN(n13417) );
  NAND2_X1 U16668 ( .A1(n14848), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13416) );
  OAI21_X1 U16669 ( .B1(n14848), .B2(n13417), .A(n13416), .ZN(n14867) );
  NAND2_X1 U16670 ( .A1(n20314), .A2(n14867), .ZN(n13476) );
  NAND2_X1 U16671 ( .A1(n13418), .A2(n13476), .ZN(P1_U2958) );
  AOI22_X1 U16672 ( .A1(n20327), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20326), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13421) );
  INV_X1 U16673 ( .A(DATAI_11_), .ZN(n13420) );
  NAND2_X1 U16674 ( .A1(n14848), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13419) );
  OAI21_X1 U16675 ( .B1(n14260), .B2(n13420), .A(n13419), .ZN(n14900) );
  NAND2_X1 U16676 ( .A1(n20314), .A2(n14900), .ZN(n13480) );
  NAND2_X1 U16677 ( .A1(n13421), .A2(n13480), .ZN(P1_U2963) );
  AOI21_X1 U16678 ( .B1(n13422), .B2(n13353), .A(n13429), .ZN(n15895) );
  INV_X1 U16679 ( .A(n15895), .ZN(n13424) );
  INV_X1 U16680 ( .A(n15487), .ZN(n13423) );
  OAI222_X1 U16681 ( .A1(n13424), .A2(n19351), .B1(n13423), .B2(n19386), .C1(
        n19400), .C2(n19349), .ZN(P2_U2910) );
  OR2_X1 U16682 ( .A1(n12927), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13426) );
  NAND2_X1 U16683 ( .A1(n13426), .A2(n13425), .ZN(n13894) );
  XOR2_X1 U16684 ( .A(n13428), .B(n13427), .Z(n13914) );
  OAI222_X1 U16685 ( .A1(n13894), .A2(n20265), .B1(n14842), .B2(n13914), .C1(
        n12877), .C2(n20270), .ZN(P1_U2872) );
  OR2_X1 U16686 ( .A1(n13430), .A2(n13429), .ZN(n13431) );
  NAND2_X1 U16687 ( .A1(n13431), .A2(n13083), .ZN(n19244) );
  INV_X1 U16688 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19398) );
  OAI222_X1 U16689 ( .A1(n19244), .A2(n19351), .B1(n15477), .B2(n19386), .C1(
        n19398), .C2(n19349), .ZN(P2_U2909) );
  NAND2_X1 U16690 ( .A1(n13434), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13435) );
  AND2_X1 U16691 ( .A1(n14450), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13439) );
  INV_X1 U16692 ( .A(n13439), .ZN(n13436) );
  NAND2_X1 U16693 ( .A1(n13437), .A2(n13436), .ZN(n13440) );
  NAND2_X1 U16694 ( .A1(n13542), .A2(n13439), .ZN(n13534) );
  OAI21_X1 U16695 ( .B1(n13441), .B2(n13440), .A(n13534), .ZN(n19357) );
  INV_X1 U16696 ( .A(n13449), .ZN(n13442) );
  AOI21_X1 U16697 ( .B1(n13444), .B2(n13443), .A(n13442), .ZN(n19427) );
  INV_X1 U16698 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13445) );
  NOR2_X1 U16699 ( .A1(n15442), .A2(n13445), .ZN(n13446) );
  AOI21_X1 U16700 ( .B1(n19427), .B2(n15442), .A(n13446), .ZN(n13447) );
  OAI21_X1 U16701 ( .B1(n19357), .B2(n15450), .A(n13447), .ZN(P2_U2883) );
  INV_X1 U16702 ( .A(n13534), .ZN(n13535) );
  XNOR2_X1 U16703 ( .A(n13535), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13452) );
  AND2_X1 U16704 ( .A1(n13449), .A2(n13448), .ZN(n13450) );
  OR2_X1 U16705 ( .A1(n13450), .A2(n9770), .ZN(n16448) );
  MUX2_X1 U16706 ( .A(n16448), .B(n10619), .S(n13273), .Z(n13451) );
  OAI21_X1 U16707 ( .B1(n13452), .B2(n15450), .A(n13451), .ZN(P2_U2882) );
  INV_X1 U16708 ( .A(n13453), .ZN(n13454) );
  OAI21_X1 U16709 ( .B1(n13456), .B2(n13455), .A(n13454), .ZN(n13952) );
  INV_X1 U16710 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13457) );
  XNOR2_X1 U16711 ( .A(n13947), .B(n14611), .ZN(n15168) );
  OAI222_X1 U16712 ( .A1(n13952), .A2(n14842), .B1(n13457), .B2(n20270), .C1(
        n20265), .C2(n15168), .ZN(P1_U2871) );
  INV_X2 U16713 ( .A(n13458), .ZN(n20327) );
  AOI22_X1 U16714 ( .A1(n20327), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U16715 ( .A1(n13718), .A2(DATAI_0_), .ZN(n13460) );
  NAND2_X1 U16716 ( .A1(n14848), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13459) );
  AND2_X1 U16717 ( .A1(n13460), .A2(n13459), .ZN(n13739) );
  INV_X1 U16718 ( .A(n13739), .ZN(n14884) );
  NAND2_X1 U16719 ( .A1(n20314), .A2(n14884), .ZN(n13484) );
  NAND2_X1 U16720 ( .A1(n13461), .A2(n13484), .ZN(P1_U2937) );
  AOI22_X1 U16721 ( .A1(n20327), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U16722 ( .A1(n13463), .A2(n13462), .ZN(P1_U2941) );
  AOI22_X1 U16723 ( .A1(n20327), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U16724 ( .A1(n13465), .A2(n13464), .ZN(P1_U2940) );
  AOI22_X1 U16725 ( .A1(n20327), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13468) );
  NAND2_X1 U16726 ( .A1(n13718), .A2(DATAI_1_), .ZN(n13467) );
  NAND2_X1 U16727 ( .A1(n14848), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13466) );
  AND2_X1 U16728 ( .A1(n13467), .A2(n13466), .ZN(n13744) );
  INV_X1 U16729 ( .A(n13744), .ZN(n16116) );
  NAND2_X1 U16730 ( .A1(n20314), .A2(n16116), .ZN(n13478) );
  NAND2_X1 U16731 ( .A1(n13468), .A2(n13478), .ZN(P1_U2938) );
  AOI22_X1 U16732 ( .A1(n20327), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U16733 ( .A1(n13718), .A2(DATAI_2_), .ZN(n13470) );
  NAND2_X1 U16734 ( .A1(n14848), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13469) );
  AND2_X1 U16735 ( .A1(n13470), .A2(n13469), .ZN(n13757) );
  INV_X1 U16736 ( .A(n13757), .ZN(n14881) );
  NAND2_X1 U16737 ( .A1(n20314), .A2(n14881), .ZN(n13474) );
  NAND2_X1 U16738 ( .A1(n13471), .A2(n13474), .ZN(P1_U2939) );
  AOI22_X1 U16739 ( .A1(n20327), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U16740 ( .A1(n13473), .A2(n13472), .ZN(P1_U2942) );
  AOI22_X1 U16741 ( .A1(n20327), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13475) );
  NAND2_X1 U16742 ( .A1(n13475), .A2(n13474), .ZN(P1_U2954) );
  AOI22_X1 U16743 ( .A1(n20327), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U16744 ( .A1(n13477), .A2(n13476), .ZN(P1_U2943) );
  AOI22_X1 U16745 ( .A1(n20327), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13479) );
  NAND2_X1 U16746 ( .A1(n13479), .A2(n13478), .ZN(P1_U2953) );
  AOI22_X1 U16747 ( .A1(n20327), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U16748 ( .A1(n13481), .A2(n13480), .ZN(P1_U2948) );
  AOI22_X1 U16749 ( .A1(n20327), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U16750 ( .A1(n13483), .A2(n13482), .ZN(P1_U2944) );
  AOI22_X1 U16751 ( .A1(n20327), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13485) );
  NAND2_X1 U16752 ( .A1(n13485), .A2(n13484), .ZN(P1_U2952) );
  AOI22_X1 U16753 ( .A1(n20327), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13487) );
  INV_X1 U16754 ( .A(DATAI_9_), .ZN(n21117) );
  NAND2_X1 U16755 ( .A1(n14848), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13486) );
  OAI21_X1 U16756 ( .B1(n14848), .B2(n21117), .A(n13486), .ZN(n14856) );
  NAND2_X1 U16757 ( .A1(n20314), .A2(n14856), .ZN(n20318) );
  NAND2_X1 U16758 ( .A1(n13487), .A2(n20318), .ZN(P1_U2946) );
  INV_X1 U16759 ( .A(n20103), .ZN(n13499) );
  INV_X1 U16760 ( .A(n16544), .ZN(n15919) );
  OR3_X1 U16761 ( .A1(n13567), .A2(n13583), .A3(n10451), .ZN(n13492) );
  INV_X1 U16762 ( .A(n13489), .ZN(n13490) );
  NAND2_X1 U16763 ( .A1(n13490), .A2(n14333), .ZN(n13569) );
  AOI22_X1 U16764 ( .A1(n13492), .A2(n13569), .B1(n13491), .B2(n10927), .ZN(
        n13497) );
  INV_X1 U16765 ( .A(n13491), .ZN(n13493) );
  NAND2_X1 U16766 ( .A1(n10927), .A2(n13493), .ZN(n13572) );
  NAND2_X1 U16767 ( .A1(n10928), .A2(n13494), .ZN(n13495) );
  NAND2_X1 U16768 ( .A1(n13495), .A2(n13570), .ZN(n13571) );
  AND3_X1 U16769 ( .A1(n13572), .A2(n13569), .A3(n13571), .ZN(n13496) );
  MUX2_X1 U16770 ( .A(n13497), .B(n13496), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13498) );
  OAI21_X1 U16771 ( .B1(n16512), .B2(n13597), .A(n13498), .ZN(n13566) );
  AOI22_X1 U16772 ( .A1(n13499), .A2(n15919), .B1(n15911), .B2(n13566), .ZN(
        n13510) );
  NOR2_X1 U16773 ( .A1(n13587), .A2(n9834), .ZN(n13501) );
  NAND2_X1 U16774 ( .A1(n13502), .A2(n13501), .ZN(n13506) );
  NAND4_X1 U16775 ( .A1(n13506), .A2(n13505), .A3(n13504), .A4(n13503), .ZN(
        n13611) );
  INV_X1 U16776 ( .A(n13611), .ZN(n13602) );
  NAND2_X1 U16777 ( .A1(n19097), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13617) );
  NOR2_X1 U16778 ( .A1(n19097), .A2(n20127), .ZN(n16535) );
  NAND2_X1 U16779 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n16535), .ZN(n13507) );
  OAI211_X1 U16780 ( .C1(n13602), .C2(n13508), .A(n13617), .B(n13507), .ZN(
        n15956) );
  INV_X1 U16781 ( .A(n15956), .ZN(n15953) );
  NAND2_X1 U16782 ( .A1(n15953), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13509) );
  OAI21_X1 U16783 ( .B1(n13510), .B2(n15953), .A(n13509), .ZN(P2_U3596) );
  INV_X1 U16784 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20300) );
  OAI222_X1 U16785 ( .A1(n14904), .A2(n13952), .B1(n14903), .B2(n20300), .C1(
        n14902), .C2(n13744), .ZN(P1_U2903) );
  INV_X1 U16786 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20304) );
  OAI222_X1 U16787 ( .A1(n14902), .A2(n13739), .B1(n14904), .B2(n13914), .C1(
        n20304), .C2(n14903), .ZN(P1_U2904) );
  OAI21_X1 U16788 ( .B1(n13513), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13512), .ZN(n13514) );
  INV_X1 U16789 ( .A(n13514), .ZN(n15179) );
  INV_X1 U16790 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13515) );
  NOR2_X1 U16791 ( .A1(n20351), .A2(n13515), .ZN(n15180) );
  INV_X1 U16792 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13516) );
  AOI21_X1 U16793 ( .B1(n15039), .B2(n13517), .A(n13516), .ZN(n13518) );
  AOI211_X1 U16794 ( .C1(n15179), .C2(n20343), .A(n15180), .B(n13518), .ZN(
        n13519) );
  OAI21_X1 U16795 ( .B1(n13914), .B2(n15054), .A(n13519), .ZN(P1_U2999) );
  INV_X1 U16796 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U16797 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20301), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16031), .ZN(n13520) );
  OAI21_X1 U16798 ( .B1(n13521), .B2(n13529), .A(n13520), .ZN(P1_U2906) );
  INV_X1 U16799 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U16800 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13522) );
  OAI21_X1 U16801 ( .B1(n13523), .B2(n13529), .A(n13522), .ZN(P1_U2919) );
  INV_X1 U16802 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U16803 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13524) );
  OAI21_X1 U16804 ( .B1(n13525), .B2(n13529), .A(n13524), .ZN(P1_U2917) );
  INV_X1 U16805 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U16806 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13526) );
  OAI21_X1 U16807 ( .B1(n13527), .B2(n13529), .A(n13526), .ZN(P1_U2918) );
  INV_X1 U16808 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U16809 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13528) );
  OAI21_X1 U16810 ( .B1(n13530), .B2(n13529), .A(n13528), .ZN(P1_U2910) );
  NOR2_X1 U16811 ( .A1(n9770), .A2(n13531), .ZN(n13532) );
  OR2_X1 U16812 ( .A1(n13561), .A2(n13532), .ZN(n19276) );
  INV_X1 U16813 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13533) );
  NOR2_X1 U16814 ( .A1(n13534), .A2(n13533), .ZN(n13536) );
  NAND3_X1 U16815 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13622) );
  OAI211_X1 U16816 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13536), .A(
        n13622), .B(n15434), .ZN(n13538) );
  NAND2_X1 U16817 ( .A1(n13273), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13537) );
  OAI211_X1 U16818 ( .C1(n19276), .C2(n13273), .A(n13538), .B(n13537), .ZN(
        P2_U2881) );
  AND4_X1 U16819 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__4__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U16820 ( .A1(n13623), .A2(n13539), .ZN(n13540) );
  NOR2_X1 U16821 ( .A1(n14429), .A2(n13540), .ZN(n13541) );
  XNOR2_X1 U16822 ( .A(n13550), .B(n13549), .ZN(n13548) );
  OR2_X1 U16823 ( .A1(n13545), .A2(n13544), .ZN(n13546) );
  AND2_X1 U16824 ( .A1(n13554), .A2(n13546), .ZN(n16425) );
  INV_X1 U16825 ( .A(n16425), .ZN(n15890) );
  MUX2_X1 U16826 ( .A(n15890), .B(n10108), .S(n13322), .Z(n13547) );
  OAI21_X1 U16827 ( .B1(n13548), .B2(n15450), .A(n13547), .ZN(P2_U2878) );
  OAI211_X1 U16828 ( .C1(n13552), .C2(n13551), .A(n13640), .B(n15434), .ZN(
        n13558) );
  AND2_X1 U16829 ( .A1(n13554), .A2(n13553), .ZN(n13555) );
  NAND2_X1 U16830 ( .A1(n9761), .A2(n15440), .ZN(n13557) );
  OAI211_X1 U16831 ( .C1(n15440), .C2(n13559), .A(n13558), .B(n13557), .ZN(
        P2_U2877) );
  XOR2_X1 U16832 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13622), .Z(n13565)
         );
  OR2_X1 U16833 ( .A1(n13561), .A2(n13560), .ZN(n13562) );
  AND2_X1 U16834 ( .A1(n13562), .A2(n13619), .ZN(n19263) );
  NOR2_X1 U16835 ( .A1(n15442), .A2(n10698), .ZN(n13563) );
  AOI21_X1 U16836 ( .B1(n19263), .B2(n15442), .A(n13563), .ZN(n13564) );
  OAI21_X1 U16837 ( .B1(n13565), .B2(n15450), .A(n13564), .ZN(P2_U2880) );
  MUX2_X1 U16838 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13566), .S(
        n13611), .Z(n13605) );
  INV_X1 U16839 ( .A(n13597), .ZN(n13577) );
  INV_X1 U16840 ( .A(n13571), .ZN(n13568) );
  AOI211_X1 U16841 ( .C1(n13568), .C2(n13569), .A(n13567), .B(n13583), .ZN(
        n13575) );
  AND3_X1 U16842 ( .A1(n13571), .A2(n13570), .A3(n13569), .ZN(n13574) );
  NOR2_X1 U16843 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13573) );
  OAI22_X1 U16844 ( .A1(n13575), .A2(n13574), .B1(n13573), .B2(n13572), .ZN(
        n13576) );
  AOI21_X1 U16845 ( .B1(n9639), .B2(n13577), .A(n13576), .ZN(n15917) );
  NOR2_X1 U16846 ( .A1(n13611), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13578) );
  AOI21_X1 U16847 ( .B1(n15917), .B2(n13611), .A(n13578), .ZN(n13604) );
  OAI22_X1 U16848 ( .A1(n13584), .A2(n13581), .B1(n13580), .B2(n13579), .ZN(
        n13582) );
  AOI21_X1 U16849 ( .B1(n13584), .B2(n13583), .A(n13582), .ZN(n20142) );
  INV_X1 U16850 ( .A(n20142), .ZN(n13590) );
  OAI21_X1 U16851 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n13585), .ZN(n13588) );
  OR3_X1 U16852 ( .A1(n13587), .A2(n13586), .A3(n14487), .ZN(n15952) );
  OAI211_X1 U16853 ( .C1(n20152), .C2(n10809), .A(n13588), .B(n15952), .ZN(
        n13589) );
  AOI211_X1 U16854 ( .C1(n13605), .C2(n13604), .A(n13590), .B(n13589), .ZN(
        n13610) );
  AOI22_X1 U16855 ( .A1(n13605), .A2(n20116), .B1(n20109), .B2(n13604), .ZN(
        n13603) );
  NOR2_X1 U16856 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19558) );
  INV_X1 U16857 ( .A(n19558), .ZN(n19535) );
  AND2_X1 U16858 ( .A1(n13592), .A2(n13591), .ZN(n13596) );
  NOR3_X1 U16859 ( .A1(n13596), .A2(n10220), .A3(n13489), .ZN(n13593) );
  AOI21_X1 U16860 ( .B1(n13594), .B2(n10927), .A(n13593), .ZN(n13595) );
  OAI21_X1 U16861 ( .B1(n13277), .B2(n13597), .A(n13595), .ZN(n15912) );
  INV_X1 U16862 ( .A(n15912), .ZN(n13599) );
  OAI22_X1 U16863 ( .A1(n19321), .A2(n13597), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13596), .ZN(n15903) );
  AOI211_X1 U16864 ( .C1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n10927), .A(
        n20135), .B(n15903), .ZN(n13598) );
  OAI21_X1 U16865 ( .B1(n13599), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13598), .ZN(n13600) );
  OAI21_X1 U16866 ( .B1(n20125), .B2(n15912), .A(n13600), .ZN(n13601) );
  AOI211_X1 U16867 ( .C1(n13603), .C2(n19535), .A(n13602), .B(n13601), .ZN(
        n13608) );
  AOI22_X1 U16868 ( .A1(n13605), .A2(n20109), .B1(n13604), .B2(n19558), .ZN(
        n13606) );
  INV_X1 U16869 ( .A(n13606), .ZN(n13607) );
  OAI21_X1 U16870 ( .B1(n13608), .B2(n13607), .A(n16037), .ZN(n13609) );
  OAI211_X1 U16871 ( .C1(n13611), .C2(n15955), .A(n13610), .B(n13609), .ZN(
        n16537) );
  OAI21_X1 U16872 ( .B1(n16537), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13615) );
  OR2_X1 U16873 ( .A1(n16539), .A2(n19884), .ZN(n20145) );
  AOI21_X1 U16874 ( .B1(n13613), .B2(n13612), .A(n20145), .ZN(n13614) );
  INV_X1 U16875 ( .A(n16540), .ZN(n13618) );
  INV_X1 U16876 ( .A(n16535), .ZN(n13616) );
  OAI211_X1 U16877 ( .C1(n13618), .C2(n19854), .A(n13617), .B(n13616), .ZN(
        P2_U3593) );
  AOI21_X1 U16878 ( .B1(n13620), .B2(n13619), .A(n13544), .ZN(n19251) );
  INV_X1 U16879 ( .A(n19251), .ZN(n15687) );
  INV_X1 U16880 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13621) );
  NOR2_X1 U16881 ( .A1(n13622), .A2(n13621), .ZN(n13624) );
  OAI211_X1 U16882 ( .C1(n13624), .C2(n13623), .A(n15434), .B(n13550), .ZN(
        n13626) );
  NAND2_X1 U16883 ( .A1(n13273), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13625) );
  OAI211_X1 U16884 ( .C1(n15687), .C2(n13273), .A(n13626), .B(n13625), .ZN(
        P2_U2879) );
  OR2_X1 U16885 ( .A1(n13627), .A2(n13084), .ZN(n13629) );
  NAND2_X1 U16886 ( .A1(n13629), .A2(n13628), .ZN(n19234) );
  INV_X1 U16887 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19395) );
  OAI222_X1 U16888 ( .A1(n19234), .A2(n19351), .B1(n15460), .B2(n19386), .C1(
        n19395), .C2(n19349), .ZN(P2_U2907) );
  INV_X1 U16889 ( .A(n13641), .ZN(n13639) );
  XNOR2_X1 U16890 ( .A(n13640), .B(n13639), .ZN(n13632) );
  MUX2_X1 U16891 ( .A(n13630), .B(n16411), .S(n15442), .Z(n13631) );
  OAI21_X1 U16892 ( .B1(n13632), .B2(n15450), .A(n13631), .ZN(P2_U2876) );
  NOR2_X1 U16893 ( .A1(n20029), .A2(n19097), .ZN(n16032) );
  AOI21_X1 U16894 ( .B1(n16032), .B2(n15911), .A(n16538), .ZN(n13634) );
  NOR2_X1 U16895 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19097), .ZN(n16534) );
  OAI211_X1 U16896 ( .C1(n16540), .C2(n16534), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20029), .ZN(n13633) );
  OAI211_X1 U16897 ( .C1(n16540), .C2(n13634), .A(n13633), .B(n19289), .ZN(
        P2_U3177) );
  NAND2_X1 U16898 ( .A1(n13637), .A2(n13636), .ZN(n13638) );
  AND2_X1 U16899 ( .A1(n13821), .A2(n13638), .ZN(n19230) );
  INV_X1 U16900 ( .A(n19230), .ZN(n13648) );
  NOR2_X1 U16901 ( .A1(n13640), .A2(n13639), .ZN(n13645) );
  NAND2_X1 U16902 ( .A1(n13642), .A2(n10210), .ZN(n13972) );
  OAI211_X1 U16903 ( .C1(n13645), .C2(n13644), .A(n15434), .B(n13643), .ZN(
        n13647) );
  NAND2_X1 U16904 ( .A1(n13273), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13646) );
  OAI211_X1 U16905 ( .C1(n13648), .C2(n13273), .A(n13647), .B(n13646), .ZN(
        P2_U2875) );
  INV_X1 U16906 ( .A(n20506), .ZN(n13711) );
  NOR2_X1 U16907 ( .A1(n11786), .A2(n13711), .ZN(n13649) );
  XOR2_X1 U16908 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n13649), .Z(
        n20228) );
  INV_X1 U16909 ( .A(n20228), .ZN(n13650) );
  NOR2_X1 U16910 ( .A1(n13650), .A2(n12449), .ZN(n16315) );
  NAND2_X1 U16911 ( .A1(n15993), .A2(n13651), .ZN(n13655) );
  NAND2_X1 U16912 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), 
        .ZN(n13654) );
  NAND2_X1 U16913 ( .A1(n13655), .A2(n13652), .ZN(n13653) );
  OAI211_X1 U16914 ( .C1(n16315), .C2(n13655), .A(n13654), .B(n13653), .ZN(
        n13681) );
  INV_X1 U16915 ( .A(n13681), .ZN(n13685) );
  INV_X1 U16916 ( .A(n13656), .ZN(n13684) );
  NOR2_X1 U16917 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13651), .ZN(n13680) );
  INV_X1 U16918 ( .A(n9689), .ZN(n13918) );
  NAND2_X1 U16919 ( .A1(n14594), .A2(n13658), .ZN(n13673) );
  INV_X1 U16920 ( .A(n13673), .ZN(n13666) );
  NOR2_X1 U16921 ( .A1(n13659), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13670) );
  NOR2_X1 U16922 ( .A1(n13670), .A2(n13660), .ZN(n15207) );
  NOR2_X1 U16923 ( .A1(n13676), .A2(n11347), .ZN(n13661) );
  NOR2_X1 U16924 ( .A1(n13676), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15196) );
  MUX2_X1 U16925 ( .A(n13661), .B(n15196), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13662) );
  INV_X1 U16926 ( .A(n13662), .ZN(n13665) );
  AND2_X1 U16927 ( .A1(n12462), .A2(n13663), .ZN(n13671) );
  NAND2_X1 U16928 ( .A1(n13671), .A2(n15207), .ZN(n13664) );
  OAI211_X1 U16929 ( .C1(n13666), .C2(n15207), .A(n13665), .B(n13664), .ZN(
        n13667) );
  AOI21_X1 U16930 ( .B1(n13918), .B2(n15197), .A(n13667), .ZN(n15210) );
  NOR2_X1 U16931 ( .A1(n15993), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13668) );
  AOI21_X1 U16932 ( .B1(n15210), .B2(n15993), .A(n13668), .ZN(n15989) );
  AOI22_X1 U16933 ( .A1(n13680), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n13651), .B2(n15989), .ZN(n13683) );
  INV_X1 U16934 ( .A(n20618), .ZN(n20254) );
  AOI21_X1 U16935 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13669), .A(
        n11358), .ZN(n13675) );
  XNOR2_X1 U16936 ( .A(n13670), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13672) );
  OAI21_X1 U16937 ( .B1(n13660), .B2(n11350), .A(n11690), .ZN(n20935) );
  AOI22_X1 U16938 ( .A1(n13673), .A2(n13672), .B1(n13671), .B2(n20935), .ZN(
        n13674) );
  OAI21_X1 U16939 ( .B1(n13676), .B2(n13675), .A(n13674), .ZN(n13677) );
  AOI21_X1 U16940 ( .B1(n15196), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13677), .ZN(n13678) );
  OAI21_X1 U16941 ( .B1(n20254), .B2(n13679), .A(n13678), .ZN(n20938) );
  MUX2_X1 U16942 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20938), .S(
        n15993), .Z(n16001) );
  AOI22_X1 U16943 ( .A1(n13680), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13651), .B2(n16001), .ZN(n13682) );
  OAI21_X1 U16944 ( .B1(n13683), .B2(n13682), .A(n13681), .ZN(n16005) );
  OAI21_X1 U16945 ( .B1(n13685), .B2(n13684), .A(n16005), .ZN(n15189) );
  INV_X1 U16946 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20168) );
  AOI21_X1 U16947 ( .B1(n15189), .B2(n20168), .A(n16322), .ZN(n13687) );
  NOR2_X1 U16948 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20958) );
  INV_X1 U16949 ( .A(n15217), .ZN(n13686) );
  INV_X1 U16950 ( .A(n20385), .ZN(n13704) );
  NOR2_X1 U16951 ( .A1(n13704), .A2(n20802), .ZN(n13703) );
  INV_X1 U16952 ( .A(n13703), .ZN(n13695) );
  NAND2_X1 U16953 ( .A1(n13688), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20806) );
  XNOR2_X1 U16954 ( .A(n13915), .B(n20806), .ZN(n13689) );
  NAND2_X1 U16955 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20689), .ZN(n15190) );
  NAND2_X1 U16956 ( .A1(n20385), .A2(n15190), .ZN(n13707) );
  OAI222_X1 U16957 ( .A1(n13695), .A2(n13689), .B1(n20385), .B2(n12290), .C1(
        n9689), .C2(n13707), .ZN(P1_U3476) );
  NAND2_X1 U16958 ( .A1(n13690), .A2(n13691), .ZN(n20807) );
  OAI22_X1 U16959 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n13916), .B1(n20807), 
        .B2(n13688), .ZN(n13693) );
  NOR2_X1 U16960 ( .A1(n20587), .A2(n20806), .ZN(n20591) );
  NOR3_X1 U16961 ( .A1(n13693), .A2(n20680), .A3(n20591), .ZN(n13694) );
  OAI222_X1 U16962 ( .A1(n20385), .A2(n20727), .B1(n13707), .B2(n20254), .C1(
        n13695), .C2(n13694), .ZN(P1_U3475) );
  AOI21_X1 U16963 ( .B1(n13697), .B2(n13773), .A(n13698), .ZN(n13699) );
  NOR2_X1 U16964 ( .A1(n9672), .A2(n13699), .ZN(n13956) );
  INV_X1 U16965 ( .A(n13956), .ZN(n20238) );
  INV_X1 U16966 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13701) );
  OR2_X1 U16967 ( .A1(n13700), .A2(n16303), .ZN(n20353) );
  OAI222_X1 U16968 ( .A1(n20238), .A2(n14842), .B1(n20270), .B2(n13701), .C1(
        n20353), .C2(n20265), .ZN(P1_U2868) );
  OAI211_X1 U16969 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n13688), .A(n13703), 
        .B(n20806), .ZN(n13706) );
  NAND2_X1 U16970 ( .A1(n13704), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13705) );
  OAI211_X1 U16971 ( .C1(n13707), .C2(n20619), .A(n13706), .B(n13705), .ZN(
        P1_U3477) );
  INV_X1 U16972 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20294) );
  INV_X1 U16973 ( .A(n14874), .ZN(n13734) );
  OAI222_X1 U16974 ( .A1(n14904), .A2(n20238), .B1(n14903), .B2(n20294), .C1(
        n14902), .C2(n13734), .ZN(P1_U2900) );
  AOI21_X1 U16975 ( .B1(n13708), .B2(n13628), .A(n9705), .ZN(n19219) );
  INV_X1 U16976 ( .A(n19219), .ZN(n13710) );
  INV_X1 U16977 ( .A(n15452), .ZN(n13709) );
  OAI222_X1 U16978 ( .A1(n13710), .A2(n19351), .B1(n13709), .B2(n19386), .C1(
        n19393), .C2(n19349), .ZN(P2_U2906) );
  NOR3_X1 U16979 ( .A1(n12290), .A2(n20727), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13722) );
  INV_X1 U16980 ( .A(n13712), .ZN(n20648) );
  NAND2_X1 U16981 ( .A1(n20800), .A2(n20648), .ZN(n13714) );
  INV_X1 U16982 ( .A(n13722), .ZN(n15216) );
  NOR2_X1 U16983 ( .A1(n20647), .A2(n15216), .ZN(n13766) );
  INV_X1 U16984 ( .A(n13766), .ZN(n13713) );
  NAND2_X1 U16985 ( .A1(n13714), .A2(n13713), .ZN(n13721) );
  INV_X1 U16986 ( .A(n13721), .ZN(n13715) );
  OAI211_X1 U16987 ( .C1(n20807), .C2(n21022), .A(n20677), .B(n13715), .ZN(
        n13716) );
  OAI211_X1 U16988 ( .C1(n20810), .C2(n13722), .A(n13716), .B(n20809), .ZN(
        n13717) );
  INV_X1 U16989 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13728) );
  INV_X1 U16990 ( .A(DATAI_23_), .ZN(n13719) );
  INV_X1 U16991 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16620) );
  OAI22_X1 U16992 ( .A1(n13719), .A2(n13763), .B1(n16620), .B2(n13764), .ZN(
        n20721) );
  NOR2_X2 U16993 ( .A1(n20807), .A2(n20653), .ZN(n20794) );
  INV_X1 U16994 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19497) );
  INV_X1 U16995 ( .A(DATAI_31_), .ZN(n21079) );
  INV_X1 U16996 ( .A(n20858), .ZN(n20676) );
  NAND2_X1 U16997 ( .A1(n13750), .A2(n11567), .ZN(n20468) );
  INV_X1 U16998 ( .A(n14863), .ZN(n13887) );
  NAND2_X1 U16999 ( .A1(n13721), .A2(n20677), .ZN(n13724) );
  NAND2_X1 U17000 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13722), .ZN(n13723) );
  NAND2_X1 U17001 ( .A1(n13724), .A2(n13723), .ZN(n13767) );
  AOI22_X1 U17002 ( .A1(n20857), .A2(n13766), .B1(n20855), .B2(n13767), .ZN(
        n13725) );
  OAI21_X1 U17003 ( .B1(n15238), .B2(n20676), .A(n13725), .ZN(n13726) );
  AOI21_X1 U17004 ( .B1(n20721), .B2(n20794), .A(n13726), .ZN(n13727) );
  OAI21_X1 U17005 ( .B1(n13772), .B2(n13728), .A(n13727), .ZN(P1_U3144) );
  INV_X1 U17006 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13733) );
  INV_X1 U17007 ( .A(DATAI_19_), .ZN(n13729) );
  INV_X1 U17008 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16627) );
  OAI22_X1 U17009 ( .A1(n13729), .A2(n13763), .B1(n16627), .B2(n13764), .ZN(
        n20704) );
  INV_X1 U17010 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16612) );
  INV_X1 U17011 ( .A(DATAI_27_), .ZN(n21085) );
  OAI22_X1 U17012 ( .A1(n16612), .A2(n13764), .B1(n21085), .B2(n13763), .ZN(
        n20830) );
  NAND2_X1 U17013 ( .A1(n13750), .A2(n11630), .ZN(n20451) );
  INV_X1 U17014 ( .A(n14877), .ZN(n13811) );
  AOI22_X1 U17015 ( .A1(n20829), .A2(n13766), .B1(n20828), .B2(n13767), .ZN(
        n13730) );
  OAI21_X1 U17016 ( .B1(n15238), .B2(n9791), .A(n13730), .ZN(n13731) );
  AOI21_X1 U17017 ( .B1(n20704), .B2(n20794), .A(n13731), .ZN(n13732) );
  OAI21_X1 U17018 ( .B1(n13772), .B2(n13733), .A(n13732), .ZN(P1_U3140) );
  INV_X1 U17019 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13738) );
  INV_X1 U17020 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16625) );
  INV_X1 U17021 ( .A(DATAI_20_), .ZN(n20972) );
  OAI22_X1 U17022 ( .A1(n16625), .A2(n13764), .B1(n20972), .B2(n13763), .ZN(
        n20708) );
  INV_X1 U17023 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19479) );
  INV_X1 U17024 ( .A(DATAI_28_), .ZN(n21090) );
  OAI22_X1 U17025 ( .A1(n19479), .A2(n13764), .B1(n21090), .B2(n13763), .ZN(
        n20836) );
  NAND2_X1 U17026 ( .A1(n13750), .A2(n11682), .ZN(n20455) );
  AOI22_X1 U17027 ( .A1(n20835), .A2(n13766), .B1(n20834), .B2(n13767), .ZN(
        n13735) );
  OAI21_X1 U17028 ( .B1(n15238), .B2(n9793), .A(n13735), .ZN(n13736) );
  AOI21_X1 U17029 ( .B1(n20708), .B2(n20794), .A(n13736), .ZN(n13737) );
  OAI21_X1 U17030 ( .B1(n13772), .B2(n13738), .A(n13737), .ZN(P1_U3141) );
  INV_X1 U17031 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13743) );
  INV_X1 U17032 ( .A(DATAI_16_), .ZN(n21088) );
  INV_X1 U17033 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16633) );
  OAI22_X1 U17034 ( .A1(n21088), .A2(n13763), .B1(n16633), .B2(n13764), .ZN(
        n20694) );
  INV_X1 U17035 ( .A(DATAI_24_), .ZN(n20965) );
  INV_X1 U17036 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16618) );
  OAI22_X2 U17037 ( .A1(n20965), .A2(n13763), .B1(n16618), .B2(n13764), .ZN(
        n20812) );
  INV_X1 U17038 ( .A(n20812), .ZN(n20657) );
  NOR2_X2 U17039 ( .A1(n13765), .A2(n11635), .ZN(n20804) );
  AOI22_X1 U17040 ( .A1(n20804), .A2(n13766), .B1(n20803), .B2(n13767), .ZN(
        n13740) );
  OAI21_X1 U17041 ( .B1(n15238), .B2(n20657), .A(n13740), .ZN(n13741) );
  AOI21_X1 U17042 ( .B1(n20694), .B2(n20794), .A(n13741), .ZN(n13742) );
  OAI21_X1 U17043 ( .B1(n13772), .B2(n13743), .A(n13742), .ZN(P1_U3137) );
  INV_X1 U17044 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13748) );
  INV_X1 U17045 ( .A(DATAI_17_), .ZN(n21073) );
  INV_X1 U17046 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16631) );
  OAI22_X1 U17047 ( .A1(n21073), .A2(n13763), .B1(n16631), .B2(n13764), .ZN(
        n20818) );
  INV_X1 U17048 ( .A(DATAI_25_), .ZN(n20998) );
  INV_X1 U17049 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16616) );
  OAI22_X1 U17050 ( .A1(n20998), .A2(n13763), .B1(n16616), .B2(n13764), .ZN(
        n20774) );
  INV_X1 U17051 ( .A(n20774), .ZN(n20821) );
  NOR2_X2 U17052 ( .A1(n13765), .A2(n9654), .ZN(n20817) );
  AOI22_X1 U17053 ( .A1(n20817), .A2(n13766), .B1(n20816), .B2(n13767), .ZN(
        n13745) );
  OAI21_X1 U17054 ( .B1(n15238), .B2(n20821), .A(n13745), .ZN(n13746) );
  AOI21_X1 U17055 ( .B1(n20818), .B2(n20794), .A(n13746), .ZN(n13747) );
  OAI21_X1 U17056 ( .B1(n13772), .B2(n13748), .A(n13747), .ZN(P1_U3138) );
  INV_X1 U17057 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13754) );
  INV_X1 U17058 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16629) );
  INV_X1 U17059 ( .A(DATAI_18_), .ZN(n21140) );
  INV_X1 U17060 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16614) );
  INV_X1 U17061 ( .A(DATAI_26_), .ZN(n21024) );
  OAI22_X1 U17062 ( .A1(n16614), .A2(n13764), .B1(n21024), .B2(n13763), .ZN(
        n20778) );
  INV_X1 U17063 ( .A(n20778), .ZN(n20827) );
  NAND2_X1 U17064 ( .A1(n13750), .A2(n13749), .ZN(n20447) );
  NOR2_X2 U17065 ( .A1(n15217), .A2(n13757), .ZN(n20822) );
  AOI22_X1 U17066 ( .A1(n20823), .A2(n13766), .B1(n20822), .B2(n13767), .ZN(
        n13751) );
  OAI21_X1 U17067 ( .B1(n15238), .B2(n20827), .A(n13751), .ZN(n13752) );
  AOI21_X1 U17068 ( .B1(n20824), .B2(n20794), .A(n13752), .ZN(n13753) );
  OAI21_X1 U17069 ( .B1(n13772), .B2(n13754), .A(n13753), .ZN(P1_U3139) );
  XOR2_X1 U17070 ( .A(n13453), .B(n13756), .Z(n20345) );
  INV_X1 U17071 ( .A(n20345), .ZN(n13796) );
  INV_X1 U17072 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20298) );
  OAI222_X1 U17073 ( .A1(n14904), .A2(n13796), .B1(n14903), .B2(n20298), .C1(
        n14902), .C2(n13757), .ZN(P1_U2902) );
  INV_X1 U17074 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13762) );
  INV_X1 U17075 ( .A(DATAI_22_), .ZN(n13758) );
  INV_X1 U17076 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16622) );
  OAI22_X1 U17077 ( .A1(n13758), .A2(n13763), .B1(n16622), .B2(n13764), .ZN(
        n20715) );
  INV_X1 U17078 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16607) );
  INV_X1 U17079 ( .A(DATAI_30_), .ZN(n21084) );
  OAI22_X1 U17080 ( .A1(n16607), .A2(n13764), .B1(n21084), .B2(n13763), .ZN(
        n20850) );
  INV_X1 U17081 ( .A(n14867), .ZN(n13831) );
  NOR2_X2 U17082 ( .A1(n13765), .A2(n9669), .ZN(n20848) );
  AOI22_X1 U17083 ( .A1(n20849), .A2(n13767), .B1(n20848), .B2(n13766), .ZN(
        n13759) );
  OAI21_X1 U17084 ( .B1(n15238), .B2(n9789), .A(n13759), .ZN(n13760) );
  AOI21_X1 U17085 ( .B1(n20715), .B2(n20794), .A(n13760), .ZN(n13761) );
  OAI21_X1 U17086 ( .B1(n13772), .B2(n13762), .A(n13761), .ZN(P1_U3143) );
  INV_X1 U17087 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13771) );
  INV_X1 U17088 ( .A(DATAI_21_), .ZN(n21120) );
  INV_X1 U17089 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19484) );
  INV_X1 U17090 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16609) );
  INV_X1 U17091 ( .A(DATAI_29_), .ZN(n21082) );
  OAI22_X1 U17092 ( .A1(n16609), .A2(n13764), .B1(n21082), .B2(n13763), .ZN(
        n20786) );
  INV_X1 U17093 ( .A(n20786), .ZN(n20847) );
  INV_X1 U17094 ( .A(n14871), .ZN(n13816) );
  NOR2_X2 U17095 ( .A1(n15217), .A2(n13816), .ZN(n20841) );
  NOR2_X2 U17096 ( .A1(n13765), .A2(n12278), .ZN(n20840) );
  AOI22_X1 U17097 ( .A1(n20841), .A2(n13767), .B1(n20840), .B2(n13766), .ZN(
        n13768) );
  OAI21_X1 U17098 ( .B1(n15238), .B2(n20847), .A(n13768), .ZN(n13769) );
  AOI21_X1 U17099 ( .B1(n20794), .B2(n20842), .A(n13769), .ZN(n13770) );
  OAI21_X1 U17100 ( .B1(n13772), .B2(n13771), .A(n13770), .ZN(P1_U3142) );
  XOR2_X1 U17101 ( .A(n13773), .B(n13697), .Z(n20334) );
  INV_X1 U17102 ( .A(n20334), .ZN(n13812) );
  AOI21_X1 U17103 ( .B1(n13795), .B2(n13775), .A(n13774), .ZN(n20361) );
  INV_X1 U17104 ( .A(n20270), .ZN(n14840) );
  AOI22_X1 U17105 ( .A1(n20361), .A2(n12975), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14840), .ZN(n13776) );
  OAI21_X1 U17106 ( .B1(n13812), .B2(n14842), .A(n13776), .ZN(P1_U2869) );
  XOR2_X1 U17107 ( .A(n20110), .B(n20111), .Z(n19370) );
  OAI21_X1 U17108 ( .B1(n13779), .B2(n13778), .A(n13777), .ZN(n20123) );
  XOR2_X1 U17109 ( .A(n20123), .B(n20121), .Z(n19375) );
  OAI21_X1 U17110 ( .B1(n13782), .B2(n13781), .A(n13780), .ZN(n19314) );
  INV_X1 U17111 ( .A(n19314), .ZN(n19383) );
  NAND2_X1 U17112 ( .A1(n19713), .A2(n19383), .ZN(n19382) );
  NAND2_X1 U17113 ( .A1(n19375), .A2(n19382), .ZN(n19374) );
  OAI21_X1 U17114 ( .B1(n20123), .B2(n20121), .A(n19374), .ZN(n19369) );
  NAND2_X1 U17115 ( .A1(n19370), .A2(n19369), .ZN(n19368) );
  OAI21_X1 U17116 ( .B1(n20111), .B2(n20110), .A(n19368), .ZN(n19363) );
  XNOR2_X1 U17117 ( .A(n13783), .B(n9765), .ZN(n19361) );
  XNOR2_X1 U17118 ( .A(n20103), .B(n19361), .ZN(n19364) );
  NAND2_X1 U17119 ( .A1(n19363), .A2(n19364), .ZN(n19362) );
  INV_X1 U17120 ( .A(n19361), .ZN(n20102) );
  NAND2_X1 U17121 ( .A1(n20103), .A2(n20102), .ZN(n13787) );
  OR2_X1 U17122 ( .A1(n13785), .A2(n13784), .ZN(n13786) );
  AND2_X1 U17123 ( .A1(n13786), .A2(n13848), .ZN(n19281) );
  AOI21_X1 U17124 ( .B1(n19362), .B2(n13787), .A(n19281), .ZN(n19358) );
  XNOR2_X1 U17125 ( .A(n19358), .B(n19357), .ZN(n13791) );
  AOI22_X1 U17126 ( .A1(n19380), .A2(n19281), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19379), .ZN(n13790) );
  INV_X1 U17127 ( .A(n19386), .ZN(n19342) );
  NAND2_X1 U17128 ( .A1(n19342), .A2(n13788), .ZN(n13789) );
  OAI211_X1 U17129 ( .C1(n13791), .C2(n19356), .A(n13790), .B(n13789), .ZN(
        P2_U2915) );
  OR2_X1 U17130 ( .A1(n13793), .A2(n13792), .ZN(n13794) );
  NAND2_X1 U17131 ( .A1(n13795), .A2(n13794), .ZN(n20366) );
  INV_X1 U17132 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13797) );
  OAI222_X1 U17133 ( .A1(n20366), .A2(n20265), .B1(n13797), .B2(n20270), .C1(
        n13796), .C2(n14842), .ZN(P1_U2870) );
  XNOR2_X1 U17134 ( .A(n13798), .B(n13799), .ZN(n16516) );
  XNOR2_X1 U17135 ( .A(n13800), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13801) );
  XNOR2_X1 U17136 ( .A(n13802), .B(n13801), .ZN(n16518) );
  NAND2_X1 U17137 ( .A1(n16518), .A2(n16450), .ZN(n13810) );
  NAND2_X1 U17138 ( .A1(n16440), .A2(n13860), .ZN(n13806) );
  NOR2_X1 U17139 ( .A1(n16466), .A2(n13804), .ZN(n16514) );
  INV_X1 U17140 ( .A(n16514), .ZN(n13805) );
  OAI211_X1 U17141 ( .C1(n13807), .C2(n16453), .A(n13806), .B(n13805), .ZN(
        n13808) );
  AOI21_X1 U17142 ( .B1(n13803), .B2(n19428), .A(n13808), .ZN(n13809) );
  OAI211_X1 U17143 ( .C1(n16516), .C2(n19423), .A(n13810), .B(n13809), .ZN(
        P2_U3011) );
  INV_X1 U17144 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20296) );
  OAI222_X1 U17145 ( .A1(n14904), .A2(n13812), .B1(n14903), .B2(n20296), .C1(
        n14902), .C2(n13811), .ZN(P1_U2901) );
  AND2_X1 U17146 ( .A1(n13696), .A2(n13814), .ZN(n13815) );
  OR2_X1 U17147 ( .A1(n13813), .A2(n13815), .ZN(n20266) );
  OAI222_X1 U17148 ( .A1(n14904), .A2(n20266), .B1(n14903), .B2(n11863), .C1(
        n14902), .C2(n13816), .ZN(P1_U2899) );
  OAI21_X1 U17149 ( .B1(n13813), .B2(n13818), .A(n13817), .ZN(n16168) );
  XOR2_X1 U17150 ( .A(n16286), .B(n16305), .Z(n20205) );
  AOI22_X1 U17151 ( .A1(n20205), .A2(n12975), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14840), .ZN(n13819) );
  OAI21_X1 U17152 ( .B1(n16168), .B2(n14842), .A(n13819), .ZN(P1_U2866) );
  INV_X1 U17153 ( .A(n13833), .ZN(n13832) );
  XNOR2_X1 U17154 ( .A(n13643), .B(n13832), .ZN(n13824) );
  NAND2_X1 U17155 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  AND2_X1 U17156 ( .A1(n13837), .A2(n13822), .ZN(n19220) );
  INV_X1 U17157 ( .A(n19220), .ZN(n16472) );
  MUX2_X1 U17158 ( .A(n10729), .B(n16472), .S(n15442), .Z(n13823) );
  OAI21_X1 U17159 ( .B1(n13824), .B2(n15450), .A(n13823), .ZN(P2_U2874) );
  INV_X1 U17160 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13825) );
  NOR2_X1 U17161 ( .A1(n20351), .A2(n13825), .ZN(n15173) );
  AOI21_X1 U17162 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15173), .ZN(n13826) );
  OAI21_X1 U17163 ( .B1(n20349), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13826), .ZN(n13827) );
  INV_X1 U17164 ( .A(n13827), .ZN(n13830) );
  OR2_X1 U17165 ( .A1(n13828), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15167) );
  NAND3_X1 U17166 ( .A1(n15167), .A2(n15166), .A3(n20343), .ZN(n13829) );
  OAI211_X1 U17167 ( .C1(n13952), .C2(n15054), .A(n13830), .B(n13829), .ZN(
        P1_U2998) );
  INV_X1 U17168 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20291) );
  OAI222_X1 U17169 ( .A1(n14904), .A2(n16168), .B1(n14903), .B2(n20291), .C1(
        n14902), .C2(n13831), .ZN(P1_U2898) );
  NOR2_X1 U17170 ( .A1(n13643), .A2(n13832), .ZN(n13835) );
  NAND2_X1 U17171 ( .A1(n13833), .A2(n13834), .ZN(n13969) );
  OR2_X1 U17172 ( .A1(n13643), .A2(n13969), .ZN(n13962) );
  OAI211_X1 U17173 ( .C1(n13835), .C2(n13834), .A(n15434), .B(n13962), .ZN(
        n13840) );
  INV_X1 U17174 ( .A(n13836), .ZN(n13964) );
  AOI21_X1 U17175 ( .B1(n13838), .B2(n13837), .A(n13836), .ZN(n19209) );
  NAND2_X1 U17176 ( .A1(n19209), .A2(n15440), .ZN(n13839) );
  OAI211_X1 U17177 ( .C1(n15442), .C2(n13841), .A(n13840), .B(n13839), .ZN(
        P2_U2873) );
  NAND2_X1 U17178 ( .A1(n19257), .A2(n13842), .ZN(n13843) );
  XNOR2_X1 U17179 ( .A(n16439), .B(n13843), .ZN(n13844) );
  NAND2_X1 U17180 ( .A1(n13844), .A2(n19306), .ZN(n13857) );
  INV_X1 U17181 ( .A(n13845), .ZN(n13849) );
  INV_X1 U17182 ( .A(n13846), .ZN(n13847) );
  AOI21_X1 U17183 ( .B1(n13849), .B2(n13848), .A(n13847), .ZN(n19354) );
  INV_X2 U17184 ( .A(n19297), .ZN(n19323) );
  AOI21_X1 U17185 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19323), .A(
        n19420), .ZN(n13851) );
  NAND2_X1 U17186 ( .A1(n19311), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13850) );
  OAI211_X1 U17187 ( .C1(n19262), .C2(n13852), .A(n13851), .B(n13850), .ZN(
        n13855) );
  NOR2_X1 U17188 ( .A1(n13853), .A2(n19302), .ZN(n13854) );
  AOI211_X1 U17189 ( .C1(n19305), .C2(n19354), .A(n13855), .B(n13854), .ZN(
        n13856) );
  OAI211_X1 U17190 ( .C1(n16448), .C2(n19320), .A(n13857), .B(n13856), .ZN(
        P2_U2850) );
  INV_X1 U17191 ( .A(n19327), .ZN(n13869) );
  NAND2_X1 U17192 ( .A1(n19257), .A2(n13858), .ZN(n13859) );
  XNOR2_X1 U17193 ( .A(n13860), .B(n13859), .ZN(n13861) );
  NAND2_X1 U17194 ( .A1(n13861), .A2(n19306), .ZN(n13868) );
  AOI22_X1 U17195 ( .A1(n19305), .A2(n19361), .B1(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19323), .ZN(n13862) );
  OAI21_X1 U17196 ( .B1(n19302), .B2(n13863), .A(n13862), .ZN(n13866) );
  OAI22_X1 U17197 ( .A1(n13864), .A2(n19180), .B1(n13804), .B2(n19262), .ZN(
        n13865) );
  AOI211_X1 U17198 ( .C1(n19285), .C2(n13803), .A(n13866), .B(n13865), .ZN(
        n13867) );
  OAI211_X1 U17199 ( .C1(n20103), .C2(n13869), .A(n13868), .B(n13867), .ZN(
        P2_U2852) );
  XNOR2_X1 U17200 ( .A(n13871), .B(n13870), .ZN(n19425) );
  XNOR2_X1 U17201 ( .A(n13872), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13873) );
  XNOR2_X1 U17202 ( .A(n13874), .B(n13873), .ZN(n19422) );
  AOI21_X1 U17203 ( .B1(n13877), .B2(n13876), .A(n13875), .ZN(n16521) );
  INV_X1 U17204 ( .A(n19434), .ZN(n15841) );
  AOI22_X1 U17205 ( .A1(n16521), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n15841), .B2(n19442), .ZN(n16501) );
  NOR2_X1 U17206 ( .A1(n16522), .A2(n16523), .ZN(n16505) );
  NOR2_X1 U17207 ( .A1(n11000), .A2(n19178), .ZN(n13878) );
  AOI221_X1 U17208 ( .B1(n16501), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n16505), .C2(n16507), .A(n13878), .ZN(n13880) );
  AOI22_X1 U17209 ( .A1(n19427), .A2(n19440), .B1(n19436), .B2(n19281), .ZN(
        n13879) );
  OAI211_X1 U17210 ( .C1(n19422), .C2(n16524), .A(n13880), .B(n13879), .ZN(
        n13881) );
  INV_X1 U17211 ( .A(n13881), .ZN(n13882) );
  OAI21_X1 U17212 ( .B1(n19425), .B2(n19449), .A(n13882), .ZN(P2_U3042) );
  INV_X1 U17213 ( .A(n13884), .ZN(n13885) );
  NAND2_X1 U17214 ( .A1(n13817), .A2(n13885), .ZN(n13886) );
  AND2_X1 U17215 ( .A1(n13883), .A2(n13886), .ZN(n20261) );
  INV_X1 U17216 ( .A(n20261), .ZN(n13888) );
  OAI222_X1 U17217 ( .A1(n14904), .A2(n13888), .B1(n14903), .B2(n11898), .C1(
        n14902), .C2(n13887), .ZN(P1_U2897) );
  NAND2_X1 U17218 ( .A1(n13889), .A2(n20952), .ZN(n13908) );
  NOR2_X1 U17219 ( .A1(n13903), .A2(n14603), .ZN(n13893) );
  OR2_X1 U17220 ( .A1(n20210), .A2(n13893), .ZN(n20247) );
  INV_X1 U17221 ( .A(n20247), .ZN(n20237) );
  NOR2_X1 U17222 ( .A1(n13903), .A2(n20955), .ZN(n20227) );
  NAND2_X1 U17223 ( .A1(n11775), .A2(n20227), .ZN(n13912) );
  INV_X1 U17224 ( .A(n13894), .ZN(n15181) );
  AND2_X1 U17225 ( .A1(n13895), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13897) );
  NAND2_X1 U17226 ( .A1(n20953), .A2(n21022), .ZN(n16010) );
  NAND2_X1 U17227 ( .A1(n13897), .A2(n16010), .ZN(n13896) );
  NOR2_X2 U17228 ( .A1(n13903), .A2(n13896), .ZN(n20257) );
  INV_X1 U17229 ( .A(n13897), .ZN(n13901) );
  INV_X1 U17230 ( .A(n16010), .ZN(n13898) );
  NAND2_X1 U17231 ( .A1(n13899), .A2(n13898), .ZN(n13904) );
  NAND3_X1 U17232 ( .A1(n13901), .A2(n13900), .A3(n13904), .ZN(n13902) );
  AOI22_X1 U17233 ( .A1(n15181), .A2(n20257), .B1(n20250), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13911) );
  NOR2_X1 U17234 ( .A1(n13904), .A2(n11635), .ZN(n13905) );
  NAND2_X1 U17235 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20958), .ZN(n16013) );
  OAI211_X1 U17236 ( .C1(n16013), .C2(n20865), .A(n20351), .B(n13908), .ZN(
        n13906) );
  NAND2_X1 U17237 ( .A1(n20220), .A2(n20198), .ZN(n20203) );
  NAND2_X1 U17238 ( .A1(n20203), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13910) );
  OAI21_X1 U17239 ( .B1(n20229), .B2(n20215), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13909) );
  AND4_X1 U17240 ( .A1(n13912), .A2(n13911), .A3(n13910), .A4(n13909), .ZN(
        n13913) );
  OAI21_X1 U17241 ( .B1(n13914), .B2(n20237), .A(n13913), .ZN(P1_U2840) );
  OAI21_X1 U17242 ( .B1(n20427), .B2(n20843), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13917) );
  NAND2_X1 U17243 ( .A1(n13917), .A2(n20677), .ZN(n13927) );
  INV_X1 U17244 ( .A(n13927), .ZN(n13921) );
  OR2_X1 U17245 ( .A1(n20618), .A2(n13918), .ZN(n20433) );
  INV_X1 U17246 ( .A(n20433), .ZN(n20478) );
  NAND2_X1 U17247 ( .A1(n20478), .A2(n20619), .ZN(n13926) );
  NOR2_X1 U17248 ( .A1(n13924), .A2(n11760), .ZN(n20560) );
  INV_X1 U17249 ( .A(n20688), .ZN(n20436) );
  NAND2_X1 U17250 ( .A1(n15214), .A2(n20683), .ZN(n20508) );
  INV_X1 U17251 ( .A(n20508), .ZN(n13919) );
  NOR3_X1 U17252 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20410) );
  INV_X1 U17253 ( .A(n20410), .ZN(n20407) );
  NOR2_X1 U17254 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20407), .ZN(
        n13922) );
  OAI22_X1 U17255 ( .A1(n13919), .A2(n11760), .B1(n13922), .B2(n20689), .ZN(
        n13920) );
  AOI211_X2 U17256 ( .C1(n13921), .C2(n13926), .A(n20436), .B(n13920), .ZN(
        n20406) );
  INV_X1 U17257 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13930) );
  INV_X1 U17258 ( .A(n13922), .ZN(n20400) );
  OAI22_X1 U17259 ( .A1(n20863), .A2(n9791), .B1(n20400), .B2(n20451), .ZN(
        n13923) );
  AOI21_X1 U17260 ( .B1(n20427), .B2(n20704), .A(n13923), .ZN(n13929) );
  INV_X1 U17261 ( .A(n13924), .ZN(n13925) );
  NOR2_X1 U17262 ( .A1(n13925), .A2(n11760), .ZN(n20685) );
  INV_X1 U17263 ( .A(n20685), .ZN(n20621) );
  NAND2_X1 U17264 ( .A1(n20402), .A2(n20828), .ZN(n13928) );
  OAI211_X1 U17265 ( .C1(n20406), .C2(n13930), .A(n13929), .B(n13928), .ZN(
        P1_U3036) );
  OAI22_X1 U17266 ( .A1(n20863), .A2(n20676), .B1(n20400), .B2(n20468), .ZN(
        n13931) );
  AOI21_X1 U17267 ( .B1(n20427), .B2(n20721), .A(n13931), .ZN(n13933) );
  NAND2_X1 U17268 ( .A1(n20402), .A2(n20855), .ZN(n13932) );
  OAI211_X1 U17269 ( .C1(n20406), .C2(n13934), .A(n13933), .B(n13932), .ZN(
        P1_U3040) );
  OAI22_X1 U17270 ( .A1(n20863), .A2(n20827), .B1(n20400), .B2(n20447), .ZN(
        n13935) );
  AOI21_X1 U17271 ( .B1(n20427), .B2(n20824), .A(n13935), .ZN(n13937) );
  NAND2_X1 U17272 ( .A1(n20402), .A2(n20822), .ZN(n13936) );
  OAI211_X1 U17273 ( .C1(n20406), .C2(n13938), .A(n13937), .B(n13936), .ZN(
        P1_U3035) );
  OAI22_X1 U17274 ( .A1(n20863), .A2(n9793), .B1(n20400), .B2(n20455), .ZN(
        n13939) );
  AOI21_X1 U17275 ( .B1(n20427), .B2(n20708), .A(n13939), .ZN(n13941) );
  NAND2_X1 U17276 ( .A1(n20402), .A2(n20834), .ZN(n13940) );
  OAI211_X1 U17277 ( .C1(n20406), .C2(n13942), .A(n13941), .B(n13940), .ZN(
        P1_U3037) );
  INV_X1 U17278 ( .A(n20227), .ZN(n20253) );
  INV_X1 U17279 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13946) );
  NAND2_X1 U17280 ( .A1(n20215), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13944) );
  INV_X1 U17281 ( .A(n20198), .ZN(n20204) );
  AOI22_X1 U17282 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n20250), .B1(n20204), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13943) );
  NAND2_X1 U17283 ( .A1(n13944), .A2(n13943), .ZN(n13945) );
  AOI21_X1 U17284 ( .B1(n20229), .B2(n13946), .A(n13945), .ZN(n13949) );
  AOI22_X1 U17285 ( .A1(n20248), .A2(n13825), .B1(n20257), .B2(n13947), .ZN(
        n13948) );
  OAI211_X1 U17286 ( .C1(n20619), .C2(n20253), .A(n13949), .B(n13948), .ZN(
        n13950) );
  INV_X1 U17287 ( .A(n13950), .ZN(n13951) );
  OAI21_X1 U17288 ( .B1(n13952), .B2(n20237), .A(n13951), .ZN(P1_U2839) );
  OAI21_X1 U17289 ( .B1(n13955), .B2(n13954), .A(n13953), .ZN(n20350) );
  NAND2_X1 U17290 ( .A1(n13956), .A2(n20344), .ZN(n13960) );
  INV_X1 U17291 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n13957) );
  OAI22_X1 U17292 ( .A1(n15039), .A2(n20235), .B1(n20351), .B2(n13957), .ZN(
        n13958) );
  AOI21_X1 U17293 ( .B1(n20230), .B2(n16152), .A(n13958), .ZN(n13959) );
  OAI211_X1 U17294 ( .C1(n20350), .C2(n20167), .A(n13960), .B(n13959), .ZN(
        P1_U2995) );
  INV_X1 U17295 ( .A(n13961), .ZN(n13970) );
  XNOR2_X1 U17296 ( .A(n13962), .B(n13970), .ZN(n13968) );
  AND2_X1 U17297 ( .A1(n13964), .A2(n13963), .ZN(n13965) );
  NOR2_X1 U17298 ( .A1(n14004), .A2(n13965), .ZN(n16461) );
  NOR2_X1 U17299 ( .A1(n15442), .A2(n10739), .ZN(n13966) );
  AOI21_X1 U17300 ( .B1(n16461), .B2(n15442), .A(n13966), .ZN(n13967) );
  OAI21_X1 U17301 ( .B1(n13968), .B2(n15450), .A(n13967), .ZN(P2_U2872) );
  NOR2_X2 U17302 ( .A1(n13972), .A2(n13971), .ZN(n13985) );
  AOI22_X1 U17303 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13976) );
  AOI22_X1 U17304 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17305 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17306 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13973) );
  NAND4_X1 U17307 ( .A1(n13976), .A2(n13975), .A3(n13974), .A4(n13973), .ZN(
        n13984) );
  AOI22_X1 U17308 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13982) );
  AOI22_X1 U17309 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13978) );
  NAND2_X1 U17310 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13977) );
  AND2_X1 U17311 ( .A1(n13978), .A2(n13977), .ZN(n13981) );
  AOI22_X1 U17312 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13980) );
  NAND2_X1 U17313 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13979) );
  NAND4_X1 U17314 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        n13983) );
  OR2_X1 U17315 ( .A1(n13984), .A2(n13983), .ZN(n13986) );
  OAI21_X1 U17316 ( .B1(n13985), .B2(n13986), .A(n9801), .ZN(n14008) );
  OR2_X1 U17317 ( .A1(n13987), .A2(n13988), .ZN(n13989) );
  NAND2_X1 U17318 ( .A1(n14060), .A2(n13989), .ZN(n19202) );
  NOR2_X2 U17319 ( .A1(n13990), .A2(n19451), .ZN(n19331) );
  AOI22_X1 U17320 ( .A1(n19331), .A2(BUF1_REG_16__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n13993) );
  AOI22_X1 U17321 ( .A1(n16364), .A2(n13991), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19379), .ZN(n13992) );
  OAI211_X1 U17322 ( .C1(n15538), .C2(n19202), .A(n13993), .B(n13992), .ZN(
        n13994) );
  INV_X1 U17323 ( .A(n13994), .ZN(n13995) );
  OAI21_X1 U17324 ( .B1(n14008), .B2(n19356), .A(n13995), .ZN(P2_U2903) );
  NAND2_X1 U17325 ( .A1(n13883), .A2(n13998), .ZN(n13999) );
  AND2_X1 U17326 ( .A1(n13997), .A2(n13999), .ZN(n20191) );
  INV_X1 U17327 ( .A(n20191), .ZN(n14012) );
  INV_X1 U17328 ( .A(DATAI_8_), .ZN(n14001) );
  NAND2_X1 U17329 ( .A1(n14848), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14000) );
  OAI21_X1 U17330 ( .B1(n14848), .B2(n14001), .A(n14000), .ZN(n20305) );
  AOI22_X1 U17331 ( .A1(n14898), .A2(n20305), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16115), .ZN(n14002) );
  OAI21_X1 U17332 ( .B1(n14012), .B2(n14904), .A(n14002), .ZN(P1_U2896) );
  OR2_X1 U17333 ( .A1(n14004), .A2(n14003), .ZN(n14005) );
  AND2_X1 U17334 ( .A1(n14005), .A2(n14068), .ZN(n19198) );
  NOR2_X1 U17335 ( .A1(n15442), .A2(n10755), .ZN(n14006) );
  AOI21_X1 U17336 ( .B1(n19198), .B2(n15442), .A(n14006), .ZN(n14007) );
  OAI21_X1 U17337 ( .B1(n14008), .B2(n15450), .A(n14007), .ZN(P2_U2871) );
  INV_X1 U17338 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14011) );
  NAND2_X1 U17339 ( .A1(n16290), .A2(n14009), .ZN(n14010) );
  NAND2_X1 U17340 ( .A1(n14016), .A2(n14010), .ZN(n20187) );
  OAI222_X1 U17341 ( .A1(n14012), .A2(n14842), .B1(n14011), .B2(n20270), .C1(
        n20265), .C2(n20187), .ZN(P1_U2864) );
  AOI21_X1 U17342 ( .B1(n14014), .B2(n13997), .A(n14013), .ZN(n14021) );
  AND2_X1 U17343 ( .A1(n14016), .A2(n14015), .ZN(n14017) );
  OR2_X1 U17344 ( .A1(n14211), .A2(n14017), .ZN(n14790) );
  INV_X1 U17345 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14018) );
  OAI22_X1 U17346 ( .A1(n14790), .A2(n20265), .B1(n14018), .B2(n20270), .ZN(
        n14019) );
  AOI21_X1 U17347 ( .B1(n14021), .B2(n12977), .A(n14019), .ZN(n14020) );
  INV_X1 U17348 ( .A(n14020), .ZN(P1_U2863) );
  INV_X1 U17349 ( .A(n14021), .ZN(n15053) );
  AOI22_X1 U17350 ( .A1(n14898), .A2(n14856), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16115), .ZN(n14022) );
  OAI21_X1 U17351 ( .B1(n15053), .B2(n14904), .A(n14022), .ZN(P1_U2895) );
  OAI21_X1 U17352 ( .B1(n14013), .B2(n14024), .A(n14023), .ZN(n14209) );
  INV_X1 U17353 ( .A(DATAI_10_), .ZN(n21132) );
  NAND2_X1 U17354 ( .A1(n14848), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14025) );
  OAI21_X1 U17355 ( .B1(n14848), .B2(n21132), .A(n14025), .ZN(n20307) );
  AOI22_X1 U17356 ( .A1(n14898), .A2(n20307), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16115), .ZN(n14026) );
  OAI21_X1 U17357 ( .B1(n14209), .B2(n14904), .A(n14026), .ZN(P1_U2894) );
  NAND2_X1 U17358 ( .A1(n9717), .A2(n14027), .ZN(n14028) );
  XNOR2_X1 U17359 ( .A(n14029), .B(n14028), .ZN(n14044) );
  NAND2_X1 U17360 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14030) );
  OR2_X1 U17361 ( .A1(n15183), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20378) );
  NAND2_X1 U17362 ( .A1(n20379), .A2(n20378), .ZN(n16250) );
  OAI21_X1 U17363 ( .B1(n14030), .B2(n16250), .A(n20369), .ZN(n16243) );
  NAND2_X1 U17364 ( .A1(n14031), .A2(n16243), .ZN(n20365) );
  INV_X1 U17365 ( .A(n20365), .ZN(n16310) );
  NAND2_X1 U17366 ( .A1(n14032), .A2(n16310), .ZN(n16301) );
  NOR2_X1 U17367 ( .A1(n14033), .A2(n16301), .ZN(n16292) );
  AOI21_X1 U17368 ( .B1(n14034), .B2(n16296), .A(n16271), .ZN(n14037) );
  NOR2_X1 U17369 ( .A1(n20369), .A2(n14031), .ZN(n20371) );
  INV_X1 U17370 ( .A(n20379), .ZN(n15144) );
  OAI21_X1 U17371 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15144), .A(
        n16268), .ZN(n20374) );
  AOI211_X1 U17372 ( .C1(n20380), .C2(n20379), .A(n20371), .B(n20374), .ZN(
        n20363) );
  OAI21_X1 U17373 ( .B1(n16269), .B2(n14032), .A(n20363), .ZN(n16307) );
  AOI21_X1 U17374 ( .B1(n14033), .B2(n15175), .A(n16307), .ZN(n16297) );
  NOR2_X1 U17375 ( .A1(n16297), .A2(n14034), .ZN(n14036) );
  NAND2_X1 U17376 ( .A1(n20377), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n14040) );
  OAI21_X1 U17377 ( .B1(n20187), .B2(n20352), .A(n14040), .ZN(n14035) );
  AOI211_X1 U17378 ( .C1(n16292), .C2(n14037), .A(n14036), .B(n14035), .ZN(
        n14038) );
  OAI21_X1 U17379 ( .B1(n14044), .B2(n16278), .A(n14038), .ZN(P1_U3023) );
  NAND2_X1 U17380 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14039) );
  OAI211_X1 U17381 ( .C1(n20349), .C2(n14041), .A(n14040), .B(n14039), .ZN(
        n14042) );
  AOI21_X1 U17382 ( .B1(n20191), .B2(n20344), .A(n14042), .ZN(n14043) );
  OAI21_X1 U17383 ( .B1(n14044), .B2(n20167), .A(n14043), .ZN(P1_U2991) );
  AOI22_X1 U17384 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14048) );
  AOI22_X1 U17385 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14047) );
  AOI22_X1 U17386 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U17387 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14045) );
  NAND4_X1 U17388 ( .A1(n14048), .A2(n14047), .A3(n14046), .A4(n14045), .ZN(
        n14056) );
  AOI22_X1 U17389 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U17390 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14358), .ZN(n14050) );
  NAND2_X1 U17391 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n14049) );
  AND2_X1 U17392 ( .A1(n14050), .A2(n14049), .ZN(n14053) );
  AOI22_X1 U17393 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14052) );
  NAND2_X1 U17394 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14051) );
  NAND4_X1 U17395 ( .A1(n14054), .A2(n14053), .A3(n14052), .A4(n14051), .ZN(
        n14055) );
  OR2_X1 U17396 ( .A1(n14056), .A2(n14055), .ZN(n14058) );
  OAI21_X1 U17397 ( .B1(n14057), .B2(n14058), .A(n14180), .ZN(n14071) );
  NAND2_X1 U17398 ( .A1(n14060), .A2(n14059), .ZN(n14061) );
  AND2_X1 U17399 ( .A1(n15532), .A2(n14061), .ZN(n19185) );
  OAI22_X1 U17400 ( .A1(n19467), .A2(n15522), .B1(n19349), .B2(n14062), .ZN(
        n14065) );
  INV_X1 U17401 ( .A(n19331), .ZN(n15525) );
  INV_X1 U17402 ( .A(n19333), .ZN(n15524) );
  INV_X1 U17403 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14063) );
  OAI22_X1 U17404 ( .A1(n15525), .A2(n16631), .B1(n15524), .B2(n14063), .ZN(
        n14064) );
  AOI211_X1 U17405 ( .C1(n19380), .C2(n19185), .A(n14065), .B(n14064), .ZN(
        n14066) );
  OAI21_X1 U17406 ( .B1(n14071), .B2(n19356), .A(n14066), .ZN(P2_U2902) );
  XNOR2_X1 U17407 ( .A(n14068), .B(n14067), .ZN(n19184) );
  NOR2_X1 U17408 ( .A1(n19184), .A2(n13322), .ZN(n14069) );
  AOI21_X1 U17409 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n13273), .A(n14069), .ZN(
        n14070) );
  OAI21_X1 U17410 ( .B1(n14071), .B2(n15450), .A(n14070), .ZN(P2_U2870) );
  AND2_X1 U17411 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17134) );
  NOR3_X1 U17412 ( .A1(n14073), .A2(n14072), .A3(n17564), .ZN(n14076) );
  INV_X1 U17413 ( .A(n18853), .ZN(n14075) );
  NOR4_X2 U17414 ( .A1(n19074), .A2(n18416), .A3(n16038), .A4(n18924), .ZN(
        n17437) );
  NAND2_X1 U17415 ( .A1(n18448), .A2(n17437), .ZN(n17439) );
  INV_X2 U17416 ( .A(n17435), .ZN(n17431) );
  INV_X1 U17417 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16824) );
  INV_X1 U17418 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17239) );
  INV_X1 U17419 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16910) );
  INV_X1 U17420 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17003) );
  INV_X1 U17421 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17404) );
  NAND4_X1 U17422 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n15933)
         );
  INV_X1 U17423 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16938) );
  INV_X1 U17424 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17305) );
  NOR2_X1 U17425 ( .A1(n16938), .A2(n17305), .ZN(n17290) );
  INV_X1 U17426 ( .A(n17290), .ZN(n14077) );
  NOR4_X1 U17427 ( .A1(n17003), .A2(n17404), .A3(n15933), .A4(n14077), .ZN(
        n17292) );
  INV_X1 U17428 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17403) );
  INV_X1 U17429 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17418) );
  INV_X1 U17430 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17079) );
  NAND3_X1 U17431 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17422) );
  NOR3_X1 U17432 ( .A1(n17079), .A2(n17423), .A3(n17422), .ZN(n17411) );
  NAND2_X1 U17433 ( .A1(n17437), .A2(n17411), .ZN(n17417) );
  NAND3_X1 U17434 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17292), .A3(n17402), 
        .ZN(n17276) );
  NAND2_X1 U17435 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17264), .ZN(n17238) );
  AND4_X1 U17436 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17135)
         );
  NAND2_X1 U17437 ( .A1(n17223), .A2(n17135), .ZN(n17180) );
  NOR2_X1 U17438 ( .A1(n16824), .A2(n17180), .ZN(n17185) );
  NAND2_X1 U17439 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17185), .ZN(n17178) );
  NAND2_X1 U17440 ( .A1(n17431), .A2(n17178), .ZN(n14078) );
  OAI21_X1 U17441 ( .B1(n17134), .B2(n17439), .A(n14078), .ZN(n17169) );
  AOI22_X1 U17442 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17443 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17444 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U17445 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14079) );
  NAND4_X1 U17446 ( .A1(n14082), .A2(n14081), .A3(n14080), .A4(n14079), .ZN(
        n14088) );
  AOI22_X1 U17447 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17448 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U17449 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U17450 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14083) );
  NAND4_X1 U17451 ( .A1(n14086), .A2(n14085), .A3(n14084), .A4(n14083), .ZN(
        n14087) );
  NOR2_X1 U17452 ( .A1(n14088), .A2(n14087), .ZN(n14153) );
  AOI22_X1 U17453 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17454 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U17455 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U17456 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14089) );
  NAND4_X1 U17457 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14098) );
  AOI22_X1 U17458 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U17459 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17460 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U17461 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14093) );
  NAND4_X1 U17462 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        n14097) );
  NOR2_X1 U17463 ( .A1(n14098), .A2(n14097), .ZN(n17176) );
  AOI22_X1 U17464 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12574), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U17465 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17367), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17369), .ZN(n14101) );
  AOI22_X1 U17466 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17385), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12550), .ZN(n14100) );
  AOI22_X1 U17467 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17387), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17386), .ZN(n14099) );
  NAND4_X1 U17468 ( .A1(n14102), .A2(n14101), .A3(n14100), .A4(n14099), .ZN(
        n14108) );
  AOI22_X1 U17469 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U17470 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17365), .ZN(n14105) );
  AOI22_X1 U17471 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17393), .ZN(n14104) );
  AOI22_X1 U17472 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14103) );
  NAND4_X1 U17473 ( .A1(n14106), .A2(n14105), .A3(n14104), .A4(n14103), .ZN(
        n14107) );
  NOR2_X1 U17474 ( .A1(n14108), .A2(n14107), .ZN(n17187) );
  AOI22_X1 U17475 ( .A1(n12581), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14119) );
  AOI22_X1 U17476 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14118) );
  INV_X1 U17477 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18495) );
  AOI22_X1 U17478 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14109) );
  OAI21_X1 U17479 ( .B1(n14110), .B2(n18495), .A(n14109), .ZN(n14116) );
  AOI22_X1 U17480 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17481 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12574), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17482 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U17483 ( .A1(n17369), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14111) );
  NAND4_X1 U17484 ( .A1(n14114), .A2(n14113), .A3(n14112), .A4(n14111), .ZN(
        n14115) );
  AOI211_X1 U17485 ( .C1(n17395), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n14116), .B(n14115), .ZN(n14117) );
  NAND3_X1 U17486 ( .A1(n14119), .A2(n14118), .A3(n14117), .ZN(n17192) );
  AOI22_X1 U17487 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U17488 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14130) );
  INV_X1 U17489 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17490 ( .A1(n12581), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14120) );
  OAI21_X1 U17491 ( .B1(n14122), .B2(n14121), .A(n14120), .ZN(n14128) );
  AOI22_X1 U17492 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17493 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17494 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14124) );
  AOI22_X1 U17495 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14123) );
  NAND4_X1 U17496 ( .A1(n14126), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        n14127) );
  AOI211_X1 U17497 ( .C1(n17366), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14128), .B(n14127), .ZN(n14129) );
  NAND3_X1 U17498 ( .A1(n14131), .A2(n14130), .A3(n14129), .ZN(n17193) );
  NAND2_X1 U17499 ( .A1(n17192), .A2(n17193), .ZN(n17191) );
  NOR2_X1 U17500 ( .A1(n17187), .A2(n17191), .ZN(n17183) );
  AOI22_X1 U17501 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14142) );
  AOI22_X1 U17502 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U17503 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14132) );
  OAI21_X1 U17504 ( .B1(n17150), .B2(n14133), .A(n14132), .ZN(n14139) );
  AOI22_X1 U17505 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17506 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U17507 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14135) );
  AOI22_X1 U17508 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14134) );
  NAND4_X1 U17509 ( .A1(n14137), .A2(n14136), .A3(n14135), .A4(n14134), .ZN(
        n14138) );
  AOI211_X1 U17510 ( .C1(n12550), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n14139), .B(n14138), .ZN(n14140) );
  NAND3_X1 U17511 ( .A1(n14142), .A2(n14141), .A3(n14140), .ZN(n17182) );
  NAND2_X1 U17512 ( .A1(n17183), .A2(n17182), .ZN(n17181) );
  NOR2_X1 U17513 ( .A1(n17176), .A2(n17181), .ZN(n17175) );
  AOI22_X1 U17514 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14152) );
  AOI22_X1 U17515 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U17516 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14143) );
  OAI21_X1 U17517 ( .B1(n17150), .B2(n17424), .A(n14143), .ZN(n14149) );
  AOI22_X1 U17518 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17519 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17520 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U17521 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14144) );
  NAND4_X1 U17522 ( .A1(n14147), .A2(n14146), .A3(n14145), .A4(n14144), .ZN(
        n14148) );
  AOI211_X1 U17523 ( .C1(n12550), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n14149), .B(n14148), .ZN(n14150) );
  NAND3_X1 U17524 ( .A1(n14152), .A2(n14151), .A3(n14150), .ZN(n17172) );
  NAND2_X1 U17525 ( .A1(n17175), .A2(n17172), .ZN(n17171) );
  NOR2_X1 U17526 ( .A1(n14153), .A2(n17171), .ZN(n17166) );
  AOI21_X1 U17527 ( .B1(n14153), .B2(n17171), .A(n17166), .ZN(n17457) );
  AOI22_X1 U17528 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17169), .B1(n17457), 
        .B2(n17435), .ZN(n14157) );
  INV_X1 U17529 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14155) );
  INV_X1 U17530 ( .A(n17178), .ZN(n14154) );
  NAND3_X1 U17531 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14155), .A3(n14154), 
        .ZN(n14156) );
  NAND2_X1 U17532 ( .A1(n14157), .A2(n14156), .ZN(P3_U2675) );
  XNOR2_X1 U17533 ( .A(n14159), .B(n14158), .ZN(n14228) );
  OAI21_X1 U17534 ( .B1(n14161), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14160), .ZN(n14162) );
  INV_X1 U17535 ( .A(n14162), .ZN(n14226) );
  OAI22_X1 U17536 ( .A1(n11007), .A2(n19178), .B1(n19432), .B2(n19271), .ZN(
        n14163) );
  INV_X1 U17537 ( .A(n14163), .ZN(n14165) );
  NAND2_X1 U17538 ( .A1(n19421), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14164) );
  OAI211_X1 U17539 ( .C1(n19276), .C2(n15688), .A(n14165), .B(n14164), .ZN(
        n14166) );
  AOI21_X1 U17540 ( .B1(n14226), .B2(n16449), .A(n14166), .ZN(n14167) );
  OAI21_X1 U17541 ( .B1(n19424), .B2(n14228), .A(n14167), .ZN(P2_U3008) );
  AOI22_X1 U17542 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U17543 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U17544 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14169) );
  AOI22_X1 U17545 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14168) );
  NAND4_X1 U17546 ( .A1(n14171), .A2(n14170), .A3(n14169), .A4(n14168), .ZN(
        n14179) );
  AOI22_X1 U17547 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14177) );
  AOI22_X1 U17548 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14358), .ZN(n14173) );
  NAND2_X1 U17549 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n14172) );
  AND2_X1 U17550 ( .A1(n14173), .A2(n14172), .ZN(n14176) );
  AOI22_X1 U17551 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14175) );
  NAND2_X1 U17552 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14174) );
  NAND4_X1 U17553 ( .A1(n14177), .A2(n14176), .A3(n14175), .A4(n14174), .ZN(
        n14178) );
  NOR2_X1 U17554 ( .A1(n14179), .A2(n14178), .ZN(n14183) );
  INV_X1 U17555 ( .A(n14183), .ZN(n14181) );
  INV_X1 U17556 ( .A(n14204), .ZN(n14182) );
  AOI21_X1 U17557 ( .B1(n14183), .B2(n14180), .A(n14182), .ZN(n15540) );
  NAND2_X1 U17558 ( .A1(n15540), .A2(n15434), .ZN(n14187) );
  AOI21_X1 U17559 ( .B1(n14185), .B2(n14184), .A(n14190), .ZN(n19170) );
  NAND2_X1 U17560 ( .A1(n19170), .A2(n15442), .ZN(n14186) );
  OAI211_X1 U17561 ( .C1(n15442), .C2(n19164), .A(n14187), .B(n14186), .ZN(
        P2_U2869) );
  OR2_X1 U17562 ( .A1(n14190), .A2(n14189), .ZN(n14191) );
  NAND2_X1 U17563 ( .A1(n14188), .A2(n14191), .ZN(n19159) );
  AOI22_X1 U17564 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14195) );
  AOI22_X1 U17565 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U17566 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14193) );
  AOI22_X1 U17567 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14192) );
  NAND4_X1 U17568 ( .A1(n14195), .A2(n14194), .A3(n14193), .A4(n14192), .ZN(
        n14203) );
  AOI22_X1 U17569 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U17570 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14358), .ZN(n14197) );
  NAND2_X1 U17571 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14196) );
  AND2_X1 U17572 ( .A1(n14197), .A2(n14196), .ZN(n14200) );
  AOI22_X1 U17573 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U17574 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14198) );
  NAND4_X1 U17575 ( .A1(n14201), .A2(n14200), .A3(n14199), .A4(n14198), .ZN(
        n14202) );
  NOR2_X1 U17576 ( .A1(n14203), .A2(n14202), .ZN(n14206) );
  AOI21_X1 U17577 ( .B1(n14206), .B2(n14204), .A(n14205), .ZN(n15517) );
  NAND2_X1 U17578 ( .A1(n15517), .A2(n15434), .ZN(n14208) );
  NAND2_X1 U17579 ( .A1(n13273), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14207) );
  OAI211_X1 U17580 ( .C1(n19159), .C2(n13273), .A(n14208), .B(n14207), .ZN(
        P2_U2868) );
  INV_X1 U17581 ( .A(n14209), .ZN(n16154) );
  OR2_X1 U17582 ( .A1(n14211), .A2(n14210), .ZN(n14212) );
  NAND2_X1 U17583 ( .A1(n14781), .A2(n14212), .ZN(n16273) );
  OAI22_X1 U17584 ( .A1(n16273), .A2(n20265), .B1(n16103), .B2(n20270), .ZN(
        n14213) );
  AOI21_X1 U17585 ( .B1(n16154), .B2(n12977), .A(n14213), .ZN(n14214) );
  INV_X1 U17586 ( .A(n14214), .ZN(P1_U2862) );
  AOI22_X1 U17587 ( .A1(n15841), .A2(n19442), .B1(n14215), .B2(n16521), .ZN(
        n16496) );
  INV_X1 U17588 ( .A(n16496), .ZN(n14217) );
  NAND2_X1 U17589 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19420), .ZN(n14216) );
  OAI221_X1 U17590 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14219), .C1(
        n14218), .C2(n14217), .A(n14216), .ZN(n14225) );
  OR2_X1 U17591 ( .A1(n14221), .A2(n14220), .ZN(n14222) );
  NAND2_X1 U17592 ( .A1(n14223), .A2(n14222), .ZN(n19350) );
  OAI22_X1 U17593 ( .A1(n19276), .A2(n16527), .B1(n16526), .B2(n19350), .ZN(
        n14224) );
  AOI211_X1 U17594 ( .C1(n14226), .C2(n19438), .A(n14225), .B(n14224), .ZN(
        n14227) );
  OAI21_X1 U17595 ( .B1(n19449), .B2(n14228), .A(n14227), .ZN(P2_U3040) );
  INV_X1 U17596 ( .A(n15674), .ZN(n14230) );
  NOR2_X1 U17597 ( .A1(n14230), .A2(n15673), .ZN(n14231) );
  XNOR2_X1 U17598 ( .A(n14229), .B(n14231), .ZN(n16434) );
  XNOR2_X1 U17599 ( .A(n14233), .B(n11192), .ZN(n14234) );
  XNOR2_X1 U17600 ( .A(n14232), .B(n14234), .ZN(n16431) );
  NOR2_X1 U17601 ( .A1(n11012), .A2(n16466), .ZN(n14235) );
  AOI221_X1 U17602 ( .B1(n16496), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n16491), .C2(n11192), .A(n14235), .ZN(n14237) );
  NAND2_X1 U17603 ( .A1(n19263), .A2(n19440), .ZN(n14236) );
  OAI211_X1 U17604 ( .C1(n16526), .C2(n19264), .A(n14237), .B(n14236), .ZN(
        n14238) );
  AOI21_X1 U17605 ( .B1(n16431), .B2(n19438), .A(n14238), .ZN(n14239) );
  OAI21_X1 U17606 ( .B1(n16434), .B2(n19449), .A(n14239), .ZN(P2_U3039) );
  NOR2_X1 U17607 ( .A1(n17422), .A2(n17439), .ZN(n17427) );
  INV_X1 U17608 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17438) );
  INV_X1 U17609 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17433) );
  NOR2_X1 U17610 ( .A1(n17438), .A2(n17433), .ZN(n14240) );
  AOI21_X1 U17611 ( .B1(n17437), .B2(n14240), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n14241) );
  NOR2_X1 U17612 ( .A1(n17427), .A2(n14241), .ZN(n14242) );
  MUX2_X1 U17613 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B(n14242), .S(n17431), 
        .Z(P3_U2701) );
  INV_X1 U17614 ( .A(n12540), .ZN(n18873) );
  AOI21_X1 U17615 ( .B1(n18873), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15950) );
  NAND2_X1 U17616 ( .A1(n15950), .A2(n17197), .ZN(n18403) );
  NOR2_X1 U17617 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18403), .ZN(n14243) );
  NAND3_X1 U17618 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19026)
         );
  OAI21_X1 U17619 ( .B1(n14243), .B2(n19026), .A(n18453), .ZN(n18409) );
  INV_X1 U17620 ( .A(n18409), .ZN(n14244) );
  NOR2_X1 U17621 ( .A1(n19068), .A2(n17907), .ZN(n15936) );
  AOI21_X1 U17622 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15936), .ZN(n15937) );
  NOR2_X1 U17623 ( .A1(n14244), .A2(n15937), .ZN(n14246) );
  INV_X1 U17624 ( .A(n18654), .ZN(n18758) );
  NOR2_X1 U17625 ( .A1(n19028), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18452) );
  OR2_X1 U17626 ( .A1(n18452), .A2(n14244), .ZN(n15935) );
  OR2_X1 U17627 ( .A1(n18758), .A2(n15935), .ZN(n14245) );
  MUX2_X1 U17628 ( .A(n14246), .B(n14245), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17629 ( .A(n14287), .ZN(n14249) );
  INV_X1 U17630 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14277) );
  NOR2_X1 U17631 ( .A1(n20351), .A2(n14277), .ZN(n15078) );
  AOI21_X1 U17632 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15078), .ZN(n14248) );
  OAI21_X1 U17633 ( .B1(n20349), .B2(n14249), .A(n14248), .ZN(n14250) );
  AOI21_X1 U17634 ( .B1(n14251), .B2(n20344), .A(n14250), .ZN(n14252) );
  INV_X1 U17635 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14255) );
  XNOR2_X1 U17636 ( .A(n14634), .B(n14254), .ZN(n15086) );
  OAI222_X1 U17637 ( .A1(n14851), .A2(n14842), .B1(n14255), .B2(n20270), .C1(
        n20265), .C2(n15086), .ZN(P1_U2844) );
  AOI22_X1 U17638 ( .A1(n12927), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14611), .ZN(n14609) );
  OAI22_X1 U17639 ( .A1(n14610), .A2(n12962), .B1(n14257), .B2(n14256), .ZN(
        n14258) );
  XOR2_X1 U17640 ( .A(n14609), .B(n14258), .Z(n15069) );
  INV_X1 U17641 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14280) );
  OAI222_X1 U17642 ( .A1(n20265), .A2(n15069), .B1(n14280), .B2(n20270), .C1(
        n14285), .C2(n14842), .ZN(P1_U2842) );
  AOI22_X1 U17643 ( .A1(n16118), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16115), .ZN(n14262) );
  INV_X1 U17644 ( .A(DATAI_14_), .ZN(n21125) );
  NAND2_X1 U17645 ( .A1(n14848), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14259) );
  OAI21_X1 U17646 ( .B1(n14260), .B2(n21125), .A(n14259), .ZN(n20313) );
  AOI22_X1 U17647 ( .A1(n16117), .A2(n20313), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n14885), .ZN(n14261) );
  OAI211_X1 U17648 ( .C1(n14285), .C2(n14904), .A(n14262), .B(n14261), .ZN(
        P1_U2874) );
  NAND3_X1 U17649 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n14274) );
  NAND3_X1 U17650 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14717) );
  NAND2_X1 U17651 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n16075) );
  INV_X1 U17652 ( .A(n16075), .ZN(n16067) );
  NAND3_X1 U17653 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n16067), .ZN(n14270) );
  INV_X1 U17654 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20894) );
  INV_X1 U17655 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20891) );
  INV_X1 U17656 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20219) );
  NAND4_X1 U17657 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20232)
         );
  NOR3_X1 U17658 ( .A1(n20891), .A2(n20219), .A3(n20232), .ZN(n20202) );
  NAND2_X1 U17659 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20202), .ZN(n20184) );
  NOR2_X1 U17660 ( .A1(n20894), .A2(n20184), .ZN(n14268) );
  NAND3_X1 U17661 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n14789), .ZN(n16074) );
  NOR2_X1 U17662 ( .A1(n14270), .A2(n16074), .ZN(n14771) );
  NAND4_X1 U17663 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .A4(n14771), .ZN(n14738) );
  NOR2_X1 U17664 ( .A1(n14717), .A2(n14738), .ZN(n14726) );
  NAND2_X1 U17665 ( .A1(n14726), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14263) );
  INV_X1 U17666 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14264) );
  NOR2_X1 U17667 ( .A1(n14718), .A2(n14264), .ZN(n14265) );
  NAND2_X1 U17668 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14265), .ZN(n14661) );
  NOR2_X1 U17669 ( .A1(n14274), .A2(n14661), .ZN(n14631) );
  NAND2_X1 U17670 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14276) );
  INV_X1 U17671 ( .A(n14276), .ZN(n14266) );
  AND2_X1 U17672 ( .A1(n14631), .A2(n14266), .ZN(n14286) );
  NAND2_X1 U17673 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14614) );
  INV_X1 U17674 ( .A(n14614), .ZN(n14267) );
  AOI21_X1 U17675 ( .B1(n14286), .B2(n14267), .A(n14788), .ZN(n14618) );
  NAND2_X1 U17676 ( .A1(n20248), .A2(n14268), .ZN(n16100) );
  NAND2_X1 U17677 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14269) );
  INV_X1 U17678 ( .A(n14270), .ZN(n14271) );
  NAND2_X1 U17679 ( .A1(n16089), .A2(n14271), .ZN(n14772) );
  INV_X1 U17680 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n16226) );
  AND2_X1 U17681 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14272) );
  NAND2_X1 U17682 ( .A1(n16044), .A2(n14272), .ZN(n14748) );
  INV_X1 U17683 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20989) );
  NAND2_X1 U17684 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14273) );
  INV_X1 U17685 ( .A(n14274), .ZN(n14275) );
  NAND2_X1 U17686 ( .A1(n14679), .A2(n14275), .ZN(n14640) );
  OAI21_X1 U17687 ( .B1(n14615), .B2(n14277), .A(n21005), .ZN(n14283) );
  AOI22_X1 U17688 ( .A1(n20229), .A2(n14278), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20215), .ZN(n14279) );
  OAI21_X1 U17689 ( .B1(n16102), .B2(n14280), .A(n14279), .ZN(n14282) );
  NOR2_X1 U17690 ( .A1(n15069), .A2(n20243), .ZN(n14281) );
  AOI211_X1 U17691 ( .C1(n14618), .C2(n14283), .A(n14282), .B(n14281), .ZN(
        n14284) );
  OAI21_X1 U17692 ( .B1(n14285), .B2(n16093), .A(n14284), .ZN(P1_U2810) );
  NOR2_X1 U17693 ( .A1(n14286), .A2(n14788), .ZN(n14627) );
  NOR2_X1 U17694 ( .A1(n14615), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14291) );
  AOI22_X1 U17695 ( .A1(n20229), .A2(n14287), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20215), .ZN(n14289) );
  NAND2_X1 U17696 ( .A1(n20250), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14288) );
  OAI211_X1 U17697 ( .C1(n15081), .C2(n20243), .A(n14289), .B(n14288), .ZN(
        n14290) );
  AOI211_X1 U17698 ( .C1(n14627), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14291), 
        .B(n14290), .ZN(n14292) );
  OAI21_X1 U17699 ( .B1(n14293), .B2(n16093), .A(n14292), .ZN(P1_U2811) );
  AOI22_X1 U17700 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U17701 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U17702 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14295) );
  AOI22_X1 U17703 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14294) );
  NAND4_X1 U17704 ( .A1(n14297), .A2(n14296), .A3(n14295), .A4(n14294), .ZN(
        n14305) );
  AOI22_X1 U17705 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U17706 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14358), .ZN(n14299) );
  NAND2_X1 U17707 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n14298) );
  AND2_X1 U17708 ( .A1(n14299), .A2(n14298), .ZN(n14302) );
  AOI22_X1 U17709 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U17710 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14300) );
  NAND4_X1 U17711 ( .A1(n14303), .A2(n14302), .A3(n14301), .A4(n14300), .ZN(
        n14304) );
  OR2_X1 U17712 ( .A1(n14305), .A2(n14304), .ZN(n15445) );
  AOI22_X1 U17713 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U17714 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14309) );
  AOI22_X1 U17715 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14308) );
  AOI22_X1 U17716 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14353), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14307) );
  NAND4_X1 U17717 ( .A1(n14310), .A2(n14309), .A3(n14308), .A4(n14307), .ZN(
        n14318) );
  AOI22_X1 U17718 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U17719 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14358), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U17720 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n14311) );
  AND2_X1 U17721 ( .A1(n14312), .A2(n14311), .ZN(n14315) );
  AOI22_X1 U17722 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U17723 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14313) );
  NAND4_X1 U17724 ( .A1(n14316), .A2(n14315), .A3(n14314), .A4(n14313), .ZN(
        n14317) );
  OR2_X1 U17725 ( .A1(n14318), .A2(n14317), .ZN(n15439) );
  AOI22_X1 U17726 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11033), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14324) );
  AOI22_X1 U17727 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17728 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14322) );
  AOI22_X1 U17729 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14353), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14321) );
  NAND4_X1 U17730 ( .A1(n14324), .A2(n14323), .A3(n14322), .A4(n14321), .ZN(
        n14332) );
  AOI22_X1 U17731 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U17732 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14358), .ZN(n14326) );
  NAND2_X1 U17733 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14325) );
  AND2_X1 U17734 ( .A1(n14326), .A2(n14325), .ZN(n14329) );
  AOI22_X1 U17735 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10659), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14328) );
  NAND2_X1 U17736 ( .A1(n14352), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n14327) );
  NAND4_X1 U17737 ( .A1(n14330), .A2(n14329), .A3(n14328), .A4(n14327), .ZN(
        n14331) );
  OR2_X1 U17738 ( .A1(n14332), .A2(n14331), .ZN(n15430) );
  NAND2_X1 U17739 ( .A1(n15431), .A2(n15430), .ZN(n14369) );
  AOI22_X1 U17740 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17741 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U17742 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9682), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14339) );
  NAND2_X1 U17743 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14337) );
  NAND2_X1 U17744 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14336) );
  NAND2_X1 U17745 ( .A1(n14333), .A2(n10275), .ZN(n14335) );
  AND2_X1 U17746 ( .A1(n14335), .A2(n14334), .ZN(n14476) );
  AND3_X1 U17747 ( .A1(n14337), .A2(n14336), .A3(n14476), .ZN(n14338) );
  NAND4_X1 U17748 ( .A1(n14341), .A2(n14340), .A3(n14339), .A4(n14338), .ZN(
        n14349) );
  AOI22_X1 U17749 ( .A1(n9647), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14347) );
  AOI22_X1 U17750 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10451), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U17751 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U17752 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14343) );
  NAND2_X1 U17753 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14342) );
  INV_X1 U17754 ( .A(n14476), .ZN(n14505) );
  AND3_X1 U17755 ( .A1(n14343), .A2(n14342), .A3(n14505), .ZN(n14344) );
  NAND4_X1 U17756 ( .A1(n14347), .A2(n14346), .A3(n14345), .A4(n14344), .ZN(
        n14348) );
  NAND2_X1 U17757 ( .A1(n14349), .A2(n14348), .ZN(n14390) );
  NOR2_X1 U17758 ( .A1(n10458), .A2(n14390), .ZN(n14368) );
  AOI22_X1 U17759 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10658), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U17760 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11033), .B1(
        n10654), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U17761 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10644), .B1(
        n14351), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U17762 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14353), .B1(
        n14352), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14354) );
  NAND4_X1 U17763 ( .A1(n14357), .A2(n14356), .A3(n14355), .A4(n14354), .ZN(
        n14367) );
  AOI22_X1 U17764 ( .A1(n11015), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10632), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14365) );
  AOI22_X1 U17765 ( .A1(n10653), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n10524), .ZN(n14364) );
  AOI22_X1 U17766 ( .A1(n14359), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14358), .ZN(n14361) );
  NAND2_X1 U17767 ( .A1(n10659), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14360) );
  AND2_X1 U17768 ( .A1(n14361), .A2(n14360), .ZN(n14363) );
  NAND2_X1 U17769 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n14362) );
  NAND4_X1 U17770 ( .A1(n14365), .A2(n14364), .A3(n14363), .A4(n14362), .ZN(
        n14366) );
  OR2_X1 U17771 ( .A1(n14367), .A2(n14366), .ZN(n14387) );
  XNOR2_X1 U17772 ( .A(n14368), .B(n14387), .ZN(n14391) );
  INV_X1 U17773 ( .A(n14390), .ZN(n14386) );
  NAND2_X1 U17774 ( .A1(n10458), .A2(n14386), .ZN(n15422) );
  INV_X1 U17775 ( .A(n14369), .ZN(n15432) );
  INV_X1 U17776 ( .A(n14391), .ZN(n14370) );
  AND2_X2 U17777 ( .A1(n15432), .A2(n14370), .ZN(n14371) );
  AOI22_X1 U17778 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U17779 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U17780 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U17781 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14373) );
  NAND2_X1 U17782 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14372) );
  AND3_X1 U17783 ( .A1(n14373), .A2(n14372), .A3(n14505), .ZN(n14374) );
  NAND4_X1 U17784 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        n14385) );
  AOI22_X1 U17785 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U17786 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U17787 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14381) );
  NAND2_X1 U17788 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14379) );
  NAND2_X1 U17789 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14378) );
  AND3_X1 U17790 ( .A1(n14379), .A2(n14378), .A3(n14476), .ZN(n14380) );
  NAND4_X1 U17791 ( .A1(n14383), .A2(n14382), .A3(n14381), .A4(n14380), .ZN(
        n14384) );
  NAND2_X1 U17792 ( .A1(n14385), .A2(n14384), .ZN(n14393) );
  NAND2_X1 U17793 ( .A1(n14387), .A2(n14386), .ZN(n14394) );
  XOR2_X1 U17794 ( .A(n14393), .B(n14394), .Z(n14388) );
  NAND2_X1 U17795 ( .A1(n14388), .A2(n14450), .ZN(n15416) );
  INV_X1 U17796 ( .A(n14393), .ZN(n14389) );
  NAND2_X1 U17797 ( .A1(n10458), .A2(n14389), .ZN(n15418) );
  NOR3_X1 U17798 ( .A1(n14391), .A2(n14390), .A3(n15418), .ZN(n14392) );
  NOR2_X1 U17799 ( .A1(n14394), .A2(n14393), .ZN(n14409) );
  AOI22_X1 U17800 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14400) );
  AOI22_X1 U17801 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U17802 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14398) );
  NAND2_X1 U17803 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14396) );
  NAND2_X1 U17804 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14395) );
  AND3_X1 U17805 ( .A1(n14396), .A2(n14395), .A3(n14505), .ZN(n14397) );
  NAND4_X1 U17806 ( .A1(n14400), .A2(n14399), .A3(n14398), .A4(n14397), .ZN(
        n14408) );
  AOI22_X1 U17807 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U17808 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U17809 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14404) );
  NAND2_X1 U17810 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14402) );
  NAND2_X1 U17811 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14401) );
  AND3_X1 U17812 ( .A1(n14402), .A2(n14401), .A3(n14476), .ZN(n14403) );
  NAND4_X1 U17813 ( .A1(n14406), .A2(n14405), .A3(n14404), .A4(n14403), .ZN(
        n14407) );
  AND2_X1 U17814 ( .A1(n14408), .A2(n14407), .ZN(n14411) );
  NAND2_X1 U17815 ( .A1(n14409), .A2(n14411), .ZN(n14430) );
  OAI211_X1 U17816 ( .C1(n14409), .C2(n14411), .A(n14450), .B(n14430), .ZN(
        n14413) );
  INV_X1 U17817 ( .A(n14411), .ZN(n14412) );
  NOR2_X1 U17818 ( .A1(n14487), .A2(n14412), .ZN(n15408) );
  NAND2_X1 U17819 ( .A1(n15406), .A2(n15408), .ZN(n15407) );
  AOI22_X1 U17820 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U17821 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14419) );
  AOI22_X1 U17822 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14418) );
  NAND2_X1 U17823 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14416) );
  NAND2_X1 U17824 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14415) );
  AND3_X1 U17825 ( .A1(n14416), .A2(n14415), .A3(n14505), .ZN(n14417) );
  NAND4_X1 U17826 ( .A1(n14420), .A2(n14419), .A3(n14418), .A4(n14417), .ZN(
        n14428) );
  AOI22_X1 U17827 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U17828 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14425) );
  AOI22_X1 U17829 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14424) );
  NAND2_X1 U17830 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14422) );
  NAND2_X1 U17831 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14421) );
  AND3_X1 U17832 ( .A1(n14422), .A2(n14421), .A3(n14476), .ZN(n14423) );
  NAND4_X1 U17833 ( .A1(n14426), .A2(n14425), .A3(n14424), .A4(n14423), .ZN(
        n14427) );
  NAND2_X1 U17834 ( .A1(n14428), .A2(n14427), .ZN(n14432) );
  AOI21_X1 U17835 ( .B1(n14430), .B2(n14432), .A(n14429), .ZN(n14431) );
  OR2_X1 U17836 ( .A1(n14430), .A2(n14432), .ZN(n14449) );
  INV_X1 U17837 ( .A(n14432), .ZN(n14433) );
  NAND2_X1 U17838 ( .A1(n10458), .A2(n14433), .ZN(n15403) );
  AOI22_X1 U17839 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U17840 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U17841 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14438) );
  NAND2_X1 U17842 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14436) );
  NAND2_X1 U17843 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14435) );
  AND3_X1 U17844 ( .A1(n14436), .A2(n14435), .A3(n14505), .ZN(n14437) );
  NAND4_X1 U17845 ( .A1(n14440), .A2(n14439), .A3(n14438), .A4(n14437), .ZN(
        n14448) );
  AOI22_X1 U17846 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U17847 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14445) );
  AOI22_X1 U17848 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14444) );
  NAND2_X1 U17849 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14442) );
  NAND2_X1 U17850 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14441) );
  AND3_X1 U17851 ( .A1(n14442), .A2(n14441), .A3(n14476), .ZN(n14443) );
  NAND4_X1 U17852 ( .A1(n14446), .A2(n14445), .A3(n14444), .A4(n14443), .ZN(
        n14447) );
  NAND2_X1 U17853 ( .A1(n14448), .A2(n14447), .ZN(n14454) );
  INV_X1 U17854 ( .A(n14454), .ZN(n14452) );
  INV_X1 U17855 ( .A(n14449), .ZN(n14451) );
  OR2_X1 U17856 ( .A1(n14449), .A2(n14454), .ZN(n14485) );
  OAI211_X1 U17857 ( .C1(n14452), .C2(n14451), .A(n14485), .B(n14450), .ZN(
        n14453) );
  NOR2_X1 U17858 ( .A1(n14487), .A2(n14454), .ZN(n15398) );
  NAND2_X1 U17859 ( .A1(n15396), .A2(n15398), .ZN(n15397) );
  AOI22_X1 U17860 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9643), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U17861 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U17862 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U17863 ( .A1(n14461), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14456) );
  NAND2_X1 U17864 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14455) );
  AND3_X1 U17865 ( .A1(n14456), .A2(n14455), .A3(n14505), .ZN(n14457) );
  NAND4_X1 U17866 ( .A1(n14460), .A2(n14459), .A3(n14458), .A4(n14457), .ZN(
        n14469) );
  AOI22_X1 U17867 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9647), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U17868 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U17869 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U17870 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14463) );
  NAND2_X1 U17871 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14462) );
  AND3_X1 U17872 ( .A1(n14463), .A2(n14462), .A3(n14476), .ZN(n14464) );
  NAND4_X1 U17873 ( .A1(n14467), .A2(n14466), .A3(n14465), .A4(n14464), .ZN(
        n14468) );
  NAND2_X1 U17874 ( .A1(n14469), .A2(n14468), .ZN(n15392) );
  AOI22_X1 U17875 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14475) );
  AOI22_X1 U17876 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14474) );
  AOI22_X1 U17877 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14473) );
  NAND2_X1 U17878 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14471) );
  NAND2_X1 U17879 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14470) );
  AND3_X1 U17880 ( .A1(n14471), .A2(n14470), .A3(n14505), .ZN(n14472) );
  NAND4_X1 U17881 ( .A1(n14475), .A2(n14474), .A3(n14473), .A4(n14472), .ZN(
        n14484) );
  AOI22_X1 U17882 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U17883 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U17884 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14480) );
  NAND2_X1 U17885 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14478) );
  NAND2_X1 U17886 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14477) );
  AND3_X1 U17887 ( .A1(n14478), .A2(n14477), .A3(n14476), .ZN(n14479) );
  NAND4_X1 U17888 ( .A1(n14482), .A2(n14481), .A3(n14480), .A4(n14479), .ZN(
        n14483) );
  NAND2_X1 U17889 ( .A1(n14484), .A2(n14483), .ZN(n14490) );
  INV_X1 U17890 ( .A(n14485), .ZN(n15390) );
  INV_X1 U17891 ( .A(n15392), .ZN(n14486) );
  AND2_X1 U17892 ( .A1(n14487), .A2(n14486), .ZN(n14488) );
  NAND2_X1 U17893 ( .A1(n15390), .A2(n14488), .ZN(n14489) );
  NOR2_X1 U17894 ( .A1(n14489), .A2(n14490), .ZN(n14491) );
  AOI21_X1 U17895 ( .B1(n14490), .B2(n14489), .A(n14491), .ZN(n15386) );
  INV_X1 U17896 ( .A(n14491), .ZN(n14492) );
  AOI22_X1 U17897 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14499), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U17898 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U17899 ( .A1(n14494), .A2(n14493), .ZN(n14512) );
  INV_X1 U17900 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14497) );
  AOI22_X1 U17901 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14496) );
  AOI21_X1 U17902 ( .B1(n14504), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14505), .ZN(n14495) );
  OAI211_X1 U17903 ( .C1(n14498), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        n14511) );
  AOI22_X1 U17904 ( .A1(n10441), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14499), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U17905 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14500), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14501) );
  NAND2_X1 U17906 ( .A1(n14502), .A2(n14501), .ZN(n14510) );
  AOI22_X1 U17907 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14503), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14508) );
  NAND2_X1 U17908 ( .A1(n14504), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14507) );
  NAND2_X1 U17909 ( .A1(n10451), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14506) );
  NAND4_X1 U17910 ( .A1(n14508), .A2(n14507), .A3(n14506), .A4(n14505), .ZN(
        n14509) );
  OAI22_X1 U17911 ( .A1(n14512), .A2(n14511), .B1(n14510), .B2(n14509), .ZN(
        n14513) );
  INV_X1 U17912 ( .A(n14513), .ZN(n14514) );
  INV_X1 U17913 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20087) );
  NAND2_X1 U17914 ( .A1(n11210), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14516) );
  AOI22_X1 U17915 ( .A1(n14561), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n14515) );
  OAI211_X1 U17916 ( .C1(n14517), .C2(n20087), .A(n14516), .B(n14515), .ZN(
        n14559) );
  NOR2_X1 U17917 ( .A1(n15699), .A2(n13322), .ZN(n14518) );
  AOI21_X1 U17918 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n13273), .A(n14518), .ZN(
        n14519) );
  OAI21_X1 U17919 ( .B1(n14526), .B2(n15450), .A(n14519), .ZN(P2_U2857) );
  INV_X1 U17920 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14521) );
  AOI22_X1 U17921 ( .A1(n16364), .A2(n19341), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19379), .ZN(n14520) );
  OAI21_X1 U17922 ( .B1(n15524), .B2(n14521), .A(n14520), .ZN(n14524) );
  AOI22_X1 U17923 ( .A1(n14577), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14522) );
  OAI21_X1 U17924 ( .B1(n14579), .B2(n20087), .A(n14522), .ZN(n14575) );
  NOR2_X1 U17925 ( .A1(n15692), .A2(n15538), .ZN(n14523) );
  AOI211_X1 U17926 ( .C1(BUF1_REG_30__SCAN_IN), .C2(n19331), .A(n14524), .B(
        n14523), .ZN(n14525) );
  OAI21_X1 U17927 ( .B1(n14526), .B2(n19356), .A(n14525), .ZN(P2_U2889) );
  AOI22_X1 U17928 ( .A1(n11777), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14531), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14536) );
  AND2_X1 U17929 ( .A1(n14533), .A2(n14532), .ZN(n14534) );
  NAND2_X1 U17930 ( .A1(n14534), .A2(n14629), .ZN(n14535) );
  INV_X1 U17931 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21004) );
  NOR2_X1 U17932 ( .A1(n20351), .A2(n21004), .ZN(n15064) );
  AOI21_X1 U17933 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15064), .ZN(n14537) );
  OAI21_X1 U17934 ( .B1(n20349), .B2(n14538), .A(n14537), .ZN(n14539) );
  AOI21_X1 U17935 ( .B1(n14844), .B2(n20344), .A(n14539), .ZN(n14540) );
  OAI21_X1 U17936 ( .B1(n15068), .B2(n20167), .A(n14540), .ZN(P1_U2968) );
  INV_X1 U17937 ( .A(n19098), .ZN(n20148) );
  INV_X1 U17938 ( .A(n19096), .ZN(n14541) );
  OAI21_X1 U17939 ( .B1(n14541), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20148), 
        .ZN(n14542) );
  OAI21_X1 U17940 ( .B1(n13122), .B2(n20148), .A(n14542), .ZN(P2_U3612) );
  NAND2_X1 U17941 ( .A1(n15542), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14544) );
  NAND2_X1 U17942 ( .A1(n14546), .A2(n14545), .ZN(n15544) );
  NAND2_X1 U17943 ( .A1(n14548), .A2(n14547), .ZN(n14553) );
  NAND2_X1 U17944 ( .A1(n14552), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14549) );
  XNOR2_X1 U17945 ( .A(n14553), .B(n14549), .ZN(n15286) );
  AOI21_X1 U17946 ( .B1(n15286), .B2(n14550), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15545) );
  INV_X1 U17947 ( .A(n15286), .ZN(n14551) );
  INV_X1 U17948 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14584) );
  OAI21_X1 U17949 ( .B1(n14553), .B2(P2_EBX_REG_30__SCAN_IN), .A(n14552), .ZN(
        n14555) );
  NAND2_X1 U17950 ( .A1(n14555), .A2(n14554), .ZN(n15273) );
  NOR2_X1 U17951 ( .A1(n15273), .A2(n10536), .ZN(n14556) );
  XOR2_X1 U17952 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14556), .Z(
        n14557) );
  XNOR2_X1 U17953 ( .A(n14558), .B(n14557), .ZN(n14574) );
  NAND2_X1 U17954 ( .A1(n14560), .A2(n14559), .ZN(n14566) );
  AOI22_X1 U17955 ( .A1(n14561), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14564) );
  NAND2_X1 U17956 ( .A1(n14562), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14563) );
  OAI211_X1 U17957 ( .C1(n10387), .C2(n14543), .A(n14564), .B(n14563), .ZN(
        n14565) );
  INV_X1 U17958 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14569) );
  NAND2_X1 U17959 ( .A1(n16440), .A2(n14567), .ZN(n14568) );
  NAND2_X1 U17960 ( .A1(n19420), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14586) );
  OAI211_X1 U17961 ( .C1(n16453), .C2(n14569), .A(n14568), .B(n14586), .ZN(
        n14570) );
  AOI21_X1 U17962 ( .B1(n15382), .B2(n19428), .A(n14570), .ZN(n14571) );
  OAI21_X1 U17963 ( .B1(n14574), .B2(n19424), .A(n14571), .ZN(n14572) );
  INV_X1 U17964 ( .A(n14572), .ZN(n14573) );
  OAI21_X1 U17965 ( .B1(n14593), .B2(n19423), .A(n14573), .ZN(P2_U2983) );
  INV_X1 U17966 ( .A(n14574), .ZN(n14592) );
  INV_X1 U17967 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U17968 ( .A1(n14577), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11032), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14578) );
  OAI21_X1 U17969 ( .B1(n14579), .B2(n15271), .A(n14578), .ZN(n14580) );
  NOR2_X1 U17970 ( .A1(n14582), .A2(n14581), .ZN(n14583) );
  NAND2_X1 U17971 ( .A1(n15705), .A2(n14583), .ZN(n15696) );
  NOR3_X1 U17972 ( .A1(n15696), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14584), .ZN(n14589) );
  OAI21_X1 U17973 ( .B1(n15841), .B2(n14583), .A(n15710), .ZN(n15693) );
  AOI21_X1 U17974 ( .B1(n14584), .B2(n19434), .A(n15693), .ZN(n14585) );
  OR2_X1 U17975 ( .A1(n14585), .A2(n14543), .ZN(n14587) );
  NAND2_X1 U17976 ( .A1(n14587), .A2(n14586), .ZN(n14588) );
  NAND3_X1 U17977 ( .A1(n9686), .A2(n14595), .A3(n14594), .ZN(n14597) );
  MUX2_X1 U17978 ( .A(n14598), .B(n14597), .S(n14596), .Z(n14599) );
  INV_X1 U17979 ( .A(n14599), .ZN(n14602) );
  NAND2_X1 U17980 ( .A1(n13002), .A2(n14600), .ZN(n14601) );
  NAND2_X1 U17981 ( .A1(n14602), .A2(n14601), .ZN(n16003) );
  NAND3_X1 U17982 ( .A1(n14611), .A2(n14603), .A3(n16029), .ZN(n14608) );
  INV_X1 U17983 ( .A(n9686), .ZN(n14606) );
  OAI22_X1 U17984 ( .A1(n14607), .A2(n14606), .B1(n14605), .B2(n14604), .ZN(
        n20163) );
  AOI21_X1 U17985 ( .B1(n20953), .B2(n14608), .A(n20163), .ZN(n16006) );
  NOR2_X1 U17986 ( .A1(n16006), .A2(n20162), .ZN(n20169) );
  MUX2_X1 U17987 ( .A(P1_MORE_REG_SCAN_IN), .B(n16003), .S(n20169), .Z(
        P1_U3484) );
  AOI22_X1 U17988 ( .A1(n12927), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14611), .ZN(n14612) );
  NAND2_X1 U17989 ( .A1(n14844), .A2(n20210), .ZN(n14620) );
  INV_X1 U17990 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14804) );
  INV_X1 U17991 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14613) );
  OAI22_X1 U17992 ( .A1(n16102), .A2(n14804), .B1(n14613), .B2(n20245), .ZN(
        n14617) );
  NOR3_X1 U17993 ( .A1(n14615), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14614), 
        .ZN(n14616) );
  AOI211_X1 U17994 ( .C1(n14618), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14617), 
        .B(n14616), .ZN(n14619) );
  OAI211_X1 U17995 ( .C1(n15059), .C2(n20243), .A(n14620), .B(n14619), .ZN(
        P1_U2809) );
  OAI22_X1 U17996 ( .A1(n20244), .A2(n14622), .B1(n14621), .B2(n20245), .ZN(
        n14624) );
  INV_X1 U17997 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21069) );
  NOR3_X1 U17998 ( .A1(n14640), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n21069), 
        .ZN(n14623) );
  AOI211_X1 U17999 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n20250), .A(n14624), .B(
        n14623), .ZN(n14625) );
  OAI21_X1 U18000 ( .B1(n15086), .B2(n20243), .A(n14625), .ZN(n14626) );
  AOI21_X1 U18001 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14627), .A(n14626), 
        .ZN(n14628) );
  OAI21_X1 U18002 ( .B1(n14851), .B2(n16093), .A(n14628), .ZN(P1_U2812) );
  NOR2_X1 U18003 ( .A1(n14631), .A2(n14788), .ZN(n14655) );
  OAI22_X1 U18004 ( .A1(n20244), .A2(n14909), .B1(n14632), .B2(n20245), .ZN(
        n14638) );
  AND2_X1 U18005 ( .A1(n14665), .A2(n14633), .ZN(n14636) );
  OAI21_X1 U18006 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n15101) );
  NOR2_X1 U18007 ( .A1(n15101), .A2(n20243), .ZN(n14637) );
  AOI211_X1 U18008 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n20250), .A(n14638), .B(
        n14637), .ZN(n14639) );
  OAI21_X1 U18009 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14640), .A(n14639), 
        .ZN(n14641) );
  AOI21_X1 U18010 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14655), .A(n14641), 
        .ZN(n14642) );
  OAI21_X1 U18011 ( .B1(n14907), .B2(n16093), .A(n14642), .ZN(P1_U2813) );
  NAND2_X1 U18012 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14643) );
  NOR2_X1 U18013 ( .A1(n14643), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14648) );
  NAND2_X1 U18014 ( .A1(n20250), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14645) );
  NAND2_X1 U18015 ( .A1(n20229), .A2(n14913), .ZN(n14644) );
  OAI211_X1 U18016 ( .C1(n20245), .C2(n14646), .A(n14645), .B(n14644), .ZN(
        n14647) );
  AOI21_X1 U18017 ( .B1(n14679), .B2(n14648), .A(n14647), .ZN(n14649) );
  OAI21_X1 U18018 ( .B1(n14806), .B2(n20243), .A(n14649), .ZN(n14654) );
  NOR2_X1 U18019 ( .A1(n14921), .A2(n16093), .ZN(n14653) );
  INV_X1 U18020 ( .A(n14656), .ZN(P1_U2814) );
  INV_X1 U18021 ( .A(n14673), .ZN(n14658) );
  NAND2_X1 U18022 ( .A1(n14657), .A2(n14658), .ZN(n14659) );
  AOI21_X1 U18023 ( .B1(n14660), .B2(n14659), .A(n14650), .ZN(n14931) );
  INV_X1 U18024 ( .A(n14931), .ZN(n14859) );
  XOR2_X1 U18025 ( .A(P1_REIP_REG_24__SCAN_IN), .B(P1_REIP_REG_25__SCAN_IN), 
        .Z(n14671) );
  NAND2_X1 U18026 ( .A1(n14661), .A2(n20203), .ZN(n14693) );
  INV_X1 U18027 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20968) );
  NOR2_X1 U18028 ( .A1(n14693), .A2(n20968), .ZN(n14670) );
  NOR2_X1 U18029 ( .A1(n14662), .A2(n14663), .ZN(n14664) );
  OR2_X1 U18030 ( .A1(n14665), .A2(n14664), .ZN(n15106) );
  INV_X1 U18031 ( .A(n14929), .ZN(n14666) );
  AOI22_X1 U18032 ( .A1(n20229), .A2(n14666), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20215), .ZN(n14668) );
  NAND2_X1 U18033 ( .A1(n20250), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n14667) );
  OAI211_X1 U18034 ( .C1(n15106), .C2(n20243), .A(n14668), .B(n14667), .ZN(
        n14669) );
  AOI211_X1 U18035 ( .C1(n14679), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        n14672) );
  OAI21_X1 U18036 ( .B1(n14859), .B2(n16093), .A(n14672), .ZN(P1_U2815) );
  INV_X1 U18037 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21087) );
  XNOR2_X1 U18038 ( .A(n14657), .B(n14673), .ZN(n14941) );
  NAND2_X1 U18039 ( .A1(n14941), .A2(n20210), .ZN(n14681) );
  NOR2_X1 U18040 ( .A1(n14687), .A2(n14674), .ZN(n14675) );
  OR2_X1 U18041 ( .A1(n14662), .A2(n14675), .ZN(n15115) );
  AOI22_X1 U18042 ( .A1(n20229), .A2(n14937), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20215), .ZN(n14677) );
  NAND2_X1 U18043 ( .A1(n20250), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14676) );
  OAI211_X1 U18044 ( .C1(n15115), .C2(n20243), .A(n14677), .B(n14676), .ZN(
        n14678) );
  AOI21_X1 U18045 ( .B1(n14679), .B2(n21087), .A(n14678), .ZN(n14680) );
  OAI211_X1 U18046 ( .C1(n21087), .C2(n14693), .A(n14681), .B(n14680), .ZN(
        P1_U2816) );
  INV_X1 U18047 ( .A(n14706), .ZN(n14682) );
  AOI21_X1 U18048 ( .B1(n14682), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14694) );
  AOI21_X1 U18049 ( .B1(n14684), .B2(n10190), .A(n14657), .ZN(n14947) );
  NAND2_X1 U18050 ( .A1(n14947), .A2(n20210), .ZN(n14692) );
  INV_X1 U18051 ( .A(n14685), .ZN(n14945) );
  OAI22_X1 U18052 ( .A1(n20244), .A2(n14945), .B1(n14686), .B2(n20245), .ZN(
        n14690) );
  AOI21_X1 U18053 ( .B1(n14688), .B2(n14699), .A(n14687), .ZN(n16178) );
  INV_X1 U18054 ( .A(n16178), .ZN(n14811) );
  NOR2_X1 U18055 ( .A1(n14811), .A2(n20243), .ZN(n14689) );
  AOI211_X1 U18056 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20250), .A(n14690), .B(
        n14689), .ZN(n14691) );
  OAI211_X1 U18057 ( .C1(n14694), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        P1_U2817) );
  AOI21_X1 U18058 ( .B1(n14696), .B2(n14695), .A(n14683), .ZN(n14956) );
  NAND2_X1 U18059 ( .A1(n14956), .A2(n20210), .ZN(n14705) );
  NAND2_X1 U18060 ( .A1(n14714), .A2(n14697), .ZN(n14698) );
  NAND2_X1 U18061 ( .A1(n14699), .A2(n14698), .ZN(n16188) );
  INV_X1 U18062 ( .A(n16188), .ZN(n14703) );
  NAND2_X1 U18063 ( .A1(n14718), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14701) );
  AOI22_X1 U18064 ( .A1(n20229), .A2(n14952), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20215), .ZN(n14700) );
  OAI211_X1 U18065 ( .C1(n14812), .C2(n16102), .A(n14701), .B(n14700), .ZN(
        n14702) );
  AOI21_X1 U18066 ( .B1(n14703), .B2(n20257), .A(n14702), .ZN(n14704) );
  OAI211_X1 U18067 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14706), .A(n14705), 
        .B(n14704), .ZN(P1_U2818) );
  OAI21_X1 U18068 ( .B1(n14707), .B2(n14708), .A(n14695), .ZN(n14962) );
  INV_X1 U18069 ( .A(n14709), .ZN(n14964) );
  OAI22_X1 U18070 ( .A1(n20244), .A2(n14964), .B1(n14710), .B2(n20245), .ZN(
        n14716) );
  NAND2_X1 U18071 ( .A1(n14711), .A2(n14712), .ZN(n14713) );
  NAND2_X1 U18072 ( .A1(n14714), .A2(n14713), .ZN(n15126) );
  NOR2_X1 U18073 ( .A1(n15126), .A2(n20243), .ZN(n14715) );
  AOI211_X1 U18074 ( .C1(n20250), .C2(P1_EBX_REG_21__SCAN_IN), .A(n14716), .B(
        n14715), .ZN(n14721) );
  NOR2_X1 U18075 ( .A1(n14748), .A2(n14717), .ZN(n14719) );
  OAI21_X1 U18076 ( .B1(n14719), .B2(P1_REIP_REG_21__SCAN_IN), .A(n14718), 
        .ZN(n14720) );
  OAI211_X1 U18077 ( .C1(n14962), .C2(n16093), .A(n14721), .B(n14720), .ZN(
        P1_U2819) );
  XNOR2_X1 U18078 ( .A(n14722), .B(n14723), .ZN(n14975) );
  OAI21_X1 U18079 ( .B1(n14737), .B2(n14724), .A(n14711), .ZN(n15139) );
  INV_X1 U18080 ( .A(n15139), .ZN(n14730) );
  INV_X1 U18081 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14816) );
  AOI22_X1 U18082 ( .A1(n20229), .A2(n14979), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20215), .ZN(n14725) );
  OAI21_X1 U18083 ( .B1(n16102), .B2(n14816), .A(n14725), .ZN(n14729) );
  INV_X1 U18084 ( .A(n14748), .ZN(n14762) );
  NAND3_X1 U18085 ( .A1(n14762), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n14727) );
  INV_X1 U18086 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21123) );
  AOI211_X1 U18087 ( .C1(n14727), .C2(n21123), .A(n14788), .B(n14726), .ZN(
        n14728) );
  AOI211_X1 U18088 ( .C1(n14730), .C2(n20257), .A(n14729), .B(n14728), .ZN(
        n14731) );
  OAI21_X1 U18089 ( .B1(n14975), .B2(n16093), .A(n14731), .ZN(P1_U2820) );
  XNOR2_X1 U18090 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14747) );
  AOI21_X1 U18091 ( .B1(n14734), .B2(n14733), .A(n14722), .ZN(n14988) );
  NAND2_X1 U18092 ( .A1(n14988), .A2(n20210), .ZN(n14746) );
  NOR2_X1 U18093 ( .A1(n14752), .A2(n14735), .ZN(n14736) );
  OR2_X1 U18094 ( .A1(n14737), .A2(n14736), .ZN(n14817) );
  INV_X1 U18095 ( .A(n14817), .ZN(n16201) );
  NAND2_X1 U18096 ( .A1(n20203), .A2(n14738), .ZN(n16054) );
  INV_X1 U18097 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14743) );
  NAND2_X1 U18098 ( .A1(n20215), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14739) );
  NAND2_X1 U18099 ( .A1(n14739), .A2(n20351), .ZN(n14740) );
  AOI21_X1 U18100 ( .B1(n14984), .B2(n20229), .A(n14740), .ZN(n14742) );
  NAND2_X1 U18101 ( .A1(n20250), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14741) );
  OAI211_X1 U18102 ( .C1(n16054), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        n14744) );
  AOI21_X1 U18103 ( .B1(n16201), .B2(n20257), .A(n14744), .ZN(n14745) );
  OAI211_X1 U18104 ( .C1(n14748), .C2(n14747), .A(n14746), .B(n14745), .ZN(
        P1_U2821) );
  OAI21_X1 U18105 ( .B1(n9660), .B2(n9780), .A(n14733), .ZN(n14997) );
  INV_X1 U18106 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14761) );
  AND2_X1 U18107 ( .A1(n9693), .A2(n14751), .ZN(n14753) );
  OR2_X1 U18108 ( .A1(n14753), .A2(n14752), .ZN(n15153) );
  INV_X1 U18109 ( .A(n16054), .ZN(n14758) );
  NAND2_X1 U18110 ( .A1(n20250), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14756) );
  NAND2_X1 U18111 ( .A1(n20229), .A2(n14995), .ZN(n14755) );
  NAND2_X1 U18112 ( .A1(n20215), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14754) );
  NAND4_X1 U18113 ( .A1(n14756), .A2(n14755), .A3(n20351), .A4(n14754), .ZN(
        n14757) );
  AOI21_X1 U18114 ( .B1(n14758), .B2(P1_REIP_REG_18__SCAN_IN), .A(n14757), 
        .ZN(n14759) );
  OAI21_X1 U18115 ( .B1(n15153), .B2(n20243), .A(n14759), .ZN(n14760) );
  AOI21_X1 U18116 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14763) );
  OAI21_X1 U18117 ( .B1(n14997), .B2(n16093), .A(n14763), .ZN(P1_U2822) );
  AOI21_X1 U18118 ( .B1(n14767), .B2(n14764), .A(n14766), .ZN(n15006) );
  INV_X1 U18119 ( .A(n15006), .ZN(n14888) );
  OAI21_X1 U18120 ( .B1(n14826), .B2(n14768), .A(n9747), .ZN(n16219) );
  AOI22_X1 U18121 ( .A1(n15002), .A2(n20229), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n20250), .ZN(n14769) );
  OAI21_X1 U18122 ( .B1(n20243), .B2(n16219), .A(n14769), .ZN(n14770) );
  AOI211_X1 U18123 ( .C1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n20215), .A(
        n20377), .B(n14770), .ZN(n14775) );
  NOR2_X1 U18124 ( .A1(n14771), .A2(n14788), .ZN(n16069) );
  INV_X1 U18125 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20906) );
  NOR2_X1 U18126 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14772), .ZN(n16058) );
  OR3_X1 U18127 ( .A1(n16069), .A2(n20906), .A3(n16058), .ZN(n14773) );
  OAI21_X1 U18128 ( .B1(n16044), .B2(P1_REIP_REG_16__SCAN_IN), .A(n14773), 
        .ZN(n14774) );
  OAI211_X1 U18129 ( .C1(n14888), .C2(n16093), .A(n14775), .B(n14774), .ZN(
        P1_U2824) );
  OAI21_X1 U18130 ( .B1(n14776), .B2(n14778), .A(n14777), .ZN(n15044) );
  INV_X1 U18131 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20899) );
  INV_X1 U18132 ( .A(n16074), .ZN(n14779) );
  NOR2_X1 U18133 ( .A1(n14788), .A2(n14779), .ZN(n16105) );
  INV_X1 U18134 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14785) );
  AOI21_X1 U18135 ( .B1(n20215), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20377), .ZN(n14784) );
  INV_X1 U18136 ( .A(n16080), .ZN(n14780) );
  AOI21_X1 U18137 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n16258) );
  AOI22_X1 U18138 ( .A1(n15041), .A2(n20229), .B1(n20257), .B2(n16258), .ZN(
        n14783) );
  OAI211_X1 U18139 ( .C1(n14785), .C2(n16102), .A(n14784), .B(n14783), .ZN(
        n14786) );
  AOI221_X1 U18140 ( .B1(n16089), .B2(n20899), .C1(n16105), .C2(
        P1_REIP_REG_11__SCAN_IN), .A(n14786), .ZN(n14787) );
  OAI21_X1 U18141 ( .B1(n15044), .B2(n16093), .A(n14787), .ZN(P1_U2829) );
  NOR2_X1 U18142 ( .A1(n14789), .A2(n14788), .ZN(n20190) );
  OAI22_X1 U18143 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n16100), .B1(n15049), 
        .B2(n20244), .ZN(n14794) );
  INV_X1 U18144 ( .A(n14790), .ZN(n16280) );
  AOI22_X1 U18145 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20250), .B1(n20257), .B2(
        n16280), .ZN(n14791) );
  OAI211_X1 U18146 ( .C1(n20245), .C2(n14792), .A(n14791), .B(n20351), .ZN(
        n14793) );
  AOI211_X1 U18147 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20190), .A(n14794), .B(
        n14793), .ZN(n14795) );
  OAI21_X1 U18148 ( .B1(n15053), .B2(n16093), .A(n14795), .ZN(P1_U2831) );
  OAI22_X1 U18149 ( .A1(n20348), .A2(n20244), .B1(n20243), .B2(n20366), .ZN(
        n14796) );
  AOI21_X1 U18150 ( .B1(n20215), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14796), .ZN(n14798) );
  NAND2_X1 U18151 ( .A1(n20250), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n14797) );
  OAI211_X1 U18152 ( .C1(n9689), .C2(n20253), .A(n14798), .B(n14797), .ZN(
        n14802) );
  INV_X1 U18153 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14800) );
  NAND2_X1 U18154 ( .A1(n20248), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14799) );
  NAND2_X1 U18155 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20231) );
  AOI21_X1 U18156 ( .B1(n20248), .B2(n20231), .A(n20204), .ZN(n20259) );
  AOI21_X1 U18157 ( .B1(n14800), .B2(n14799), .A(n20259), .ZN(n14801) );
  AOI211_X1 U18158 ( .C1(n20345), .C2(n20247), .A(n14802), .B(n14801), .ZN(
        n14803) );
  INV_X1 U18159 ( .A(n14803), .ZN(P1_U2838) );
  OAI22_X1 U18160 ( .A1(n15059), .A2(n20265), .B1(n20270), .B2(n14804), .ZN(
        P1_U2841) );
  OAI222_X1 U18161 ( .A1(n14907), .A2(n14842), .B1(n14805), .B2(n20270), .C1(
        n15101), .C2(n20265), .ZN(P1_U2845) );
  INV_X1 U18162 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14807) );
  OAI222_X1 U18163 ( .A1(n14842), .A2(n14921), .B1(n14807), .B2(n20270), .C1(
        n20265), .C2(n14806), .ZN(P1_U2846) );
  OAI222_X1 U18164 ( .A1(n14859), .A2(n14842), .B1(n14808), .B2(n20270), .C1(
        n15106), .C2(n20265), .ZN(P1_U2847) );
  INV_X1 U18165 ( .A(n14941), .ZN(n14862) );
  INV_X1 U18166 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14809) );
  OAI222_X1 U18167 ( .A1(n14862), .A2(n14842), .B1(n14809), .B2(n20270), .C1(
        n15115), .C2(n20265), .ZN(P1_U2848) );
  INV_X1 U18168 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14810) );
  INV_X1 U18169 ( .A(n14947), .ZN(n14866) );
  OAI222_X1 U18170 ( .A1(n14811), .A2(n20265), .B1(n14810), .B2(n20270), .C1(
        n14866), .C2(n14842), .ZN(P1_U2849) );
  INV_X1 U18171 ( .A(n14956), .ZN(n14870) );
  OAI222_X1 U18172 ( .A1(n16188), .A2(n20265), .B1(n14812), .B2(n20270), .C1(
        n14870), .C2(n14842), .ZN(P1_U2850) );
  INV_X1 U18173 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14813) );
  OAI22_X1 U18174 ( .A1(n15126), .A2(n20265), .B1(n14813), .B2(n20270), .ZN(
        n14814) );
  INV_X1 U18175 ( .A(n14814), .ZN(n14815) );
  OAI21_X1 U18176 ( .B1(n14962), .B2(n14842), .A(n14815), .ZN(P1_U2851) );
  OAI222_X1 U18177 ( .A1(n14975), .A2(n14842), .B1(n14816), .B2(n20270), .C1(
        n15139), .C2(n20265), .ZN(P1_U2852) );
  INV_X1 U18178 ( .A(n14988), .ZN(n14880) );
  OAI222_X1 U18179 ( .A1(n14880), .A2(n14842), .B1(n14818), .B2(n20270), .C1(
        n14817), .C2(n20265), .ZN(P1_U2853) );
  INV_X1 U18180 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14819) );
  OAI222_X1 U18181 ( .A1(n15153), .A2(n20265), .B1(n20270), .B2(n14819), .C1(
        n14997), .C2(n14842), .ZN(P1_U2854) );
  INV_X1 U18182 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14820) );
  OAI222_X1 U18183 ( .A1(n14888), .A2(n14842), .B1(n20270), .B2(n14820), .C1(
        n16219), .C2(n20265), .ZN(P1_U2856) );
  INV_X1 U18184 ( .A(n14764), .ZN(n14822) );
  AOI21_X1 U18185 ( .B1(n14823), .B2(n14821), .A(n14822), .ZN(n16142) );
  INV_X1 U18186 ( .A(n16142), .ZN(n14891) );
  NOR2_X1 U18187 ( .A1(n14832), .A2(n14824), .ZN(n14825) );
  OR2_X1 U18188 ( .A1(n14826), .A2(n14825), .ZN(n16056) );
  OAI222_X1 U18189 ( .A1(n14891), .A2(n14842), .B1(n14827), .B2(n20270), .C1(
        n20265), .C2(n16056), .ZN(P1_U2857) );
  NAND2_X1 U18190 ( .A1(n14829), .A2(n14830), .ZN(n14831) );
  AND2_X1 U18191 ( .A1(n14821), .A2(n14831), .ZN(n16070) );
  INV_X1 U18192 ( .A(n16070), .ZN(n14893) );
  AOI21_X1 U18193 ( .B1(n14833), .B2(n16081), .A(n14832), .ZN(n16065) );
  AOI22_X1 U18194 ( .A1(n16065), .A2(n12975), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14840), .ZN(n14834) );
  OAI21_X1 U18195 ( .B1(n14893), .B2(n14842), .A(n14834), .ZN(P1_U2858) );
  NAND3_X1 U18196 ( .A1(n14777), .A2(n10182), .A3(n14837), .ZN(n14838) );
  NAND2_X1 U18197 ( .A1(n14835), .A2(n14838), .ZN(n16094) );
  XNOR2_X1 U18198 ( .A(n16080), .B(n16076), .ZN(n16245) );
  AOI22_X1 U18199 ( .A1(n16245), .A2(n12975), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14840), .ZN(n14839) );
  OAI21_X1 U18200 ( .B1(n16094), .B2(n14842), .A(n14839), .ZN(P1_U2860) );
  AOI22_X1 U18201 ( .A1(n16258), .A2(n12975), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14840), .ZN(n14841) );
  OAI21_X1 U18202 ( .B1(n15044), .B2(n14842), .A(n14841), .ZN(P1_U2861) );
  NAND3_X1 U18203 ( .A1(n14844), .A2(n14843), .A3(n14903), .ZN(n14846) );
  AOI22_X1 U18204 ( .A1(n16118), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16115), .ZN(n14845) );
  OAI211_X1 U18205 ( .C1(n16122), .C2(n19497), .A(n14846), .B(n14845), .ZN(
        P1_U2873) );
  AOI22_X1 U18206 ( .A1(n16118), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16115), .ZN(n14850) );
  INV_X1 U18207 ( .A(DATAI_12_), .ZN(n21074) );
  NAND2_X1 U18208 ( .A1(n14848), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14847) );
  OAI21_X1 U18209 ( .B1(n14848), .B2(n21074), .A(n14847), .ZN(n20309) );
  AOI22_X1 U18210 ( .A1(n16117), .A2(n20309), .B1(BUF1_REG_28__SCAN_IN), .B2(
        n14885), .ZN(n14849) );
  OAI211_X1 U18211 ( .C1(n14851), .C2(n14904), .A(n14850), .B(n14849), .ZN(
        P1_U2876) );
  AOI22_X1 U18212 ( .A1(n16118), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16115), .ZN(n14853) );
  AOI22_X1 U18213 ( .A1(n16117), .A2(n14900), .B1(n14885), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14852) );
  OAI211_X1 U18214 ( .C1(n14907), .C2(n14904), .A(n14853), .B(n14852), .ZN(
        P1_U2877) );
  AOI22_X1 U18215 ( .A1(n16118), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n16115), .ZN(n14855) );
  AOI22_X1 U18216 ( .A1(n16117), .A2(n20307), .B1(n14885), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14854) );
  OAI211_X1 U18217 ( .C1(n14921), .C2(n14904), .A(n14855), .B(n14854), .ZN(
        P1_U2878) );
  AOI22_X1 U18218 ( .A1(n16118), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16115), .ZN(n14858) );
  AOI22_X1 U18219 ( .A1(n16117), .A2(n14856), .B1(n14885), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14857) );
  OAI211_X1 U18220 ( .C1(n14859), .C2(n14904), .A(n14858), .B(n14857), .ZN(
        P1_U2879) );
  AOI22_X1 U18221 ( .A1(n16118), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16115), .ZN(n14861) );
  AOI22_X1 U18222 ( .A1(n16117), .A2(n20305), .B1(n14885), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14860) );
  OAI211_X1 U18223 ( .C1(n14862), .C2(n14904), .A(n14861), .B(n14860), .ZN(
        P1_U2880) );
  AOI22_X1 U18224 ( .A1(n16118), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16115), .ZN(n14865) );
  AOI22_X1 U18225 ( .A1(n16117), .A2(n14863), .B1(n14885), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14864) );
  OAI211_X1 U18226 ( .C1(n14866), .C2(n14904), .A(n14865), .B(n14864), .ZN(
        P1_U2881) );
  AOI22_X1 U18227 ( .A1(n16118), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16115), .ZN(n14869) );
  AOI22_X1 U18228 ( .A1(n16117), .A2(n14867), .B1(n14885), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14868) );
  OAI211_X1 U18229 ( .C1(n14870), .C2(n14904), .A(n14869), .B(n14868), .ZN(
        P1_U2882) );
  AOI22_X1 U18230 ( .A1(n16118), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16115), .ZN(n14873) );
  AOI22_X1 U18231 ( .A1(n16117), .A2(n14871), .B1(n14885), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14872) );
  OAI211_X1 U18232 ( .C1(n14962), .C2(n14904), .A(n14873), .B(n14872), .ZN(
        P1_U2883) );
  AOI22_X1 U18233 ( .A1(n16118), .A2(DATAI_20_), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16115), .ZN(n14876) );
  AOI22_X1 U18234 ( .A1(n16117), .A2(n14874), .B1(n14885), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14875) );
  OAI211_X1 U18235 ( .C1(n14975), .C2(n14904), .A(n14876), .B(n14875), .ZN(
        P1_U2884) );
  AOI22_X1 U18236 ( .A1(n16118), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16115), .ZN(n14879) );
  AOI22_X1 U18237 ( .A1(n16117), .A2(n14877), .B1(n14885), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14878) );
  OAI211_X1 U18238 ( .C1(n14880), .C2(n14904), .A(n14879), .B(n14878), .ZN(
        P1_U2885) );
  AOI22_X1 U18239 ( .A1(n16117), .A2(n14881), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16115), .ZN(n14883) );
  AOI22_X1 U18240 ( .A1(n16118), .A2(DATAI_18_), .B1(n14885), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14882) );
  OAI211_X1 U18241 ( .C1(n14997), .C2(n14904), .A(n14883), .B(n14882), .ZN(
        P1_U2886) );
  AOI22_X1 U18242 ( .A1(n16117), .A2(n14884), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16115), .ZN(n14887) );
  AOI22_X1 U18243 ( .A1(n16118), .A2(DATAI_16_), .B1(n14885), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14886) );
  OAI211_X1 U18244 ( .C1(n14888), .C2(n14904), .A(n14887), .B(n14886), .ZN(
        P1_U2888) );
  OAI222_X1 U18245 ( .A1(n14904), .A2(n14891), .B1(n14903), .B2(n14890), .C1(
        n14902), .C2(n14889), .ZN(P1_U2889) );
  AOI22_X1 U18246 ( .A1(n14898), .A2(n20313), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16115), .ZN(n14892) );
  OAI21_X1 U18247 ( .B1(n14893), .B2(n14904), .A(n14892), .ZN(P1_U2890) );
  NAND2_X1 U18248 ( .A1(n14835), .A2(n14894), .ZN(n14895) );
  AND2_X1 U18249 ( .A1(n14829), .A2(n14895), .ZN(n16112) );
  INV_X1 U18250 ( .A(n16112), .ZN(n14897) );
  AOI22_X1 U18251 ( .A1(n14898), .A2(n20311), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16115), .ZN(n14896) );
  OAI21_X1 U18252 ( .B1(n14897), .B2(n14904), .A(n14896), .ZN(P1_U2891) );
  AOI22_X1 U18253 ( .A1(n14898), .A2(n20309), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16115), .ZN(n14899) );
  OAI21_X1 U18254 ( .B1(n16094), .B2(n14904), .A(n14899), .ZN(P1_U2892) );
  INV_X1 U18255 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20282) );
  INV_X1 U18256 ( .A(n14900), .ZN(n14901) );
  OAI222_X1 U18257 ( .A1(n15044), .A2(n14904), .B1(n20282), .B2(n14903), .C1(
        n14902), .C2(n14901), .ZN(P1_U2893) );
  NOR2_X1 U18258 ( .A1(n14905), .A2(n13016), .ZN(n14906) );
  XNOR2_X1 U18259 ( .A(n14906), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15105) );
  INV_X1 U18260 ( .A(n14907), .ZN(n14911) );
  NOR2_X1 U18261 ( .A1(n20351), .A2(n21069), .ZN(n15097) );
  AOI21_X1 U18262 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15097), .ZN(n14908) );
  OAI21_X1 U18263 ( .B1(n20349), .B2(n14909), .A(n14908), .ZN(n14910) );
  OAI21_X1 U18264 ( .B1(n20167), .B2(n15105), .A(n14912), .ZN(P1_U2972) );
  INV_X1 U18265 ( .A(n14913), .ZN(n14918) );
  NAND3_X1 U18266 ( .A1(n12992), .A2(n14914), .A3(n20343), .ZN(n14917) );
  AOI21_X1 U18267 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14915), .ZN(n14916) );
  OAI211_X1 U18268 ( .C1(n20349), .C2(n14918), .A(n14917), .B(n14916), .ZN(
        n14919) );
  INV_X1 U18269 ( .A(n14919), .ZN(n14920) );
  OAI21_X1 U18270 ( .B1(n14921), .B2(n15054), .A(n14920), .ZN(P1_U2973) );
  AOI21_X1 U18271 ( .B1(n14922), .B2(n15046), .A(n16183), .ZN(n14935) );
  MUX2_X1 U18272 ( .A(n16183), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .S(
        n16146), .Z(n14923) );
  OAI211_X1 U18273 ( .C1(n14935), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        n14927) );
  XNOR2_X1 U18274 ( .A(n14927), .B(n14926), .ZN(n15114) );
  NOR2_X1 U18275 ( .A1(n20351), .A2(n20968), .ZN(n15108) );
  AOI21_X1 U18276 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15108), .ZN(n14928) );
  OAI21_X1 U18277 ( .B1(n20349), .B2(n14929), .A(n14928), .ZN(n14930) );
  AOI21_X1 U18278 ( .B1(n14931), .B2(n20344), .A(n14930), .ZN(n14932) );
  OAI21_X1 U18279 ( .B1(n20167), .B2(n15114), .A(n14932), .ZN(P1_U2974) );
  NOR2_X1 U18280 ( .A1(n14935), .A2(n12491), .ZN(n14934) );
  MUX2_X1 U18281 ( .A(n14935), .B(n14934), .S(n14933), .Z(n14936) );
  XNOR2_X1 U18282 ( .A(n14936), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15124) );
  INV_X1 U18283 ( .A(n14937), .ZN(n14939) );
  NOR2_X1 U18284 ( .A1(n20351), .A2(n21087), .ZN(n15118) );
  AOI21_X1 U18285 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15118), .ZN(n14938) );
  OAI21_X1 U18286 ( .B1(n20349), .B2(n14939), .A(n14938), .ZN(n14940) );
  AOI21_X1 U18287 ( .B1(n14941), .B2(n20344), .A(n14940), .ZN(n14942) );
  OAI21_X1 U18288 ( .B1(n20167), .B2(n15124), .A(n14942), .ZN(P1_U2975) );
  XNOR2_X1 U18289 ( .A(n15046), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14943) );
  XNOR2_X1 U18290 ( .A(n12491), .B(n14943), .ZN(n16177) );
  AOI22_X1 U18291 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14944) );
  OAI21_X1 U18292 ( .B1(n20349), .B2(n14945), .A(n14944), .ZN(n14946) );
  AOI21_X1 U18293 ( .B1(n14947), .B2(n20344), .A(n14946), .ZN(n14948) );
  OAI21_X1 U18294 ( .B1(n16177), .B2(n20167), .A(n14948), .ZN(P1_U2976) );
  NAND2_X1 U18295 ( .A1(n14949), .A2(n14950), .ZN(n14951) );
  XNOR2_X1 U18296 ( .A(n14951), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16192) );
  INV_X1 U18297 ( .A(n16192), .ZN(n14958) );
  INV_X1 U18298 ( .A(n14952), .ZN(n14954) );
  AOI22_X1 U18299 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n14953) );
  OAI21_X1 U18300 ( .B1(n20349), .B2(n14954), .A(n14953), .ZN(n14955) );
  AOI21_X1 U18301 ( .B1(n14956), .B2(n20344), .A(n14955), .ZN(n14957) );
  OAI21_X1 U18302 ( .B1(n20167), .B2(n14958), .A(n14957), .ZN(P1_U2977) );
  NOR2_X1 U18303 ( .A1(n15035), .A2(n15125), .ZN(n14960) );
  OR3_X1 U18304 ( .A1(n15046), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14969) );
  NOR3_X1 U18305 ( .A1(n14992), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n14969), .ZN(n14959) );
  AOI21_X1 U18306 ( .B1(n15154), .B2(n14960), .A(n14959), .ZN(n14961) );
  XNOR2_X1 U18307 ( .A(n14961), .B(n15127), .ZN(n15128) );
  INV_X1 U18308 ( .A(n14962), .ZN(n14966) );
  NOR2_X1 U18309 ( .A1(n20351), .A2(n20989), .ZN(n15130) );
  AOI21_X1 U18310 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15130), .ZN(n14963) );
  OAI21_X1 U18311 ( .B1(n20349), .B2(n14964), .A(n14963), .ZN(n14965) );
  AOI21_X1 U18312 ( .B1(n14966), .B2(n20344), .A(n14965), .ZN(n14967) );
  OAI21_X1 U18313 ( .B1(n15128), .B2(n20167), .A(n14967), .ZN(P1_U2978) );
  AND2_X1 U18314 ( .A1(n16146), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14968) );
  NAND2_X1 U18315 ( .A1(n15154), .A2(n14968), .ZN(n14973) );
  INV_X1 U18316 ( .A(n14992), .ZN(n14971) );
  INV_X1 U18317 ( .A(n14969), .ZN(n14970) );
  NAND2_X1 U18318 ( .A1(n14971), .A2(n14970), .ZN(n14972) );
  NAND2_X1 U18319 ( .A1(n14973), .A2(n14972), .ZN(n14974) );
  XNOR2_X1 U18320 ( .A(n14974), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15137) );
  INV_X1 U18321 ( .A(n14975), .ZN(n14976) );
  NAND2_X1 U18322 ( .A1(n14976), .A2(n20344), .ZN(n14981) );
  NOR2_X1 U18323 ( .A1(n20351), .A2(n21123), .ZN(n15141) );
  INV_X1 U18324 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14977) );
  NOR2_X1 U18325 ( .A1(n15039), .A2(n14977), .ZN(n14978) );
  AOI211_X1 U18326 ( .C1(n16152), .C2(n14979), .A(n15141), .B(n14978), .ZN(
        n14980) );
  OAI211_X1 U18327 ( .C1(n15137), .C2(n20167), .A(n14981), .B(n14980), .ZN(
        P1_U2979) );
  NOR2_X1 U18328 ( .A1(n16146), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14982) );
  MUX2_X1 U18329 ( .A(n14982), .B(n16146), .S(n15154), .Z(n14983) );
  XNOR2_X1 U18330 ( .A(n14983), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16200) );
  INV_X1 U18331 ( .A(n14984), .ZN(n14986) );
  AOI22_X1 U18332 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14985) );
  OAI21_X1 U18333 ( .B1(n20349), .B2(n14986), .A(n14985), .ZN(n14987) );
  AOI21_X1 U18334 ( .B1(n14988), .B2(n20344), .A(n14987), .ZN(n14989) );
  OAI21_X1 U18335 ( .B1(n20167), .B2(n16200), .A(n14989), .ZN(P1_U2980) );
  INV_X1 U18336 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14990) );
  NAND2_X1 U18337 ( .A1(n20377), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15152) );
  OAI21_X1 U18338 ( .B1(n15039), .B2(n14990), .A(n15152), .ZN(n14994) );
  NOR2_X1 U18339 ( .A1(n14992), .A2(n14991), .ZN(n15155) );
  NOR3_X1 U18340 ( .A1(n15155), .A2(n15154), .A3(n20167), .ZN(n14993) );
  AOI211_X1 U18341 ( .C1(n16152), .C2(n14995), .A(n14994), .B(n14993), .ZN(
        n14996) );
  OAI21_X1 U18342 ( .B1(n14997), .B2(n15054), .A(n14996), .ZN(P1_U2981) );
  NOR2_X1 U18343 ( .A1(n10157), .A2(n15018), .ZN(n16123) );
  NOR2_X1 U18344 ( .A1(n16123), .A2(n14999), .ZN(n16136) );
  OAI21_X1 U18345 ( .B1(n16136), .B2(n16125), .A(n16137), .ZN(n15000) );
  XOR2_X1 U18346 ( .A(n15001), .B(n15000), .Z(n16216) );
  INV_X1 U18347 ( .A(n15002), .ZN(n15004) );
  AOI22_X1 U18348 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15003) );
  OAI21_X1 U18349 ( .B1(n15004), .B2(n20349), .A(n15003), .ZN(n15005) );
  AOI21_X1 U18350 ( .B1(n15006), .B2(n20344), .A(n15005), .ZN(n15007) );
  OAI21_X1 U18351 ( .B1(n16216), .B2(n20167), .A(n15007), .ZN(P1_U2983) );
  MUX2_X1 U18352 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n12923), .S(
        n16146), .Z(n15011) );
  OAI21_X1 U18353 ( .B1(n16123), .B2(n15009), .A(n15008), .ZN(n15010) );
  XOR2_X1 U18354 ( .A(n15011), .B(n15010), .Z(n15165) );
  INV_X1 U18355 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15012) );
  NOR2_X1 U18356 ( .A1(n20351), .A2(n15012), .ZN(n15163) );
  AOI21_X1 U18357 ( .B1(n20338), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15163), .ZN(n15013) );
  OAI21_X1 U18358 ( .B1(n20349), .B2(n15014), .A(n15013), .ZN(n15015) );
  AOI21_X1 U18359 ( .B1(n16070), .B2(n20344), .A(n15015), .ZN(n15016) );
  OAI21_X1 U18360 ( .B1(n15165), .B2(n20167), .A(n15016), .ZN(P1_U2985) );
  NOR2_X1 U18361 ( .A1(n14998), .A2(n15017), .ZN(n15025) );
  OAI21_X1 U18362 ( .B1(n15025), .B2(n15018), .A(n9740), .ZN(n15020) );
  XNOR2_X1 U18363 ( .A(n15020), .B(n15019), .ZN(n16236) );
  AOI22_X1 U18364 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15021) );
  OAI21_X1 U18365 ( .B1(n20349), .B2(n15022), .A(n15021), .ZN(n15023) );
  AOI21_X1 U18366 ( .B1(n16112), .B2(n20344), .A(n15023), .ZN(n15024) );
  OAI21_X1 U18367 ( .B1(n16236), .B2(n20167), .A(n15024), .ZN(P1_U2986) );
  INV_X1 U18368 ( .A(n15025), .ZN(n15027) );
  NAND2_X1 U18369 ( .A1(n15027), .A2(n15026), .ZN(n15030) );
  NAND2_X1 U18370 ( .A1(n9740), .A2(n15028), .ZN(n15029) );
  XNOR2_X1 U18371 ( .A(n15030), .B(n15029), .ZN(n16251) );
  NAND2_X1 U18372 ( .A1(n16251), .A2(n20343), .ZN(n15034) );
  INV_X1 U18373 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15031) );
  NOR2_X1 U18374 ( .A1(n20351), .A2(n15031), .ZN(n16244) );
  NOR2_X1 U18375 ( .A1(n20349), .A2(n16092), .ZN(n15032) );
  AOI211_X1 U18376 ( .C1(n20338), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16244), .B(n15032), .ZN(n15033) );
  OAI211_X1 U18377 ( .C1(n15054), .C2(n16094), .A(n15034), .B(n15033), .ZN(
        P1_U2987) );
  NOR3_X1 U18378 ( .A1(n14998), .A2(n15035), .A3(n12908), .ZN(n16149) );
  NOR3_X1 U18379 ( .A1(n16145), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15046), .ZN(n15036) );
  NOR2_X1 U18380 ( .A1(n16149), .A2(n15036), .ZN(n15037) );
  XNOR2_X1 U18381 ( .A(n15037), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16260) );
  NAND2_X1 U18382 ( .A1(n16260), .A2(n20343), .ZN(n15043) );
  NAND2_X1 U18383 ( .A1(n20377), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n16256) );
  OAI21_X1 U18384 ( .B1(n15039), .B2(n15038), .A(n16256), .ZN(n15040) );
  AOI21_X1 U18385 ( .B1(n16152), .B2(n15041), .A(n15040), .ZN(n15042) );
  OAI211_X1 U18386 ( .C1(n15054), .C2(n15044), .A(n15043), .B(n15042), .ZN(
        P1_U2988) );
  XNOR2_X1 U18387 ( .A(n15046), .B(n16272), .ZN(n15047) );
  XNOR2_X1 U18388 ( .A(n15045), .B(n15047), .ZN(n16282) );
  NAND2_X1 U18389 ( .A1(n16282), .A2(n20343), .ZN(n15052) );
  INV_X1 U18390 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U18391 ( .A1(n20351), .A2(n15048), .ZN(n16279) );
  NOR2_X1 U18392 ( .A1(n20349), .A2(n15049), .ZN(n15050) );
  AOI211_X1 U18393 ( .C1(n20338), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16279), .B(n15050), .ZN(n15051) );
  OAI211_X1 U18394 ( .C1(n15054), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        P1_U2990) );
  INV_X1 U18395 ( .A(n15055), .ZN(n15120) );
  NAND2_X1 U18396 ( .A1(n15120), .A2(n16269), .ZN(n15056) );
  INV_X1 U18397 ( .A(n15056), .ZN(n15058) );
  NAND3_X1 U18398 ( .A1(n15110), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15057) );
  NAND2_X1 U18399 ( .A1(n15057), .A2(n15056), .ZN(n15093) );
  OAI21_X1 U18400 ( .B1(n15087), .B2(n15058), .A(n15093), .ZN(n15083) );
  AOI211_X1 U18401 ( .C1(n14247), .C2(n15175), .A(n14528), .B(n15083), .ZN(
        n15071) );
  INV_X1 U18402 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15198) );
  NOR3_X1 U18403 ( .A1(n15071), .A2(n15058), .A3(n15198), .ZN(n15066) );
  INV_X1 U18404 ( .A(n15060), .ZN(n15062) );
  NOR3_X1 U18405 ( .A1(n15116), .A2(n15062), .A3(n15061), .ZN(n15099) );
  NAND3_X1 U18406 ( .A1(n15099), .A2(n15087), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15072) );
  NOR3_X1 U18407 ( .A1(n15072), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14528), .ZN(n15063) );
  NOR4_X1 U18408 ( .A1(n15066), .A2(n15065), .A3(n15064), .A4(n15063), .ZN(
        n15067) );
  OAI21_X1 U18409 ( .B1(n15068), .B2(n16278), .A(n15067), .ZN(P1_U3000) );
  INV_X1 U18410 ( .A(n15069), .ZN(n15075) );
  INV_X1 U18411 ( .A(n15070), .ZN(n15074) );
  AOI21_X1 U18412 ( .B1(n14528), .B2(n15072), .A(n15071), .ZN(n15073) );
  AOI211_X1 U18413 ( .C1(n20372), .C2(n15075), .A(n15074), .B(n15073), .ZN(
        n15076) );
  OAI21_X1 U18414 ( .B1(n15077), .B2(n16278), .A(n15076), .ZN(P1_U3001) );
  INV_X1 U18415 ( .A(n15078), .ZN(n15080) );
  NAND3_X1 U18416 ( .A1(n15099), .A2(n15087), .A3(n14247), .ZN(n15079) );
  OAI211_X1 U18417 ( .C1(n15081), .C2(n20352), .A(n15080), .B(n15079), .ZN(
        n15082) );
  AOI21_X1 U18418 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15083), .A(
        n15082), .ZN(n15084) );
  OAI21_X1 U18419 ( .B1(n15085), .B2(n16278), .A(n15084), .ZN(P1_U3002) );
  INV_X1 U18420 ( .A(n15086), .ZN(n15092) );
  INV_X1 U18421 ( .A(n15099), .ZN(n15089) );
  NOR3_X1 U18422 ( .A1(n15089), .A2(n15088), .A3(n15087), .ZN(n15090) );
  AOI211_X1 U18423 ( .C1(n15092), .C2(n20372), .A(n15091), .B(n15090), .ZN(
        n15095) );
  INV_X1 U18424 ( .A(n15093), .ZN(n15103) );
  NAND2_X1 U18425 ( .A1(n15103), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15094) );
  OAI211_X1 U18426 ( .C1(n15096), .C2(n16278), .A(n15095), .B(n15094), .ZN(
        P1_U3003) );
  INV_X1 U18427 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15098) );
  AOI21_X1 U18428 ( .B1(n15099), .B2(n15098), .A(n15097), .ZN(n15100) );
  OAI21_X1 U18429 ( .B1(n15101), .B2(n20352), .A(n15100), .ZN(n15102) );
  AOI21_X1 U18430 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15103), .A(
        n15102), .ZN(n15104) );
  OAI21_X1 U18431 ( .B1(n15105), .B2(n16278), .A(n15104), .ZN(P1_U3004) );
  INV_X1 U18432 ( .A(n15106), .ZN(n15109) );
  AOI211_X1 U18433 ( .C1(n15109), .C2(n20372), .A(n15108), .B(n15107), .ZN(
        n15113) );
  INV_X1 U18434 ( .A(n15110), .ZN(n15111) );
  NAND2_X1 U18435 ( .A1(n15111), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15112) );
  OAI211_X1 U18436 ( .C1(n15114), .C2(n16278), .A(n15113), .B(n15112), .ZN(
        P1_U3006) );
  INV_X1 U18437 ( .A(n15115), .ZN(n15119) );
  NOR3_X1 U18438 ( .A1(n15116), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16183), .ZN(n15117) );
  AOI211_X1 U18439 ( .C1(n15119), .C2(n20372), .A(n15118), .B(n15117), .ZN(
        n15123) );
  OAI21_X1 U18440 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16250), .A(
        n15120), .ZN(n15121) );
  NAND2_X1 U18441 ( .A1(n15121), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15122) );
  OAI211_X1 U18442 ( .C1(n15124), .C2(n16278), .A(n15123), .B(n15122), .ZN(
        P1_U3007) );
  NOR3_X1 U18443 ( .A1(n16198), .A2(n16197), .A3(n15125), .ZN(n16187) );
  INV_X1 U18444 ( .A(n16187), .ZN(n15133) );
  INV_X1 U18445 ( .A(n15126), .ZN(n15131) );
  OAI22_X1 U18446 ( .A1(n15128), .A2(n16278), .B1(n15127), .B2(n16190), .ZN(
        n15129) );
  AOI211_X1 U18447 ( .C1(n15131), .C2(n20372), .A(n15130), .B(n15129), .ZN(
        n15132) );
  OAI21_X1 U18448 ( .B1(n15133), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15132), .ZN(P1_U3010) );
  AOI221_X1 U18449 ( .B1(n15183), .B2(n15138), .C1(n15134), .C2(n15138), .A(
        n16199), .ZN(n15136) );
  OAI22_X1 U18450 ( .A1(n15137), .A2(n16278), .B1(n15136), .B2(n15135), .ZN(
        n15143) );
  NOR4_X1 U18451 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16198), .A3(
        n15138), .A4(n16197), .ZN(n15142) );
  NOR2_X1 U18452 ( .A1(n15139), .A2(n20352), .ZN(n15140) );
  OR4_X1 U18453 ( .A1(n15143), .A2(n15142), .A3(n15141), .A4(n15140), .ZN(
        P1_U3011) );
  AOI21_X1 U18454 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15145), .A(
        n15144), .ZN(n15146) );
  INV_X1 U18455 ( .A(n16268), .ZN(n16247) );
  AOI211_X1 U18456 ( .C1(n15169), .C2(n15147), .A(n15146), .B(n16247), .ZN(
        n16242) );
  OAI21_X1 U18457 ( .B1(n16269), .B2(n15148), .A(n16242), .ZN(n16211) );
  INV_X1 U18458 ( .A(n15148), .ZN(n15149) );
  NOR2_X1 U18459 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15149), .ZN(
        n15150) );
  NAND2_X1 U18460 ( .A1(n15150), .A2(n16206), .ZN(n15151) );
  OAI211_X1 U18461 ( .C1(n15153), .C2(n20352), .A(n15152), .B(n15151), .ZN(
        n15157) );
  NOR3_X1 U18462 ( .A1(n15155), .A2(n15154), .A3(n16278), .ZN(n15156) );
  AOI211_X1 U18463 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n16211), .A(
        n15157), .B(n15156), .ZN(n15158) );
  INV_X1 U18464 ( .A(n15158), .ZN(P1_U3013) );
  NOR2_X1 U18465 ( .A1(n15159), .A2(n16301), .ZN(n16259) );
  NAND3_X1 U18466 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16259), .A3(
        n12923), .ZN(n15160) );
  OAI22_X1 U18467 ( .A1(n16242), .A2(n12923), .B1(n15161), .B2(n15160), .ZN(
        n15162) );
  AOI211_X1 U18468 ( .C1(n20372), .C2(n16065), .A(n15163), .B(n15162), .ZN(
        n15164) );
  OAI21_X1 U18469 ( .B1(n15165), .B2(n16278), .A(n15164), .ZN(P1_U3017) );
  NAND3_X1 U18470 ( .A1(n15167), .A2(n15166), .A3(n20375), .ZN(n15178) );
  INV_X1 U18471 ( .A(n15168), .ZN(n15174) );
  OAI21_X1 U18472 ( .B1(n15170), .B2(n15169), .A(n20368), .ZN(n15185) );
  AOI21_X1 U18473 ( .B1(n15171), .B2(n15185), .A(n20367), .ZN(n15172) );
  AOI211_X1 U18474 ( .C1(n20372), .C2(n15174), .A(n15173), .B(n15172), .ZN(
        n15177) );
  NAND3_X1 U18475 ( .A1(n15175), .A2(n20367), .A3(n20378), .ZN(n15176) );
  NAND3_X1 U18476 ( .A1(n15178), .A2(n15177), .A3(n15176), .ZN(P1_U3030) );
  NAND2_X1 U18477 ( .A1(n15179), .A2(n20375), .ZN(n15187) );
  AOI21_X1 U18478 ( .B1(n20372), .B2(n15181), .A(n15180), .ZN(n15186) );
  OAI21_X1 U18479 ( .B1(n15183), .B2(n15182), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15184) );
  NAND4_X1 U18480 ( .A1(n15187), .A2(n15186), .A3(n15185), .A4(n15184), .ZN(
        P1_U3031) );
  NAND2_X1 U18481 ( .A1(n15189), .A2(n15188), .ZN(n16019) );
  AOI22_X1 U18482 ( .A1(n15191), .A2(n20810), .B1(n11775), .B2(n15190), .ZN(
        n15192) );
  NAND2_X1 U18483 ( .A1(n16019), .A2(n15192), .ZN(n15193) );
  MUX2_X1 U18484 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15193), .S(
        n20385), .Z(P1_U3478) );
  NOR3_X1 U18485 ( .A1(n15194), .A2(n13656), .A3(n13659), .ZN(n15195) );
  AOI211_X1 U18486 ( .C1(n11751), .C2(n15197), .A(n15196), .B(n15195), .ZN(
        n15996) );
  INV_X1 U18487 ( .A(n20937), .ZN(n15209) );
  OAI22_X1 U18488 ( .A1(n15198), .A2(n20367), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15204) );
  NOR2_X1 U18489 ( .A1(n13651), .A2(n20368), .ZN(n15206) );
  NOR3_X1 U18490 ( .A1(n13656), .A2(n13659), .A3(n15199), .ZN(n15200) );
  AOI21_X1 U18491 ( .B1(n15204), .B2(n15206), .A(n15200), .ZN(n15201) );
  OAI21_X1 U18492 ( .B1(n15996), .B2(n15209), .A(n15201), .ZN(n15202) );
  MUX2_X1 U18493 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15202), .S(
        n16317), .Z(P1_U3473) );
  INV_X1 U18494 ( .A(n15204), .ZN(n15205) );
  AOI22_X1 U18495 ( .A1(n15207), .A2(n20936), .B1(n15206), .B2(n15205), .ZN(
        n15208) );
  OAI21_X1 U18496 ( .B1(n15210), .B2(n15209), .A(n15208), .ZN(n15211) );
  MUX2_X1 U18497 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15211), .S(
        n16317), .Z(P1_U3472) );
  INV_X1 U18498 ( .A(n20586), .ZN(n15212) );
  OAI21_X1 U18499 ( .B1(n15240), .B2(n20758), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15213) );
  NAND2_X1 U18500 ( .A1(n15213), .A2(n20677), .ZN(n15218) );
  NAND2_X1 U18501 ( .A1(n20800), .A2(n20619), .ZN(n15219) );
  INV_X1 U18502 ( .A(n15214), .ZN(n15215) );
  NAND2_X1 U18503 ( .A1(n15215), .A2(n20683), .ZN(n20620) );
  INV_X1 U18504 ( .A(n20560), .ZN(n20766) );
  OAI22_X1 U18505 ( .A1(n15218), .A2(n15219), .B1(n20620), .B2(n20766), .ZN(
        n20759) );
  INV_X1 U18506 ( .A(n20803), .ZN(n20697) );
  INV_X1 U18507 ( .A(n20694), .ZN(n20815) );
  NOR2_X1 U18508 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15216), .ZN(
        n20757) );
  INV_X1 U18509 ( .A(n15218), .ZN(n15220) );
  AOI22_X1 U18510 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20620), .B1(n15220), 
        .B2(n15219), .ZN(n15221) );
  AOI22_X1 U18511 ( .A1(n20804), .A2(n20757), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n20760), .ZN(n15222) );
  OAI21_X1 U18512 ( .B1(n15238), .B2(n20815), .A(n15222), .ZN(n15223) );
  AOI21_X1 U18513 ( .B1(n15240), .B2(n20812), .A(n15223), .ZN(n15224) );
  OAI21_X1 U18514 ( .B1(n15242), .B2(n20697), .A(n15224), .ZN(P1_U3129) );
  INV_X1 U18515 ( .A(n20816), .ZN(n20700) );
  INV_X1 U18516 ( .A(n20818), .ZN(n20777) );
  AOI22_X1 U18517 ( .A1(n20817), .A2(n20757), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n20760), .ZN(n15225) );
  OAI21_X1 U18518 ( .B1(n15238), .B2(n20777), .A(n15225), .ZN(n15226) );
  AOI21_X1 U18519 ( .B1(n15240), .B2(n20774), .A(n15226), .ZN(n15227) );
  OAI21_X1 U18520 ( .B1(n15242), .B2(n20700), .A(n15227), .ZN(P1_U3130) );
  INV_X1 U18521 ( .A(n20828), .ZN(n20707) );
  INV_X1 U18522 ( .A(n20704), .ZN(n20833) );
  AOI22_X1 U18523 ( .A1(n20829), .A2(n20757), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n20760), .ZN(n15228) );
  OAI21_X1 U18524 ( .B1(n15238), .B2(n20833), .A(n15228), .ZN(n15229) );
  AOI21_X1 U18525 ( .B1(n9792), .B2(n15240), .A(n15229), .ZN(n15230) );
  OAI21_X1 U18526 ( .B1(n15242), .B2(n20707), .A(n15230), .ZN(P1_U3132) );
  INV_X1 U18527 ( .A(n20834), .ZN(n20711) );
  INV_X1 U18528 ( .A(n20708), .ZN(n20839) );
  AOI22_X1 U18529 ( .A1(n20835), .A2(n20757), .B1(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n20760), .ZN(n15231) );
  OAI21_X1 U18530 ( .B1(n15238), .B2(n20839), .A(n15231), .ZN(n15232) );
  AOI21_X1 U18531 ( .B1(n9794), .B2(n15240), .A(n15232), .ZN(n15233) );
  OAI21_X1 U18532 ( .B1(n15242), .B2(n20711), .A(n15233), .ZN(P1_U3133) );
  INV_X1 U18533 ( .A(n20849), .ZN(n20718) );
  INV_X1 U18534 ( .A(n20715), .ZN(n20853) );
  AOI22_X1 U18535 ( .A1(n20848), .A2(n20757), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n20760), .ZN(n15234) );
  OAI21_X1 U18536 ( .B1(n15238), .B2(n20853), .A(n15234), .ZN(n15235) );
  AOI21_X1 U18537 ( .B1(n15240), .B2(n9790), .A(n15235), .ZN(n15236) );
  OAI21_X1 U18538 ( .B1(n15242), .B2(n20718), .A(n15236), .ZN(P1_U3135) );
  INV_X1 U18539 ( .A(n20855), .ZN(n20725) );
  INV_X1 U18540 ( .A(n20721), .ZN(n20864) );
  AOI22_X1 U18541 ( .A1(n20857), .A2(n20757), .B1(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n20760), .ZN(n15237) );
  OAI21_X1 U18542 ( .B1(n15238), .B2(n20864), .A(n15237), .ZN(n15239) );
  AOI21_X1 U18543 ( .B1(n20858), .B2(n15240), .A(n15239), .ZN(n15241) );
  OAI21_X1 U18544 ( .B1(n15242), .B2(n20725), .A(n15241), .ZN(P1_U3136) );
  INV_X1 U18545 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15550) );
  XNOR2_X1 U18546 ( .A(n13071), .B(n15550), .ZN(n15552) );
  OAI21_X1 U18547 ( .B1(n15246), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15244), .ZN(n15560) );
  INV_X1 U18548 ( .A(n15560), .ZN(n16341) );
  NOR2_X1 U18549 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n15247), .ZN(
        n15245) );
  NOR2_X1 U18550 ( .A1(n15246), .A2(n15245), .ZN(n15566) );
  OAI21_X1 U18551 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n15250), .A(
        n15248), .ZN(n15249) );
  INV_X1 U18552 ( .A(n15249), .ZN(n15579) );
  AOI21_X1 U18553 ( .B1(n16349), .B2(n15251), .A(n15250), .ZN(n16357) );
  OAI21_X1 U18554 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15254), .A(
        n15251), .ZN(n15601) );
  INV_X1 U18555 ( .A(n15601), .ZN(n15320) );
  NOR2_X1 U18556 ( .A1(n15252), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15253) );
  NOR2_X1 U18557 ( .A1(n15254), .A2(n15253), .ZN(n15608) );
  INV_X1 U18558 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15255) );
  AOI21_X1 U18559 ( .B1(n15263), .B2(n15255), .A(n15265), .ZN(n19136) );
  AOI21_X1 U18560 ( .B1(n15642), .B2(n15262), .A(n15264), .ZN(n19154) );
  AOI21_X1 U18561 ( .B1(n15260), .B2(n15661), .A(n9739), .ZN(n19176) );
  AOI21_X1 U18562 ( .B1(n16381), .B2(n15258), .A(n15261), .ZN(n16370) );
  AOI21_X1 U18563 ( .B1(n16399), .B2(n15256), .A(n15259), .ZN(n19215) );
  OAI21_X1 U18564 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15257), .A(
        n15256), .ZN(n19228) );
  NAND2_X1 U18565 ( .A1(n19227), .A2(n19228), .ZN(n19213) );
  NOR2_X1 U18566 ( .A1(n19215), .A2(n19213), .ZN(n19206) );
  OAI21_X1 U18567 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15259), .A(
        n15258), .ZN(n19207) );
  NAND2_X1 U18568 ( .A1(n19206), .A2(n19207), .ZN(n15347) );
  NOR2_X1 U18569 ( .A1(n16370), .A2(n15347), .ZN(n19195) );
  OAI21_X1 U18570 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15261), .A(
        n15260), .ZN(n19196) );
  NAND2_X1 U18571 ( .A1(n19195), .A2(n19196), .ZN(n19177) );
  OAI21_X1 U18572 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9739), .A(
        n15262), .ZN(n19168) );
  NAND2_X1 U18573 ( .A1(n19175), .A2(n19168), .ZN(n19152) );
  NOR2_X1 U18574 ( .A1(n19154), .A2(n19152), .ZN(n19139) );
  OAI21_X1 U18575 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15264), .A(
        n15263), .ZN(n19143) );
  NAND2_X1 U18576 ( .A1(n19139), .A2(n19143), .ZN(n19125) );
  INV_X1 U18577 ( .A(n15252), .ZN(n15269) );
  INV_X1 U18578 ( .A(n15265), .ZN(n15267) );
  INV_X1 U18579 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15266) );
  NAND2_X1 U18580 ( .A1(n15267), .A2(n15266), .ZN(n15268) );
  NAND2_X1 U18581 ( .A1(n15269), .A2(n15268), .ZN(n15976) );
  NOR2_X1 U18582 ( .A1(n15320), .A2(n15319), .ZN(n15318) );
  NOR2_X1 U18583 ( .A1(n19288), .A2(n15318), .ZN(n16356) );
  NOR2_X1 U18584 ( .A1(n16357), .A2(n16356), .ZN(n16355) );
  NOR2_X1 U18585 ( .A1(n19288), .A2(n16355), .ZN(n15304) );
  NOR2_X1 U18586 ( .A1(n19288), .A2(n15303), .ZN(n15298) );
  NOR2_X1 U18587 ( .A1(n15566), .A2(n15298), .ZN(n15297) );
  NOR2_X1 U18588 ( .A1(n19288), .A2(n15297), .ZN(n16340) );
  INV_X1 U18589 ( .A(n19329), .ZN(n19123) );
  NAND2_X1 U18590 ( .A1(n15382), .A2(n19285), .ZN(n15275) );
  AOI22_X1 U18591 ( .A1(n19311), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19323), .ZN(n15270) );
  OAI21_X1 U18592 ( .B1(n15271), .B2(n19262), .A(n15270), .ZN(n15272) );
  AOI21_X1 U18593 ( .B1(n15278), .B2(n19123), .A(n15276), .ZN(n15277) );
  INV_X1 U18594 ( .A(n15277), .ZN(P2_U2824) );
  INV_X1 U18595 ( .A(n15278), .ZN(n15281) );
  NAND2_X1 U18596 ( .A1(n15281), .A2(n15280), .ZN(n15288) );
  NAND2_X1 U18597 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19323), .ZN(
        n15283) );
  NAND2_X1 U18598 ( .A1(n19311), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15282) );
  OAI211_X1 U18599 ( .C1(n19262), .C2(n20087), .A(n15283), .B(n15282), .ZN(
        n15285) );
  NOR2_X1 U18600 ( .A1(n15692), .A2(n19315), .ZN(n15284) );
  AOI211_X1 U18601 ( .C1(n19317), .C2(n15286), .A(n15285), .B(n15284), .ZN(
        n15287) );
  OAI211_X1 U18602 ( .C1(n15699), .C2(n19320), .A(n15288), .B(n15287), .ZN(
        P2_U2825) );
  OR2_X1 U18603 ( .A1(n15311), .A2(n15289), .ZN(n15290) );
  AND2_X1 U18604 ( .A1(n15291), .A2(n15290), .ZN(n15712) );
  INV_X1 U18605 ( .A(n15712), .ZN(n15302) );
  NOR2_X1 U18606 ( .A1(n15306), .A2(n15292), .ZN(n15293) );
  OR2_X1 U18607 ( .A1(n12858), .A2(n15293), .ZN(n15706) );
  INV_X1 U18608 ( .A(n19262), .ZN(n19312) );
  AOI22_X1 U18609 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19311), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19312), .ZN(n15296) );
  AOI22_X1 U18610 ( .A1(n15294), .A2(n19317), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19323), .ZN(n15295) );
  OAI211_X1 U18611 ( .C1(n15706), .C2(n19315), .A(n15296), .B(n15295), .ZN(
        n15300) );
  AOI211_X1 U18612 ( .C1(n15566), .C2(n15298), .A(n15297), .B(n19289), .ZN(
        n15299) );
  NOR2_X1 U18613 ( .A1(n15300), .A2(n15299), .ZN(n15301) );
  OAI21_X1 U18614 ( .B1(n15302), .B2(n19320), .A(n15301), .ZN(P2_U2828) );
  AOI211_X1 U18615 ( .C1(n15579), .C2(n15304), .A(n15303), .B(n19289), .ZN(
        n15305) );
  INV_X1 U18616 ( .A(n15305), .ZN(n15316) );
  AOI21_X1 U18617 ( .B1(n15307), .B2(n15482), .A(n15306), .ZN(n15723) );
  INV_X1 U18618 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15309) );
  AOI22_X1 U18619 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19311), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19312), .ZN(n15308) );
  OAI21_X1 U18620 ( .B1(n15309), .B2(n19297), .A(n15308), .ZN(n15314) );
  AND2_X1 U18621 ( .A1(n15412), .A2(n15310), .ZN(n15312) );
  OR2_X1 U18622 ( .A1(n15312), .A2(n15311), .ZN(n15718) );
  NOR2_X1 U18623 ( .A1(n15718), .A2(n19320), .ZN(n15313) );
  AOI211_X1 U18624 ( .C1(n19305), .C2(n15723), .A(n15314), .B(n15313), .ZN(
        n15315) );
  OAI211_X1 U18625 ( .C1(n19302), .C2(n15317), .A(n15316), .B(n15315), .ZN(
        P2_U2829) );
  AOI211_X1 U18626 ( .C1(n15320), .C2(n15319), .A(n15318), .B(n19289), .ZN(
        n15321) );
  INV_X1 U18627 ( .A(n15321), .ZN(n15330) );
  AOI21_X1 U18628 ( .B1(n15322), .B2(n9696), .A(n10013), .ZN(n15751) );
  NAND2_X1 U18629 ( .A1(n15323), .A2(n15324), .ZN(n15325) );
  NAND2_X1 U18630 ( .A1(n15483), .A2(n15325), .ZN(n15749) );
  AOI22_X1 U18631 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19311), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19312), .ZN(n15327) );
  NAND2_X1 U18632 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19323), .ZN(
        n15326) );
  OAI211_X1 U18633 ( .C1(n15749), .C2(n19315), .A(n15327), .B(n15326), .ZN(
        n15328) );
  AOI21_X1 U18634 ( .B1(n15751), .B2(n19285), .A(n15328), .ZN(n15329) );
  OAI211_X1 U18635 ( .C1(n19302), .C2(n15331), .A(n15330), .B(n15329), .ZN(
        P2_U2831) );
  AOI211_X1 U18636 ( .C1(n15608), .C2(n15333), .A(n15332), .B(n19289), .ZN(
        n15334) );
  INV_X1 U18637 ( .A(n15334), .ZN(n15345) );
  OR2_X1 U18638 ( .A1(n15336), .A2(n15335), .ZN(n15337) );
  AND2_X1 U18639 ( .A1(n15323), .A2(n15337), .ZN(n15760) );
  NAND2_X1 U18640 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19323), .ZN(
        n15339) );
  NAND2_X1 U18641 ( .A1(n19311), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15338) );
  OAI211_X1 U18642 ( .C1(n19262), .C2(n20074), .A(n15339), .B(n15338), .ZN(
        n15343) );
  OR2_X1 U18643 ( .A1(n15429), .A2(n15340), .ZN(n15341) );
  NAND2_X1 U18644 ( .A1(n9696), .A2(n15341), .ZN(n15763) );
  NOR2_X1 U18645 ( .A1(n15763), .A2(n19320), .ZN(n15342) );
  AOI211_X1 U18646 ( .C1(n19305), .C2(n15760), .A(n15343), .B(n15342), .ZN(
        n15344) );
  OAI211_X1 U18647 ( .C1(n19302), .C2(n15346), .A(n15345), .B(n15344), .ZN(
        P2_U2832) );
  AOI211_X1 U18648 ( .C1(n16370), .C2(n15347), .A(n19195), .B(n19329), .ZN(
        n15358) );
  NOR2_X1 U18649 ( .A1(n15348), .A2(n15349), .ZN(n15350) );
  OR2_X1 U18650 ( .A1(n13987), .A2(n15350), .ZN(n19337) );
  NOR2_X1 U18651 ( .A1(n19315), .A2(n19337), .ZN(n15353) );
  AOI22_X1 U18652 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19323), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n19311), .ZN(n15351) );
  OAI211_X1 U18653 ( .C1(n19262), .C2(n11140), .A(n15351), .B(n19178), .ZN(
        n15352) );
  AOI211_X1 U18654 ( .C1(n16370), .C2(n19322), .A(n15353), .B(n15352), .ZN(
        n15355) );
  NAND2_X1 U18655 ( .A1(n16461), .A2(n19285), .ZN(n15354) );
  OAI211_X1 U18656 ( .C1(n15356), .C2(n19302), .A(n15355), .B(n15354), .ZN(
        n15357) );
  OR2_X1 U18657 ( .A1(n15358), .A2(n15357), .ZN(P2_U2840) );
  NAND2_X1 U18658 ( .A1(n19257), .A2(n15359), .ZN(n15360) );
  XNOR2_X1 U18659 ( .A(n16424), .B(n15360), .ZN(n15361) );
  NAND2_X1 U18660 ( .A1(n15361), .A2(n19306), .ZN(n15367) );
  AOI22_X1 U18661 ( .A1(n15362), .A2(n19317), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19323), .ZN(n15363) );
  OAI211_X1 U18662 ( .C1(n10108), .C2(n19180), .A(n15363), .B(n19178), .ZN(
        n15364) );
  AOI21_X1 U18663 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n19312), .A(n15364), .ZN(
        n15366) );
  AOI22_X1 U18664 ( .A1(n16425), .A2(n19285), .B1(n19305), .B2(n15895), .ZN(
        n15365) );
  NAND3_X1 U18665 ( .A1(n15367), .A2(n15366), .A3(n15365), .ZN(P2_U2846) );
  NAND2_X1 U18666 ( .A1(n19317), .A2(n15368), .ZN(n15370) );
  AOI22_X1 U18667 ( .A1(n19311), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19323), .ZN(n15369) );
  OAI211_X1 U18668 ( .C1(n19262), .C2(n15371), .A(n15370), .B(n15369), .ZN(
        n15372) );
  AOI21_X1 U18669 ( .B1(n20110), .B2(n19305), .A(n15372), .ZN(n15373) );
  OAI21_X1 U18670 ( .B1(n15374), .B2(n19320), .A(n15373), .ZN(n15380) );
  INV_X1 U18671 ( .A(n15376), .ZN(n15378) );
  NOR2_X1 U18672 ( .A1(n19288), .A2(n15907), .ZN(n15377) );
  INV_X1 U18673 ( .A(n15377), .ZN(n15375) );
  AOI221_X1 U18674 ( .B1(n15378), .B2(n15377), .C1(n15376), .C2(n15375), .A(
        n19289), .ZN(n15379) );
  AOI211_X1 U18675 ( .C1(n19327), .C2(n20111), .A(n15380), .B(n15379), .ZN(
        n15381) );
  INV_X1 U18676 ( .A(n15381), .ZN(P2_U2853) );
  NAND2_X1 U18677 ( .A1(n15382), .A2(n15442), .ZN(n15383) );
  OAI21_X1 U18678 ( .B1(n15440), .B2(n15384), .A(n15383), .ZN(P2_U2856) );
  INV_X1 U18679 ( .A(n15385), .ZN(n16332) );
  NAND3_X1 U18680 ( .A1(n15451), .A2(n15387), .A3(n15434), .ZN(n15389) );
  NAND2_X1 U18681 ( .A1(n13273), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15388) );
  OAI211_X1 U18682 ( .C1(n16332), .C2(n13273), .A(n15389), .B(n15388), .ZN(
        P2_U2858) );
  NOR2_X1 U18683 ( .A1(n15391), .A2(n15390), .ZN(n15393) );
  XNOR2_X1 U18684 ( .A(n15393), .B(n15392), .ZN(n15467) );
  NAND2_X1 U18685 ( .A1(n13273), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15395) );
  NAND2_X1 U18686 ( .A1(n16338), .A2(n15442), .ZN(n15394) );
  OAI211_X1 U18687 ( .C1(n15467), .C2(n15450), .A(n15395), .B(n15394), .ZN(
        P2_U2859) );
  OAI21_X1 U18688 ( .B1(n15396), .B2(n15398), .A(n15397), .ZN(n15474) );
  NAND2_X1 U18689 ( .A1(n13273), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15400) );
  NAND2_X1 U18690 ( .A1(n15712), .A2(n15440), .ZN(n15399) );
  OAI211_X1 U18691 ( .C1(n15474), .C2(n15450), .A(n15400), .B(n15399), .ZN(
        P2_U2860) );
  AOI21_X1 U18692 ( .B1(n15401), .B2(n15403), .A(n15402), .ZN(n15475) );
  NAND2_X1 U18693 ( .A1(n15475), .A2(n15434), .ZN(n15405) );
  NAND2_X1 U18694 ( .A1(n13273), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15404) );
  OAI211_X1 U18695 ( .C1(n15718), .C2(n13322), .A(n15405), .B(n15404), .ZN(
        P2_U2861) );
  OAI21_X1 U18696 ( .B1(n15406), .B2(n15408), .A(n15407), .ZN(n15490) );
  NAND2_X1 U18697 ( .A1(n15410), .A2(n15409), .ZN(n15411) );
  NAND2_X1 U18698 ( .A1(n15412), .A2(n15411), .ZN(n16352) );
  NOR2_X1 U18699 ( .A1(n16352), .A2(n13322), .ZN(n15413) );
  AOI21_X1 U18700 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n13273), .A(n15413), .ZN(
        n15414) );
  OAI21_X1 U18701 ( .B1(n15490), .B2(n15450), .A(n15414), .ZN(P2_U2862) );
  AOI21_X1 U18702 ( .B1(n9749), .B2(n15416), .A(n15415), .ZN(n15417) );
  XOR2_X1 U18703 ( .A(n15418), .B(n15417), .Z(n15497) );
  NAND2_X1 U18704 ( .A1(n13273), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15420) );
  NAND2_X1 U18705 ( .A1(n15751), .A2(n15442), .ZN(n15419) );
  OAI211_X1 U18706 ( .C1(n15497), .C2(n15450), .A(n15420), .B(n15419), .ZN(
        P2_U2863) );
  AOI21_X1 U18707 ( .B1(n15423), .B2(n15422), .A(n15421), .ZN(n15498) );
  NAND2_X1 U18708 ( .A1(n15498), .A2(n15434), .ZN(n15425) );
  NAND2_X1 U18709 ( .A1(n13273), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15424) );
  OAI211_X1 U18710 ( .C1(n15763), .C2(n13322), .A(n15425), .B(n15424), .ZN(
        P2_U2864) );
  NOR2_X1 U18711 ( .A1(n15427), .A2(n15426), .ZN(n15428) );
  OR2_X1 U18712 ( .A1(n15429), .A2(n15428), .ZN(n15983) );
  INV_X1 U18713 ( .A(n15430), .ZN(n15433) );
  INV_X1 U18714 ( .A(n15431), .ZN(n15438) );
  AOI21_X1 U18715 ( .B1(n15433), .B2(n15438), .A(n15432), .ZN(n16366) );
  NAND2_X1 U18716 ( .A1(n16366), .A2(n15434), .ZN(n15436) );
  NAND2_X1 U18717 ( .A1(n13273), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15435) );
  OAI211_X1 U18718 ( .C1(n15983), .C2(n13322), .A(n15436), .B(n15435), .ZN(
        P2_U2865) );
  OAI21_X1 U18719 ( .B1(n15444), .B2(n15439), .A(n15438), .ZN(n15508) );
  NOR2_X1 U18720 ( .A1(n15440), .A2(n10783), .ZN(n15441) );
  AOI21_X1 U18721 ( .B1(n19128), .B2(n15442), .A(n15441), .ZN(n15443) );
  OAI21_X1 U18722 ( .B1(n15508), .B2(n15450), .A(n15443), .ZN(P2_U2866) );
  OAI21_X1 U18723 ( .B1(n14205), .B2(n15445), .A(n15437), .ZN(n15516) );
  NAND2_X1 U18724 ( .A1(n14188), .A2(n15446), .ZN(n15447) );
  AND2_X1 U18725 ( .A1(n15448), .A2(n15447), .ZN(n19148) );
  INV_X1 U18726 ( .A(n19148), .ZN(n15785) );
  MUX2_X1 U18727 ( .A(n15785), .B(n10781), .S(n13273), .Z(n15449) );
  OAI21_X1 U18728 ( .B1(n15516), .B2(n15450), .A(n15449), .ZN(P2_U2867) );
  NAND3_X1 U18729 ( .A1(n15451), .A2(n15387), .A3(n19381), .ZN(n15457) );
  INV_X1 U18730 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n15454) );
  AOI22_X1 U18731 ( .A1(n16364), .A2(n15452), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19379), .ZN(n15453) );
  OAI21_X1 U18732 ( .B1(n15524), .B2(n15454), .A(n15453), .ZN(n15455) );
  AOI21_X1 U18733 ( .B1(n19331), .B2(BUF1_REG_29__SCAN_IN), .A(n15455), .ZN(
        n15456) );
  OAI211_X1 U18734 ( .C1(n15458), .C2(n15538), .A(n15457), .B(n15456), .ZN(
        P2_U2890) );
  NAND2_X1 U18735 ( .A1(n19379), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n15459) );
  OAI21_X1 U18736 ( .B1(n15522), .B2(n15460), .A(n15459), .ZN(n15461) );
  AOI21_X1 U18737 ( .B1(n19333), .B2(BUF2_REG_28__SCAN_IN), .A(n15461), .ZN(
        n15463) );
  NAND2_X1 U18738 ( .A1(n19331), .A2(BUF1_REG_28__SCAN_IN), .ZN(n15462) );
  OAI211_X1 U18739 ( .C1(n15464), .C2(n15538), .A(n15463), .B(n15462), .ZN(
        n15465) );
  INV_X1 U18740 ( .A(n15465), .ZN(n15466) );
  OAI21_X1 U18741 ( .B1(n15467), .B2(n19356), .A(n15466), .ZN(P2_U2891) );
  NAND2_X1 U18742 ( .A1(n19379), .A2(P2_EAX_REG_27__SCAN_IN), .ZN(n15468) );
  OAI21_X1 U18743 ( .B1(n15522), .B2(n19347), .A(n15468), .ZN(n15469) );
  AOI21_X1 U18744 ( .B1(n19333), .B2(BUF2_REG_27__SCAN_IN), .A(n15469), .ZN(
        n15471) );
  NAND2_X1 U18745 ( .A1(n19331), .A2(BUF1_REG_27__SCAN_IN), .ZN(n15470) );
  OAI211_X1 U18746 ( .C1(n15706), .C2(n15538), .A(n15471), .B(n15470), .ZN(
        n15472) );
  INV_X1 U18747 ( .A(n15472), .ZN(n15473) );
  OAI21_X1 U18748 ( .B1(n15474), .B2(n19356), .A(n15473), .ZN(P2_U2892) );
  INV_X1 U18749 ( .A(n15475), .ZN(n15481) );
  OAI22_X1 U18750 ( .A1(n15477), .A2(n15522), .B1(n19349), .B2(n15476), .ZN(
        n15478) );
  AOI21_X1 U18751 ( .B1(n15723), .B2(n19380), .A(n15478), .ZN(n15480) );
  AOI22_X1 U18752 ( .A1(n19331), .A2(BUF1_REG_26__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15479) );
  OAI211_X1 U18753 ( .C1(n15481), .C2(n19356), .A(n15480), .B(n15479), .ZN(
        P2_U2893) );
  AOI21_X1 U18754 ( .B1(n15484), .B2(n15483), .A(n10103), .ZN(n16353) );
  INV_X1 U18755 ( .A(n16353), .ZN(n15485) );
  OAI22_X1 U18756 ( .A1(n15485), .A2(n15538), .B1(n19349), .B2(n13226), .ZN(
        n15486) );
  AOI21_X1 U18757 ( .B1(n16364), .B2(n15487), .A(n15486), .ZN(n15489) );
  AOI22_X1 U18758 ( .A1(n19331), .A2(BUF1_REG_25__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15488) );
  OAI211_X1 U18759 ( .C1(n15490), .C2(n19356), .A(n15489), .B(n15488), .ZN(
        P2_U2894) );
  INV_X1 U18760 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n15491) );
  OAI22_X1 U18761 ( .A1(n15525), .A2(n16618), .B1(n15524), .B2(n15491), .ZN(
        n15494) );
  OAI22_X1 U18762 ( .A1(n15749), .A2(n15538), .B1(n19349), .B2(n15492), .ZN(
        n15493) );
  AOI211_X1 U18763 ( .C1(n16364), .C2(n15495), .A(n15494), .B(n15493), .ZN(
        n15496) );
  OAI21_X1 U18764 ( .B1(n15497), .B2(n19356), .A(n15496), .ZN(P2_U2895) );
  NAND2_X1 U18765 ( .A1(n15498), .A2(n19381), .ZN(n15503) );
  AOI22_X1 U18766 ( .A1(n16364), .A2(n15499), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n19379), .ZN(n15502) );
  AOI22_X1 U18767 ( .A1(n19331), .A2(BUF1_REG_23__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15501) );
  NAND2_X1 U18768 ( .A1(n15760), .A2(n19380), .ZN(n15500) );
  NAND4_X1 U18769 ( .A1(n15503), .A2(n15502), .A3(n15501), .A4(n15500), .ZN(
        P2_U2896) );
  OAI22_X1 U18770 ( .A1(n19486), .A2(n15522), .B1(n19349), .B2(n15504), .ZN(
        n15505) );
  AOI21_X1 U18771 ( .B1(n19133), .B2(n19380), .A(n15505), .ZN(n15507) );
  AOI22_X1 U18772 ( .A1(n19331), .A2(BUF1_REG_21__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15506) );
  OAI211_X1 U18773 ( .C1(n15508), .C2(n19356), .A(n15507), .B(n15506), .ZN(
        P2_U2898) );
  OR2_X1 U18774 ( .A1(n15520), .A2(n15509), .ZN(n15510) );
  NAND2_X1 U18775 ( .A1(n11243), .A2(n15510), .ZN(n19151) );
  INV_X1 U18776 ( .A(n19151), .ZN(n15513) );
  OAI22_X1 U18777 ( .A1(n19480), .A2(n15522), .B1(n19349), .B2(n15511), .ZN(
        n15512) );
  AOI21_X1 U18778 ( .B1(n19380), .B2(n15513), .A(n15512), .ZN(n15515) );
  AOI22_X1 U18779 ( .A1(n19331), .A2(BUF1_REG_20__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15514) );
  OAI211_X1 U18780 ( .C1(n15516), .C2(n19356), .A(n15515), .B(n15514), .ZN(
        P2_U2899) );
  INV_X1 U18781 ( .A(n15517), .ZN(n15530) );
  NOR2_X1 U18782 ( .A1(n15534), .A2(n15518), .ZN(n15519) );
  OR2_X1 U18783 ( .A1(n15520), .A2(n15519), .ZN(n19158) );
  INV_X1 U18784 ( .A(n19158), .ZN(n15528) );
  OAI22_X1 U18785 ( .A1(n19475), .A2(n15522), .B1(n19349), .B2(n15521), .ZN(
        n15527) );
  INV_X1 U18786 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15523) );
  OAI22_X1 U18787 ( .A1(n15525), .A2(n16627), .B1(n15524), .B2(n15523), .ZN(
        n15526) );
  AOI211_X1 U18788 ( .C1(n19380), .C2(n15528), .A(n15527), .B(n15526), .ZN(
        n15529) );
  OAI21_X1 U18789 ( .B1(n15530), .B2(n19356), .A(n15529), .ZN(P2_U2900) );
  AND2_X1 U18790 ( .A1(n15532), .A2(n15531), .ZN(n15533) );
  OR2_X1 U18791 ( .A1(n15534), .A2(n15533), .ZN(n19174) );
  AOI22_X1 U18792 ( .A1(n19331), .A2(BUF1_REG_18__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n15537) );
  INV_X1 U18793 ( .A(n19471), .ZN(n15535) );
  AOI22_X1 U18794 ( .A1(n16364), .A2(n15535), .B1(n19379), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15536) );
  OAI211_X1 U18795 ( .C1(n15538), .C2(n19174), .A(n15537), .B(n15536), .ZN(
        n15539) );
  AOI21_X1 U18796 ( .B1(n15540), .B2(n19381), .A(n15539), .ZN(n15541) );
  INV_X1 U18797 ( .A(n15541), .ZN(P2_U2901) );
  NAND2_X1 U18798 ( .A1(n15544), .A2(n15543), .ZN(n15549) );
  INV_X1 U18799 ( .A(n15545), .ZN(n15547) );
  NAND2_X1 U18800 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  NAND2_X1 U18801 ( .A1(n19420), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15695) );
  OAI21_X1 U18802 ( .B1(n16453), .B2(n15550), .A(n15695), .ZN(n15551) );
  AOI21_X1 U18803 ( .B1(n16440), .B2(n15552), .A(n15551), .ZN(n15553) );
  OAI21_X1 U18804 ( .B1(n15699), .B2(n15688), .A(n15553), .ZN(n15554) );
  AOI21_X1 U18805 ( .B1(n15701), .B2(n16450), .A(n15554), .ZN(n15555) );
  OAI21_X1 U18806 ( .B1(n19423), .B2(n15703), .A(n15555), .ZN(P2_U2984) );
  INV_X1 U18807 ( .A(n15556), .ZN(n15562) );
  NAND2_X1 U18808 ( .A1(n16338), .A2(n19428), .ZN(n15559) );
  AOI21_X1 U18809 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15557), .ZN(n15558) );
  OAI211_X1 U18810 ( .C1(n19432), .C2(n15560), .A(n15559), .B(n15558), .ZN(
        n15561) );
  OAI21_X1 U18811 ( .B1(n15564), .B2(n19424), .A(n15563), .ZN(P2_U2986) );
  OAI21_X1 U18812 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n9694), .A(
        n9933), .ZN(n15717) );
  NOR2_X1 U18813 ( .A1(n16466), .A2(n20082), .ZN(n15704) );
  AOI21_X1 U18814 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15704), .ZN(n15568) );
  NAND2_X1 U18815 ( .A1(n16440), .A2(n15566), .ZN(n15567) );
  NAND2_X1 U18816 ( .A1(n15568), .A2(n15567), .ZN(n15569) );
  AOI21_X1 U18817 ( .B1(n15712), .B2(n19428), .A(n15569), .ZN(n15572) );
  OR2_X1 U18818 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15714) );
  NAND3_X1 U18819 ( .A1(n15714), .A2(n15713), .A3(n16450), .ZN(n15571) );
  OAI211_X1 U18820 ( .C1(n15717), .C2(n19423), .A(n15572), .B(n15571), .ZN(
        P2_U2987) );
  INV_X1 U18821 ( .A(n15597), .ZN(n15574) );
  NAND2_X1 U18822 ( .A1(n15574), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15575) );
  AOI22_X1 U18823 ( .A1(n15575), .A2(n15595), .B1(n15597), .B2(n15745), .ZN(
        n15590) );
  AOI21_X1 U18824 ( .B1(n15590), .B2(n15587), .A(n15586), .ZN(n15576) );
  XOR2_X1 U18825 ( .A(n15577), .B(n15576), .Z(n15729) );
  INV_X1 U18826 ( .A(n15578), .ZN(n15585) );
  AOI21_X1 U18827 ( .B1(n9930), .B2(n15585), .A(n9694), .ZN(n15727) );
  NOR2_X1 U18828 ( .A1(n16466), .A2(n20079), .ZN(n15722) );
  AOI21_X1 U18829 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15722), .ZN(n15581) );
  NAND2_X1 U18830 ( .A1(n16440), .A2(n15579), .ZN(n15580) );
  OAI211_X1 U18831 ( .C1(n15718), .C2(n15688), .A(n15581), .B(n15580), .ZN(
        n15582) );
  AOI21_X1 U18832 ( .B1(n15727), .B2(n16449), .A(n15582), .ZN(n15583) );
  OAI21_X1 U18833 ( .B1(n15729), .B2(n19424), .A(n15583), .ZN(P2_U2988) );
  INV_X1 U18834 ( .A(n15584), .ZN(n15599) );
  OAI21_X1 U18835 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15599), .A(
        n15585), .ZN(n15740) );
  INV_X1 U18836 ( .A(n15586), .ZN(n15588) );
  NAND2_X1 U18837 ( .A1(n15588), .A2(n15587), .ZN(n15589) );
  XNOR2_X1 U18838 ( .A(n15590), .B(n15589), .ZN(n15738) );
  NAND2_X1 U18839 ( .A1(n19420), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15730) );
  OAI21_X1 U18840 ( .B1(n16453), .B2(n16349), .A(n15730), .ZN(n15591) );
  AOI21_X1 U18841 ( .B1(n16440), .B2(n16357), .A(n15591), .ZN(n15592) );
  OAI21_X1 U18842 ( .B1(n16352), .B2(n15688), .A(n15592), .ZN(n15593) );
  AOI21_X1 U18843 ( .B1(n15738), .B2(n16450), .A(n15593), .ZN(n15594) );
  OAI21_X1 U18844 ( .B1(n19423), .B2(n15740), .A(n15594), .ZN(P2_U2989) );
  XNOR2_X1 U18845 ( .A(n15595), .B(n15745), .ZN(n15596) );
  XNOR2_X1 U18846 ( .A(n15597), .B(n15596), .ZN(n15754) );
  AOI21_X1 U18847 ( .B1(n15745), .B2(n15598), .A(n15599), .ZN(n15741) );
  NAND2_X1 U18848 ( .A1(n15741), .A2(n16449), .ZN(n15604) );
  NOR2_X1 U18849 ( .A1(n16466), .A2(n20076), .ZN(n15744) );
  AOI21_X1 U18850 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15744), .ZN(n15600) );
  OAI21_X1 U18851 ( .B1(n19432), .B2(n15601), .A(n15600), .ZN(n15602) );
  AOI21_X1 U18852 ( .B1(n15751), .B2(n19428), .A(n15602), .ZN(n15603) );
  OAI211_X1 U18853 ( .C1(n15754), .C2(n19424), .A(n15604), .B(n15603), .ZN(
        P2_U2990) );
  INV_X1 U18854 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15756) );
  NOR2_X1 U18855 ( .A1(n15605), .A2(n15756), .ZN(n15613) );
  OAI21_X1 U18856 ( .B1(n15613), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15598), .ZN(n15767) );
  XOR2_X1 U18857 ( .A(n15607), .B(n15606), .Z(n15765) );
  NOR2_X1 U18858 ( .A1(n16466), .A2(n20074), .ZN(n15759) );
  AOI21_X1 U18859 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15759), .ZN(n15610) );
  NAND2_X1 U18860 ( .A1(n16440), .A2(n15608), .ZN(n15609) );
  OAI211_X1 U18861 ( .C1(n15763), .C2(n15688), .A(n15610), .B(n15609), .ZN(
        n15611) );
  AOI21_X1 U18862 ( .B1(n15765), .B2(n16450), .A(n15611), .ZN(n15612) );
  OAI21_X1 U18863 ( .B1(n15767), .B2(n19423), .A(n15612), .ZN(P2_U2991) );
  INV_X1 U18864 ( .A(n15613), .ZN(n15614) );
  OAI21_X1 U18865 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n11205), .A(
        n15614), .ZN(n15778) );
  INV_X1 U18866 ( .A(n15615), .ZN(n15616) );
  NOR2_X1 U18867 ( .A1(n15617), .A2(n15616), .ZN(n15618) );
  XNOR2_X1 U18868 ( .A(n15619), .B(n15618), .ZN(n15776) );
  NOR2_X1 U18869 ( .A1(n16466), .A2(n20072), .ZN(n15771) );
  NOR2_X1 U18870 ( .A1(n19432), .A2(n15976), .ZN(n15620) );
  AOI211_X1 U18871 ( .C1(n19421), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15771), .B(n15620), .ZN(n15621) );
  OAI21_X1 U18872 ( .B1(n15983), .B2(n15688), .A(n15621), .ZN(n15622) );
  AOI21_X1 U18873 ( .B1(n15776), .B2(n16450), .A(n15622), .ZN(n15623) );
  OAI21_X1 U18874 ( .B1(n15778), .B2(n19423), .A(n15623), .ZN(P2_U2992) );
  INV_X1 U18875 ( .A(n19136), .ZN(n19124) );
  AOI21_X1 U18876 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15624), .ZN(n15625) );
  OAI21_X1 U18877 ( .B1(n19432), .B2(n19124), .A(n15625), .ZN(n15628) );
  NOR2_X1 U18878 ( .A1(n15626), .A2(n19423), .ZN(n15627) );
  AOI211_X1 U18879 ( .C1(n19428), .C2(n19128), .A(n15628), .B(n15627), .ZN(
        n15629) );
  OAI21_X1 U18880 ( .B1(n15630), .B2(n19424), .A(n15629), .ZN(P2_U2993) );
  INV_X1 U18881 ( .A(n15631), .ZN(n15641) );
  NOR2_X1 U18882 ( .A1(n15641), .A2(n15791), .ZN(n15640) );
  OAI21_X1 U18883 ( .B1(n15640), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11199), .ZN(n15790) );
  NAND3_X1 U18884 ( .A1(n15780), .A2(n15779), .A3(n16450), .ZN(n15635) );
  NOR2_X1 U18885 ( .A1(n19178), .A2(n20068), .ZN(n15781) );
  AOI21_X1 U18886 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15781), .ZN(n15632) );
  OAI21_X1 U18887 ( .B1(n19432), .B2(n19143), .A(n15632), .ZN(n15633) );
  AOI21_X1 U18888 ( .B1(n19148), .B2(n19428), .A(n15633), .ZN(n15634) );
  OAI211_X1 U18889 ( .C1(n19423), .C2(n15790), .A(n15635), .B(n15634), .ZN(
        P2_U2994) );
  NOR2_X1 U18890 ( .A1(n15651), .A2(n15638), .ZN(n15639) );
  AOI21_X1 U18891 ( .B1(n15791), .B2(n15641), .A(n15640), .ZN(n15797) );
  NAND2_X1 U18892 ( .A1(n19420), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15794) );
  OAI21_X1 U18893 ( .B1(n16453), .B2(n15642), .A(n15794), .ZN(n15643) );
  AOI21_X1 U18894 ( .B1(n16440), .B2(n19154), .A(n15643), .ZN(n15644) );
  OAI21_X1 U18895 ( .B1(n19159), .B2(n15688), .A(n15644), .ZN(n15645) );
  AOI21_X1 U18896 ( .B1(n15797), .B2(n16449), .A(n15645), .ZN(n15646) );
  OAI21_X1 U18897 ( .B1(n15800), .B2(n19424), .A(n15646), .ZN(P2_U2995) );
  AOI21_X1 U18898 ( .B1(n15650), .B2(n15648), .A(n15647), .ZN(n15649) );
  AOI21_X1 U18899 ( .B1(n15651), .B2(n15650), .A(n15649), .ZN(n15811) );
  AOI21_X1 U18900 ( .B1(n15802), .B2(n15652), .A(n15631), .ZN(n15808) );
  NAND2_X1 U18901 ( .A1(n19170), .A2(n19428), .ZN(n15654) );
  NOR2_X1 U18902 ( .A1(n19178), .A2(n20065), .ZN(n15801) );
  AOI21_X1 U18903 ( .B1(n19421), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15801), .ZN(n15653) );
  OAI211_X1 U18904 ( .C1(n19168), .C2(n19432), .A(n15654), .B(n15653), .ZN(
        n15655) );
  AOI21_X1 U18905 ( .B1(n15808), .B2(n16449), .A(n15655), .ZN(n15656) );
  OAI21_X1 U18906 ( .B1(n15811), .B2(n19424), .A(n15656), .ZN(P2_U2996) );
  NAND2_X1 U18907 ( .A1(n15658), .A2(n15657), .ZN(n15660) );
  XOR2_X1 U18908 ( .A(n15660), .B(n15659), .Z(n15825) );
  NAND2_X1 U18909 ( .A1(n19420), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15820) );
  OAI21_X1 U18910 ( .B1(n16453), .B2(n15661), .A(n15820), .ZN(n15663) );
  NOR2_X1 U18911 ( .A1(n19184), .A2(n15688), .ZN(n15662) );
  AOI211_X1 U18912 ( .C1(n16440), .C2(n19176), .A(n15663), .B(n15662), .ZN(
        n15666) );
  INV_X1 U18913 ( .A(n15664), .ZN(n15813) );
  OAI211_X1 U18914 ( .C1(n15813), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16449), .B(n15652), .ZN(n15665) );
  OAI211_X1 U18915 ( .C1(n15825), .C2(n19424), .A(n15666), .B(n15665), .ZN(
        P2_U2997) );
  OAI21_X1 U18916 ( .B1(n10214), .B2(n10750), .A(n15668), .ZN(n15833) );
  NOR2_X1 U18917 ( .A1(n20062), .A2(n19178), .ZN(n15670) );
  OAI22_X1 U18918 ( .A1(n10035), .A2(n16453), .B1(n19432), .B2(n19196), .ZN(
        n15669) );
  AOI211_X1 U18919 ( .C1(n19428), .C2(n19198), .A(n15670), .B(n15669), .ZN(
        n15672) );
  OAI211_X1 U18920 ( .C1(n9725), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16449), .B(n15664), .ZN(n15671) );
  OAI211_X1 U18921 ( .C1(n15833), .C2(n19424), .A(n15672), .B(n15671), .ZN(
        P2_U2998) );
  AOI21_X1 U18922 ( .B1(n14229), .B2(n15674), .A(n15673), .ZN(n15679) );
  INV_X1 U18923 ( .A(n15675), .ZN(n15677) );
  NAND2_X1 U18924 ( .A1(n15677), .A2(n15676), .ZN(n15678) );
  XNOR2_X1 U18925 ( .A(n15679), .B(n15678), .ZN(n16500) );
  NAND2_X1 U18926 ( .A1(n15680), .A2(n15681), .ZN(n15683) );
  NAND2_X1 U18927 ( .A1(n15683), .A2(n15682), .ZN(n15684) );
  OAI22_X1 U18928 ( .A1(n11030), .A2(n19178), .B1(n19432), .B2(n19249), .ZN(
        n15690) );
  INV_X1 U18929 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15686) );
  OAI22_X1 U18930 ( .A1(n15688), .A2(n15687), .B1(n16453), .B2(n15686), .ZN(
        n15689) );
  AOI211_X1 U18931 ( .C1(n16497), .C2(n16449), .A(n15690), .B(n15689), .ZN(
        n15691) );
  OAI21_X1 U18932 ( .B1(n16500), .B2(n19424), .A(n15691), .ZN(P2_U3006) );
  INV_X1 U18933 ( .A(n15693), .ZN(n15694) );
  NOR2_X1 U18934 ( .A1(n15694), .A2(n14584), .ZN(n15698) );
  OAI21_X1 U18935 ( .B1(n15696), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15695), .ZN(n15697) );
  OAI21_X1 U18936 ( .B1(n16524), .B2(n15703), .A(n15702), .ZN(P2_U3016) );
  AOI21_X1 U18937 ( .B1(n15705), .B2(n11318), .A(n15704), .ZN(n15709) );
  INV_X1 U18938 ( .A(n15706), .ZN(n15707) );
  NAND2_X1 U18939 ( .A1(n15707), .A2(n19436), .ZN(n15708) );
  OAI211_X1 U18940 ( .C1(n15710), .C2(n11318), .A(n15709), .B(n15708), .ZN(
        n15711) );
  AOI21_X1 U18941 ( .B1(n15712), .B2(n19440), .A(n15711), .ZN(n15716) );
  NAND3_X1 U18942 ( .A1(n15714), .A2(n15713), .A3(n16519), .ZN(n15715) );
  OAI211_X1 U18943 ( .C1(n15717), .C2(n16524), .A(n15716), .B(n15715), .ZN(
        P2_U3019) );
  NOR2_X1 U18944 ( .A1(n15718), .A2(n16527), .ZN(n15726) );
  INV_X1 U18945 ( .A(n15719), .ZN(n15731) );
  AOI211_X1 U18946 ( .C1(n9930), .C2(n15732), .A(n15720), .B(n15731), .ZN(
        n15721) );
  AOI211_X1 U18947 ( .C1(n15723), .C2(n19436), .A(n15722), .B(n15721), .ZN(
        n15724) );
  OAI21_X1 U18948 ( .B1(n15733), .B2(n9930), .A(n15724), .ZN(n15725) );
  AOI211_X1 U18949 ( .C1(n15727), .C2(n19438), .A(n15726), .B(n15725), .ZN(
        n15728) );
  OAI21_X1 U18950 ( .B1(n15729), .B2(n19449), .A(n15728), .ZN(P2_U3020) );
  OAI21_X1 U18951 ( .B1(n15731), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15730), .ZN(n15735) );
  NOR2_X1 U18952 ( .A1(n15733), .A2(n15732), .ZN(n15734) );
  AOI211_X1 U18953 ( .C1(n19436), .C2(n16353), .A(n15735), .B(n15734), .ZN(
        n15736) );
  OAI21_X1 U18954 ( .B1(n16527), .B2(n16352), .A(n15736), .ZN(n15737) );
  AOI21_X1 U18955 ( .B1(n15738), .B2(n16519), .A(n15737), .ZN(n15739) );
  OAI21_X1 U18956 ( .B1(n16524), .B2(n15740), .A(n15739), .ZN(P2_U3021) );
  NAND2_X1 U18957 ( .A1(n15741), .A2(n19438), .ZN(n15753) );
  NAND2_X1 U18958 ( .A1(n15742), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15748) );
  INV_X1 U18959 ( .A(n15743), .ZN(n15746) );
  AOI21_X1 U18960 ( .B1(n15746), .B2(n15745), .A(n15744), .ZN(n15747) );
  OAI211_X1 U18961 ( .C1(n16526), .C2(n15749), .A(n15748), .B(n15747), .ZN(
        n15750) );
  AOI21_X1 U18962 ( .B1(n15751), .B2(n19440), .A(n15750), .ZN(n15752) );
  OAI211_X1 U18963 ( .C1(n15754), .C2(n19449), .A(n15753), .B(n15752), .ZN(
        P2_U3022) );
  AOI211_X1 U18964 ( .C1(n15757), .C2(n15756), .A(n15755), .B(n15769), .ZN(
        n15758) );
  AOI211_X1 U18965 ( .C1(n15760), .C2(n19436), .A(n15759), .B(n15758), .ZN(
        n15762) );
  NAND2_X1 U18966 ( .A1(n15772), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15761) );
  OAI211_X1 U18967 ( .C1(n15763), .C2(n16527), .A(n15762), .B(n15761), .ZN(
        n15764) );
  AOI21_X1 U18968 ( .B1(n15765), .B2(n16519), .A(n15764), .ZN(n15766) );
  OAI21_X1 U18969 ( .B1(n15767), .B2(n16524), .A(n15766), .ZN(P2_U3023) );
  XNOR2_X1 U18970 ( .A(n15768), .B(n9778), .ZN(n16365) );
  NOR2_X1 U18971 ( .A1(n15769), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15770) );
  AOI211_X1 U18972 ( .C1(n19436), .C2(n16365), .A(n15771), .B(n15770), .ZN(
        n15774) );
  NAND2_X1 U18973 ( .A1(n15772), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15773) );
  OAI211_X1 U18974 ( .C1(n15983), .C2(n16527), .A(n15774), .B(n15773), .ZN(
        n15775) );
  AOI21_X1 U18975 ( .B1(n15776), .B2(n16519), .A(n15775), .ZN(n15777) );
  OAI21_X1 U18976 ( .B1(n15778), .B2(n16524), .A(n15777), .ZN(P2_U3024) );
  NAND3_X1 U18977 ( .A1(n15780), .A2(n15779), .A3(n16519), .ZN(n15789) );
  INV_X1 U18978 ( .A(n15781), .ZN(n15784) );
  OAI211_X1 U18979 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15792), .B(n15782), .ZN(
        n15783) );
  OAI211_X1 U18980 ( .C1(n16526), .C2(n19151), .A(n15784), .B(n15783), .ZN(
        n15787) );
  NOR2_X1 U18981 ( .A1(n15785), .A2(n16527), .ZN(n15786) );
  AOI211_X1 U18982 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15807), .A(
        n15787), .B(n15786), .ZN(n15788) );
  OAI211_X1 U18983 ( .C1(n15790), .C2(n16524), .A(n15789), .B(n15788), .ZN(
        P2_U3026) );
  NAND2_X1 U18984 ( .A1(n15792), .A2(n15791), .ZN(n15793) );
  OAI211_X1 U18985 ( .C1(n16526), .C2(n19158), .A(n15794), .B(n15793), .ZN(
        n15796) );
  NOR2_X1 U18986 ( .A1(n19159), .A2(n16527), .ZN(n15795) );
  AOI211_X1 U18987 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15807), .A(
        n15796), .B(n15795), .ZN(n15799) );
  NAND2_X1 U18988 ( .A1(n15797), .A2(n19438), .ZN(n15798) );
  OAI211_X1 U18989 ( .C1(n15800), .C2(n19449), .A(n15799), .B(n15798), .ZN(
        P2_U3027) );
  NAND2_X1 U18990 ( .A1(n19170), .A2(n19440), .ZN(n15805) );
  AOI21_X1 U18991 ( .B1(n15803), .B2(n15802), .A(n15801), .ZN(n15804) );
  OAI211_X1 U18992 ( .C1(n16526), .C2(n19174), .A(n15805), .B(n15804), .ZN(
        n15806) );
  AOI21_X1 U18993 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15807), .A(
        n15806), .ZN(n15810) );
  NAND2_X1 U18994 ( .A1(n15808), .A2(n19438), .ZN(n15809) );
  OAI211_X1 U18995 ( .C1(n15811), .C2(n19449), .A(n15810), .B(n15809), .ZN(
        P2_U3028) );
  INV_X1 U18996 ( .A(n15812), .ZN(n15816) );
  AOI21_X1 U18997 ( .B1(n16524), .B2(n15814), .A(n15813), .ZN(n15815) );
  INV_X1 U18998 ( .A(n15817), .ZN(n16456) );
  NOR3_X1 U18999 ( .A1(n15829), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15818), .ZN(n15822) );
  NAND2_X1 U19000 ( .A1(n19436), .A2(n19185), .ZN(n15819) );
  OAI211_X1 U19001 ( .C1(n19184), .C2(n16527), .A(n15820), .B(n15819), .ZN(
        n15821) );
  OAI21_X1 U19002 ( .B1(n15825), .B2(n19449), .A(n15824), .ZN(P2_U3029) );
  INV_X1 U19003 ( .A(n19202), .ZN(n15826) );
  AOI22_X1 U19004 ( .A1(n19436), .A2(n15826), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19420), .ZN(n15828) );
  NAND2_X1 U19005 ( .A1(n19198), .A2(n19440), .ZN(n15827) );
  OAI211_X1 U19006 ( .C1(n15829), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15828), .B(n15827), .ZN(n15830) );
  AOI21_X1 U19007 ( .B1(n15831), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15830), .ZN(n15832) );
  OAI21_X1 U19008 ( .B1(n19449), .B2(n15833), .A(n15832), .ZN(P2_U3030) );
  NAND2_X1 U19009 ( .A1(n15834), .A2(n16371), .ZN(n15836) );
  XOR2_X1 U19010 ( .A(n15836), .B(n15835), .Z(n16383) );
  OR2_X1 U19011 ( .A1(n15838), .A2(n15846), .ZN(n16388) );
  NAND2_X1 U19012 ( .A1(n16388), .A2(n15842), .ZN(n15839) );
  NAND2_X1 U19013 ( .A1(n9999), .A2(n15839), .ZN(n16382) );
  INV_X1 U19014 ( .A(n16382), .ZN(n15852) );
  NAND2_X1 U19015 ( .A1(n16479), .A2(n15877), .ZN(n15840) );
  NOR2_X1 U19016 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15840), .ZN(
        n15860) );
  OAI21_X1 U19017 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15841), .A(
        n15892), .ZN(n15876) );
  INV_X1 U19018 ( .A(n15876), .ZN(n16489) );
  OAI21_X1 U19019 ( .B1(n16479), .B2(n15841), .A(n16489), .ZN(n15861) );
  NOR2_X1 U19020 ( .A1(n15860), .A2(n15861), .ZN(n16469) );
  NAND3_X1 U19021 ( .A1(n16479), .A2(n15877), .A3(n16468), .ZN(n16467) );
  AOI21_X1 U19022 ( .B1(n16469), .B2(n16467), .A(n15842), .ZN(n15851) );
  INV_X1 U19023 ( .A(n15348), .ZN(n15843) );
  OAI21_X1 U19024 ( .B1(n9705), .B2(n15844), .A(n15843), .ZN(n19344) );
  OAI22_X1 U19025 ( .A1(n16526), .A2(n19344), .B1(n15845), .B2(n19178), .ZN(
        n15848) );
  NOR3_X1 U19026 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15846), .A3(
        n16478), .ZN(n15847) );
  AOI211_X1 U19027 ( .C1(n19440), .C2(n19209), .A(n15848), .B(n15847), .ZN(
        n15849) );
  INV_X1 U19028 ( .A(n15849), .ZN(n15850) );
  AOI211_X1 U19029 ( .C1(n15852), .C2(n19438), .A(n15851), .B(n15850), .ZN(
        n15853) );
  OAI21_X1 U19030 ( .B1(n16383), .B2(n19449), .A(n15853), .ZN(P2_U3032) );
  INV_X1 U19031 ( .A(n16479), .ZN(n15854) );
  OR2_X1 U19032 ( .A1(n15838), .A2(n15854), .ZN(n16413) );
  XNOR2_X1 U19033 ( .A(n16413), .B(n16387), .ZN(n16401) );
  NOR2_X1 U19034 ( .A1(n15856), .A2(n15855), .ZN(n15857) );
  XNOR2_X1 U19035 ( .A(n15858), .B(n15857), .ZN(n16400) );
  NOR2_X1 U19036 ( .A1(n11094), .A2(n19178), .ZN(n15859) );
  AOI211_X1 U19037 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15861), .A(
        n15860), .B(n15859), .ZN(n15864) );
  INV_X1 U19038 ( .A(n19234), .ZN(n15862) );
  AOI22_X1 U19039 ( .A1(n19440), .A2(n19230), .B1(n19436), .B2(n15862), .ZN(
        n15863) );
  OAI211_X1 U19040 ( .C1(n16400), .C2(n19449), .A(n15864), .B(n15863), .ZN(
        n15865) );
  INV_X1 U19041 ( .A(n15865), .ZN(n15866) );
  OAI21_X1 U19042 ( .B1(n16401), .B2(n16524), .A(n15866), .ZN(P2_U3034) );
  XNOR2_X1 U19043 ( .A(n15838), .B(n15867), .ZN(n16420) );
  NAND2_X1 U19044 ( .A1(n15869), .A2(n15868), .ZN(n15888) );
  INV_X1 U19045 ( .A(n15886), .ZN(n15870) );
  OAI21_X1 U19046 ( .B1(n15888), .B2(n15870), .A(n15885), .ZN(n15874) );
  AND2_X1 U19047 ( .A1(n15872), .A2(n15871), .ZN(n15873) );
  XNOR2_X1 U19048 ( .A(n15874), .B(n15873), .ZN(n16419) );
  NOR2_X1 U19049 ( .A1(n11063), .A2(n16466), .ZN(n15875) );
  AOI221_X1 U19050 ( .B1(n15877), .B2(n15867), .C1(n15876), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15875), .ZN(n15880) );
  INV_X1 U19051 ( .A(n19244), .ZN(n15878) );
  AOI22_X1 U19052 ( .A1(n19440), .A2(n9761), .B1(n19436), .B2(n15878), .ZN(
        n15879) );
  OAI211_X1 U19053 ( .C1(n16419), .C2(n19449), .A(n15880), .B(n15879), .ZN(
        n15881) );
  INV_X1 U19054 ( .A(n15881), .ZN(n15882) );
  OAI21_X1 U19055 ( .B1(n16420), .B2(n16524), .A(n15882), .ZN(P2_U3036) );
  INV_X1 U19056 ( .A(n15883), .ZN(n15884) );
  INV_X1 U19057 ( .A(n15838), .ZN(n16412) );
  AOI21_X1 U19058 ( .B1(n15884), .B2(n15891), .A(n16412), .ZN(n16427) );
  INV_X1 U19059 ( .A(n16427), .ZN(n15900) );
  AND2_X1 U19060 ( .A1(n15886), .A2(n15885), .ZN(n15887) );
  XNOR2_X1 U19061 ( .A(n15888), .B(n15887), .ZN(n16426) );
  NAND2_X1 U19062 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19420), .ZN(n15889) );
  OAI21_X1 U19063 ( .B1(n16527), .B2(n15890), .A(n15889), .ZN(n15894) );
  NOR2_X1 U19064 ( .A1(n15892), .A2(n15891), .ZN(n15893) );
  AOI211_X1 U19065 ( .C1(n19436), .C2(n15895), .A(n15894), .B(n15893), .ZN(
        n15896) );
  OAI21_X1 U19066 ( .B1(n15897), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15896), .ZN(n15898) );
  AOI21_X1 U19067 ( .B1(n16426), .B2(n16519), .A(n15898), .ZN(n15899) );
  OAI21_X1 U19068 ( .B1(n15900), .B2(n16524), .A(n15899), .ZN(P2_U3037) );
  NOR2_X1 U19069 ( .A1(n13314), .A2(n16544), .ZN(n15902) );
  AOI22_X1 U19070 ( .A1(n19288), .A2(n10375), .B1(n19330), .B2(n19257), .ZN(
        n15906) );
  NOR2_X1 U19071 ( .A1(n15906), .A2(n16035), .ZN(n15901) );
  AOI211_X1 U19072 ( .C1(n15911), .C2(n15903), .A(n15902), .B(n15901), .ZN(
        n15905) );
  AOI21_X1 U19073 ( .B1(n10927), .B2(n15911), .A(n15953), .ZN(n15904) );
  OAI22_X1 U19074 ( .A1(n15905), .A2(n15953), .B1(n15904), .B2(n10222), .ZN(
        P2_U3601) );
  NAND2_X1 U19075 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15906), .ZN(n15916) );
  INV_X1 U19076 ( .A(n15916), .ZN(n15910) );
  AOI211_X1 U19077 ( .C1(n15909), .C2(n15908), .A(n19288), .B(n15907), .ZN(
        n19307) );
  AOI21_X1 U19078 ( .B1(n19288), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19307), .ZN(n15915) );
  AOI22_X1 U19079 ( .A1(n15912), .A2(n15911), .B1(n15910), .B2(n15915), .ZN(
        n15913) );
  OAI21_X1 U19080 ( .B1(n20099), .B2(n16544), .A(n15913), .ZN(n15914) );
  MUX2_X1 U19081 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15914), .S(
        n15956), .Z(P2_U3600) );
  OAI22_X1 U19082 ( .A1(n15917), .A2(n20100), .B1(n15916), .B2(n15915), .ZN(
        n15918) );
  AOI21_X1 U19083 ( .B1(n20111), .B2(n15919), .A(n15918), .ZN(n15921) );
  NAND2_X1 U19084 ( .A1(n15953), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15920) );
  OAI21_X1 U19085 ( .B1(n15921), .B2(n15953), .A(n15920), .ZN(P2_U3599) );
  AOI22_X1 U19086 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15925) );
  AOI22_X1 U19087 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15924) );
  AOI22_X1 U19088 ( .A1(n17368), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15923) );
  AOI22_X1 U19089 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15922) );
  NAND4_X1 U19090 ( .A1(n15925), .A2(n15924), .A3(n15923), .A4(n15922), .ZN(
        n15931) );
  AOI22_X1 U19091 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15929) );
  AOI22_X1 U19092 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12584), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15928) );
  AOI22_X1 U19093 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15927) );
  AOI22_X1 U19094 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15926) );
  NAND4_X1 U19095 ( .A1(n15929), .A2(n15928), .A3(n15927), .A4(n15926), .ZN(
        n15930) );
  NOR2_X1 U19096 ( .A1(n15931), .A2(n15930), .ZN(n17537) );
  NAND3_X1 U19097 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .ZN(n15932) );
  NAND3_X1 U19098 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17402), .ZN(n17381) );
  NOR2_X1 U19099 ( .A1(n15932), .A2(n17381), .ZN(n17333) );
  NOR2_X1 U19100 ( .A1(n15933), .A2(n17381), .ZN(n17318) );
  INV_X1 U19101 ( .A(n17318), .ZN(n17304) );
  OAI21_X1 U19102 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17333), .A(n17304), .ZN(
        n15934) );
  AOI22_X1 U19103 ( .A1(n17435), .A2(n17537), .B1(n15934), .B2(n17431), .ZN(
        P3_U2690) );
  NAND2_X1 U19104 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18630) );
  AOI221_X1 U19105 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18630), .C1(n15936), 
        .C2(n18630), .A(n15935), .ZN(n18408) );
  NOR2_X1 U19106 ( .A1(n15937), .A2(n18679), .ZN(n15938) );
  OAI21_X1 U19107 ( .B1(n15938), .B2(n18758), .A(n18409), .ZN(n18406) );
  AOI22_X1 U19108 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18408), .B1(
        n18406), .B2(n18906), .ZN(P3_U2865) );
  NAND2_X1 U19109 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19075) );
  NAND2_X1 U19110 ( .A1(n18856), .A2(n19075), .ZN(n15947) );
  INV_X2 U19111 ( .A(n19084), .ZN(n19083) );
  OAI211_X1 U19112 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18952), .B(n19017), .ZN(n19072) );
  INV_X1 U19113 ( .A(n19072), .ZN(n16732) );
  NAND2_X1 U19114 ( .A1(n16731), .A2(n16732), .ZN(n17599) );
  INV_X1 U19115 ( .A(n19075), .ZN(n18943) );
  INV_X1 U19116 ( .A(n18879), .ZN(n18863) );
  NOR3_X4 U19117 ( .A1(n18943), .A2(n15939), .A3(n16710), .ZN(n16040) );
  NOR2_X1 U19118 ( .A1(n15941), .A2(n15940), .ZN(n15944) );
  OAI21_X1 U19119 ( .B1(n15944), .B2(n15943), .A(n15942), .ZN(n15959) );
  NOR3_X1 U19120 ( .A1(n16040), .A2(n15945), .A3(n15959), .ZN(n15946) );
  NOR2_X1 U19121 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19028), .ZN(n18415) );
  INV_X1 U19122 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18404) );
  NOR2_X1 U19123 ( .A1(n18404), .A2(n19026), .ZN(n15948) );
  AOI211_X1 U19124 ( .C1(n19069), .C2(n18900), .A(n18415), .B(n15948), .ZN(
        n19056) );
  INV_X1 U19125 ( .A(n19056), .ZN(n19054) );
  INV_X1 U19126 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18862) );
  INV_X1 U19127 ( .A(n19032), .ZN(n19087) );
  INV_X1 U19128 ( .A(n18885), .ZN(n15949) );
  NOR2_X1 U19129 ( .A1(n15950), .A2(n15949), .ZN(n18915) );
  NAND3_X1 U19130 ( .A1(n19054), .A2(n19087), .A3(n18915), .ZN(n15951) );
  OAI21_X1 U19131 ( .B1(n19054), .B2(n18862), .A(n15951), .ZN(P3_U3284) );
  OR3_X1 U19132 ( .A1(n15953), .A2(n20100), .A3(n15952), .ZN(n15954) );
  OAI21_X1 U19133 ( .B1(n15956), .B2(n15955), .A(n15954), .ZN(P2_U3595) );
  INV_X1 U19134 ( .A(n18857), .ZN(n15964) );
  OAI21_X1 U19135 ( .B1(n18423), .B2(n16733), .A(n19072), .ZN(n15957) );
  OAI21_X1 U19136 ( .B1(n15958), .B2(n15957), .A(n19075), .ZN(n16709) );
  NOR3_X1 U19137 ( .A1(n15961), .A2(n16710), .A3(n16709), .ZN(n15960) );
  AOI211_X1 U19138 ( .C1(n15961), .C2(n18853), .A(n15960), .B(n15959), .ZN(
        n15963) );
  AOI221_X4 U19139 ( .B1(n15964), .B2(n15963), .C1(n15962), .C2(n15963), .A(
        n18924), .ZN(n18382) );
  INV_X1 U19140 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19036) );
  NAND3_X1 U19141 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18191) );
  NAND2_X1 U19142 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18307) );
  NOR2_X1 U19143 ( .A1(n9664), .A2(n18307), .ZN(n18192) );
  INV_X1 U19144 ( .A(n18192), .ZN(n18255) );
  NOR4_X1 U19145 ( .A1(n18380), .A2(n19036), .A3(n18191), .A4(n18255), .ZN(
        n18206) );
  NAND2_X1 U19146 ( .A1(n17863), .A2(n18206), .ZN(n15972) );
  INV_X1 U19147 ( .A(n15972), .ZN(n18143) );
  NAND2_X1 U19148 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18206), .ZN(
        n18275) );
  INV_X1 U19149 ( .A(n18275), .ZN(n18230) );
  NAND2_X1 U19150 ( .A1(n17863), .A2(n18230), .ZN(n18207) );
  NAND2_X1 U19151 ( .A1(n18081), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16589) );
  INV_X1 U19152 ( .A(n18191), .ZN(n18306) );
  OAI21_X1 U19153 ( .B1(n18385), .B2(n19036), .A(n18380), .ZN(n18362) );
  NAND2_X1 U19154 ( .A1(n18306), .A2(n18362), .ZN(n18304) );
  NOR2_X1 U19155 ( .A1(n18304), .A2(n18255), .ZN(n18232) );
  NAND2_X1 U19156 ( .A1(n17863), .A2(n18232), .ZN(n18145) );
  NAND2_X1 U19157 ( .A1(n18881), .A2(n18145), .ZN(n18183) );
  OAI21_X1 U19158 ( .B1(n18081), .B2(n18363), .A(n18183), .ZN(n18086) );
  AOI221_X1 U19159 ( .B1(n18207), .B2(n18864), .C1(n16589), .C2(n18864), .A(
        n18086), .ZN(n15965) );
  OAI221_X1 U19160 ( .B1(n18872), .B2(n18081), .C1(n18872), .C2(n18143), .A(
        n15965), .ZN(n16024) );
  AOI21_X1 U19161 ( .B1(n18248), .B2(n9991), .A(n16024), .ZN(n16596) );
  OAI21_X1 U19162 ( .B1(n18345), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16596), .ZN(n15968) );
  INV_X1 U19163 ( .A(n15969), .ZN(n18858) );
  NOR2_X1 U19164 ( .A1(n18858), .A2(n18399), .ZN(n18398) );
  NAND2_X1 U19165 ( .A1(n17565), .A2(n18398), .ZN(n18310) );
  NOR2_X1 U19166 ( .A1(n18249), .A2(n18399), .ZN(n18396) );
  OAI22_X1 U19167 ( .A1(n16561), .A2(n18310), .B1(n16558), .B2(n18374), .ZN(
        n15966) );
  NOR2_X1 U19168 ( .A1(n18359), .A2(n15966), .ZN(n16025) );
  INV_X1 U19169 ( .A(n16025), .ZN(n15967) );
  AOI21_X1 U19170 ( .B1(n18382), .B2(n15968), .A(n15967), .ZN(n15975) );
  NAND3_X1 U19171 ( .A1(n16594), .A2(n15969), .A3(n18382), .ZN(n18312) );
  OAI21_X1 U19172 ( .B1(n15971), .B2(n16563), .A(n15970), .ZN(n16566) );
  OAI21_X1 U19173 ( .B1(n18385), .B2(n18894), .A(n18872), .ZN(n18190) );
  INV_X1 U19174 ( .A(n18190), .ZN(n18364) );
  OAI22_X1 U19175 ( .A1(n18363), .A2(n18145), .B1(n15972), .B2(n18364), .ZN(
        n18104) );
  NOR2_X1 U19176 ( .A1(n18858), .A2(n16594), .ZN(n18277) );
  AOI22_X1 U19177 ( .A1(n18852), .A2(n17885), .B1(n17886), .B2(n18277), .ZN(
        n18194) );
  INV_X1 U19178 ( .A(n18194), .ZN(n15973) );
  NOR2_X1 U19179 ( .A1(n18399), .A2(n18152), .ZN(n16591) );
  INV_X1 U19180 ( .A(n16591), .ZN(n18156) );
  NOR3_X1 U19181 ( .A1(n16587), .A2(n16589), .A3(n18156), .ZN(n16027) );
  AOI22_X1 U19182 ( .A1(n18299), .A2(n16566), .B1(n16027), .B2(n16563), .ZN(
        n15974) );
  NAND2_X1 U19183 ( .A1(n18393), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16573) );
  OAI211_X1 U19184 ( .C1(n15975), .C2(n16563), .A(n15974), .B(n16573), .ZN(
        P3_U2833) );
  OAI21_X1 U19185 ( .B1(n15977), .B2(n15976), .A(n19306), .ZN(n15987) );
  INV_X1 U19186 ( .A(n15978), .ZN(n15980) );
  OAI222_X1 U19187 ( .A1(n19302), .A2(n15980), .B1(n19262), .B2(n20072), .C1(
        n15979), .C2(n19180), .ZN(n15981) );
  AOI21_X1 U19188 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19323), .A(
        n15981), .ZN(n15986) );
  INV_X1 U19189 ( .A(n16365), .ZN(n15982) );
  OAI22_X1 U19190 ( .A1(n15983), .A2(n19320), .B1(n15982), .B2(n19315), .ZN(
        n15984) );
  INV_X1 U19191 ( .A(n15984), .ZN(n15985) );
  OAI211_X1 U19192 ( .C1(n15988), .C2(n15987), .A(n15986), .B(n15985), .ZN(
        P2_U2833) );
  INV_X1 U19193 ( .A(n15989), .ZN(n16000) );
  AOI21_X1 U19194 ( .B1(n15990), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20647), .ZN(n15991) );
  AND2_X1 U19195 ( .A1(n15992), .A2(n15991), .ZN(n15994) );
  INV_X1 U19196 ( .A(n15994), .ZN(n15998) );
  INV_X1 U19197 ( .A(n15993), .ZN(n15995) );
  OAI22_X1 U19198 ( .A1(n15996), .A2(n15995), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15994), .ZN(n15997) );
  OAI21_X1 U19199 ( .B1(n15998), .B2(n20686), .A(n15997), .ZN(n15999) );
  AOI222_X1 U19200 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16000), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15999), .C1(n16000), 
        .C2(n15999), .ZN(n16002) );
  AOI222_X1 U19201 ( .A1(n16002), .A2(n20727), .B1(n16002), .B2(n16001), .C1(
        n20727), .C2(n16001), .ZN(n16009) );
  NOR3_X1 U19202 ( .A1(n16005), .A2(n16004), .A3(n16003), .ZN(n16008) );
  OAI21_X1 U19203 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16006), .ZN(n16007) );
  OAI211_X1 U19204 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n16009), .A(
        n16008), .B(n16007), .ZN(n16014) );
  NOR3_X1 U19205 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11760), .A3(n20953), 
        .ZN(n16012) );
  OAI22_X1 U19206 ( .A1(n16015), .A2(n16012), .B1(n16011), .B2(n16010), .ZN(
        n16320) );
  AOI221_X1 U19207 ( .B1(n20865), .B2(n13651), .C1(n16014), .C2(n13651), .A(
        n16320), .ZN(n16016) );
  NOR2_X1 U19208 ( .A1(n16016), .A2(n20865), .ZN(n16323) );
  OAI211_X1 U19209 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20953), .A(n16323), 
        .B(n16013), .ZN(n16321) );
  AOI21_X1 U19210 ( .B1(n16015), .B2(n16014), .A(n16321), .ZN(n16020) );
  AOI21_X1 U19211 ( .B1(n20958), .B2(n20936), .A(n16016), .ZN(n16017) );
  INV_X1 U19212 ( .A(n16017), .ZN(n16018) );
  AOI22_X1 U19213 ( .A1(n16020), .A2(n16019), .B1(n20865), .B2(n16018), .ZN(
        P1_U3161) );
  NAND2_X1 U19214 ( .A1(n16022), .A2(n16021), .ZN(n16023) );
  XOR2_X1 U19215 ( .A(n16023), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16557) );
  NOR2_X1 U19216 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16578), .ZN(
        n16553) );
  INV_X1 U19217 ( .A(n18345), .ZN(n18210) );
  OAI211_X1 U19218 ( .C1(n16024), .C2(n16578), .A(n18210), .B(n18382), .ZN(
        n16575) );
  INV_X1 U19219 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16577) );
  AOI21_X1 U19220 ( .B1(n16575), .B2(n16025), .A(n16577), .ZN(n16026) );
  AOI21_X1 U19221 ( .B1(n16027), .B2(n16553), .A(n16026), .ZN(n16028) );
  INV_X2 U19222 ( .A(n9655), .ZN(n18393) );
  NAND2_X1 U19223 ( .A1(n18393), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16548) );
  OAI211_X1 U19224 ( .C1(n18312), .C2(n16557), .A(n16028), .B(n16548), .ZN(
        P3_U2832) );
  INV_X1 U19225 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20874) );
  INV_X1 U19226 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21122) );
  NOR2_X1 U19227 ( .A1(n12994), .A2(n21122), .ZN(n20870) );
  INV_X1 U19228 ( .A(HOLD), .ZN(n21071) );
  INV_X1 U19229 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20883) );
  OAI222_X1 U19230 ( .A1(n20870), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n20870), 
        .B2(HOLD), .C1(n21071), .C2(n20883), .ZN(n16030) );
  OAI211_X1 U19231 ( .C1(n20953), .C2(n20874), .A(n16030), .B(n16029), .ZN(
        P1_U3195) );
  AND2_X1 U19232 ( .A1(n16031), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U19233 ( .A1(n16032), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16034) );
  AOI21_X1 U19234 ( .B1(n20117), .B2(n19097), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16033) );
  AOI21_X1 U19235 ( .B1(n16034), .B2(n16033), .A(n16535), .ZN(P2_U3178) );
  AOI21_X1 U19236 ( .B1(n19884), .B2(n16035), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20149) );
  NAND2_X1 U19237 ( .A1(n20149), .A2(n20127), .ZN(n16036) );
  INV_X1 U19238 ( .A(n20133), .ZN(n20134) );
  NOR2_X1 U19239 ( .A1(n16037), .A2(n20134), .ZN(P2_U3047) );
  NAND2_X1 U19240 ( .A1(n18448), .A2(n17591), .ZN(n17522) );
  INV_X1 U19241 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17672) );
  NOR2_X1 U19242 ( .A1(n16041), .A2(n17563), .ZN(n17595) );
  AOI22_X1 U19243 ( .A1(n17595), .A2(BUF2_REG_0__SCAN_IN), .B1(n17594), .B2(
        n16042), .ZN(n16043) );
  OAI221_X1 U19244 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17522), .C1(n17672), 
        .C2(n17591), .A(n16043), .ZN(P3_U2735) );
  AOI21_X1 U19245 ( .B1(n16044), .B2(P1_REIP_REG_16__SCAN_IN), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16055) );
  INV_X1 U19246 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16111) );
  OAI22_X1 U19247 ( .A1(n16045), .A2(n20245), .B1(n16111), .B2(n16102), .ZN(
        n16046) );
  AOI211_X1 U19248 ( .C1(n20229), .C2(n16130), .A(n20377), .B(n16046), .ZN(
        n16053) );
  OR2_X1 U19249 ( .A1(n14766), .A2(n16047), .ZN(n16048) );
  AND2_X1 U19250 ( .A1(n16048), .A2(n14749), .ZN(n16131) );
  NAND2_X1 U19251 ( .A1(n9747), .A2(n16049), .ZN(n16050) );
  NAND2_X1 U19252 ( .A1(n9693), .A2(n16050), .ZN(n16208) );
  NOR2_X1 U19253 ( .A1(n16208), .A2(n20243), .ZN(n16051) );
  AOI21_X1 U19254 ( .B1(n16131), .B2(n20210), .A(n16051), .ZN(n16052) );
  OAI211_X1 U19255 ( .C1(n16055), .C2(n16054), .A(n16053), .B(n16052), .ZN(
        P1_U2823) );
  INV_X1 U19256 ( .A(n16056), .ZN(n16230) );
  AOI22_X1 U19257 ( .A1(n16141), .A2(n20229), .B1(n20257), .B2(n16230), .ZN(
        n16064) );
  NOR2_X1 U19258 ( .A1(n20245), .A2(n16057), .ZN(n16062) );
  AOI22_X1 U19259 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(n20250), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n16069), .ZN(n16060) );
  INV_X1 U19260 ( .A(n16058), .ZN(n16059) );
  NAND3_X1 U19261 ( .A1(n20351), .A2(n16060), .A3(n16059), .ZN(n16061) );
  AOI211_X1 U19262 ( .C1(n16142), .C2(n20210), .A(n16062), .B(n16061), .ZN(
        n16063) );
  NAND2_X1 U19263 ( .A1(n16064), .A2(n16063), .ZN(P1_U2825) );
  AOI22_X1 U19264 ( .A1(n16066), .A2(n20229), .B1(n20257), .B2(n16065), .ZN(
        n16073) );
  AOI22_X1 U19265 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20215), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n20250), .ZN(n16072) );
  INV_X1 U19266 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20901) );
  NAND2_X1 U19267 ( .A1(n16089), .A2(n16067), .ZN(n16088) );
  OAI21_X1 U19268 ( .B1(n20901), .B2(n16088), .A(n15012), .ZN(n16068) );
  AOI22_X1 U19269 ( .A1(n16070), .A2(n20210), .B1(n16069), .B2(n16068), .ZN(
        n16071) );
  NAND4_X1 U19270 ( .A1(n16073), .A2(n16072), .A3(n16071), .A4(n20351), .ZN(
        P1_U2826) );
  OAI21_X1 U19271 ( .B1(n16075), .B2(n16074), .A(n20203), .ZN(n16098) );
  INV_X1 U19272 ( .A(n16076), .ZN(n16079) );
  INV_X1 U19273 ( .A(n16077), .ZN(n16078) );
  OAI21_X1 U19274 ( .B1(n16080), .B2(n16079), .A(n16078), .ZN(n16082) );
  AND2_X1 U19275 ( .A1(n16082), .A2(n16081), .ZN(n16234) );
  AOI22_X1 U19276 ( .A1(n16083), .A2(n20229), .B1(n20257), .B2(n16234), .ZN(
        n16085) );
  AOI21_X1 U19277 ( .B1(n20215), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20377), .ZN(n16084) );
  OAI211_X1 U19278 ( .C1(n16102), .C2(n16114), .A(n16085), .B(n16084), .ZN(
        n16086) );
  AOI21_X1 U19279 ( .B1(n16112), .B2(n20210), .A(n16086), .ZN(n16087) );
  OAI221_X1 U19280 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n16088), .C1(n20901), 
        .C2(n16098), .A(n16087), .ZN(P1_U2827) );
  AOI21_X1 U19281 ( .B1(n16089), .B2(P1_REIP_REG_11__SCAN_IN), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16099) );
  AOI22_X1 U19282 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20215), .B1(
        n20257), .B2(n16245), .ZN(n16090) );
  INV_X1 U19283 ( .A(n16090), .ZN(n16091) );
  AOI211_X1 U19284 ( .C1(n20250), .C2(P1_EBX_REG_12__SCAN_IN), .A(n20377), .B(
        n16091), .ZN(n16097) );
  OAI22_X1 U19285 ( .A1(n16094), .A2(n16093), .B1(n16092), .B2(n20244), .ZN(
        n16095) );
  INV_X1 U19286 ( .A(n16095), .ZN(n16096) );
  OAI211_X1 U19287 ( .C1(n16099), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        P1_U2828) );
  NOR2_X1 U19288 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n16100), .ZN(n16101) );
  AOI22_X1 U19289 ( .A1(n16153), .A2(n20229), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n16101), .ZN(n16108) );
  OAI22_X1 U19290 ( .A1(n16103), .A2(n16102), .B1(n20243), .B2(n16273), .ZN(
        n16104) );
  AOI211_X1 U19291 ( .C1(n20215), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20377), .B(n16104), .ZN(n16107) );
  AOI22_X1 U19292 ( .A1(n16154), .A2(n20210), .B1(n16105), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n16106) );
  NAND3_X1 U19293 ( .A1(n16108), .A2(n16107), .A3(n16106), .ZN(P1_U2830) );
  NOR2_X1 U19294 ( .A1(n16208), .A2(n20265), .ZN(n16109) );
  AOI21_X1 U19295 ( .B1(n16131), .B2(n12977), .A(n16109), .ZN(n16110) );
  OAI21_X1 U19296 ( .B1(n20270), .B2(n16111), .A(n16110), .ZN(P1_U2855) );
  AOI22_X1 U19297 ( .A1(n16112), .A2(n12977), .B1(n12975), .B2(n16234), .ZN(
        n16113) );
  OAI21_X1 U19298 ( .B1(n20270), .B2(n16114), .A(n16113), .ZN(P1_U2859) );
  AOI22_X1 U19299 ( .A1(n16117), .A2(n16116), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16115), .ZN(n16121) );
  AOI22_X1 U19300 ( .A1(n16131), .A2(n16119), .B1(n16118), .B2(DATAI_17_), 
        .ZN(n16120) );
  OAI211_X1 U19301 ( .C1(n16122), .C2(n16631), .A(n16121), .B(n16120), .ZN(
        P1_U2887) );
  NOR2_X1 U19302 ( .A1(n12396), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16128) );
  INV_X1 U19303 ( .A(n16123), .ZN(n16126) );
  OAI21_X1 U19304 ( .B1(n16126), .B2(n16125), .A(n16124), .ZN(n16127) );
  MUX2_X1 U19305 ( .A(n16146), .B(n16128), .S(n16127), .Z(n16129) );
  XNOR2_X1 U19306 ( .A(n16129), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16214) );
  AOI22_X1 U19307 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16133) );
  AOI22_X1 U19308 ( .A1(n16131), .A2(n20344), .B1(n16130), .B2(n16152), .ZN(
        n16132) );
  OAI211_X1 U19309 ( .C1(n20167), .C2(n16214), .A(n16133), .B(n16132), .ZN(
        P1_U2982) );
  INV_X1 U19310 ( .A(n16134), .ZN(n16135) );
  NOR2_X1 U19311 ( .A1(n16136), .A2(n16135), .ZN(n16140) );
  NAND2_X1 U19312 ( .A1(n16138), .A2(n16137), .ZN(n16139) );
  XNOR2_X1 U19313 ( .A(n16140), .B(n16139), .ZN(n16227) );
  AOI22_X1 U19314 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16144) );
  AOI22_X1 U19315 ( .A1(n16142), .A2(n20344), .B1(n16141), .B2(n16152), .ZN(
        n16143) );
  OAI211_X1 U19316 ( .C1(n16227), .C2(n20167), .A(n16144), .B(n16143), .ZN(
        P1_U2984) );
  XOR2_X1 U19317 ( .A(n16145), .B(n12908), .Z(n16148) );
  NAND2_X1 U19318 ( .A1(n14998), .A2(n12908), .ZN(n16147) );
  MUX2_X1 U19319 ( .A(n16148), .B(n16147), .S(n16146), .Z(n16151) );
  INV_X1 U19320 ( .A(n16149), .ZN(n16150) );
  NAND2_X1 U19321 ( .A1(n16151), .A2(n16150), .ZN(n16277) );
  AOI22_X1 U19322 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n16156) );
  AOI22_X1 U19323 ( .A1(n16154), .A2(n20344), .B1(n16153), .B2(n16152), .ZN(
        n16155) );
  OAI211_X1 U19324 ( .C1(n20167), .C2(n16277), .A(n16156), .B(n16155), .ZN(
        P1_U2989) );
  AOI22_X1 U19325 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16163) );
  INV_X1 U19326 ( .A(n16157), .ZN(n16159) );
  NAND2_X1 U19327 ( .A1(n16159), .A2(n16158), .ZN(n16160) );
  XNOR2_X1 U19328 ( .A(n16161), .B(n16160), .ZN(n16293) );
  AOI22_X1 U19329 ( .A1(n16293), .A2(n20343), .B1(n20344), .B2(n20261), .ZN(
        n16162) );
  OAI211_X1 U19330 ( .C1(n20349), .C2(n20195), .A(n16163), .B(n16162), .ZN(
        P1_U2992) );
  AOI22_X1 U19331 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16170) );
  OAI21_X1 U19332 ( .B1(n16166), .B2(n16165), .A(n16164), .ZN(n16167) );
  INV_X1 U19333 ( .A(n16167), .ZN(n16298) );
  INV_X1 U19334 ( .A(n16168), .ZN(n20211) );
  AOI22_X1 U19335 ( .A1(n16298), .A2(n20343), .B1(n20344), .B2(n20211), .ZN(
        n16169) );
  OAI211_X1 U19336 ( .C1(n20349), .C2(n20207), .A(n16170), .B(n16169), .ZN(
        P1_U2993) );
  AOI22_X1 U19337 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16176) );
  OAI21_X1 U19338 ( .B1(n16173), .B2(n16172), .A(n16171), .ZN(n16174) );
  INV_X1 U19339 ( .A(n16174), .ZN(n16308) );
  INV_X1 U19340 ( .A(n20266), .ZN(n20223) );
  AOI22_X1 U19341 ( .A1(n16308), .A2(n20343), .B1(n20344), .B2(n20223), .ZN(
        n16175) );
  OAI211_X1 U19342 ( .C1(n20349), .C2(n20226), .A(n16176), .B(n16175), .ZN(
        P1_U2994) );
  INV_X1 U19343 ( .A(n16177), .ZN(n16179) );
  AOI22_X1 U19344 ( .A1(n16179), .A2(n20375), .B1(n20372), .B2(n16178), .ZN(
        n16186) );
  INV_X1 U19345 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n16180) );
  NOR2_X1 U19346 ( .A1(n20351), .A2(n16180), .ZN(n16181) );
  AOI221_X1 U19347 ( .B1(n16184), .B2(n16183), .C1(n16182), .C2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16181), .ZN(n16185) );
  NAND2_X1 U19348 ( .A1(n16186), .A2(n16185), .ZN(P1_U3008) );
  OAI21_X1 U19349 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16187), .ZN(n16195) );
  OAI22_X1 U19350 ( .A1(n16190), .A2(n16189), .B1(n20352), .B2(n16188), .ZN(
        n16191) );
  AOI21_X1 U19351 ( .B1(n20375), .B2(n16192), .A(n16191), .ZN(n16194) );
  NAND2_X1 U19352 ( .A1(n20377), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16193) );
  OAI211_X1 U19353 ( .C1(n16196), .C2(n16195), .A(n16194), .B(n16193), .ZN(
        P1_U3009) );
  OR2_X1 U19354 ( .A1(n16198), .A2(n16197), .ZN(n16205) );
  AOI22_X1 U19355 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16199), .B1(
        n20377), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16204) );
  INV_X1 U19356 ( .A(n16200), .ZN(n16202) );
  AOI22_X1 U19357 ( .A1(n16202), .A2(n20375), .B1(n20372), .B2(n16201), .ZN(
        n16203) );
  OAI211_X1 U19358 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16205), .A(
        n16204), .B(n16203), .ZN(P1_U3012) );
  NAND2_X1 U19359 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16206), .ZN(
        n16225) );
  OAI21_X1 U19360 ( .B1(n16217), .B2(n16225), .A(n16207), .ZN(n16210) );
  INV_X1 U19361 ( .A(n16208), .ZN(n16209) );
  AOI22_X1 U19362 ( .A1(n16211), .A2(n16210), .B1(n20372), .B2(n16209), .ZN(
        n16213) );
  NAND2_X1 U19363 ( .A1(n20377), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16212) );
  OAI211_X1 U19364 ( .C1(n16214), .C2(n16278), .A(n16213), .B(n16212), .ZN(
        P1_U3014) );
  OAI21_X1 U19365 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16269), .A(
        n16242), .ZN(n16215) );
  INV_X1 U19366 ( .A(n16215), .ZN(n16233) );
  INV_X1 U19367 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16224) );
  INV_X1 U19368 ( .A(n16216), .ZN(n16222) );
  INV_X1 U19369 ( .A(n16217), .ZN(n16218) );
  AOI211_X1 U19370 ( .C1(n16232), .C2(n16224), .A(n16218), .B(n16225), .ZN(
        n16221) );
  OAI22_X1 U19371 ( .A1(n16219), .A2(n20352), .B1(n20906), .B2(n20351), .ZN(
        n16220) );
  AOI211_X1 U19372 ( .C1(n16222), .C2(n20375), .A(n16221), .B(n16220), .ZN(
        n16223) );
  OAI21_X1 U19373 ( .B1(n16233), .B2(n16224), .A(n16223), .ZN(P1_U3015) );
  OAI22_X1 U19374 ( .A1(n20351), .A2(n16226), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16225), .ZN(n16229) );
  NOR2_X1 U19375 ( .A1(n16227), .A2(n16278), .ZN(n16228) );
  AOI211_X1 U19376 ( .C1(n20372), .C2(n16230), .A(n16229), .B(n16228), .ZN(
        n16231) );
  OAI21_X1 U19377 ( .B1(n16233), .B2(n16232), .A(n16231), .ZN(P1_U3016) );
  INV_X1 U19378 ( .A(n16234), .ZN(n16235) );
  OAI22_X1 U19379 ( .A1(n16235), .A2(n20352), .B1(n20901), .B2(n20351), .ZN(
        n16238) );
  NOR2_X1 U19380 ( .A1(n16236), .A2(n16278), .ZN(n16237) );
  AOI211_X1 U19381 ( .C1(n16241), .C2(n16239), .A(n16238), .B(n16237), .ZN(
        n16240) );
  OAI21_X1 U19382 ( .B1(n16242), .B2(n16241), .A(n16240), .ZN(P1_U3018) );
  NAND3_X1 U19383 ( .A1(n16246), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16243), .ZN(n16255) );
  AOI21_X1 U19384 ( .B1(n16245), .B2(n20372), .A(n16244), .ZN(n16254) );
  AOI21_X1 U19385 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16246), .A(
        n20369), .ZN(n16248) );
  AOI211_X1 U19386 ( .C1(n20379), .C2(n16249), .A(n16248), .B(n16247), .ZN(
        n16264) );
  OAI21_X1 U19387 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16250), .A(
        n16264), .ZN(n16252) );
  AOI22_X1 U19388 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16252), .B1(
        n20375), .B2(n16251), .ZN(n16253) );
  OAI211_X1 U19389 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16255), .A(
        n16254), .B(n16253), .ZN(P1_U3019) );
  INV_X1 U19390 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16263) );
  INV_X1 U19391 ( .A(n16256), .ZN(n16257) );
  AOI21_X1 U19392 ( .B1(n16258), .B2(n20372), .A(n16257), .ZN(n16262) );
  AOI22_X1 U19393 ( .A1(n16260), .A2(n20375), .B1(n16259), .B2(n16263), .ZN(
        n16261) );
  OAI211_X1 U19394 ( .C1(n16264), .C2(n16263), .A(n16262), .B(n16261), .ZN(
        P1_U3020) );
  AOI211_X1 U19395 ( .C1(n16267), .C2(n20379), .A(n16266), .B(n16265), .ZN(
        n16270) );
  OAI21_X1 U19396 ( .B1(n16270), .B2(n16269), .A(n16268), .ZN(n16281) );
  NAND2_X1 U19397 ( .A1(n16271), .A2(n16292), .ZN(n16285) );
  AOI221_X1 U19398 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12908), .C2(n16272), .A(
        n16285), .ZN(n16275) );
  INV_X1 U19399 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20896) );
  OAI22_X1 U19400 ( .A1(n16273), .A2(n20352), .B1(n20896), .B2(n20351), .ZN(
        n16274) );
  AOI211_X1 U19401 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16281), .A(
        n16275), .B(n16274), .ZN(n16276) );
  OAI21_X1 U19402 ( .B1(n16278), .B2(n16277), .A(n16276), .ZN(P1_U3021) );
  AOI21_X1 U19403 ( .B1(n16280), .B2(n20372), .A(n16279), .ZN(n16284) );
  AOI22_X1 U19404 ( .A1(n16282), .A2(n20375), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16281), .ZN(n16283) );
  OAI211_X1 U19405 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16285), .A(
        n16284), .B(n16283), .ZN(P1_U3022) );
  NAND2_X1 U19406 ( .A1(n16305), .A2(n16286), .ZN(n16289) );
  INV_X1 U19407 ( .A(n16287), .ZN(n16288) );
  NAND2_X1 U19408 ( .A1(n16289), .A2(n16288), .ZN(n16291) );
  AND2_X1 U19409 ( .A1(n16291), .A2(n16290), .ZN(n20260) );
  AOI22_X1 U19410 ( .A1(n20260), .A2(n20372), .B1(n20377), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16295) );
  AOI22_X1 U19411 ( .A1(n16293), .A2(n20375), .B1(n16296), .B2(n16292), .ZN(
        n16294) );
  OAI211_X1 U19412 ( .C1(n16297), .C2(n16296), .A(n16295), .B(n16294), .ZN(
        P1_U3024) );
  AOI22_X1 U19413 ( .A1(n20205), .A2(n20372), .B1(n20377), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16300) );
  AOI22_X1 U19414 ( .A1(n16298), .A2(n20375), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16307), .ZN(n16299) );
  OAI211_X1 U19415 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16301), .A(
        n16300), .B(n16299), .ZN(P1_U3025) );
  NOR2_X1 U19416 ( .A1(n16303), .A2(n16302), .ZN(n16304) );
  OR2_X1 U19417 ( .A1(n16305), .A2(n16304), .ZN(n20264) );
  OAI22_X1 U19418 ( .A1(n20264), .A2(n20352), .B1(n20351), .B2(n20219), .ZN(
        n16306) );
  INV_X1 U19419 ( .A(n16306), .ZN(n16313) );
  AOI22_X1 U19420 ( .A1(n16308), .A2(n20375), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16307), .ZN(n16312) );
  NAND3_X1 U19421 ( .A1(n20354), .A2(n16310), .A3(n16309), .ZN(n16311) );
  NAND3_X1 U19422 ( .A1(n16313), .A2(n16312), .A3(n16311), .ZN(P1_U3026) );
  NAND3_X1 U19423 ( .A1(n16315), .A2(n20937), .A3(n16314), .ZN(n16316) );
  OAI21_X1 U19424 ( .B1(n16317), .B2(n13652), .A(n16316), .ZN(P1_U3468) );
  OAI221_X1 U19425 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20865), .C2(n20953), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20866) );
  NAND2_X1 U19426 ( .A1(n20866), .A2(n16318), .ZN(n16319) );
  AOI22_X1 U19427 ( .A1(n13651), .A2(n16321), .B1(n16320), .B2(n16319), .ZN(
        P1_U3162) );
  OAI21_X1 U19428 ( .B1(n16323), .B2(n20689), .A(n16322), .ZN(P1_U3466) );
  AOI211_X1 U19429 ( .C1(n16326), .C2(n16325), .A(n16324), .B(n19289), .ZN(
        n16334) );
  AOI22_X1 U19430 ( .A1(n19311), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19323), .ZN(n16327) );
  OAI21_X1 U19431 ( .B1(n16328), .B2(n19262), .A(n16327), .ZN(n16329) );
  AOI21_X1 U19432 ( .B1(n16330), .B2(n19317), .A(n16329), .ZN(n16331) );
  OAI21_X1 U19433 ( .B1(n16332), .B2(n19320), .A(n16331), .ZN(n16333) );
  AOI211_X1 U19434 ( .C1(n19305), .C2(n16335), .A(n16334), .B(n16333), .ZN(
        n16336) );
  INV_X1 U19435 ( .A(n16336), .ZN(P2_U2826) );
  AOI22_X1 U19436 ( .A1(n16338), .A2(n19285), .B1(n16337), .B2(n19305), .ZN(
        n16348) );
  AOI211_X1 U19437 ( .C1(n16341), .C2(n16340), .A(n16339), .B(n19289), .ZN(
        n16346) );
  INV_X1 U19438 ( .A(n16342), .ZN(n16344) );
  OAI222_X1 U19439 ( .A1(n19302), .A2(n16344), .B1(n19262), .B2(n20083), .C1(
        n16343), .C2(n19180), .ZN(n16345) );
  AOI211_X1 U19440 ( .C1(n19323), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16346), .B(n16345), .ZN(n16347) );
  NAND2_X1 U19441 ( .A1(n16348), .A2(n16347), .ZN(P2_U2827) );
  AOI22_X1 U19442 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19311), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19312), .ZN(n16362) );
  OAI22_X1 U19443 ( .A1(n16350), .A2(n19302), .B1(n19297), .B2(n16349), .ZN(
        n16351) );
  INV_X1 U19444 ( .A(n16351), .ZN(n16361) );
  INV_X1 U19445 ( .A(n16352), .ZN(n16354) );
  AOI22_X1 U19446 ( .A1(n16354), .A2(n19285), .B1(n16353), .B2(n19305), .ZN(
        n16360) );
  AOI21_X1 U19447 ( .B1(n16357), .B2(n16356), .A(n16355), .ZN(n16358) );
  NAND2_X1 U19448 ( .A1(n19306), .A2(n16358), .ZN(n16359) );
  NAND4_X1 U19449 ( .A1(n16362), .A2(n16361), .A3(n16360), .A4(n16359), .ZN(
        P2_U2830) );
  AOI22_X1 U19450 ( .A1(n16364), .A2(n16363), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19379), .ZN(n16369) );
  AOI22_X1 U19451 ( .A1(n19331), .A2(BUF1_REG_22__SCAN_IN), .B1(n19333), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16368) );
  AOI22_X1 U19452 ( .A1(n16366), .A2(n19381), .B1(n19380), .B2(n16365), .ZN(
        n16367) );
  NAND3_X1 U19453 ( .A1(n16369), .A2(n16368), .A3(n16367), .ZN(P2_U2897) );
  AOI22_X1 U19454 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19420), .B1(n16440), 
        .B2(n16370), .ZN(n16380) );
  NAND2_X1 U19455 ( .A1(n16372), .A2(n16371), .ZN(n16376) );
  AND2_X1 U19456 ( .A1(n16374), .A2(n16373), .ZN(n16375) );
  XNOR2_X1 U19457 ( .A(n16376), .B(n16375), .ZN(n16465) );
  OR2_X1 U19458 ( .A1(n16465), .A2(n19424), .ZN(n16378) );
  XNOR2_X1 U19459 ( .A(n15837), .B(n16455), .ZN(n16462) );
  AOI22_X1 U19460 ( .A1(n16462), .A2(n16449), .B1(n19428), .B2(n16461), .ZN(
        n16377) );
  AND2_X1 U19461 ( .A1(n16378), .A2(n16377), .ZN(n16379) );
  OAI211_X1 U19462 ( .C1(n16381), .C2(n16453), .A(n16380), .B(n16379), .ZN(
        P2_U2999) );
  AOI22_X1 U19463 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19421), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19420), .ZN(n16386) );
  OAI22_X1 U19464 ( .A1(n16383), .A2(n19424), .B1(n19423), .B2(n16382), .ZN(
        n16384) );
  AOI21_X1 U19465 ( .B1(n19428), .B2(n19209), .A(n16384), .ZN(n16385) );
  OAI211_X1 U19466 ( .C1(n19432), .C2(n19207), .A(n16386), .B(n16385), .ZN(
        P2_U3000) );
  AOI22_X1 U19467 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19420), .B1(n16440), 
        .B2(n19215), .ZN(n16398) );
  OAI21_X1 U19468 ( .B1(n16413), .B2(n16387), .A(n16468), .ZN(n16389) );
  NAND2_X1 U19469 ( .A1(n16389), .A2(n16388), .ZN(n16473) );
  NAND2_X1 U19470 ( .A1(n16391), .A2(n16390), .ZN(n16392) );
  XNOR2_X1 U19471 ( .A(n16393), .B(n16392), .ZN(n16477) );
  OR2_X1 U19472 ( .A1(n16477), .A2(n19424), .ZN(n16395) );
  NAND2_X1 U19473 ( .A1(n19220), .A2(n19428), .ZN(n16394) );
  OAI211_X1 U19474 ( .C1(n16473), .C2(n19423), .A(n16395), .B(n16394), .ZN(
        n16396) );
  INV_X1 U19475 ( .A(n16396), .ZN(n16397) );
  OAI211_X1 U19476 ( .C1(n16399), .C2(n16453), .A(n16398), .B(n16397), .ZN(
        P2_U3001) );
  AOI22_X1 U19477 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19421), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19420), .ZN(n16404) );
  OAI22_X1 U19478 ( .A1(n16401), .A2(n19423), .B1(n16400), .B2(n19424), .ZN(
        n16402) );
  AOI21_X1 U19479 ( .B1(n19428), .B2(n19230), .A(n16402), .ZN(n16403) );
  OAI211_X1 U19480 ( .C1(n19432), .C2(n19228), .A(n16404), .B(n16403), .ZN(
        P2_U3002) );
  AOI22_X1 U19481 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19420), .B1(n16440), 
        .B2(n16405), .ZN(n16417) );
  NOR2_X1 U19482 ( .A1(n9729), .A2(n16406), .ZN(n16410) );
  NOR2_X1 U19483 ( .A1(n16408), .A2(n16407), .ZN(n16409) );
  XNOR2_X1 U19484 ( .A(n16410), .B(n16409), .ZN(n16485) );
  INV_X1 U19485 ( .A(n16411), .ZN(n16484) );
  AOI21_X1 U19486 ( .B1(n16412), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16415) );
  INV_X1 U19487 ( .A(n16413), .ZN(n16414) );
  NOR2_X1 U19488 ( .A1(n16415), .A2(n16414), .ZN(n16483) );
  AOI222_X1 U19489 ( .A1(n16485), .A2(n16450), .B1(n19428), .B2(n16484), .C1(
        n16449), .C2(n16483), .ZN(n16416) );
  OAI211_X1 U19490 ( .C1(n16418), .C2(n16453), .A(n16417), .B(n16416), .ZN(
        P2_U3003) );
  AOI22_X1 U19491 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19421), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19420), .ZN(n16423) );
  OAI22_X1 U19492 ( .A1(n16420), .A2(n19423), .B1(n16419), .B2(n19424), .ZN(
        n16421) );
  AOI21_X1 U19493 ( .B1(n19428), .B2(n9761), .A(n16421), .ZN(n16422) );
  OAI211_X1 U19494 ( .C1(n19432), .C2(n19239), .A(n16423), .B(n16422), .ZN(
        P2_U3004) );
  AOI22_X1 U19495 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19420), .B1(n16440), 
        .B2(n16424), .ZN(n16429) );
  AOI222_X1 U19496 ( .A1(n16427), .A2(n16449), .B1(n16450), .B2(n16426), .C1(
        n19428), .C2(n16425), .ZN(n16428) );
  OAI211_X1 U19497 ( .C1(n16430), .C2(n16453), .A(n16429), .B(n16428), .ZN(
        P2_U3005) );
  AOI22_X1 U19498 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19420), .B1(n16440), 
        .B2(n19258), .ZN(n16437) );
  NAND2_X1 U19499 ( .A1(n16431), .A2(n16449), .ZN(n16433) );
  NAND2_X1 U19500 ( .A1(n19263), .A2(n19428), .ZN(n16432) );
  OAI211_X1 U19501 ( .C1(n16434), .C2(n19424), .A(n16433), .B(n16432), .ZN(
        n16435) );
  INV_X1 U19502 ( .A(n16435), .ZN(n16436) );
  OAI211_X1 U19503 ( .C1(n16438), .C2(n16453), .A(n16437), .B(n16436), .ZN(
        P2_U3007) );
  AOI22_X1 U19504 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19420), .B1(n16440), 
        .B2(n16439), .ZN(n16452) );
  XOR2_X1 U19505 ( .A(n16442), .B(n16441), .Z(n16504) );
  INV_X1 U19506 ( .A(n16443), .ZN(n16447) );
  AOI21_X1 U19507 ( .B1(n11176), .B2(n16445), .A(n16444), .ZN(n16446) );
  AOI21_X1 U19508 ( .B1(n16447), .B2(n11176), .A(n16446), .ZN(n16503) );
  INV_X1 U19509 ( .A(n16448), .ZN(n16502) );
  AOI222_X1 U19510 ( .A1(n16504), .A2(n16450), .B1(n16503), .B2(n16449), .C1(
        n19428), .C2(n16502), .ZN(n16451) );
  OAI211_X1 U19511 ( .C1(n16454), .C2(n16453), .A(n16452), .B(n16451), .ZN(
        P2_U3009) );
  NAND2_X1 U19512 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19420), .ZN(n16458) );
  NAND2_X1 U19513 ( .A1(n16456), .A2(n16455), .ZN(n16457) );
  OAI211_X1 U19514 ( .C1(n16526), .C2(n19337), .A(n16458), .B(n16457), .ZN(
        n16459) );
  AOI21_X1 U19515 ( .B1(n16460), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16459), .ZN(n16464) );
  AOI22_X1 U19516 ( .A1(n16462), .A2(n19438), .B1(n19440), .B2(n16461), .ZN(
        n16463) );
  OAI211_X1 U19517 ( .C1(n16465), .C2(n19449), .A(n16464), .B(n16463), .ZN(
        P2_U3031) );
  NOR2_X1 U19518 ( .A1(n16466), .A2(n11095), .ZN(n16471) );
  OAI22_X1 U19519 ( .A1(n16469), .A2(n16468), .B1(n16387), .B2(n16467), .ZN(
        n16470) );
  AOI211_X1 U19520 ( .C1(n19436), .C2(n19219), .A(n16471), .B(n16470), .ZN(
        n16476) );
  OAI22_X1 U19521 ( .A1(n16473), .A2(n16524), .B1(n16527), .B2(n16472), .ZN(
        n16474) );
  INV_X1 U19522 ( .A(n16474), .ZN(n16475) );
  OAI211_X1 U19523 ( .C1(n19449), .C2(n16477), .A(n16476), .B(n16475), .ZN(
        P2_U3033) );
  AOI211_X1 U19524 ( .C1(n15867), .C2(n16488), .A(n16479), .B(n16478), .ZN(
        n16482) );
  NAND2_X1 U19525 ( .A1(n19436), .A2(n19345), .ZN(n16480) );
  OAI21_X1 U19526 ( .B1(n11064), .B2(n19178), .A(n16480), .ZN(n16481) );
  NOR2_X1 U19527 ( .A1(n16482), .A2(n16481), .ZN(n16487) );
  AOI222_X1 U19528 ( .A1(n16485), .A2(n16519), .B1(n19440), .B2(n16484), .C1(
        n19438), .C2(n16483), .ZN(n16486) );
  OAI211_X1 U19529 ( .C1(n16489), .C2(n16488), .A(n16487), .B(n16486), .ZN(
        P2_U3035) );
  NAND2_X1 U19530 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16490) );
  OAI211_X1 U19531 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16491), .B(n16490), .ZN(n16494) );
  INV_X1 U19532 ( .A(n19255), .ZN(n16492) );
  AOI22_X1 U19533 ( .A1(n19436), .A2(n16492), .B1(n19420), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n16493) );
  NAND2_X1 U19534 ( .A1(n16494), .A2(n16493), .ZN(n16495) );
  AOI21_X1 U19535 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16496), .A(
        n16495), .ZN(n16499) );
  AOI22_X1 U19536 ( .A1(n16497), .A2(n19438), .B1(n19440), .B2(n19251), .ZN(
        n16498) );
  OAI211_X1 U19537 ( .C1(n16500), .C2(n19449), .A(n16499), .B(n16498), .ZN(
        P2_U3038) );
  AOI22_X1 U19538 ( .A1(n16501), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19436), .B2(n19354), .ZN(n16511) );
  AOI222_X1 U19539 ( .A1(n16504), .A2(n16519), .B1(n16503), .B2(n19438), .C1(
        n19440), .C2(n16502), .ZN(n16510) );
  NAND2_X1 U19540 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19420), .ZN(n16509) );
  OAI221_X1 U19541 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n16507), .C2(n16506), .A(
        n16505), .ZN(n16508) );
  NAND4_X1 U19542 ( .A1(n16511), .A2(n16510), .A3(n16509), .A4(n16508), .ZN(
        P2_U3041) );
  NOR2_X1 U19543 ( .A1(n16512), .A2(n16527), .ZN(n16513) );
  AOI211_X1 U19544 ( .C1(n19436), .C2(n19361), .A(n16514), .B(n16513), .ZN(
        n16515) );
  OAI21_X1 U19545 ( .B1(n16516), .B2(n16524), .A(n16515), .ZN(n16517) );
  AOI21_X1 U19546 ( .B1(n16519), .B2(n16518), .A(n16517), .ZN(n16520) );
  OAI221_X1 U19547 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16523), .C1(
        n16522), .C2(n16521), .A(n16520), .ZN(P2_U3043) );
  OAI22_X1 U19548 ( .A1(n16526), .A2(n19314), .B1(n16525), .B2(n16524), .ZN(
        n16529) );
  OAI22_X1 U19549 ( .A1(n16527), .A2(n19321), .B1(n19442), .B2(n10375), .ZN(
        n16528) );
  AOI211_X1 U19550 ( .C1(n10375), .C2(n19434), .A(n16529), .B(n16528), .ZN(
        n16531) );
  OAI211_X1 U19551 ( .C1(n19449), .C2(n16532), .A(n16531), .B(n16530), .ZN(
        P2_U3046) );
  AOI21_X1 U19552 ( .B1(n20029), .B2(n16534), .A(n16533), .ZN(n16547) );
  INV_X1 U19553 ( .A(n20140), .ZN(n16536) );
  AOI22_X1 U19554 ( .A1(n16538), .A2(n16537), .B1(n16536), .B2(n16535), .ZN(
        n16546) );
  NAND2_X1 U19555 ( .A1(n16539), .A2(n19884), .ZN(n16543) );
  NAND2_X1 U19556 ( .A1(n16540), .A2(n20029), .ZN(n16541) );
  MUX2_X1 U19557 ( .A(n16541), .B(n16540), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16542) );
  OAI21_X1 U19558 ( .B1(n16544), .B2(n16543), .A(n16542), .ZN(n16545) );
  NAND3_X1 U19559 ( .A1(n16547), .A2(n16546), .A3(n16545), .ZN(P2_U3176) );
  INV_X1 U19560 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16764) );
  XNOR2_X1 U19561 ( .A(n16764), .B(n16567), .ZN(n16763) );
  OAI221_X1 U19562 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16550), .C1(
        n16764), .C2(n16549), .A(n16548), .ZN(n16551) );
  AOI21_X1 U19563 ( .B1(n17927), .B2(n16763), .A(n16551), .ZN(n16556) );
  OAI22_X1 U19565 ( .A1(n16558), .A2(n18080), .B1(n16561), .B2(n17986), .ZN(
        n16554) );
  OAI22_X2 U19566 ( .A1(n18080), .A2(n18274), .B1(n17986), .B2(n18276), .ZN(
        n17944) );
  NAND2_X1 U19567 ( .A1(n17944), .A2(n17863), .ZN(n17875) );
  NOR2_X1 U19568 ( .A1(n18135), .A2(n17875), .ZN(n17768) );
  INV_X1 U19569 ( .A(n17768), .ZN(n17787) );
  NOR2_X1 U19570 ( .A1(n16552), .A2(n17787), .ZN(n17736) );
  AOI22_X1 U19571 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16554), .B1(
        n16553), .B2(n17736), .ZN(n16555) );
  OAI211_X1 U19572 ( .C1(n17991), .C2(n16557), .A(n16556), .B(n16555), .ZN(
        P3_U2800) );
  NAND2_X1 U19573 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16560) );
  NOR2_X1 U19574 ( .A1(n18087), .A2(n16560), .ZN(n16597) );
  INV_X1 U19575 ( .A(n16597), .ZN(n16559) );
  AOI211_X1 U19576 ( .C1(n16563), .C2(n16559), .A(n16558), .B(n18080), .ZN(
        n16565) );
  NOR2_X1 U19577 ( .A1(n16560), .A2(n18090), .ZN(n16595) );
  INV_X1 U19578 ( .A(n16595), .ZN(n16562) );
  AOI211_X1 U19579 ( .C1(n16563), .C2(n16562), .A(n16561), .B(n17986), .ZN(
        n16564) );
  AOI211_X1 U19580 ( .C1(n17973), .C2(n16566), .A(n16565), .B(n16564), .ZN(
        n16574) );
  AOI21_X1 U19581 ( .B1(n9968), .B2(n16568), .A(n16567), .ZN(n16773) );
  OAI21_X1 U19582 ( .B1(n16569), .B2(n17927), .A(n16773), .ZN(n16572) );
  OAI221_X1 U19583 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n9777), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18798), .A(n16570), .ZN(
        n16571) );
  NAND4_X1 U19584 ( .A1(n16574), .A2(n16573), .A3(n16572), .A4(n16571), .ZN(
        P3_U2801) );
  NOR2_X1 U19585 ( .A1(n18399), .A2(n18345), .ZN(n18308) );
  INV_X1 U19586 ( .A(n18308), .ZN(n18384) );
  OAI211_X1 U19587 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18384), .A(
        n16575), .B(n18383), .ZN(n16581) );
  NAND3_X1 U19588 ( .A1(n18382), .A2(n18081), .A3(n18104), .ZN(n16576) );
  NOR4_X1 U19589 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16578), .A3(
        n16577), .A4(n16576), .ZN(n16579) );
  AOI211_X1 U19590 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16581), .A(
        n16580), .B(n16579), .ZN(n16585) );
  INV_X1 U19591 ( .A(n18310), .ZN(n18116) );
  AOI22_X1 U19592 ( .A1(n16583), .A2(n18116), .B1(n16582), .B2(n18299), .ZN(
        n16584) );
  OAI211_X1 U19593 ( .C1(n16586), .C2(n18374), .A(n16585), .B(n16584), .ZN(
        P3_U2831) );
  NAND4_X1 U19594 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17955), .A3(
        n16588), .A4(n16587), .ZN(n16602) );
  INV_X1 U19595 ( .A(n18398), .ZN(n18391) );
  NOR2_X1 U19596 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16589), .ZN(
        n17717) );
  INV_X1 U19597 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19010) );
  NOR2_X1 U19598 ( .A1(n9655), .A2(n19010), .ZN(n17716) );
  NOR3_X1 U19599 ( .A1(n17721), .A2(n17725), .A3(n18312), .ZN(n16590) );
  AOI211_X1 U19600 ( .C1(n16591), .C2(n17717), .A(n17716), .B(n16590), .ZN(
        n16601) );
  NAND3_X1 U19601 ( .A1(n17955), .A2(n17726), .A3(n17725), .ZN(n17727) );
  NAND2_X1 U19602 ( .A1(n17725), .A2(n17727), .ZN(n17720) );
  NAND2_X1 U19603 ( .A1(n17721), .A2(n17720), .ZN(n17719) );
  NAND2_X1 U19604 ( .A1(n16592), .A2(n17719), .ZN(n16593) );
  AOI221_X1 U19605 ( .B1(n17565), .B2(n16595), .C1(n16594), .C2(n16593), .A(
        n18858), .ZN(n16599) );
  OAI211_X1 U19606 ( .C1(n16597), .C2(n18249), .A(n18382), .B(n16596), .ZN(
        n16598) );
  OAI211_X1 U19607 ( .C1(n16599), .C2(n16598), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n9655), .ZN(n16600) );
  OAI211_X1 U19608 ( .C1(n16602), .C2(n18391), .A(n16601), .B(n16600), .ZN(
        P3_U2834) );
  NOR3_X1 U19609 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16604) );
  NOR4_X1 U19610 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16603) );
  INV_X2 U19611 ( .A(n16698), .ZN(U215) );
  NAND4_X1 U19612 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16604), .A3(n16603), .A4(
        U215), .ZN(U213) );
  INV_X1 U19613 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16700) );
  INV_X2 U19614 ( .A(U214), .ZN(n16661) );
  INV_X1 U19615 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16701) );
  OAI222_X1 U19616 ( .A1(U212), .A2(n16700), .B1(n16663), .B2(n19497), .C1(
        U214), .C2(n16701), .ZN(U216) );
  AOI22_X1 U19617 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16660), .ZN(n16606) );
  OAI21_X1 U19618 ( .B1(n16607), .B2(n16663), .A(n16606), .ZN(U217) );
  AOI22_X1 U19619 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16660), .ZN(n16608) );
  OAI21_X1 U19620 ( .B1(n16609), .B2(n16663), .A(n16608), .ZN(U218) );
  AOI22_X1 U19621 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16660), .ZN(n16610) );
  OAI21_X1 U19622 ( .B1(n19479), .B2(n16663), .A(n16610), .ZN(U219) );
  AOI22_X1 U19623 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16660), .ZN(n16611) );
  OAI21_X1 U19624 ( .B1(n16612), .B2(n16663), .A(n16611), .ZN(U220) );
  AOI22_X1 U19625 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16660), .ZN(n16613) );
  OAI21_X1 U19626 ( .B1(n16614), .B2(n16663), .A(n16613), .ZN(U221) );
  AOI22_X1 U19627 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16660), .ZN(n16615) );
  OAI21_X1 U19628 ( .B1(n16616), .B2(n16663), .A(n16615), .ZN(U222) );
  AOI22_X1 U19629 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16660), .ZN(n16617) );
  OAI21_X1 U19630 ( .B1(n16618), .B2(n16663), .A(n16617), .ZN(U223) );
  AOI22_X1 U19631 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16660), .ZN(n16619) );
  OAI21_X1 U19632 ( .B1(n16620), .B2(n16663), .A(n16619), .ZN(U224) );
  AOI22_X1 U19633 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16660), .ZN(n16621) );
  OAI21_X1 U19634 ( .B1(n16622), .B2(n16663), .A(n16621), .ZN(U225) );
  AOI22_X1 U19635 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16660), .ZN(n16623) );
  OAI21_X1 U19636 ( .B1(n19484), .B2(n16663), .A(n16623), .ZN(U226) );
  AOI22_X1 U19637 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16660), .ZN(n16624) );
  OAI21_X1 U19638 ( .B1(n16625), .B2(n16663), .A(n16624), .ZN(U227) );
  AOI22_X1 U19639 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16660), .ZN(n16626) );
  OAI21_X1 U19640 ( .B1(n16627), .B2(n16663), .A(n16626), .ZN(U228) );
  AOI22_X1 U19641 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16660), .ZN(n16628) );
  OAI21_X1 U19642 ( .B1(n16629), .B2(n16663), .A(n16628), .ZN(U229) );
  AOI22_X1 U19643 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16660), .ZN(n16630) );
  OAI21_X1 U19644 ( .B1(n16631), .B2(n16663), .A(n16630), .ZN(U230) );
  AOI22_X1 U19645 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16660), .ZN(n16632) );
  OAI21_X1 U19646 ( .B1(n16633), .B2(n16663), .A(n16632), .ZN(U231) );
  AOI22_X1 U19647 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16660), .ZN(n16634) );
  OAI21_X1 U19648 ( .B1(n13297), .B2(n16663), .A(n16634), .ZN(U232) );
  AOI22_X1 U19649 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16660), .ZN(n16635) );
  OAI21_X1 U19650 ( .B1(n16636), .B2(n16663), .A(n16635), .ZN(U233) );
  AOI22_X1 U19651 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16660), .ZN(n16637) );
  OAI21_X1 U19652 ( .B1(n16638), .B2(n16663), .A(n16637), .ZN(U234) );
  INV_X1 U19653 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16640) );
  AOI22_X1 U19654 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16660), .ZN(n16639) );
  OAI21_X1 U19655 ( .B1(n16640), .B2(n16663), .A(n16639), .ZN(U235) );
  AOI22_X1 U19656 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16660), .ZN(n16641) );
  OAI21_X1 U19657 ( .B1(n13183), .B2(n16663), .A(n16641), .ZN(U236) );
  AOI22_X1 U19658 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16660), .ZN(n16642) );
  OAI21_X1 U19659 ( .B1(n16643), .B2(n16663), .A(n16642), .ZN(U237) );
  AOI22_X1 U19660 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16660), .ZN(n16644) );
  OAI21_X1 U19661 ( .B1(n16645), .B2(n16663), .A(n16644), .ZN(U238) );
  AOI22_X1 U19662 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16660), .ZN(n16646) );
  OAI21_X1 U19663 ( .B1(n13165), .B2(n16663), .A(n16646), .ZN(U239) );
  AOI22_X1 U19664 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16660), .ZN(n16647) );
  OAI21_X1 U19665 ( .B1(n13160), .B2(n16663), .A(n16647), .ZN(U240) );
  INV_X1 U19666 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16649) );
  AOI22_X1 U19667 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16660), .ZN(n16648) );
  OAI21_X1 U19668 ( .B1(n16649), .B2(n16663), .A(n16648), .ZN(U241) );
  INV_X1 U19669 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16651) );
  AOI22_X1 U19670 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16660), .ZN(n16650) );
  OAI21_X1 U19671 ( .B1(n16651), .B2(n16663), .A(n16650), .ZN(U242) );
  AOI22_X1 U19672 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16660), .ZN(n16652) );
  OAI21_X1 U19673 ( .B1(n16653), .B2(n16663), .A(n16652), .ZN(U243) );
  INV_X1 U19674 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16655) );
  AOI22_X1 U19675 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16660), .ZN(n16654) );
  OAI21_X1 U19676 ( .B1(n16655), .B2(n16663), .A(n16654), .ZN(U244) );
  INV_X1 U19677 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16657) );
  AOI22_X1 U19678 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16660), .ZN(n16656) );
  OAI21_X1 U19679 ( .B1(n16657), .B2(n16663), .A(n16656), .ZN(U245) );
  INV_X1 U19680 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16659) );
  AOI22_X1 U19681 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16660), .ZN(n16658) );
  OAI21_X1 U19682 ( .B1(n16659), .B2(n16663), .A(n16658), .ZN(U246) );
  INV_X1 U19683 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16664) );
  AOI22_X1 U19684 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16661), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16660), .ZN(n16662) );
  OAI21_X1 U19685 ( .B1(n16664), .B2(n16663), .A(n16662), .ZN(U247) );
  OAI22_X1 U19686 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16698), .ZN(n16665) );
  INV_X1 U19687 ( .A(n16665), .ZN(U251) );
  OAI22_X1 U19688 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16698), .ZN(n16666) );
  INV_X1 U19689 ( .A(n16666), .ZN(U252) );
  OAI22_X1 U19690 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16698), .ZN(n16667) );
  INV_X1 U19691 ( .A(n16667), .ZN(U253) );
  OAI22_X1 U19692 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16698), .ZN(n16668) );
  INV_X1 U19693 ( .A(n16668), .ZN(U254) );
  OAI22_X1 U19694 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16698), .ZN(n16669) );
  INV_X1 U19695 ( .A(n16669), .ZN(U255) );
  OAI22_X1 U19696 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16698), .ZN(n16670) );
  INV_X1 U19697 ( .A(n16670), .ZN(U256) );
  OAI22_X1 U19698 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16698), .ZN(n16671) );
  INV_X1 U19699 ( .A(n16671), .ZN(U257) );
  OAI22_X1 U19700 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16698), .ZN(n16672) );
  INV_X1 U19701 ( .A(n16672), .ZN(U258) );
  OAI22_X1 U19702 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16698), .ZN(n16673) );
  INV_X1 U19703 ( .A(n16673), .ZN(U259) );
  OAI22_X1 U19704 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16692), .ZN(n16674) );
  INV_X1 U19705 ( .A(n16674), .ZN(U260) );
  OAI22_X1 U19706 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16692), .ZN(n16675) );
  INV_X1 U19707 ( .A(n16675), .ZN(U261) );
  OAI22_X1 U19708 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16698), .ZN(n16676) );
  INV_X1 U19709 ( .A(n16676), .ZN(U262) );
  OAI22_X1 U19710 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16698), .ZN(n16677) );
  INV_X1 U19711 ( .A(n16677), .ZN(U263) );
  OAI22_X1 U19712 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16698), .ZN(n16678) );
  INV_X1 U19713 ( .A(n16678), .ZN(U264) );
  OAI22_X1 U19714 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16698), .ZN(n16679) );
  INV_X1 U19715 ( .A(n16679), .ZN(U265) );
  OAI22_X1 U19716 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16692), .ZN(n16680) );
  INV_X1 U19717 ( .A(n16680), .ZN(U266) );
  OAI22_X1 U19718 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16692), .ZN(n16681) );
  INV_X1 U19719 ( .A(n16681), .ZN(U267) );
  OAI22_X1 U19720 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16692), .ZN(n16682) );
  INV_X1 U19721 ( .A(n16682), .ZN(U268) );
  OAI22_X1 U19722 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16692), .ZN(n16683) );
  INV_X1 U19723 ( .A(n16683), .ZN(U269) );
  OAI22_X1 U19724 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16692), .ZN(n16684) );
  INV_X1 U19725 ( .A(n16684), .ZN(U270) );
  OAI22_X1 U19726 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16692), .ZN(n16685) );
  INV_X1 U19727 ( .A(n16685), .ZN(U271) );
  OAI22_X1 U19728 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16698), .ZN(n16686) );
  INV_X1 U19729 ( .A(n16686), .ZN(U272) );
  OAI22_X1 U19730 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16698), .ZN(n16687) );
  INV_X1 U19731 ( .A(n16687), .ZN(U273) );
  OAI22_X1 U19732 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16692), .ZN(n16688) );
  INV_X1 U19733 ( .A(n16688), .ZN(U274) );
  OAI22_X1 U19734 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16698), .ZN(n16689) );
  INV_X1 U19735 ( .A(n16689), .ZN(U275) );
  OAI22_X1 U19736 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16698), .ZN(n16690) );
  INV_X1 U19737 ( .A(n16690), .ZN(U276) );
  OAI22_X1 U19738 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16698), .ZN(n16691) );
  INV_X1 U19739 ( .A(n16691), .ZN(U277) );
  OAI22_X1 U19740 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16692), .ZN(n16693) );
  INV_X1 U19741 ( .A(n16693), .ZN(U278) );
  OAI22_X1 U19742 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16698), .ZN(n16694) );
  INV_X1 U19743 ( .A(n16694), .ZN(U279) );
  OAI22_X1 U19744 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16698), .ZN(n16695) );
  INV_X1 U19745 ( .A(n16695), .ZN(U280) );
  OAI22_X1 U19746 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16698), .ZN(n16697) );
  INV_X1 U19747 ( .A(n16697), .ZN(U281) );
  INV_X1 U19748 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19495) );
  AOI22_X1 U19749 ( .A1(n16698), .A2(n16700), .B1(n19495), .B2(U215), .ZN(U282) );
  INV_X1 U19750 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16699) );
  AOI222_X1 U19751 ( .A1(n16701), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16700), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16699), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16702) );
  INV_X2 U19752 ( .A(n16704), .ZN(n16703) );
  INV_X1 U19753 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18974) );
  INV_X1 U19754 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20056) );
  AOI22_X1 U19755 ( .A1(n16703), .A2(n18974), .B1(n20056), .B2(n16704), .ZN(
        U347) );
  INV_X1 U19756 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18972) );
  INV_X1 U19757 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20055) );
  AOI22_X1 U19758 ( .A1(n16703), .A2(n18972), .B1(n20055), .B2(n16704), .ZN(
        U348) );
  INV_X1 U19759 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18969) );
  INV_X1 U19760 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20054) );
  AOI22_X1 U19761 ( .A1(n16703), .A2(n18969), .B1(n20054), .B2(n16704), .ZN(
        U349) );
  INV_X1 U19762 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18968) );
  INV_X1 U19763 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20053) );
  AOI22_X1 U19764 ( .A1(n16703), .A2(n18968), .B1(n20053), .B2(n16704), .ZN(
        U350) );
  INV_X1 U19765 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18966) );
  INV_X1 U19766 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20052) );
  AOI22_X1 U19767 ( .A1(n16703), .A2(n18966), .B1(n20052), .B2(n16704), .ZN(
        U351) );
  INV_X1 U19768 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18963) );
  INV_X1 U19769 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20051) );
  AOI22_X1 U19770 ( .A1(n16703), .A2(n18963), .B1(n20051), .B2(n16704), .ZN(
        U352) );
  INV_X1 U19771 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18962) );
  INV_X1 U19772 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20050) );
  AOI22_X1 U19773 ( .A1(n16703), .A2(n18962), .B1(n20050), .B2(n16704), .ZN(
        U353) );
  INV_X1 U19774 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18960) );
  AOI22_X1 U19775 ( .A1(n16703), .A2(n18960), .B1(n20049), .B2(n16704), .ZN(
        U354) );
  INV_X1 U19776 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19012) );
  INV_X1 U19777 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20085) );
  AOI22_X1 U19778 ( .A1(n16703), .A2(n19012), .B1(n20085), .B2(n16704), .ZN(
        U356) );
  INV_X1 U19779 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19009) );
  INV_X1 U19780 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20084) );
  AOI22_X1 U19781 ( .A1(n16703), .A2(n19009), .B1(n20084), .B2(n16704), .ZN(
        U357) );
  INV_X1 U19782 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19008) );
  INV_X1 U19783 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20081) );
  AOI22_X1 U19784 ( .A1(n16703), .A2(n19008), .B1(n20081), .B2(n16704), .ZN(
        U358) );
  INV_X1 U19785 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19006) );
  INV_X1 U19786 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20080) );
  AOI22_X1 U19787 ( .A1(n16703), .A2(n19006), .B1(n20080), .B2(n16704), .ZN(
        U359) );
  INV_X1 U19788 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19004) );
  INV_X1 U19789 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20078) );
  AOI22_X1 U19790 ( .A1(n16703), .A2(n19004), .B1(n20078), .B2(n16704), .ZN(
        U360) );
  INV_X1 U19791 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19002) );
  INV_X1 U19792 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20077) );
  AOI22_X1 U19793 ( .A1(n16703), .A2(n19002), .B1(n20077), .B2(n16704), .ZN(
        U361) );
  INV_X1 U19794 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18999) );
  INV_X1 U19795 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20075) );
  AOI22_X1 U19796 ( .A1(n16703), .A2(n18999), .B1(n20075), .B2(n16704), .ZN(
        U362) );
  INV_X1 U19797 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18998) );
  INV_X1 U19798 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20073) );
  AOI22_X1 U19799 ( .A1(n16703), .A2(n18998), .B1(n20073), .B2(n16704), .ZN(
        U363) );
  INV_X1 U19800 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18995) );
  INV_X1 U19801 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20071) );
  AOI22_X1 U19802 ( .A1(n16703), .A2(n18995), .B1(n20071), .B2(n16704), .ZN(
        U364) );
  INV_X1 U19803 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18958) );
  INV_X1 U19804 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20048) );
  AOI22_X1 U19805 ( .A1(n16703), .A2(n18958), .B1(n20048), .B2(n16704), .ZN(
        U365) );
  INV_X1 U19806 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18994) );
  INV_X1 U19807 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20069) );
  AOI22_X1 U19808 ( .A1(n16703), .A2(n18994), .B1(n20069), .B2(n16704), .ZN(
        U366) );
  INV_X1 U19809 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18992) );
  INV_X1 U19810 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20067) );
  AOI22_X1 U19811 ( .A1(n16703), .A2(n18992), .B1(n20067), .B2(n16704), .ZN(
        U367) );
  INV_X1 U19812 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18990) );
  INV_X1 U19813 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20066) );
  AOI22_X1 U19814 ( .A1(n16703), .A2(n18990), .B1(n20066), .B2(n16704), .ZN(
        U368) );
  INV_X1 U19815 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18987) );
  INV_X1 U19816 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20064) );
  AOI22_X1 U19817 ( .A1(n16703), .A2(n18987), .B1(n20064), .B2(n16704), .ZN(
        U369) );
  INV_X1 U19818 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18986) );
  INV_X1 U19819 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20063) );
  AOI22_X1 U19820 ( .A1(n16703), .A2(n18986), .B1(n20063), .B2(n16704), .ZN(
        U370) );
  INV_X1 U19821 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18984) );
  INV_X1 U19822 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20061) );
  AOI22_X1 U19823 ( .A1(n16703), .A2(n18984), .B1(n20061), .B2(n16704), .ZN(
        U371) );
  INV_X1 U19824 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18981) );
  INV_X1 U19825 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20060) );
  AOI22_X1 U19826 ( .A1(n16703), .A2(n18981), .B1(n20060), .B2(n16704), .ZN(
        U372) );
  INV_X1 U19827 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18980) );
  INV_X1 U19828 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20059) );
  AOI22_X1 U19829 ( .A1(n16703), .A2(n18980), .B1(n20059), .B2(n16704), .ZN(
        U373) );
  INV_X1 U19830 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18978) );
  INV_X1 U19831 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20058) );
  AOI22_X1 U19832 ( .A1(n16703), .A2(n18978), .B1(n20058), .B2(n16704), .ZN(
        U374) );
  INV_X1 U19833 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18976) );
  INV_X1 U19834 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U19835 ( .A1(n16703), .A2(n18976), .B1(n20057), .B2(n16704), .ZN(
        U375) );
  INV_X1 U19836 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18955) );
  INV_X1 U19837 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U19838 ( .A1(n16703), .A2(n18955), .B1(n20047), .B2(n16704), .ZN(
        U376) );
  INV_X1 U19839 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18954) );
  NAND2_X1 U19840 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18954), .ZN(n18946) );
  AOI22_X1 U19841 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18946), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18952), .ZN(n19025) );
  AOI21_X1 U19842 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19025), .ZN(n16705) );
  INV_X1 U19843 ( .A(n16705), .ZN(P3_U2633) );
  OAI21_X1 U19844 ( .B1(n16712), .B2(n17638), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16706) );
  OAI21_X1 U19845 ( .B1(n16707), .B2(n18929), .A(n16706), .ZN(P3_U2634) );
  AOI21_X1 U19846 ( .B1(n18952), .B2(n18954), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16708) );
  AOI22_X1 U19847 ( .A1(n19083), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16708), 
        .B2(n19084), .ZN(P3_U2635) );
  NOR2_X1 U19848 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18939) );
  OAI21_X1 U19849 ( .B1(n18939), .B2(BS16), .A(n19025), .ZN(n19023) );
  OAI21_X1 U19850 ( .B1(n19025), .B2(n19073), .A(n19023), .ZN(P3_U2636) );
  INV_X1 U19851 ( .A(n16709), .ZN(n16711) );
  NOR3_X1 U19852 ( .A1(n16712), .A2(n16711), .A3(n16710), .ZN(n18859) );
  NOR2_X1 U19853 ( .A1(n18859), .A2(n18924), .ZN(n19065) );
  OAI21_X1 U19854 ( .B1(n19065), .B2(n18404), .A(n16713), .ZN(P3_U2637) );
  NOR4_X1 U19855 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16717) );
  NOR4_X1 U19856 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16716) );
  NOR4_X1 U19857 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16715) );
  NOR4_X1 U19858 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16714) );
  NAND4_X1 U19859 ( .A1(n16717), .A2(n16716), .A3(n16715), .A4(n16714), .ZN(
        n16723) );
  NOR4_X1 U19860 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16721) );
  AOI211_X1 U19861 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16720) );
  NOR4_X1 U19862 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16719) );
  NOR4_X1 U19863 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16718) );
  NAND4_X1 U19864 ( .A1(n16721), .A2(n16720), .A3(n16719), .A4(n16718), .ZN(
        n16722) );
  NOR2_X1 U19865 ( .A1(n16723), .A2(n16722), .ZN(n19063) );
  INV_X1 U19866 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16725) );
  NOR3_X1 U19867 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16726) );
  OAI21_X1 U19868 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16726), .A(n19063), .ZN(
        n16724) );
  OAI21_X1 U19869 ( .B1(n19063), .B2(n16725), .A(n16724), .ZN(P3_U2638) );
  INV_X1 U19870 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18956) );
  INV_X1 U19871 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19024) );
  AOI21_X1 U19872 ( .B1(n18956), .B2(n19024), .A(n16726), .ZN(n16728) );
  INV_X1 U19873 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16727) );
  INV_X1 U19874 ( .A(n19063), .ZN(n19060) );
  AOI22_X1 U19875 ( .A1(n19063), .A2(n16728), .B1(n16727), .B2(n19060), .ZN(
        P3_U2639) );
  NAND4_X1 U19876 ( .A1(n19086), .A2(n18926), .A3(n19073), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18933) );
  NAND2_X1 U19877 ( .A1(n19086), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18792) );
  OR2_X1 U19878 ( .A1(n18929), .A2(n18792), .ZN(n18922) );
  INV_X1 U19879 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n17138) );
  OAI211_X1 U19880 ( .C1(n16733), .C2(n16732), .A(n19075), .B(n19073), .ZN(
        n18918) );
  OAI211_X2 U19881 ( .C1(n17138), .C2(n19074), .A(n18918), .B(n16737), .ZN(
        n17127) );
  INV_X1 U19882 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19016) );
  INV_X1 U19883 ( .A(n18918), .ZN(n16734) );
  INV_X1 U19884 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19001) );
  INV_X1 U19885 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19000) );
  INV_X1 U19886 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18996) );
  INV_X1 U19887 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18997) );
  INV_X1 U19888 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18982) );
  INV_X1 U19889 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18979) );
  INV_X1 U19890 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18975) );
  INV_X1 U19891 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18964) );
  INV_X1 U19892 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18957) );
  NOR2_X1 U19893 ( .A1(n18956), .A2(n18957), .ZN(n17104) );
  NAND2_X1 U19894 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17104), .ZN(n17064) );
  INV_X1 U19895 ( .A(n17064), .ZN(n17071) );
  NAND2_X1 U19896 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17071), .ZN(n17054) );
  NOR2_X1 U19897 ( .A1(n18964), .A2(n17054), .ZN(n17025) );
  NAND4_X1 U19898 ( .A1(n17025), .A2(P3_REIP_REG_8__SCAN_IN), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n16997) );
  NAND2_X1 U19899 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16979) );
  NOR3_X1 U19900 ( .A1(n18975), .A2(n16997), .A3(n16979), .ZN(n16975) );
  NAND2_X1 U19901 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16975), .ZN(n16945) );
  NOR3_X1 U19902 ( .A1(n18982), .A2(n18979), .A3(n16945), .ZN(n16882) );
  INV_X1 U19903 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18993) );
  NAND3_X1 U19904 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16883) );
  NAND2_X1 U19905 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16874) );
  NOR3_X1 U19906 ( .A1(n18993), .A2(n16883), .A3(n16874), .ZN(n16855) );
  NAND2_X1 U19907 ( .A1(n16882), .A2(n16855), .ZN(n16854) );
  NOR2_X1 U19908 ( .A1(n19000), .A2(n16845), .ZN(n16831) );
  INV_X1 U19909 ( .A(n16831), .ZN(n16816) );
  NOR2_X1 U19910 ( .A1(n19001), .A2(n16816), .ZN(n16803) );
  NAND3_X1 U19911 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16803), .ZN(n16750) );
  NOR2_X1 U19912 ( .A1(n17118), .A2(n16750), .ZN(n16782) );
  NAND4_X1 U19913 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16782), .ZN(n16753) );
  NOR3_X1 U19914 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19016), .A3(n16753), 
        .ZN(n16735) );
  AOI21_X1 U19915 ( .B1(n17116), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16735), .ZN(
        n16759) );
  NOR2_X1 U19916 ( .A1(n17138), .A2(n19074), .ZN(n16736) );
  OAI211_X2 U19917 ( .C1(P3_STATEBS16_REG_SCAN_IN), .C2(n18943), .A(n16737), 
        .B(n16736), .ZN(n17126) );
  NOR3_X1 U19918 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17107) );
  NAND2_X1 U19919 ( .A1(n17107), .A2(n17423), .ZN(n17090) );
  NOR2_X1 U19920 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17090), .ZN(n17063) );
  NAND2_X1 U19921 ( .A1(n17063), .A2(n17418), .ZN(n17057) );
  NAND2_X1 U19922 ( .A1(n17041), .A2(n17403), .ZN(n17031) );
  NAND2_X1 U19923 ( .A1(n17010), .A2(n17003), .ZN(n16994) );
  INV_X1 U19924 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17345) );
  NAND2_X1 U19925 ( .A1(n16993), .A2(n17345), .ZN(n16986) );
  NOR2_X1 U19926 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16986), .ZN(n16971) );
  INV_X1 U19927 ( .A(n16971), .ZN(n16955) );
  NAND2_X1 U19928 ( .A1(n16944), .A2(n16938), .ZN(n16934) );
  NAND2_X1 U19929 ( .A1(n16918), .A2(n16910), .ZN(n16909) );
  NAND2_X1 U19930 ( .A1(n16893), .A2(n17239), .ZN(n16890) );
  INV_X1 U19931 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17222) );
  NAND2_X1 U19932 ( .A1(n16872), .A2(n17222), .ZN(n16866) );
  INV_X1 U19933 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17186) );
  NAND2_X1 U19934 ( .A1(n16852), .A2(n17186), .ZN(n16848) );
  NOR2_X1 U19935 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16848), .ZN(n16819) );
  NAND2_X1 U19936 ( .A1(n16819), .A2(n16824), .ZN(n16805) );
  NOR2_X1 U19937 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16805), .ZN(n16804) );
  INV_X1 U19938 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16796) );
  NAND2_X1 U19939 ( .A1(n16804), .A2(n16796), .ZN(n16799) );
  NOR2_X1 U19940 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16799), .ZN(n16783) );
  INV_X1 U19941 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17136) );
  NAND2_X1 U19942 ( .A1(n16783), .A2(n17136), .ZN(n16761) );
  NOR2_X1 U19943 ( .A1(n17126), .A2(n16761), .ZN(n16768) );
  INV_X1 U19944 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16757) );
  INV_X1 U19945 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16739) );
  NOR2_X1 U19946 ( .A1(n18070), .A2(n17711), .ZN(n16741) );
  NAND2_X1 U19947 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16741), .ZN(
        n16740) );
  AOI21_X1 U19948 ( .B1(n16739), .B2(n16740), .A(n16738), .ZN(n17710) );
  OAI21_X1 U19949 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16741), .A(
        n16740), .ZN(n17730) );
  INV_X1 U19950 ( .A(n17730), .ZN(n16795) );
  NOR2_X1 U19951 ( .A1(n18070), .A2(n17795), .ZN(n16747) );
  INV_X1 U19952 ( .A(n16747), .ZN(n16748) );
  NOR2_X1 U19953 ( .A1(n17796), .A2(n16748), .ZN(n17779) );
  NAND2_X1 U19954 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17779), .ZN(
        n16744) );
  NOR2_X1 U19955 ( .A1(n17758), .A2(n16744), .ZN(n17708) );
  INV_X1 U19956 ( .A(n16741), .ZN(n16742) );
  OAI21_X1 U19957 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17708), .A(
        n16742), .ZN(n17742) );
  INV_X1 U19958 ( .A(n17742), .ZN(n16808) );
  INV_X1 U19959 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16829) );
  INV_X1 U19960 ( .A(n16744), .ZN(n17749) );
  NAND2_X1 U19961 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17749), .ZN(
        n16743) );
  AOI21_X1 U19962 ( .B1(n16829), .B2(n16743), .A(n17708), .ZN(n17750) );
  OAI21_X1 U19963 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17749), .A(
        n16743), .ZN(n17771) );
  INV_X1 U19964 ( .A(n17771), .ZN(n16835) );
  OAI21_X1 U19965 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17779), .A(
        n16744), .ZN(n17783) );
  INV_X1 U19966 ( .A(n17783), .ZN(n16843) );
  INV_X1 U19967 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17807) );
  NOR2_X1 U19968 ( .A1(n17807), .A2(n16748), .ZN(n16746) );
  INV_X1 U19969 ( .A(n17779), .ZN(n16745) );
  OAI21_X1 U19970 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16746), .A(
        n16745), .ZN(n17799) );
  INV_X1 U19971 ( .A(n17799), .ZN(n16858) );
  OAI22_X1 U19972 ( .A1(n17807), .A2(n16747), .B1(n16748), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17803) );
  AND2_X1 U19973 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17818), .ZN(
        n17793) );
  OAI21_X1 U19974 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17793), .A(
        n16748), .ZN(n16749) );
  INV_X1 U19975 ( .A(n16749), .ZN(n17822) );
  NOR2_X1 U19976 ( .A1(n18070), .A2(n17867), .ZN(n17866) );
  NAND2_X1 U19977 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17866), .ZN(
        n16932) );
  NOR2_X1 U19978 ( .A1(n16932), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16912) );
  NOR2_X1 U19979 ( .A1(n9975), .A2(n16912), .ZN(n16923) );
  INV_X1 U19980 ( .A(n16923), .ZN(n16921) );
  OAI21_X1 U19981 ( .B1(n17793), .B2(n9975), .A(n16921), .ZN(n16876) );
  NOR2_X1 U19982 ( .A1(n16858), .A2(n16857), .ZN(n16856) );
  NOR2_X1 U19983 ( .A1(n16856), .A2(n9975), .ZN(n16842) );
  NOR2_X1 U19984 ( .A1(n16843), .A2(n16842), .ZN(n16841) );
  NOR2_X1 U19985 ( .A1(n16841), .A2(n9975), .ZN(n16834) );
  NOR2_X1 U19986 ( .A1(n16835), .A2(n16834), .ZN(n16833) );
  NOR2_X1 U19987 ( .A1(n16833), .A2(n9975), .ZN(n16822) );
  NOR2_X1 U19988 ( .A1(n17750), .A2(n16822), .ZN(n16821) );
  NOR2_X1 U19989 ( .A1(n16821), .A2(n9975), .ZN(n16807) );
  NOR2_X1 U19990 ( .A1(n16808), .A2(n16807), .ZN(n16806) );
  NOR2_X1 U19991 ( .A1(n16806), .A2(n9975), .ZN(n16794) );
  NOR2_X1 U19992 ( .A1(n16795), .A2(n16794), .ZN(n16793) );
  NOR2_X1 U19993 ( .A1(n16793), .A2(n9975), .ZN(n16785) );
  NOR2_X1 U19994 ( .A1(n9975), .A2(n18933), .ZN(n17120) );
  INV_X1 U19995 ( .A(n17120), .ZN(n17029) );
  NOR3_X1 U19996 ( .A1(n16763), .A2(n16762), .A3(n17029), .ZN(n16756) );
  NAND3_X1 U19997 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16752) );
  AOI21_X1 U19998 ( .B1(n16750), .B2(n17106), .A(n17115), .ZN(n16814) );
  INV_X1 U19999 ( .A(n16814), .ZN(n16751) );
  AOI21_X1 U20000 ( .B1(n17106), .B2(n16752), .A(n16751), .ZN(n16781) );
  NOR2_X1 U20001 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16753), .ZN(n16766) );
  INV_X1 U20002 ( .A(n16766), .ZN(n16754) );
  AOI21_X1 U20003 ( .B1(n16781), .B2(n16754), .A(n19014), .ZN(n16755) );
  AOI211_X1 U20004 ( .C1(n16768), .C2(n16757), .A(n16756), .B(n16755), .ZN(
        n16758) );
  OAI211_X1 U20005 ( .C1(n16760), .C2(n17095), .A(n16759), .B(n16758), .ZN(
        P3_U2640) );
  NAND2_X1 U20006 ( .A1(n17091), .A2(n16761), .ZN(n16777) );
  XOR2_X1 U20007 ( .A(n16763), .B(n16762), .Z(n16767) );
  INV_X1 U20008 ( .A(n18933), .ZN(n17084) );
  OAI22_X1 U20009 ( .A1(n16781), .A2(n19016), .B1(n16764), .B2(n17095), .ZN(
        n16765) );
  AOI211_X1 U20010 ( .C1(n16767), .C2(n17084), .A(n16766), .B(n16765), .ZN(
        n16770) );
  OAI21_X1 U20011 ( .B1(n17116), .B2(n16768), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16769) );
  INV_X1 U20012 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19011) );
  AOI211_X1 U20013 ( .C1(n16773), .C2(n16772), .A(n16771), .B(n18933), .ZN(
        n16776) );
  NAND3_X1 U20014 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16782), .ZN(n16774) );
  OAI22_X1 U20015 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16774), .B1(n9968), 
        .B2(n17095), .ZN(n16775) );
  AOI211_X1 U20016 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17116), .A(n16776), .B(
        n16775), .ZN(n16780) );
  INV_X1 U20017 ( .A(n16777), .ZN(n16778) );
  OAI21_X1 U20018 ( .B1(n16783), .B2(n17136), .A(n16778), .ZN(n16779) );
  OAI211_X1 U20019 ( .C1(n16781), .C2(n19011), .A(n16780), .B(n16779), .ZN(
        P3_U2642) );
  NAND2_X1 U20020 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16782), .ZN(n16791) );
  AOI22_X1 U20021 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17121), .B1(
        n17116), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16790) );
  INV_X1 U20022 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19007) );
  NAND2_X1 U20023 ( .A1(n16782), .A2(n19007), .ZN(n16801) );
  NAND2_X1 U20024 ( .A1(n16814), .A2(n16801), .ZN(n16788) );
  AOI211_X1 U20025 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16799), .A(n16783), .B(
        n17126), .ZN(n16787) );
  AOI211_X1 U20026 ( .C1(n17710), .C2(n16785), .A(n16784), .B(n18933), .ZN(
        n16786) );
  AOI211_X1 U20027 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16788), .A(n16787), 
        .B(n16786), .ZN(n16789) );
  OAI211_X1 U20028 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16791), .A(n16790), 
        .B(n16789), .ZN(P3_U2643) );
  OAI21_X1 U20029 ( .B1(n16796), .B2(n16804), .A(n17091), .ZN(n16792) );
  INV_X1 U20030 ( .A(n16792), .ZN(n16800) );
  AOI211_X1 U20031 ( .C1(n16795), .C2(n16794), .A(n16793), .B(n18933), .ZN(
        n16798) );
  INV_X1 U20032 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17733) );
  OAI22_X1 U20033 ( .A1(n17733), .A2(n17095), .B1(n17127), .B2(n16796), .ZN(
        n16797) );
  AOI211_X1 U20034 ( .C1(n16800), .C2(n16799), .A(n16798), .B(n16797), .ZN(
        n16802) );
  OAI211_X1 U20035 ( .C1(n16814), .C2(n19007), .A(n16802), .B(n16801), .ZN(
        P3_U2644) );
  AND2_X1 U20036 ( .A1(n17106), .A2(n16803), .ZN(n16815) );
  AOI21_X1 U20037 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16815), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16813) );
  AOI22_X1 U20038 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17121), .B1(
        n17116), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16812) );
  AOI211_X1 U20039 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16805), .A(n16804), .B(
        n17126), .ZN(n16810) );
  AOI211_X1 U20040 ( .C1(n16808), .C2(n16807), .A(n16806), .B(n18933), .ZN(
        n16809) );
  NOR2_X1 U20041 ( .A1(n16810), .A2(n16809), .ZN(n16811) );
  OAI211_X1 U20042 ( .C1(n16814), .C2(n16813), .A(n16812), .B(n16811), .ZN(
        P3_U2645) );
  INV_X1 U20043 ( .A(n16815), .ZN(n16818) );
  NOR2_X1 U20044 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17118), .ZN(n16830) );
  NAND2_X1 U20045 ( .A1(n17106), .A2(n16816), .ZN(n16844) );
  NAND2_X1 U20046 ( .A1(n17130), .A2(n16844), .ZN(n16840) );
  NOR2_X1 U20047 ( .A1(n16830), .A2(n16840), .ZN(n16817) );
  MUX2_X1 U20048 ( .A(n16818), .B(n16817), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n16828) );
  INV_X1 U20049 ( .A(n16819), .ZN(n16820) );
  OAI21_X1 U20050 ( .B1(n17126), .B2(n16820), .A(n17127), .ZN(n16826) );
  NAND2_X1 U20051 ( .A1(n16820), .A2(n17091), .ZN(n16832) );
  INV_X1 U20052 ( .A(n16832), .ZN(n16825) );
  AOI211_X1 U20053 ( .C1(n17750), .C2(n16822), .A(n16821), .B(n18933), .ZN(
        n16823) );
  AOI221_X1 U20054 ( .B1(n16826), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n16825), 
        .C2(n16824), .A(n16823), .ZN(n16827) );
  OAI211_X1 U20055 ( .C1(n16829), .C2(n17095), .A(n16828), .B(n16827), .ZN(
        P3_U2646) );
  INV_X1 U20056 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17762) );
  AOI22_X1 U20057 ( .A1(n17116), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16831), 
        .B2(n16830), .ZN(n16839) );
  AOI21_X1 U20058 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16848), .A(n16832), .ZN(
        n16837) );
  AOI211_X1 U20059 ( .C1(n16835), .C2(n16834), .A(n16833), .B(n18933), .ZN(
        n16836) );
  AOI211_X1 U20060 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16840), .A(n16837), 
        .B(n16836), .ZN(n16838) );
  OAI211_X1 U20061 ( .C1(n17762), .C2(n17095), .A(n16839), .B(n16838), .ZN(
        P3_U2647) );
  INV_X1 U20062 ( .A(n16840), .ZN(n16851) );
  AOI211_X1 U20063 ( .C1(n16843), .C2(n16842), .A(n16841), .B(n18933), .ZN(
        n16847) );
  OAI22_X1 U20064 ( .A1(n17127), .A2(n17186), .B1(n16845), .B2(n16844), .ZN(
        n16846) );
  AOI211_X1 U20065 ( .C1(n17121), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16847), .B(n16846), .ZN(n16850) );
  OAI211_X1 U20066 ( .C1(n16852), .C2(n17186), .A(n17091), .B(n16848), .ZN(
        n16849) );
  OAI211_X1 U20067 ( .C1(n16851), .C2(n19000), .A(n16850), .B(n16849), .ZN(
        P3_U2648) );
  INV_X1 U20068 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16864) );
  AOI211_X1 U20069 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16866), .A(n16852), .B(
        n17126), .ZN(n16853) );
  AOI21_X1 U20070 ( .B1(n17121), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16853), .ZN(n16863) );
  AOI21_X1 U20071 ( .B1(n16854), .B2(n17106), .A(n17115), .ZN(n16881) );
  INV_X1 U20072 ( .A(n16881), .ZN(n16861) );
  NAND2_X1 U20073 ( .A1(n17106), .A2(n16882), .ZN(n16943) );
  INV_X1 U20074 ( .A(n16943), .ZN(n16929) );
  NAND2_X1 U20075 ( .A1(n16855), .A2(n16929), .ZN(n16871) );
  AOI221_X1 U20076 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(P3_REIP_REG_22__SCAN_IN), .C1(n18996), .C2(n18997), .A(n16871), .ZN(n16860) );
  AOI211_X1 U20077 ( .C1(n16858), .C2(n16857), .A(n16856), .B(n18933), .ZN(
        n16859) );
  AOI211_X1 U20078 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16861), .A(n16860), 
        .B(n16859), .ZN(n16862) );
  OAI211_X1 U20079 ( .C1(n17127), .C2(n16864), .A(n16863), .B(n16862), .ZN(
        P3_U2649) );
  AOI211_X1 U20080 ( .C1(n17803), .C2(n16865), .A(n9768), .B(n18933), .ZN(
        n16869) );
  OAI211_X1 U20081 ( .C1(n16872), .C2(n17222), .A(n17091), .B(n16866), .ZN(
        n16867) );
  OAI21_X1 U20082 ( .B1(n17222), .B2(n17127), .A(n16867), .ZN(n16868) );
  AOI211_X1 U20083 ( .C1(n17121), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16869), .B(n16868), .ZN(n16870) );
  OAI221_X1 U20084 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16871), .C1(n18996), 
        .C2(n16881), .A(n16870), .ZN(P3_U2650) );
  AOI211_X1 U20085 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16890), .A(n16872), .B(
        n17126), .ZN(n16873) );
  AOI21_X1 U20086 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17116), .A(n16873), .ZN(
        n16880) );
  OR2_X1 U20087 ( .A1(n16883), .A2(n16943), .ZN(n16895) );
  NOR3_X1 U20088 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16874), .A3(n16895), 
        .ZN(n16878) );
  AOI211_X1 U20089 ( .C1(n17822), .C2(n16876), .A(n16875), .B(n18933), .ZN(
        n16877) );
  AOI211_X1 U20090 ( .C1(n17121), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16878), .B(n16877), .ZN(n16879) );
  OAI211_X1 U20091 ( .C1(n18993), .C2(n16881), .A(n16880), .B(n16879), .ZN(
        P3_U2651) );
  NAND2_X1 U20092 ( .A1(n16882), .A2(n17130), .ZN(n16946) );
  NOR2_X1 U20093 ( .A1(n16883), .A2(n16946), .ZN(n16904) );
  NAND2_X1 U20094 ( .A1(n17130), .A2(n17118), .ZN(n17128) );
  INV_X1 U20095 ( .A(n17128), .ZN(n16905) );
  AOI21_X1 U20096 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16904), .A(n16905), 
        .ZN(n16901) );
  INV_X1 U20097 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18989) );
  NOR3_X1 U20098 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18989), .A3(n16895), 
        .ZN(n16889) );
  INV_X1 U20099 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16887) );
  INV_X1 U20100 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16911) );
  NAND2_X1 U20101 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17851), .ZN(
        n16919) );
  NOR2_X1 U20102 ( .A1(n16911), .A2(n16919), .ZN(n17828) );
  NAND2_X1 U20103 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17828), .ZN(
        n16896) );
  INV_X1 U20104 ( .A(n16912), .ZN(n16936) );
  OAI21_X1 U20105 ( .B1(n16896), .B2(n16936), .A(n17083), .ZN(n16898) );
  AOI21_X1 U20106 ( .B1(n16887), .B2(n16896), .A(n17793), .ZN(n16884) );
  INV_X1 U20107 ( .A(n16884), .ZN(n17832) );
  AOI21_X1 U20108 ( .B1(n16898), .B2(n17832), .A(n18933), .ZN(n16885) );
  OAI21_X1 U20109 ( .B1(n16898), .B2(n17832), .A(n16885), .ZN(n16886) );
  OAI211_X1 U20110 ( .C1(n16887), .C2(n17095), .A(n9655), .B(n16886), .ZN(
        n16888) );
  AOI211_X1 U20111 ( .C1(n16901), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16889), 
        .B(n16888), .ZN(n16892) );
  OAI211_X1 U20112 ( .C1(n16893), .C2(n17239), .A(n17091), .B(n16890), .ZN(
        n16891) );
  OAI211_X1 U20113 ( .C1(n17239), .C2(n17127), .A(n16892), .B(n16891), .ZN(
        P3_U2652) );
  INV_X1 U20114 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17845) );
  AOI211_X1 U20115 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16909), .A(n16893), .B(
        n17126), .ZN(n16894) );
  AOI21_X1 U20116 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17116), .A(n16894), .ZN(
        n16903) );
  NAND2_X1 U20117 ( .A1(n18989), .A2(n16895), .ZN(n16900) );
  OAI21_X1 U20118 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17828), .A(
        n16896), .ZN(n17842) );
  NAND2_X1 U20119 ( .A1(n9975), .A2(n17084), .ZN(n17101) );
  OAI221_X1 U20120 ( .B1(n17842), .B2(n16912), .C1(n17842), .C2(n17845), .A(
        n17084), .ZN(n16897) );
  AOI22_X1 U20121 ( .A1(n16898), .A2(n17842), .B1(n17101), .B2(n16897), .ZN(
        n16899) );
  AOI211_X1 U20122 ( .C1(n16901), .C2(n16900), .A(n18393), .B(n16899), .ZN(
        n16902) );
  OAI211_X1 U20123 ( .C1(n17845), .C2(n17095), .A(n16903), .B(n16902), .ZN(
        P3_U2653) );
  NAND2_X1 U20124 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16928) );
  NOR2_X1 U20125 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16928), .ZN(n16908) );
  INV_X1 U20126 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18988) );
  NOR3_X1 U20127 ( .A1(n16905), .A2(n16904), .A3(n18988), .ZN(n16907) );
  OAI22_X1 U20128 ( .A1(n16911), .A2(n17095), .B1(n17127), .B2(n16910), .ZN(
        n16906) );
  AOI211_X1 U20129 ( .C1(n16929), .C2(n16908), .A(n16907), .B(n16906), .ZN(
        n16917) );
  OAI211_X1 U20130 ( .C1(n16918), .C2(n16910), .A(n17091), .B(n16909), .ZN(
        n16916) );
  AOI21_X1 U20131 ( .B1(n16911), .B2(n16919), .A(n17828), .ZN(n17855) );
  AOI21_X1 U20132 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16912), .A(
        n9975), .ZN(n16914) );
  AOI21_X1 U20133 ( .B1(n17855), .B2(n16914), .A(n18933), .ZN(n16913) );
  OAI21_X1 U20134 ( .B1(n17855), .B2(n16914), .A(n16913), .ZN(n16915) );
  NAND4_X1 U20135 ( .A1(n16917), .A2(n9655), .A3(n16916), .A4(n16915), .ZN(
        P3_U2654) );
  NAND2_X1 U20136 ( .A1(n17128), .A2(n16946), .ZN(n16951) );
  INV_X1 U20137 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18985) );
  AOI211_X1 U20138 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16934), .A(n16918), .B(
        n17126), .ZN(n16927) );
  INV_X1 U20139 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16925) );
  INV_X1 U20140 ( .A(n16932), .ZN(n16920) );
  OAI21_X1 U20141 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16920), .A(
        n16919), .ZN(n17871) );
  INV_X1 U20142 ( .A(n17871), .ZN(n16922) );
  OAI221_X1 U20143 ( .B1(n16923), .B2(n16922), .C1(n16921), .C2(n17871), .A(
        n17084), .ZN(n16924) );
  OAI211_X1 U20144 ( .C1(n16925), .C2(n17095), .A(n9655), .B(n16924), .ZN(
        n16926) );
  AOI211_X1 U20145 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17116), .A(n16927), .B(
        n16926), .ZN(n16931) );
  OAI211_X1 U20146 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16929), .B(n16928), .ZN(n16930) );
  OAI211_X1 U20147 ( .C1(n16951), .C2(n18985), .A(n16931), .B(n16930), .ZN(
        P3_U2655) );
  INV_X1 U20148 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18983) );
  INV_X1 U20149 ( .A(n17866), .ZN(n16933) );
  INV_X1 U20150 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17053) );
  OAI21_X1 U20151 ( .B1(n9975), .B2(n17053), .A(n17084), .ZN(n17113) );
  OAI21_X1 U20152 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17866), .A(
        n16932), .ZN(n17880) );
  AOI211_X1 U20153 ( .C1(n17083), .C2(n16933), .A(n17113), .B(n17880), .ZN(
        n16941) );
  INV_X1 U20154 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17883) );
  OAI211_X1 U20155 ( .C1(n16944), .C2(n16938), .A(n17091), .B(n16934), .ZN(
        n16935) );
  OAI21_X1 U20156 ( .B1(n17095), .B2(n17883), .A(n16935), .ZN(n16940) );
  NAND2_X1 U20157 ( .A1(n16936), .A2(n17880), .ZN(n16937) );
  OAI22_X1 U20158 ( .A1(n17127), .A2(n16938), .B1(n17029), .B2(n16937), .ZN(
        n16939) );
  NOR4_X1 U20159 ( .A1(n18393), .A2(n16941), .A3(n16940), .A4(n16939), .ZN(
        n16942) );
  OAI221_X1 U20160 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16943), .C1(n18983), 
        .C2(n16951), .A(n16942), .ZN(P3_U2656) );
  AOI211_X1 U20161 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16956), .A(n16944), .B(
        n17126), .ZN(n16953) );
  NOR2_X1 U20162 ( .A1(n17118), .A2(n16945), .ZN(n16960) );
  NAND3_X1 U20163 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16960), .A3(n16946), 
        .ZN(n16950) );
  INV_X1 U20164 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16947) );
  INV_X1 U20165 ( .A(n17994), .ZN(n17939) );
  NAND2_X1 U20166 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17939), .ZN(
        n17026) );
  NOR2_X1 U20167 ( .A1(n17906), .A2(n17026), .ZN(n17909) );
  NAND2_X1 U20168 ( .A1(n17914), .A2(n17909), .ZN(n16958) );
  AOI21_X1 U20169 ( .B1(n16947), .B2(n16958), .A(n17866), .ZN(n17901) );
  INV_X1 U20170 ( .A(n17925), .ZN(n17891) );
  NOR2_X1 U20171 ( .A1(n18070), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17015) );
  INV_X1 U20172 ( .A(n17015), .ZN(n17099) );
  OAI21_X1 U20173 ( .B1(n17891), .B2(n17099), .A(n17083), .ZN(n16970) );
  OAI21_X1 U20174 ( .B1(n17914), .B2(n9975), .A(n16970), .ZN(n16963) );
  AOI21_X1 U20175 ( .B1(n17901), .B2(n16963), .A(n18933), .ZN(n16948) );
  OAI21_X1 U20176 ( .B1(n17901), .B2(n16963), .A(n16948), .ZN(n16949) );
  OAI211_X1 U20177 ( .C1(n16951), .C2(n18982), .A(n16950), .B(n16949), .ZN(
        n16952) );
  AOI211_X1 U20178 ( .C1(n17121), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16953), .B(n16952), .ZN(n16954) );
  OAI211_X1 U20179 ( .C1(n17127), .C2(n17305), .A(n16954), .B(n9655), .ZN(
        P3_U2657) );
  AOI21_X1 U20180 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16955), .A(n17126), .ZN(
        n16957) );
  AOI22_X1 U20181 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17121), .B1(
        n16957), .B2(n16956), .ZN(n16967) );
  INV_X1 U20182 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16969) );
  INV_X1 U20183 ( .A(n17909), .ZN(n16980) );
  NOR2_X1 U20184 ( .A1(n16969), .A2(n16980), .ZN(n16968) );
  OAI21_X1 U20185 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16968), .A(
        n16958), .ZN(n17912) );
  AOI211_X1 U20186 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17101), .A(
        n17113), .B(n17912), .ZN(n16959) );
  AOI211_X1 U20187 ( .C1(n17116), .C2(P3_EBX_REG_13__SCAN_IN), .A(n18393), .B(
        n16959), .ZN(n16966) );
  INV_X1 U20188 ( .A(n16960), .ZN(n16962) );
  NOR2_X1 U20189 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17118), .ZN(n16974) );
  OAI21_X1 U20190 ( .B1(n16975), .B2(n17118), .A(n17130), .ZN(n16984) );
  NOR2_X1 U20191 ( .A1(n16974), .A2(n16984), .ZN(n16961) );
  MUX2_X1 U20192 ( .A(n16962), .B(n16961), .S(P3_REIP_REG_13__SCAN_IN), .Z(
        n16965) );
  NAND3_X1 U20193 ( .A1(n17084), .A2(n17912), .A3(n16963), .ZN(n16964) );
  NAND4_X1 U20194 ( .A1(n16967), .A2(n16966), .A3(n16965), .A4(n16964), .ZN(
        P3_U2658) );
  AOI22_X1 U20195 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17121), .B1(
        n17116), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16978) );
  AOI21_X1 U20196 ( .B1(n16969), .B2(n16980), .A(n16968), .ZN(n17926) );
  XNOR2_X1 U20197 ( .A(n17926), .B(n16970), .ZN(n16973) );
  AOI211_X1 U20198 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16986), .A(n16971), .B(
        n17126), .ZN(n16972) );
  AOI211_X1 U20199 ( .C1(n17084), .C2(n16973), .A(n18393), .B(n16972), .ZN(
        n16977) );
  AOI22_X1 U20200 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16984), .B1(n16975), 
        .B2(n16974), .ZN(n16976) );
  NAND3_X1 U20201 ( .A1(n16978), .A2(n16977), .A3(n16976), .ZN(P3_U2659) );
  AOI22_X1 U20202 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17121), .B1(
        n17116), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n16989) );
  NOR3_X1 U20203 ( .A1(n17118), .A2(n18964), .A3(n17054), .ZN(n17042) );
  NAND4_X1 U20204 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .A4(n17042), .ZN(n16998) );
  OAI21_X1 U20205 ( .B1(n16979), .B2(n16998), .A(n18975), .ZN(n16985) );
  INV_X1 U20206 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17950) );
  NOR2_X1 U20207 ( .A1(n17979), .A2(n17026), .ZN(n17014) );
  NAND2_X1 U20208 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17014), .ZN(
        n17002) );
  NOR2_X1 U20209 ( .A1(n17950), .A2(n17002), .ZN(n16990) );
  OAI21_X1 U20210 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16990), .A(
        n16980), .ZN(n17940) );
  NOR2_X1 U20211 ( .A1(n17994), .A2(n17099), .ZN(n17030) );
  NAND3_X1 U20212 ( .A1(n17938), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17030), .ZN(n16991) );
  OAI21_X1 U20213 ( .B1(n17950), .B2(n16991), .A(n17083), .ZN(n16982) );
  OAI21_X1 U20214 ( .B1(n17940), .B2(n16982), .A(n17084), .ZN(n16981) );
  AOI21_X1 U20215 ( .B1(n17940), .B2(n16982), .A(n16981), .ZN(n16983) );
  AOI211_X1 U20216 ( .C1(n16985), .C2(n16984), .A(n18393), .B(n16983), .ZN(
        n16988) );
  OAI211_X1 U20217 ( .C1(n16993), .C2(n17345), .A(n17091), .B(n16986), .ZN(
        n16987) );
  NAND3_X1 U20218 ( .A1(n16989), .A2(n16988), .A3(n16987), .ZN(P3_U2660) );
  AOI21_X1 U20219 ( .B1(n17950), .B2(n17002), .A(n16990), .ZN(n17953) );
  NAND2_X1 U20220 ( .A1(n17083), .A2(n16991), .ZN(n17007) );
  XNOR2_X1 U20221 ( .A(n17953), .B(n17007), .ZN(n16992) );
  AOI22_X1 U20222 ( .A1(n17116), .A2(P3_EBX_REG_10__SCAN_IN), .B1(n17084), 
        .B2(n16992), .ZN(n17001) );
  INV_X1 U20223 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18971) );
  NOR3_X1 U20224 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18971), .A3(n16998), 
        .ZN(n16996) );
  AOI211_X1 U20225 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16994), .A(n16993), .B(
        n17126), .ZN(n16995) );
  AOI211_X1 U20226 ( .C1(n17121), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16996), .B(n16995), .ZN(n17000) );
  AOI21_X1 U20227 ( .B1(n16997), .B2(n17106), .A(n17115), .ZN(n17013) );
  INV_X1 U20228 ( .A(n17013), .ZN(n17021) );
  NOR2_X1 U20229 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16998), .ZN(n17009) );
  OAI21_X1 U20230 ( .B1(n17021), .B2(n17009), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16999) );
  NAND4_X1 U20231 ( .A1(n17001), .A2(n17000), .A3(n9655), .A4(n16999), .ZN(
        P3_U2661) );
  OAI21_X1 U20232 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17014), .A(
        n17002), .ZN(n17969) );
  OAI221_X1 U20233 ( .B1(n17969), .B2(n17938), .C1(n17969), .C2(n17030), .A(
        n17084), .ZN(n17006) );
  INV_X1 U20234 ( .A(n17101), .ZN(n17066) );
  INV_X1 U20235 ( .A(n17969), .ZN(n17004) );
  NOR2_X1 U20236 ( .A1(n17010), .A2(n17126), .ZN(n17018) );
  AOI22_X1 U20237 ( .A1(n17066), .A2(n17004), .B1(n17018), .B2(n17003), .ZN(
        n17005) );
  OAI211_X1 U20238 ( .C1(n17007), .C2(n17006), .A(n17005), .B(n9655), .ZN(
        n17008) );
  AOI211_X1 U20239 ( .C1(n17121), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17009), .B(n17008), .ZN(n17012) );
  OAI221_X1 U20240 ( .B1(n17116), .B2(n17091), .C1(n17116), .C2(n17010), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n17011) );
  OAI211_X1 U20241 ( .C1(n17013), .C2(n18971), .A(n17012), .B(n17011), .ZN(
        P3_U2662) );
  AOI22_X1 U20242 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17121), .B1(
        n17116), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n17024) );
  INV_X1 U20243 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17982) );
  INV_X1 U20244 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17995) );
  NOR2_X1 U20245 ( .A1(n17994), .A2(n17995), .ZN(n17980) );
  NAND2_X1 U20246 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17980), .ZN(
        n17027) );
  AOI21_X1 U20247 ( .B1(n17982), .B2(n17027), .A(n17014), .ZN(n17989) );
  AOI21_X1 U20248 ( .B1(n17980), .B2(n17015), .A(n9975), .ZN(n17016) );
  XOR2_X1 U20249 ( .A(n17989), .B(n17016), .Z(n17019) );
  NAND2_X1 U20250 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17031), .ZN(n17017) );
  AOI22_X1 U20251 ( .A1(n17084), .A2(n17019), .B1(n17018), .B2(n17017), .ZN(
        n17023) );
  INV_X1 U20252 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18967) );
  INV_X1 U20253 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18965) );
  NOR3_X1 U20254 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18967), .A3(n18965), .ZN(
        n17020) );
  AOI22_X1 U20255 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17021), .B1(n17042), 
        .B2(n17020), .ZN(n17022) );
  NAND4_X1 U20256 ( .A1(n17024), .A2(n17023), .A3(n17022), .A4(n9655), .ZN(
        P3_U2663) );
  NAND2_X1 U20257 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17042), .ZN(n17037) );
  NAND2_X1 U20258 ( .A1(n17025), .A2(n17130), .ZN(n17055) );
  OAI21_X1 U20259 ( .B1(n18965), .B2(n17055), .A(n17128), .ZN(n17044) );
  OAI22_X1 U20260 ( .A1(n17995), .A2(n17095), .B1(n17127), .B2(n17403), .ZN(
        n17035) );
  INV_X1 U20261 ( .A(n17026), .ZN(n17038) );
  OAI21_X1 U20262 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17038), .A(
        n17027), .ZN(n17028) );
  INV_X1 U20263 ( .A(n17028), .ZN(n18002) );
  OR2_X1 U20264 ( .A1(n17030), .A2(n17029), .ZN(n17050) );
  OAI211_X1 U20265 ( .C1(n17030), .C2(n9975), .A(n17084), .B(n18002), .ZN(
        n17033) );
  OAI211_X1 U20266 ( .C1(n17041), .C2(n17403), .A(n17091), .B(n17031), .ZN(
        n17032) );
  OAI211_X1 U20267 ( .C1(n18002), .C2(n17050), .A(n17033), .B(n17032), .ZN(
        n17034) );
  NOR3_X1 U20268 ( .A1(n18393), .A2(n17035), .A3(n17034), .ZN(n17036) );
  OAI221_X1 U20269 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n17037), .C1(n18967), 
        .C2(n17044), .A(n17036), .ZN(P3_U2664) );
  NAND2_X1 U20270 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18013), .ZN(
        n17051) );
  AOI21_X1 U20271 ( .B1(n9982), .B2(n17051), .A(n17038), .ZN(n18014) );
  NAND2_X1 U20272 ( .A1(n17084), .A2(n17053), .ZN(n17039) );
  OAI21_X1 U20273 ( .B1(n17051), .B2(n17039), .A(n17101), .ZN(n17040) );
  AOI21_X1 U20274 ( .B1(n18014), .B2(n17040), .A(n18393), .ZN(n17049) );
  AOI211_X1 U20275 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17057), .A(n17041), .B(
        n17126), .ZN(n17047) );
  NOR2_X1 U20276 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17042), .ZN(n17045) );
  INV_X1 U20277 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17043) );
  OAI22_X1 U20278 ( .A1(n17045), .A2(n17044), .B1(n17127), .B2(n17043), .ZN(
        n17046) );
  AOI211_X1 U20279 ( .C1(n17121), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17047), .B(n17046), .ZN(n17048) );
  OAI211_X1 U20280 ( .C1(n18014), .C2(n17050), .A(n17049), .B(n17048), .ZN(
        P3_U2665) );
  NOR2_X1 U20281 ( .A1(n18070), .A2(n18021), .ZN(n17065) );
  OAI21_X1 U20282 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17065), .A(
        n17051), .ZN(n18025) );
  AOI21_X1 U20283 ( .B1(n17053), .B2(n17065), .A(n9975), .ZN(n17073) );
  XNOR2_X1 U20284 ( .A(n18025), .B(n17073), .ZN(n17061) );
  NOR2_X1 U20285 ( .A1(n17118), .A2(n17054), .ZN(n17056) );
  OAI211_X1 U20286 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n17056), .A(n17055), .B(
        n17128), .ZN(n17059) );
  OAI211_X1 U20287 ( .C1(n17063), .C2(n17418), .A(n17091), .B(n17057), .ZN(
        n17058) );
  OAI211_X1 U20288 ( .C1(n17418), .C2(n17127), .A(n17059), .B(n17058), .ZN(
        n17060) );
  AOI211_X1 U20289 ( .C1(n17084), .C2(n17061), .A(n18393), .B(n17060), .ZN(
        n17062) );
  OAI21_X1 U20290 ( .B1(n18020), .B2(n17095), .A(n17062), .ZN(P3_U2666) );
  NOR2_X1 U20291 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17118), .ZN(n17072) );
  AOI211_X1 U20292 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17090), .A(n17063), .B(
        n17126), .ZN(n17070) );
  AOI21_X1 U20293 ( .B1(n17106), .B2(n17064), .A(n17115), .ZN(n17086) );
  INV_X1 U20294 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18961) );
  INV_X1 U20295 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17074) );
  NAND2_X1 U20296 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18047), .ZN(
        n17081) );
  AOI21_X1 U20297 ( .B1(n17074), .B2(n17081), .A(n17065), .ZN(n18037) );
  AOI22_X1 U20298 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17121), .B1(
        n18037), .B2(n17066), .ZN(n17068) );
  NAND2_X1 U20299 ( .A1(n18416), .A2(n19089), .ZN(n17133) );
  INV_X1 U20300 ( .A(n17133), .ZN(n19091) );
  OAI21_X1 U20301 ( .B1(n12550), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19091), .ZN(n17067) );
  OAI211_X1 U20302 ( .C1(n17086), .C2(n18961), .A(n17068), .B(n17067), .ZN(
        n17069) );
  AOI211_X1 U20303 ( .C1(n17072), .C2(n17071), .A(n17070), .B(n17069), .ZN(
        n17078) );
  INV_X1 U20304 ( .A(n17073), .ZN(n17075) );
  NAND2_X1 U20305 ( .A1(n18047), .A2(n17074), .ZN(n18035) );
  OAI22_X1 U20306 ( .A1(n18037), .A2(n17075), .B1(n17099), .B2(n18035), .ZN(
        n17076) );
  AOI21_X1 U20307 ( .B1(n17084), .B2(n17076), .A(n18393), .ZN(n17077) );
  OAI211_X1 U20308 ( .C1(n17079), .C2(n17127), .A(n17078), .B(n17077), .ZN(
        P3_U2667) );
  AOI21_X1 U20309 ( .B1(n17096), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n17385), .ZN(n17080) );
  INV_X1 U20310 ( .A(n17080), .ZN(n19029) );
  NOR2_X1 U20311 ( .A1(n18070), .A2(n17097), .ZN(n17082) );
  OAI21_X1 U20312 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17082), .A(
        n17081), .ZN(n18054) );
  OAI21_X1 U20313 ( .B1(n17097), .B2(n17099), .A(n17083), .ZN(n17098) );
  OAI21_X1 U20314 ( .B1(n18054), .B2(n17098), .A(n17084), .ZN(n17085) );
  AOI21_X1 U20315 ( .B1(n18054), .B2(n17098), .A(n17085), .ZN(n17089) );
  AOI21_X1 U20316 ( .B1(n17106), .B2(n17104), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n17087) );
  OAI22_X1 U20317 ( .A1(n17087), .A2(n17086), .B1(n17127), .B2(n17423), .ZN(
        n17088) );
  AOI211_X1 U20318 ( .C1(n19091), .C2(n19029), .A(n17089), .B(n17088), .ZN(
        n17093) );
  OAI211_X1 U20319 ( .C1(n17107), .C2(n17423), .A(n17091), .B(n17090), .ZN(
        n17092) );
  OAI211_X1 U20320 ( .C1(n17095), .C2(n17094), .A(n17093), .B(n17092), .ZN(
        P3_U2668) );
  NAND2_X1 U20321 ( .A1(n12678), .A2(n18875), .ZN(n18866) );
  NAND2_X1 U20322 ( .A1(n17096), .A2(n18866), .ZN(n18880) );
  INV_X1 U20323 ( .A(n18880), .ZN(n19038) );
  AOI22_X1 U20324 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17121), .B1(
        n19038), .B2(n19091), .ZN(n17112) );
  OAI22_X1 U20325 ( .A1(n18070), .A2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n17097), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17100) );
  AOI211_X1 U20326 ( .C1(n17100), .C2(n17099), .A(n18933), .B(n17098), .ZN(
        n17103) );
  INV_X1 U20327 ( .A(n17100), .ZN(n18061) );
  OAI22_X1 U20328 ( .A1(n17130), .A2(n18957), .B1(n18061), .B2(n17101), .ZN(
        n17102) );
  AOI211_X1 U20329 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17116), .A(n17103), .B(
        n17102), .ZN(n17111) );
  INV_X1 U20330 ( .A(n17104), .ZN(n17105) );
  OAI211_X1 U20331 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17106), .B(n17105), .ZN(n17110) );
  NAND2_X1 U20332 ( .A1(n17438), .A2(n17433), .ZN(n17117) );
  AOI211_X1 U20333 ( .C1(n17117), .C2(P3_EBX_REG_2__SCAN_IN), .A(n17126), .B(
        n17107), .ZN(n17108) );
  INV_X1 U20334 ( .A(n17108), .ZN(n17109) );
  NAND4_X1 U20335 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        P3_U2669) );
  OAI21_X1 U20336 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18875), .ZN(n18892) );
  OAI22_X1 U20337 ( .A1(n17133), .A2(n18892), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17113), .ZN(n17114) );
  INV_X1 U20338 ( .A(n17114), .ZN(n17125) );
  AOI22_X1 U20339 ( .A1(n17116), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n17115), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17124) );
  OAI21_X1 U20340 ( .B1(n17433), .B2(n17438), .A(n17117), .ZN(n17434) );
  OAI22_X1 U20341 ( .A1(n17126), .A2(n17434), .B1(n17118), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17119) );
  INV_X1 U20342 ( .A(n17119), .ZN(n17123) );
  OAI221_X1 U20343 ( .B1(n17121), .B2(n17120), .C1(n17121), .C2(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17122) );
  NAND4_X1 U20344 ( .A1(n17125), .A2(n17124), .A3(n17123), .A4(n17122), .ZN(
        P3_U2670) );
  NAND2_X1 U20345 ( .A1(n17127), .A2(n17126), .ZN(n17129) );
  AOI22_X1 U20346 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17129), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17128), .ZN(n17132) );
  NAND3_X1 U20347 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19032), .A3(
        n17130), .ZN(n17131) );
  OAI211_X1 U20348 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17133), .A(
        n17132), .B(n17131), .ZN(P3_U2671) );
  NAND4_X1 U20349 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17135), .A4(n17134), .ZN(n17167) );
  NAND2_X1 U20350 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17252), .ZN(n17221) );
  NOR3_X1 U20351 ( .A1(n17136), .A2(n17167), .A3(n17221), .ZN(n17162) );
  NAND2_X1 U20352 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17162), .ZN(n17161) );
  INV_X1 U20353 ( .A(n17161), .ZN(n17137) );
  OAI33_X1 U20354 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17161), .A3(n17564), 
        .B1(n17138), .B2(n17435), .B3(n17137), .ZN(P3_U2672) );
  AOI22_X1 U20355 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20356 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20357 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20358 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17139) );
  NAND4_X1 U20359 ( .A1(n17142), .A2(n17141), .A3(n17140), .A4(n17139), .ZN(
        n17148) );
  AOI22_X1 U20360 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20361 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17145) );
  AOI22_X1 U20362 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20363 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17143) );
  NAND4_X1 U20364 ( .A1(n17146), .A2(n17145), .A3(n17144), .A4(n17143), .ZN(
        n17147) );
  NOR2_X1 U20365 ( .A1(n17148), .A2(n17147), .ZN(n17160) );
  AOI22_X1 U20366 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20367 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20368 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17149) );
  OAI21_X1 U20369 ( .B1(n17150), .B2(n17415), .A(n17149), .ZN(n17156) );
  AOI22_X1 U20370 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20371 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17153) );
  AOI22_X1 U20372 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20373 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17151) );
  NAND4_X1 U20374 ( .A1(n17154), .A2(n17153), .A3(n17152), .A4(n17151), .ZN(
        n17155) );
  AOI211_X1 U20375 ( .C1(n17350), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n17156), .B(n17155), .ZN(n17157) );
  NAND3_X1 U20376 ( .A1(n17159), .A2(n17158), .A3(n17157), .ZN(n17165) );
  NAND2_X1 U20377 ( .A1(n17166), .A2(n17165), .ZN(n17164) );
  XNOR2_X1 U20378 ( .A(n17160), .B(n17164), .ZN(n17452) );
  OAI211_X1 U20379 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17162), .A(n17161), .B(
        n17431), .ZN(n17163) );
  OAI21_X1 U20380 ( .B1(n17452), .B2(n17431), .A(n17163), .ZN(P3_U2673) );
  OAI21_X1 U20381 ( .B1(n17166), .B2(n17165), .A(n17164), .ZN(n17456) );
  NOR2_X1 U20382 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17167), .ZN(n17168) );
  AOI22_X1 U20383 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17169), .B1(n17223), 
        .B2(n17168), .ZN(n17170) );
  OAI21_X1 U20384 ( .B1(n17456), .B2(n17431), .A(n17170), .ZN(P3_U2674) );
  OAI21_X1 U20385 ( .B1(n17175), .B2(n17172), .A(n17171), .ZN(n17465) );
  NAND3_X1 U20386 ( .A1(n17178), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17431), 
        .ZN(n17173) );
  OAI221_X1 U20387 ( .B1(n17178), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17431), 
        .C2(n17465), .A(n17173), .ZN(P3_U2676) );
  AOI21_X1 U20388 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17431), .A(n17185), .ZN(
        n17174) );
  INV_X1 U20389 ( .A(n17174), .ZN(n17177) );
  AOI21_X1 U20390 ( .B1(n17176), .B2(n17181), .A(n17175), .ZN(n17466) );
  AOI22_X1 U20391 ( .A1(n17178), .A2(n17177), .B1(n17466), .B2(n17435), .ZN(
        n17179) );
  INV_X1 U20392 ( .A(n17179), .ZN(P3_U2677) );
  INV_X1 U20393 ( .A(n17180), .ZN(n17189) );
  AOI21_X1 U20394 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17431), .A(n17189), .ZN(
        n17184) );
  OAI21_X1 U20395 ( .B1(n17183), .B2(n17182), .A(n17181), .ZN(n17475) );
  OAI22_X1 U20396 ( .A1(n17185), .A2(n17184), .B1(n17431), .B2(n17475), .ZN(
        P3_U2678) );
  NAND3_X1 U20397 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17223), .ZN(n17190) );
  NOR2_X1 U20398 ( .A1(n17186), .A2(n17190), .ZN(n17195) );
  AOI21_X1 U20399 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17431), .A(n17195), .ZN(
        n17188) );
  XNOR2_X1 U20400 ( .A(n17187), .B(n17191), .ZN(n17480) );
  OAI22_X1 U20401 ( .A1(n17189), .A2(n17188), .B1(n17431), .B2(n17480), .ZN(
        P3_U2679) );
  INV_X1 U20402 ( .A(n17190), .ZN(n17209) );
  AOI21_X1 U20403 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17431), .A(n17209), .ZN(
        n17194) );
  OAI21_X1 U20404 ( .B1(n17193), .B2(n17192), .A(n17191), .ZN(n17485) );
  OAI22_X1 U20405 ( .A1(n17195), .A2(n17194), .B1(n17431), .B2(n17485), .ZN(
        P3_U2680) );
  AOI22_X1 U20406 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17431), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n17223), .ZN(n17208) );
  AOI22_X1 U20407 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U20408 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17205) );
  AOI22_X1 U20409 ( .A1(n12581), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17196) );
  OAI21_X1 U20410 ( .B1(n17197), .B2(n17415), .A(n17196), .ZN(n17203) );
  AOI22_X1 U20411 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20412 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20413 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17199) );
  AOI22_X1 U20414 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17198) );
  NAND4_X1 U20415 ( .A1(n17201), .A2(n17200), .A3(n17199), .A4(n17198), .ZN(
        n17202) );
  AOI211_X1 U20416 ( .C1(n17384), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17203), .B(n17202), .ZN(n17204) );
  NAND3_X1 U20417 ( .A1(n17206), .A2(n17205), .A3(n17204), .ZN(n17486) );
  INV_X1 U20418 ( .A(n17486), .ZN(n17207) );
  OAI22_X1 U20419 ( .A1(n17209), .A2(n17208), .B1(n17207), .B2(n17431), .ZN(
        P3_U2681) );
  AOI22_X1 U20420 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20421 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20422 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20423 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17210) );
  NAND4_X1 U20424 ( .A1(n17213), .A2(n17212), .A3(n17211), .A4(n17210), .ZN(
        n17220) );
  AOI22_X1 U20425 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20426 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20427 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20428 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17215) );
  NAND4_X1 U20429 ( .A1(n17218), .A2(n17217), .A3(n17216), .A4(n17215), .ZN(
        n17219) );
  NOR2_X1 U20430 ( .A1(n17220), .A2(n17219), .ZN(n17492) );
  AND2_X1 U20431 ( .A1(n17431), .A2(n17221), .ZN(n17235) );
  AOI22_X1 U20432 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17235), .B1(n17223), 
        .B2(n17222), .ZN(n17224) );
  OAI21_X1 U20433 ( .B1(n17492), .B2(n17431), .A(n17224), .ZN(P3_U2682) );
  AOI22_X1 U20434 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20435 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20436 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20437 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17225) );
  NAND4_X1 U20438 ( .A1(n17228), .A2(n17227), .A3(n17226), .A4(n17225), .ZN(
        n17234) );
  AOI22_X1 U20439 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U20440 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20441 ( .A1(n12581), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20442 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17229) );
  NAND4_X1 U20443 ( .A1(n17232), .A2(n17231), .A3(n17230), .A4(n17229), .ZN(
        n17233) );
  NOR2_X1 U20444 ( .A1(n17234), .A2(n17233), .ZN(n17499) );
  OAI21_X1 U20445 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17236), .A(n17235), .ZN(
        n17237) );
  OAI21_X1 U20446 ( .B1(n17499), .B2(n17431), .A(n17237), .ZN(P3_U2683) );
  AOI21_X1 U20447 ( .B1(n17239), .B2(n17238), .A(n17435), .ZN(n17240) );
  INV_X1 U20448 ( .A(n17240), .ZN(n17251) );
  AOI22_X1 U20449 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17244) );
  AOI22_X1 U20450 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20451 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20452 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17241) );
  NAND4_X1 U20453 ( .A1(n17244), .A2(n17243), .A3(n17242), .A4(n17241), .ZN(
        n17250) );
  AOI22_X1 U20454 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20455 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20456 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U20457 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17245) );
  NAND4_X1 U20458 ( .A1(n17248), .A2(n17247), .A3(n17246), .A4(n17245), .ZN(
        n17249) );
  NOR2_X1 U20459 ( .A1(n17250), .A2(n17249), .ZN(n17504) );
  OAI22_X1 U20460 ( .A1(n17252), .A2(n17251), .B1(n17504), .B2(n17431), .ZN(
        P3_U2684) );
  AOI22_X1 U20461 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20462 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20463 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20464 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17253) );
  NAND4_X1 U20465 ( .A1(n17256), .A2(n17255), .A3(n17254), .A4(n17253), .ZN(
        n17262) );
  AOI22_X1 U20466 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20467 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20468 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20469 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17257) );
  NAND4_X1 U20470 ( .A1(n17260), .A2(n17259), .A3(n17258), .A4(n17257), .ZN(
        n17261) );
  NOR2_X1 U20471 ( .A1(n17262), .A2(n17261), .ZN(n17508) );
  NOR2_X1 U20472 ( .A1(n17435), .A2(n17264), .ZN(n17277) );
  NOR2_X1 U20473 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17564), .ZN(n17263) );
  AOI22_X1 U20474 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17277), .B1(n17264), 
        .B2(n17263), .ZN(n17265) );
  OAI21_X1 U20475 ( .B1(n17508), .B2(n17431), .A(n17265), .ZN(P3_U2685) );
  AOI22_X1 U20476 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17355), .ZN(n17269) );
  AOI22_X1 U20477 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17387), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17385), .ZN(n17268) );
  AOI22_X1 U20478 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17367), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12550), .ZN(n17267) );
  AOI22_X1 U20479 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17266) );
  NAND4_X1 U20480 ( .A1(n17269), .A2(n17268), .A3(n17267), .A4(n17266), .ZN(
        n17275) );
  AOI22_X1 U20481 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17349), .ZN(n17273) );
  AOI22_X1 U20482 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n12563), .ZN(n17272) );
  AOI22_X1 U20483 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17384), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20484 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17270) );
  NAND4_X1 U20485 ( .A1(n17273), .A2(n17272), .A3(n17271), .A4(n17270), .ZN(
        n17274) );
  NOR2_X1 U20486 ( .A1(n17275), .A2(n17274), .ZN(n17514) );
  INV_X1 U20487 ( .A(n17276), .ZN(n17278) );
  OAI21_X1 U20488 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17278), .A(n17277), .ZN(
        n17279) );
  OAI21_X1 U20489 ( .B1(n17514), .B2(n17431), .A(n17279), .ZN(P3_U2686) );
  AOI22_X1 U20490 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20491 ( .A1(n12576), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20492 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20493 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17280) );
  NAND4_X1 U20494 ( .A1(n17283), .A2(n17282), .A3(n17281), .A4(n17280), .ZN(
        n17289) );
  AOI22_X1 U20495 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20496 ( .A1(n12585), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12581), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20497 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20498 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17284) );
  NAND4_X1 U20499 ( .A1(n17287), .A2(n17286), .A3(n17285), .A4(n17284), .ZN(
        n17288) );
  NOR2_X1 U20500 ( .A1(n17289), .A2(n17288), .ZN(n17521) );
  AOI21_X1 U20501 ( .B1(n17290), .B2(n17318), .A(n17435), .ZN(n17306) );
  NOR4_X1 U20502 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17564), .A3(n17403), .A4(
        n17413), .ZN(n17291) );
  AOI22_X1 U20503 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17306), .B1(n17292), 
        .B2(n17291), .ZN(n17293) );
  OAI21_X1 U20504 ( .B1(n17521), .B2(n17431), .A(n17293), .ZN(P3_U2687) );
  AOI22_X1 U20505 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20506 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20507 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20508 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17294) );
  NAND4_X1 U20509 ( .A1(n17297), .A2(n17296), .A3(n17295), .A4(n17294), .ZN(
        n17303) );
  AOI22_X1 U20510 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20511 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20512 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20513 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17298) );
  NAND4_X1 U20514 ( .A1(n17301), .A2(n17300), .A3(n17299), .A4(n17298), .ZN(
        n17302) );
  NOR2_X1 U20515 ( .A1(n17303), .A2(n17302), .ZN(n17526) );
  NOR2_X1 U20516 ( .A1(n17305), .A2(n17304), .ZN(n17320) );
  OAI21_X1 U20517 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17320), .A(n17306), .ZN(
        n17307) );
  OAI21_X1 U20518 ( .B1(n17526), .B2(n17431), .A(n17307), .ZN(P3_U2688) );
  AOI22_X1 U20519 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U20520 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U20521 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17308) );
  OAI21_X1 U20522 ( .B1(n12541), .B2(n17415), .A(n17308), .ZN(n17314) );
  AOI22_X1 U20523 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U20524 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U20525 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20526 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17368), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17309) );
  NAND4_X1 U20527 ( .A1(n17312), .A2(n17311), .A3(n17310), .A4(n17309), .ZN(
        n17313) );
  AOI211_X1 U20528 ( .C1(n17394), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17314), .B(n17313), .ZN(n17315) );
  NAND3_X1 U20529 ( .A1(n17317), .A2(n17316), .A3(n17315), .ZN(n17532) );
  INV_X1 U20530 ( .A(n17532), .ZN(n17321) );
  OAI21_X1 U20531 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17318), .A(n17431), .ZN(
        n17319) );
  OAI22_X1 U20532 ( .A1(n17321), .A2(n17431), .B1(n17320), .B2(n17319), .ZN(
        P3_U2689) );
  AOI22_X1 U20533 ( .A1(n12583), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20534 ( .A1(n17387), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U20535 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12550), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20536 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17322) );
  NAND4_X1 U20537 ( .A1(n17325), .A2(n17324), .A3(n17323), .A4(n17322), .ZN(
        n17331) );
  AOI22_X1 U20538 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20539 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20540 ( .A1(n12574), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12697), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U20541 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17326) );
  NAND4_X1 U20542 ( .A1(n17329), .A2(n17328), .A3(n17327), .A4(n17326), .ZN(
        n17330) );
  NOR2_X1 U20543 ( .A1(n17331), .A2(n17330), .ZN(n17542) );
  INV_X1 U20544 ( .A(n17381), .ZN(n17363) );
  NAND2_X1 U20545 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17363), .ZN(n17362) );
  NOR2_X1 U20546 ( .A1(n17345), .A2(n17362), .ZN(n17344) );
  OAI21_X1 U20547 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17344), .A(n17431), .ZN(
        n17332) );
  OAI22_X1 U20548 ( .A1(n17542), .A2(n17431), .B1(n17333), .B2(n17332), .ZN(
        P3_U2691) );
  AOI22_X1 U20549 ( .A1(n12697), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U20550 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17342) );
  INV_X1 U20551 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20552 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9648), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17334) );
  OAI21_X1 U20553 ( .B1(n12541), .B2(n17428), .A(n17334), .ZN(n17340) );
  AOI22_X1 U20554 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20555 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U20556 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20557 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17386), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17335) );
  NAND4_X1 U20558 ( .A1(n17338), .A2(n17337), .A3(n17336), .A4(n17335), .ZN(
        n17339) );
  AOI211_X1 U20559 ( .C1(n17366), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n17340), .B(n17339), .ZN(n17341) );
  NAND3_X1 U20560 ( .A1(n17343), .A2(n17342), .A3(n17341), .ZN(n17546) );
  INV_X1 U20561 ( .A(n17344), .ZN(n17347) );
  AOI21_X1 U20562 ( .B1(n17345), .B2(n17362), .A(n17435), .ZN(n17346) );
  AOI22_X1 U20563 ( .A1(n17546), .A2(n17435), .B1(n17347), .B2(n17346), .ZN(
        n17348) );
  INV_X1 U20564 ( .A(n17348), .ZN(P3_U2692) );
  AOI22_X1 U20565 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17349), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17354) );
  AOI22_X1 U20566 ( .A1(n17350), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20567 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20568 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17367), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17351) );
  NAND4_X1 U20569 ( .A1(n17354), .A2(n17353), .A3(n17352), .A4(n17351), .ZN(
        n17361) );
  AOI22_X1 U20570 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20571 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U20572 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20573 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17356) );
  NAND4_X1 U20574 ( .A1(n17359), .A2(n17358), .A3(n17357), .A4(n17356), .ZN(
        n17360) );
  NOR2_X1 U20575 ( .A1(n17361), .A2(n17360), .ZN(n17549) );
  OAI21_X1 U20576 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17363), .A(n17362), .ZN(
        n17364) );
  AOI22_X1 U20577 ( .A1(n17435), .A2(n17549), .B1(n17364), .B2(n17431), .ZN(
        P3_U2693) );
  AOI22_X1 U20578 ( .A1(n17366), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17365), .ZN(n17373) );
  AOI22_X1 U20579 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12550), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17367), .ZN(n17372) );
  AOI22_X1 U20580 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17368), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17386), .ZN(n17371) );
  AOI22_X1 U20581 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17369), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17387), .ZN(n17370) );
  NAND4_X1 U20582 ( .A1(n17373), .A2(n17372), .A3(n17371), .A4(n17370), .ZN(
        n17380) );
  AOI22_X1 U20583 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12574), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17384), .ZN(n17378) );
  AOI22_X1 U20584 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17355), .ZN(n17377) );
  AOI22_X1 U20585 ( .A1(n12583), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17393), .ZN(n17376) );
  AOI22_X1 U20586 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17395), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17375) );
  NAND4_X1 U20587 ( .A1(n17378), .A2(n17377), .A3(n17376), .A4(n17375), .ZN(
        n17379) );
  NOR2_X1 U20588 ( .A1(n17380), .A2(n17379), .ZN(n17554) );
  AND2_X1 U20589 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17402), .ZN(n17382) );
  OAI21_X1 U20590 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17382), .A(n17381), .ZN(
        n17383) );
  AOI22_X1 U20591 ( .A1(n17435), .A2(n17554), .B1(n17383), .B2(n17431), .ZN(
        P3_U2694) );
  AOI22_X1 U20592 ( .A1(n12563), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20593 ( .A1(n17386), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20594 ( .A1(n12602), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17387), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20595 ( .A1(n12550), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17388), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17389) );
  NAND4_X1 U20596 ( .A1(n17392), .A2(n17391), .A3(n17390), .A4(n17389), .ZN(
        n17401) );
  AOI22_X1 U20597 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20598 ( .A1(n17349), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U20599 ( .A1(n9650), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12574), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20600 ( .A1(n17395), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17365), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17396) );
  NAND4_X1 U20601 ( .A1(n17399), .A2(n17398), .A3(n17397), .A4(n17396), .ZN(
        n17400) );
  NOR2_X1 U20602 ( .A1(n17401), .A2(n17400), .ZN(n17562) );
  NOR2_X1 U20603 ( .A1(n17435), .A2(n17402), .ZN(n17407) );
  NOR3_X1 U20604 ( .A1(n17564), .A2(n17403), .A3(n17413), .ZN(n17405) );
  AOI22_X1 U20605 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17407), .B1(n17405), .B2(
        n17404), .ZN(n17406) );
  OAI21_X1 U20606 ( .B1(n17562), .B2(n17431), .A(n17406), .ZN(P3_U2695) );
  INV_X1 U20607 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17410) );
  INV_X1 U20608 ( .A(n17413), .ZN(n17408) );
  OAI21_X1 U20609 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17408), .A(n17407), .ZN(
        n17409) );
  OAI21_X1 U20610 ( .B1(n17431), .B2(n17410), .A(n17409), .ZN(P3_U2696) );
  INV_X1 U20611 ( .A(n17411), .ZN(n17412) );
  NOR2_X1 U20612 ( .A1(n17412), .A2(n17439), .ZN(n17426) );
  OAI221_X1 U20613 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(P3_EBX_REG_5__SCAN_IN), 
        .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17426), .A(n17413), .ZN(n17414) );
  AOI22_X1 U20614 ( .A1(n17435), .A2(n17415), .B1(n17414), .B2(n17431), .ZN(
        P3_U2697) );
  INV_X1 U20615 ( .A(n17416), .ZN(n17420) );
  AOI21_X1 U20616 ( .B1(n17418), .B2(n17417), .A(n17435), .ZN(n17419) );
  AOI22_X1 U20617 ( .A1(n17420), .A2(n17419), .B1(
        P3_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n17435), .ZN(n17421) );
  INV_X1 U20618 ( .A(n17421), .ZN(P3_U2698) );
  NOR3_X1 U20619 ( .A1(n17423), .A2(n17422), .A3(n17439), .ZN(n17430) );
  AOI21_X1 U20620 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17431), .A(n17430), .ZN(
        n17425) );
  OAI22_X1 U20621 ( .A1(n17426), .A2(n17425), .B1(n17424), .B2(n17431), .ZN(
        P3_U2699) );
  AOI21_X1 U20622 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17431), .A(n17427), .ZN(
        n17429) );
  OAI22_X1 U20623 ( .A1(n17430), .A2(n17429), .B1(n17428), .B2(n17431), .ZN(
        P3_U2700) );
  INV_X1 U20624 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17432) );
  OAI222_X1 U20625 ( .A1(n17434), .A2(n17439), .B1(n17433), .B2(n17437), .C1(
        n17432), .C2(n17431), .ZN(P3_U2702) );
  NAND2_X1 U20626 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17435), .ZN(
        n17436) );
  OAI221_X1 U20627 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17439), .C1(n17438), 
        .C2(n17437), .A(n17436), .ZN(P3_U2703) );
  INV_X1 U20628 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17666) );
  INV_X1 U20629 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17662) );
  INV_X1 U20630 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17707) );
  INV_X1 U20631 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17682) );
  INV_X1 U20632 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17680) );
  NAND4_X1 U20633 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n17440) );
  NOR3_X1 U20634 ( .A1(n17682), .A2(n17680), .A3(n17440), .ZN(n17441) );
  NAND3_X1 U20635 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(n17441), .ZN(n17523) );
  INV_X1 U20636 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17688) );
  NAND2_X1 U20637 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n17530) );
  NAND4_X1 U20638 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .A4(P3_EAX_REG_11__SCAN_IN), .ZN(n17442)
         );
  NOR3_X1 U20639 ( .A1(n17688), .A2(n17530), .A3(n17442), .ZN(n17524) );
  NAND2_X1 U20640 ( .A1(n17559), .A2(n17524), .ZN(n17525) );
  INV_X1 U20641 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17654) );
  INV_X1 U20642 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17652) );
  NAND4_X1 U20643 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17443)
         );
  NAND2_X1 U20644 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17482), .ZN(n17481) );
  NAND2_X1 U20645 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17477), .ZN(n17476) );
  NAND2_X1 U20646 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17458), .ZN(n17453) );
  NAND2_X1 U20647 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17449), .ZN(n17448) );
  NAND2_X1 U20648 ( .A1(n17448), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17446) );
  NAND2_X1 U20649 ( .A1(n17444), .A2(n17598), .ZN(n17491) );
  NAND2_X1 U20650 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17515), .ZN(n17445) );
  OAI221_X1 U20651 ( .B1(n17448), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17446), 
        .C2(n17598), .A(n17445), .ZN(P3_U2704) );
  NOR2_X2 U20652 ( .A1(n17447), .A2(n17585), .ZN(n17516) );
  AOI22_X1 U20653 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17515), .ZN(n17451) );
  OAI211_X1 U20654 ( .C1(n17449), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17585), .B(
        n17448), .ZN(n17450) );
  OAI211_X1 U20655 ( .C1(n17452), .C2(n17587), .A(n17451), .B(n17450), .ZN(
        P3_U2705) );
  AOI22_X1 U20656 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17515), .ZN(n17455) );
  OAI211_X1 U20657 ( .C1(n17458), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17585), .B(
        n17453), .ZN(n17454) );
  OAI211_X1 U20658 ( .C1(n17456), .C2(n17587), .A(n17455), .B(n17454), .ZN(
        P3_U2706) );
  INV_X1 U20659 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19478) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17516), .B1(n17594), .B2(
        n17457), .ZN(n17461) );
  AOI211_X1 U20661 ( .C1(n17666), .C2(n17462), .A(n17458), .B(n17598), .ZN(
        n17459) );
  INV_X1 U20662 ( .A(n17459), .ZN(n17460) );
  OAI211_X1 U20663 ( .C1(n17491), .C2(n19478), .A(n17461), .B(n17460), .ZN(
        P3_U2707) );
  AOI22_X1 U20664 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17515), .ZN(n17464) );
  OAI211_X1 U20665 ( .C1(n17467), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17585), .B(
        n17462), .ZN(n17463) );
  OAI211_X1 U20666 ( .C1(n17465), .C2(n17587), .A(n17464), .B(n17463), .ZN(
        P3_U2708) );
  INV_X1 U20667 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18421) );
  AOI22_X1 U20668 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17516), .B1(n17594), .B2(
        n17466), .ZN(n17470) );
  AOI211_X1 U20669 ( .C1(n17662), .C2(n17471), .A(n17467), .B(n17598), .ZN(
        n17468) );
  INV_X1 U20670 ( .A(n17468), .ZN(n17469) );
  OAI211_X1 U20671 ( .C1(n17491), .C2(n18421), .A(n17470), .B(n17469), .ZN(
        P3_U2709) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17515), .ZN(n17474) );
  OAI211_X1 U20673 ( .C1(n17472), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17585), .B(
        n17471), .ZN(n17473) );
  OAI211_X1 U20674 ( .C1(n17475), .C2(n17587), .A(n17474), .B(n17473), .ZN(
        P3_U2710) );
  AOI22_X1 U20675 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17515), .ZN(n17479) );
  OAI211_X1 U20676 ( .C1(n17477), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17585), .B(
        n17476), .ZN(n17478) );
  OAI211_X1 U20677 ( .C1(n17480), .C2(n17587), .A(n17479), .B(n17478), .ZN(
        P3_U2711) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17515), .ZN(n17484) );
  OAI211_X1 U20679 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17482), .A(n17585), .B(
        n17481), .ZN(n17483) );
  OAI211_X1 U20680 ( .C1(n17485), .C2(n17587), .A(n17484), .B(n17483), .ZN(
        P3_U2712) );
  INV_X1 U20681 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17648) );
  INV_X1 U20682 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17644) );
  NAND2_X1 U20683 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17509), .ZN(n17505) );
  NAND2_X1 U20684 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17500), .ZN(n17496) );
  NAND2_X1 U20685 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17654), .ZN(n17490) );
  AOI22_X1 U20686 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17515), .B1(n17594), .B2(
        n17486), .ZN(n17489) );
  NAND2_X1 U20687 ( .A1(n17585), .A2(n17496), .ZN(n17495) );
  OAI21_X1 U20688 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17522), .A(n17495), .ZN(
        n17487) );
  AOI22_X1 U20689 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17516), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17487), .ZN(n17488) );
  OAI211_X1 U20690 ( .C1(n17496), .C2(n17490), .A(n17489), .B(n17488), .ZN(
        P3_U2713) );
  INV_X1 U20691 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19483) );
  OAI22_X1 U20692 ( .A1(n17492), .A2(n17587), .B1(n19483), .B2(n17491), .ZN(
        n17493) );
  AOI21_X1 U20693 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17516), .A(n17493), .ZN(
        n17494) );
  OAI221_X1 U20694 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17496), .C1(n17652), 
        .C2(n17495), .A(n17494), .ZN(P3_U2714) );
  AOI22_X1 U20695 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17515), .ZN(n17498) );
  OAI211_X1 U20696 ( .C1(n17500), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17585), .B(
        n17496), .ZN(n17497) );
  OAI211_X1 U20697 ( .C1(n17499), .C2(n17587), .A(n17498), .B(n17497), .ZN(
        P3_U2715) );
  AOI22_X1 U20698 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17515), .ZN(n17503) );
  AOI211_X1 U20699 ( .C1(n17648), .C2(n17505), .A(n17500), .B(n17598), .ZN(
        n17501) );
  INV_X1 U20700 ( .A(n17501), .ZN(n17502) );
  OAI211_X1 U20701 ( .C1(n17504), .C2(n17587), .A(n17503), .B(n17502), .ZN(
        P3_U2716) );
  AOI22_X1 U20702 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17515), .ZN(n17507) );
  OAI211_X1 U20703 ( .C1(n17509), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17585), .B(
        n17505), .ZN(n17506) );
  OAI211_X1 U20704 ( .C1(n17508), .C2(n17587), .A(n17507), .B(n17506), .ZN(
        P3_U2717) );
  AOI22_X1 U20705 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17515), .ZN(n17513) );
  INV_X1 U20706 ( .A(n17517), .ZN(n17511) );
  INV_X1 U20707 ( .A(n17509), .ZN(n17510) );
  OAI211_X1 U20708 ( .C1(n17511), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17585), .B(
        n17510), .ZN(n17512) );
  OAI211_X1 U20709 ( .C1(n17514), .C2(n17587), .A(n17513), .B(n17512), .ZN(
        P3_U2718) );
  AOI22_X1 U20710 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17516), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17515), .ZN(n17520) );
  OAI211_X1 U20711 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17518), .A(n17585), .B(
        n17517), .ZN(n17519) );
  OAI211_X1 U20712 ( .C1(n17521), .C2(n17587), .A(n17520), .B(n17519), .ZN(
        P3_U2719) );
  NAND2_X1 U20713 ( .A1(n17524), .A2(n17567), .ZN(n17529) );
  NAND2_X1 U20714 ( .A1(n17585), .A2(n17525), .ZN(n17534) );
  INV_X1 U20715 ( .A(n17526), .ZN(n17527) );
  AOI22_X1 U20716 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17595), .B1(n17594), .B2(
        n17527), .ZN(n17528) );
  OAI221_X1 U20717 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17529), .C1(n17707), 
        .C2(n17534), .A(n17528), .ZN(P3_U2720) );
  NAND2_X1 U20718 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n17531) );
  INV_X1 U20719 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17694) );
  NAND2_X1 U20720 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17567), .ZN(n17558) );
  NOR2_X1 U20721 ( .A1(n17694), .A2(n17548), .ZN(n17541) );
  INV_X1 U20722 ( .A(n17541), .ZN(n17536) );
  NOR2_X1 U20723 ( .A1(n17531), .A2(n17536), .ZN(n17538) );
  INV_X1 U20724 ( .A(n17538), .ZN(n17535) );
  INV_X1 U20725 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17702) );
  AOI22_X1 U20726 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17595), .B1(n17594), .B2(
        n17532), .ZN(n17533) );
  OAI221_X1 U20727 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17535), .C1(n17702), 
        .C2(n17534), .A(n17533), .ZN(P3_U2721) );
  INV_X1 U20728 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17540) );
  INV_X1 U20729 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17698) );
  NOR2_X1 U20730 ( .A1(n17698), .A2(n17536), .ZN(n17544) );
  AOI21_X1 U20731 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17585), .A(n17544), .ZN(
        n17539) );
  OAI222_X1 U20732 ( .A1(n17590), .A2(n17540), .B1(n17539), .B2(n17538), .C1(
        n17587), .C2(n17537), .ZN(P3_U2722) );
  INV_X1 U20733 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17545) );
  AOI21_X1 U20734 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17585), .A(n17541), .ZN(
        n17543) );
  OAI222_X1 U20735 ( .A1(n17590), .A2(n17545), .B1(n17544), .B2(n17543), .C1(
        n17587), .C2(n17542), .ZN(P3_U2723) );
  NAND2_X1 U20736 ( .A1(n17585), .A2(n17548), .ZN(n17551) );
  AOI22_X1 U20737 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17595), .B1(n17594), .B2(
        n17546), .ZN(n17547) );
  OAI221_X1 U20738 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17548), .C1(n17694), 
        .C2(n17551), .A(n17547), .ZN(P3_U2724) );
  INV_X1 U20739 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17552) );
  INV_X1 U20740 ( .A(n17558), .ZN(n17553) );
  AOI21_X1 U20741 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17553), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n17550) );
  OAI222_X1 U20742 ( .A1(n17590), .A2(n17552), .B1(n17551), .B2(n17550), .C1(
        n17587), .C2(n17549), .ZN(P3_U2725) );
  INV_X1 U20743 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17557) );
  INV_X1 U20744 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17690) );
  NOR2_X1 U20745 ( .A1(n17690), .A2(n17558), .ZN(n17556) );
  AOI21_X1 U20746 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17585), .A(n17553), .ZN(
        n17555) );
  OAI222_X1 U20747 ( .A1(n17590), .A2(n17557), .B1(n17556), .B2(n17555), .C1(
        n17587), .C2(n17554), .ZN(P3_U2726) );
  NAND2_X1 U20748 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17595), .ZN(n17561) );
  OAI211_X1 U20749 ( .C1(n17559), .C2(P3_EAX_REG_8__SCAN_IN), .A(n17585), .B(
        n17558), .ZN(n17560) );
  OAI211_X1 U20750 ( .C1(n17562), .C2(n17587), .A(n17561), .B(n17560), .ZN(
        P3_U2727) );
  INV_X1 U20751 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18445) );
  INV_X1 U20752 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17684) );
  INV_X1 U20753 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17674) );
  NOR4_X1 U20754 ( .A1(n17564), .A2(n17563), .A3(n17674), .A4(n17672), .ZN(
        n17584) );
  AND2_X1 U20755 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17584), .ZN(n17589) );
  NAND2_X1 U20756 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17589), .ZN(n17576) );
  NOR2_X1 U20757 ( .A1(n17680), .A2(n17576), .ZN(n17580) );
  NAND2_X1 U20758 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17580), .ZN(n17568) );
  NOR2_X1 U20759 ( .A1(n17684), .A2(n17568), .ZN(n17572) );
  AOI21_X1 U20760 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17585), .A(n17572), .ZN(
        n17566) );
  OAI222_X1 U20761 ( .A1(n17590), .A2(n18445), .B1(n17567), .B2(n17566), .C1(
        n17587), .C2(n17565), .ZN(P3_U2728) );
  INV_X1 U20762 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18440) );
  INV_X1 U20763 ( .A(n17568), .ZN(n17575) );
  AOI21_X1 U20764 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17585), .A(n17575), .ZN(
        n17571) );
  INV_X1 U20765 ( .A(n17569), .ZN(n17570) );
  OAI222_X1 U20766 ( .A1(n18440), .A2(n17590), .B1(n17572), .B2(n17571), .C1(
        n17587), .C2(n17570), .ZN(P3_U2729) );
  INV_X1 U20767 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18435) );
  AOI21_X1 U20768 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17585), .A(n17580), .ZN(
        n17574) );
  OAI222_X1 U20769 ( .A1(n18435), .A2(n17590), .B1(n17575), .B2(n17574), .C1(
        n17587), .C2(n17573), .ZN(P3_U2730) );
  INV_X1 U20770 ( .A(n17576), .ZN(n17583) );
  AOI21_X1 U20771 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17585), .A(n17583), .ZN(
        n17579) );
  INV_X1 U20772 ( .A(n17577), .ZN(n17578) );
  OAI222_X1 U20773 ( .A1(n18431), .A2(n17590), .B1(n17580), .B2(n17579), .C1(
        n17587), .C2(n17578), .ZN(P3_U2731) );
  INV_X1 U20774 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18426) );
  AOI21_X1 U20775 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17585), .A(n17589), .ZN(
        n17582) );
  OAI222_X1 U20776 ( .A1(n18426), .A2(n17590), .B1(n17583), .B2(n17582), .C1(
        n17587), .C2(n17581), .ZN(P3_U2732) );
  INV_X1 U20777 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18422) );
  AOI21_X1 U20778 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17585), .A(n17584), .ZN(
        n17588) );
  OAI222_X1 U20779 ( .A1(n18422), .A2(n17590), .B1(n17589), .B2(n17588), .C1(
        n17587), .C2(n17586), .ZN(P3_U2733) );
  NAND2_X1 U20780 ( .A1(n17591), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17592) );
  XNOR2_X1 U20781 ( .A(n17674), .B(n17592), .ZN(n17597) );
  AOI22_X1 U20782 ( .A1(n17595), .A2(BUF2_REG_1__SCAN_IN), .B1(n17594), .B2(
        n17593), .ZN(n17596) );
  OAI21_X1 U20783 ( .B1(n17598), .B2(n17597), .A(n17596), .ZN(P3_U2734) );
  NOR2_X1 U20784 ( .A1(n19049), .A2(n18937), .ZN(n19071) );
  AND2_X1 U20785 ( .A1(n17615), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20786 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17670) );
  NAND2_X1 U20787 ( .A1(n17618), .A2(n17600), .ZN(n17617) );
  AOI22_X1 U20788 ( .A1(n19071), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17634), .ZN(n17601) );
  OAI21_X1 U20789 ( .B1(n17670), .B2(n17617), .A(n17601), .ZN(P3_U2737) );
  INV_X1 U20790 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U20791 ( .A1(n19071), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17602) );
  OAI21_X1 U20792 ( .B1(n17668), .B2(n17617), .A(n17602), .ZN(P3_U2738) );
  AOI22_X1 U20793 ( .A1(n19071), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17603) );
  OAI21_X1 U20794 ( .B1(n17666), .B2(n17617), .A(n17603), .ZN(P3_U2739) );
  INV_X1 U20795 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U20796 ( .A1(n19071), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17604) );
  OAI21_X1 U20797 ( .B1(n17664), .B2(n17617), .A(n17604), .ZN(P3_U2740) );
  AOI22_X1 U20798 ( .A1(n19071), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17605) );
  OAI21_X1 U20799 ( .B1(n17662), .B2(n17617), .A(n17605), .ZN(P3_U2741) );
  INV_X1 U20800 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17660) );
  AOI22_X1 U20801 ( .A1(n19071), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17606) );
  OAI21_X1 U20802 ( .B1(n17660), .B2(n17617), .A(n17606), .ZN(P3_U2742) );
  INV_X1 U20803 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17658) );
  AOI22_X1 U20804 ( .A1(n19071), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17607) );
  OAI21_X1 U20805 ( .B1(n17658), .B2(n17617), .A(n17607), .ZN(P3_U2743) );
  INV_X1 U20806 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17656) );
  CLKBUF_X1 U20807 ( .A(n19071), .Z(n17635) );
  AOI22_X1 U20808 ( .A1(n17635), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17608) );
  OAI21_X1 U20809 ( .B1(n17656), .B2(n17617), .A(n17608), .ZN(P3_U2744) );
  AOI22_X1 U20810 ( .A1(n17635), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17609) );
  OAI21_X1 U20811 ( .B1(n17654), .B2(n17617), .A(n17609), .ZN(P3_U2745) );
  AOI22_X1 U20812 ( .A1(n17635), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17610) );
  OAI21_X1 U20813 ( .B1(n17652), .B2(n17617), .A(n17610), .ZN(P3_U2746) );
  INV_X1 U20814 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U20815 ( .A1(n17635), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17611) );
  OAI21_X1 U20816 ( .B1(n17650), .B2(n17617), .A(n17611), .ZN(P3_U2747) );
  AOI22_X1 U20817 ( .A1(n17635), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17612) );
  OAI21_X1 U20818 ( .B1(n17648), .B2(n17617), .A(n17612), .ZN(P3_U2748) );
  INV_X1 U20819 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17646) );
  AOI22_X1 U20820 ( .A1(n17635), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17613) );
  OAI21_X1 U20821 ( .B1(n17646), .B2(n17617), .A(n17613), .ZN(P3_U2749) );
  AOI22_X1 U20822 ( .A1(n17635), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17614) );
  OAI21_X1 U20823 ( .B1(n17644), .B2(n17617), .A(n17614), .ZN(P3_U2750) );
  INV_X1 U20824 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17642) );
  AOI22_X1 U20825 ( .A1(n17635), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17615), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17616) );
  OAI21_X1 U20826 ( .B1(n17642), .B2(n17617), .A(n17616), .ZN(P3_U2751) );
  AOI22_X1 U20827 ( .A1(n17635), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U20828 ( .B1(n17707), .B2(n17637), .A(n17619), .ZN(P3_U2752) );
  AOI22_X1 U20829 ( .A1(n17635), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17620) );
  OAI21_X1 U20830 ( .B1(n17702), .B2(n17637), .A(n17620), .ZN(P3_U2753) );
  INV_X1 U20831 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17700) );
  AOI22_X1 U20832 ( .A1(n17635), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17621) );
  OAI21_X1 U20833 ( .B1(n17700), .B2(n17637), .A(n17621), .ZN(P3_U2754) );
  AOI22_X1 U20834 ( .A1(n17635), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17622) );
  OAI21_X1 U20835 ( .B1(n17698), .B2(n17637), .A(n17622), .ZN(P3_U2755) );
  AOI22_X1 U20836 ( .A1(n17635), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17623) );
  OAI21_X1 U20837 ( .B1(n17694), .B2(n17637), .A(n17623), .ZN(P3_U2756) );
  INV_X1 U20838 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17692) );
  AOI22_X1 U20839 ( .A1(n17635), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17624) );
  OAI21_X1 U20840 ( .B1(n17692), .B2(n17637), .A(n17624), .ZN(P3_U2757) );
  AOI22_X1 U20841 ( .A1(n17635), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17625) );
  OAI21_X1 U20842 ( .B1(n17690), .B2(n17637), .A(n17625), .ZN(P3_U2758) );
  AOI22_X1 U20843 ( .A1(n17635), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17626) );
  OAI21_X1 U20844 ( .B1(n17688), .B2(n17637), .A(n17626), .ZN(P3_U2759) );
  INV_X1 U20845 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U20846 ( .A1(n17635), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17627) );
  OAI21_X1 U20847 ( .B1(n17686), .B2(n17637), .A(n17627), .ZN(P3_U2760) );
  AOI22_X1 U20848 ( .A1(n17635), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17628) );
  OAI21_X1 U20849 ( .B1(n17684), .B2(n17637), .A(n17628), .ZN(P3_U2761) );
  AOI22_X1 U20850 ( .A1(n17635), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17629) );
  OAI21_X1 U20851 ( .B1(n17682), .B2(n17637), .A(n17629), .ZN(P3_U2762) );
  AOI22_X1 U20852 ( .A1(n17635), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17630) );
  OAI21_X1 U20853 ( .B1(n17680), .B2(n17637), .A(n17630), .ZN(P3_U2763) );
  INV_X1 U20854 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U20855 ( .A1(n17635), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17631) );
  OAI21_X1 U20856 ( .B1(n17678), .B2(n17637), .A(n17631), .ZN(P3_U2764) );
  INV_X1 U20857 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17676) );
  AOI22_X1 U20858 ( .A1(n17635), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17632) );
  OAI21_X1 U20859 ( .B1(n17676), .B2(n17637), .A(n17632), .ZN(P3_U2765) );
  AOI22_X1 U20860 ( .A1(n17635), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17633) );
  OAI21_X1 U20861 ( .B1(n17674), .B2(n17637), .A(n17633), .ZN(P3_U2766) );
  AOI22_X1 U20862 ( .A1(n17635), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17634), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17636) );
  OAI21_X1 U20863 ( .B1(n17672), .B2(n17637), .A(n17636), .ZN(P3_U2767) );
  NAND2_X1 U20864 ( .A1(n19074), .A2(n17640), .ZN(n18917) );
  AOI22_X1 U20865 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17695), .ZN(n17641) );
  OAI21_X1 U20866 ( .B1(n17642), .B2(n17706), .A(n17641), .ZN(P3_U2768) );
  AOI22_X1 U20867 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17695), .ZN(n17643) );
  OAI21_X1 U20868 ( .B1(n17644), .B2(n17706), .A(n17643), .ZN(P3_U2769) );
  AOI22_X1 U20869 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17695), .ZN(n17645) );
  OAI21_X1 U20870 ( .B1(n17646), .B2(n17706), .A(n17645), .ZN(P3_U2770) );
  AOI22_X1 U20871 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17695), .ZN(n17647) );
  OAI21_X1 U20872 ( .B1(n17648), .B2(n17706), .A(n17647), .ZN(P3_U2771) );
  AOI22_X1 U20873 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17695), .ZN(n17649) );
  OAI21_X1 U20874 ( .B1(n17650), .B2(n17706), .A(n17649), .ZN(P3_U2772) );
  AOI22_X1 U20875 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17695), .ZN(n17651) );
  OAI21_X1 U20876 ( .B1(n17652), .B2(n17706), .A(n17651), .ZN(P3_U2773) );
  AOI22_X1 U20877 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17695), .ZN(n17653) );
  OAI21_X1 U20878 ( .B1(n17654), .B2(n17706), .A(n17653), .ZN(P3_U2774) );
  AOI22_X1 U20879 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17695), .ZN(n17655) );
  OAI21_X1 U20880 ( .B1(n17656), .B2(n17706), .A(n17655), .ZN(P3_U2775) );
  AOI22_X1 U20881 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17695), .ZN(n17657) );
  OAI21_X1 U20882 ( .B1(n17658), .B2(n17706), .A(n17657), .ZN(P3_U2776) );
  AOI22_X1 U20883 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17695), .ZN(n17659) );
  OAI21_X1 U20884 ( .B1(n17660), .B2(n17706), .A(n17659), .ZN(P3_U2777) );
  AOI22_X1 U20885 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17695), .ZN(n17661) );
  OAI21_X1 U20886 ( .B1(n17662), .B2(n17706), .A(n17661), .ZN(P3_U2778) );
  AOI22_X1 U20887 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17696), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17703), .ZN(n17663) );
  OAI21_X1 U20888 ( .B1(n17664), .B2(n17706), .A(n17663), .ZN(P3_U2779) );
  AOI22_X1 U20889 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17695), .ZN(n17665) );
  OAI21_X1 U20890 ( .B1(n17666), .B2(n17706), .A(n17665), .ZN(P3_U2780) );
  AOI22_X1 U20891 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17695), .ZN(n17667) );
  OAI21_X1 U20892 ( .B1(n17668), .B2(n17706), .A(n17667), .ZN(P3_U2781) );
  AOI22_X1 U20893 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17695), .ZN(n17669) );
  OAI21_X1 U20894 ( .B1(n17670), .B2(n17706), .A(n17669), .ZN(P3_U2782) );
  AOI22_X1 U20895 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17695), .ZN(n17671) );
  OAI21_X1 U20896 ( .B1(n17672), .B2(n17706), .A(n17671), .ZN(P3_U2783) );
  AOI22_X1 U20897 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17695), .ZN(n17673) );
  OAI21_X1 U20898 ( .B1(n17674), .B2(n17706), .A(n17673), .ZN(P3_U2784) );
  AOI22_X1 U20899 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17695), .ZN(n17675) );
  OAI21_X1 U20900 ( .B1(n17676), .B2(n17706), .A(n17675), .ZN(P3_U2785) );
  AOI22_X1 U20901 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17695), .ZN(n17677) );
  OAI21_X1 U20902 ( .B1(n17678), .B2(n17706), .A(n17677), .ZN(P3_U2786) );
  AOI22_X1 U20903 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17695), .ZN(n17679) );
  OAI21_X1 U20904 ( .B1(n17680), .B2(n17706), .A(n17679), .ZN(P3_U2787) );
  AOI22_X1 U20905 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17703), .ZN(n17681) );
  OAI21_X1 U20906 ( .B1(n17682), .B2(n17706), .A(n17681), .ZN(P3_U2788) );
  AOI22_X1 U20907 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17703), .ZN(n17683) );
  OAI21_X1 U20908 ( .B1(n17684), .B2(n17706), .A(n17683), .ZN(P3_U2789) );
  AOI22_X1 U20909 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17703), .ZN(n17685) );
  OAI21_X1 U20910 ( .B1(n17686), .B2(n17706), .A(n17685), .ZN(P3_U2790) );
  AOI22_X1 U20911 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17703), .ZN(n17687) );
  OAI21_X1 U20912 ( .B1(n17688), .B2(n17706), .A(n17687), .ZN(P3_U2791) );
  AOI22_X1 U20913 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17703), .ZN(n17689) );
  OAI21_X1 U20914 ( .B1(n17690), .B2(n17706), .A(n17689), .ZN(P3_U2792) );
  AOI22_X1 U20915 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17696), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17695), .ZN(n17691) );
  OAI21_X1 U20916 ( .B1(n17692), .B2(n17706), .A(n17691), .ZN(P3_U2793) );
  AOI22_X1 U20917 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17703), .ZN(n17693) );
  OAI21_X1 U20918 ( .B1(n17694), .B2(n17706), .A(n17693), .ZN(P3_U2794) );
  AOI22_X1 U20919 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17696), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17695), .ZN(n17697) );
  OAI21_X1 U20920 ( .B1(n17698), .B2(n17706), .A(n17697), .ZN(P3_U2795) );
  AOI22_X1 U20921 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17703), .ZN(n17699) );
  OAI21_X1 U20922 ( .B1(n17700), .B2(n17706), .A(n17699), .ZN(P3_U2796) );
  AOI22_X1 U20923 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17703), .ZN(n17701) );
  OAI21_X1 U20924 ( .B1(n17702), .B2(n17706), .A(n17701), .ZN(P3_U2797) );
  AOI22_X1 U20925 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17703), .ZN(n17705) );
  OAI21_X1 U20926 ( .B1(n17707), .B2(n17706), .A(n17705), .ZN(P3_U2798) );
  INV_X1 U20927 ( .A(n17875), .ZN(n17858) );
  OAI21_X1 U20928 ( .B1(n17708), .B2(n18937), .A(n9676), .ZN(n17709) );
  AOI21_X1 U20929 ( .B1(n17907), .B2(n17711), .A(n17709), .ZN(n17741) );
  OAI21_X1 U20930 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17817), .A(
        n17741), .ZN(n17732) );
  AOI22_X1 U20931 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17732), .B1(
        n17927), .B2(n17710), .ZN(n17714) );
  NOR2_X1 U20932 ( .A1(n17910), .A2(n17711), .ZN(n17734) );
  OAI211_X1 U20933 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17734), .B(n17712), .ZN(n17713) );
  NAND2_X1 U20934 ( .A1(n17714), .A2(n17713), .ZN(n17715) );
  AOI211_X1 U20935 ( .C1(n17858), .C2(n17717), .A(n17716), .B(n17715), .ZN(
        n17724) );
  NOR2_X1 U20936 ( .A1(n18069), .A2(n17945), .ZN(n17823) );
  INV_X1 U20937 ( .A(n17823), .ZN(n17718) );
  AOI22_X1 U20938 ( .A1(n18069), .A2(n18087), .B1(n17945), .B2(n18090), .ZN(
        n17748) );
  NAND2_X1 U20939 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17748), .ZN(
        n17735) );
  NAND3_X1 U20940 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17718), .A3(
        n17735), .ZN(n17723) );
  OAI211_X1 U20941 ( .C1(n17721), .C2(n17720), .A(n17973), .B(n17719), .ZN(
        n17722) );
  NAND3_X1 U20942 ( .A1(n17724), .A2(n17723), .A3(n17722), .ZN(P3_U2802) );
  NAND2_X1 U20943 ( .A1(n17726), .A2(n17725), .ZN(n17729) );
  INV_X1 U20944 ( .A(n17727), .ZN(n17728) );
  AOI21_X1 U20945 ( .B1(n17978), .B2(n17729), .A(n17728), .ZN(n18095) );
  OAI22_X1 U20946 ( .A1(n9655), .A2(n19007), .B1(n17911), .B2(n17730), .ZN(
        n17731) );
  AOI221_X1 U20947 ( .B1(n17734), .B2(n17733), .C1(n17732), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17731), .ZN(n17738) );
  OAI21_X1 U20948 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17736), .A(
        n17735), .ZN(n17737) );
  OAI211_X1 U20949 ( .C1(n18095), .C2(n17991), .A(n17738), .B(n17737), .ZN(
        P3_U2803) );
  NOR2_X1 U20950 ( .A1(n17927), .A2(n17780), .ZN(n18062) );
  AOI21_X1 U20951 ( .B1(n17739), .B2(n18798), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17740) );
  OAI22_X1 U20952 ( .A1(n18062), .A2(n17742), .B1(n17741), .B2(n17740), .ZN(
        n17746) );
  AOI21_X1 U20953 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17744), .A(
        n17743), .ZN(n18101) );
  NAND3_X1 U20954 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18106), .A3(
        n9990), .ZN(n18097) );
  OAI22_X1 U20955 ( .A1(n18101), .A2(n17991), .B1(n17787), .B2(n18097), .ZN(
        n17745) );
  AOI211_X1 U20956 ( .C1(n18393), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17746), 
        .B(n17745), .ZN(n17747) );
  OAI21_X1 U20957 ( .B1(n17748), .B2(n9990), .A(n17747), .ZN(P3_U2804) );
  NAND2_X1 U20958 ( .A1(n18798), .A2(n17757), .ZN(n17775) );
  OAI211_X1 U20959 ( .C1(n17749), .C2(n18937), .A(n9676), .B(n17775), .ZN(
        n17778) );
  AOI22_X1 U20960 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17778), .B1(
        n17927), .B2(n17750), .ZN(n17761) );
  NAND3_X1 U20961 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17764), .A3(
        n17886), .ZN(n17751) );
  XOR2_X1 U20962 ( .A(n17751), .B(n18107), .Z(n18115) );
  NAND3_X1 U20963 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17764), .A3(
        n17885), .ZN(n17752) );
  XOR2_X1 U20964 ( .A(n17752), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18118) );
  OAI21_X1 U20965 ( .B1(n17978), .B2(n17754), .A(n17753), .ZN(n17755) );
  XOR2_X1 U20966 ( .A(n17755), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18113) );
  OAI22_X1 U20967 ( .A1(n18080), .A2(n18118), .B1(n17991), .B2(n18113), .ZN(
        n17756) );
  AOI21_X1 U20968 ( .B1(n17945), .B2(n18115), .A(n17756), .ZN(n17760) );
  NAND2_X1 U20969 ( .A1(n18393), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18111) );
  NOR2_X1 U20970 ( .A1(n17910), .A2(n17757), .ZN(n17763) );
  OAI211_X1 U20971 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17763), .B(n17758), .ZN(n17759) );
  NAND4_X1 U20972 ( .A1(n17761), .A2(n17760), .A3(n18111), .A4(n17759), .ZN(
        P3_U2805) );
  NOR2_X1 U20973 ( .A1(n9655), .A2(n19001), .ZN(n18130) );
  AOI221_X1 U20974 ( .B1(n17763), .B2(n17762), .C1(n17778), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18130), .ZN(n17770) );
  NOR2_X1 U20975 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18139), .ZN(
        n18132) );
  NAND2_X1 U20976 ( .A1(n17885), .A2(n17764), .ZN(n18120) );
  NAND2_X1 U20977 ( .A1(n17886), .A2(n17764), .ZN(n18119) );
  AOI22_X1 U20978 ( .A1(n18069), .A2(n18120), .B1(n17945), .B2(n18119), .ZN(
        n17786) );
  INV_X1 U20979 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18127) );
  AOI21_X1 U20980 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17766), .A(
        n17765), .ZN(n18134) );
  OAI22_X1 U20981 ( .A1(n17786), .A2(n18127), .B1(n18134), .B2(n17991), .ZN(
        n17767) );
  AOI21_X1 U20982 ( .B1(n17768), .B2(n18132), .A(n17767), .ZN(n17769) );
  OAI211_X1 U20983 ( .C1(n17911), .C2(n17771), .A(n17770), .B(n17769), .ZN(
        P3_U2806) );
  AOI22_X1 U20984 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17978), .B1(
        n17772), .B2(n17789), .ZN(n17773) );
  NAND2_X1 U20985 ( .A1(n17824), .A2(n17773), .ZN(n17774) );
  XOR2_X1 U20986 ( .A(n17774), .B(n18139), .Z(n18136) );
  INV_X1 U20987 ( .A(n17775), .ZN(n17776) );
  AOI22_X1 U20988 ( .A1(n18393), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17777), 
        .B2(n17776), .ZN(n17782) );
  OAI221_X1 U20989 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17780), .C1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n17779), .A(n17778), .ZN(
        n17781) );
  OAI211_X1 U20990 ( .C1(n17783), .C2(n17911), .A(n17782), .B(n17781), .ZN(
        n17784) );
  AOI21_X1 U20991 ( .B1(n17973), .B2(n18136), .A(n17784), .ZN(n17785) );
  OAI221_X1 U20992 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17787), 
        .C1(n18139), .C2(n17786), .A(n17785), .ZN(P3_U2807) );
  INV_X1 U20993 ( .A(n17824), .ZN(n17788) );
  AOI221_X1 U20994 ( .B1(n17790), .B2(n17789), .C1(n17809), .C2(n17789), .A(
        n17788), .ZN(n17791) );
  XOR2_X1 U20995 ( .A(n18151), .B(n17791), .Z(n18155) );
  AOI22_X1 U20996 ( .A1(n18069), .A2(n18142), .B1(n17945), .B2(n18217), .ZN(
        n17874) );
  OAI21_X1 U20997 ( .B1(n18146), .B2(n17823), .A(n17874), .ZN(n17814) );
  AOI21_X1 U20998 ( .B1(n17795), .B2(n17907), .A(n18022), .ZN(n17792) );
  OAI21_X1 U20999 ( .B1(n18937), .B2(n17793), .A(n17792), .ZN(n17794) );
  INV_X1 U21000 ( .A(n17794), .ZN(n17820) );
  OAI21_X1 U21001 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17817), .A(
        n17820), .ZN(n17806) );
  AOI22_X1 U21002 ( .A1(n18393), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17806), .ZN(n17798) );
  NOR2_X1 U21003 ( .A1(n17910), .A2(n17795), .ZN(n17808) );
  OAI211_X1 U21004 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17808), .B(n17796), .ZN(n17797) );
  OAI211_X1 U21005 ( .C1(n17911), .C2(n17799), .A(n17798), .B(n17797), .ZN(
        n17800) );
  AOI21_X1 U21006 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17814), .A(
        n17800), .ZN(n17802) );
  NAND3_X1 U21007 ( .A1(n18146), .A2(n17858), .A3(n18151), .ZN(n17801) );
  OAI211_X1 U21008 ( .C1(n17991), .C2(n18155), .A(n17802), .B(n17801), .ZN(
        P3_U2808) );
  NAND2_X1 U21009 ( .A1(n18160), .A2(n18149), .ZN(n18164) );
  NAND2_X1 U21010 ( .A1(n18184), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18158) );
  OR2_X1 U21011 ( .A1(n17875), .A2(n18158), .ZN(n17839) );
  AOI22_X1 U21012 ( .A1(n18393), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17927), 
        .B2(n17803), .ZN(n17804) );
  INV_X1 U21013 ( .A(n17804), .ZN(n17805) );
  AOI221_X1 U21014 ( .B1(n17808), .B2(n17807), .C1(n17806), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17805), .ZN(n17816) );
  INV_X1 U21015 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17810) );
  NOR3_X1 U21016 ( .A1(n17810), .A2(n17978), .A3(n17809), .ZN(n17834) );
  AOI22_X1 U21017 ( .A1(n18160), .A2(n17834), .B1(n17811), .B2(n17812), .ZN(
        n17813) );
  XOR2_X1 U21018 ( .A(n18149), .B(n17813), .Z(n18157) );
  AOI22_X1 U21019 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17814), .B1(
        n17973), .B2(n18157), .ZN(n17815) );
  OAI211_X1 U21020 ( .C1(n18164), .C2(n17839), .A(n17816), .B(n17815), .ZN(
        P3_U2809) );
  NAND2_X1 U21021 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18148), .ZN(
        n18176) );
  AOI21_X1 U21022 ( .B1(n17818), .B2(n18798), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17819) );
  OAI22_X1 U21023 ( .A1(n17820), .A2(n17819), .B1(n9655), .B2(n18993), .ZN(
        n17821) );
  AOI221_X1 U21024 ( .B1(n17927), .B2(n17822), .C1(n17780), .C2(n17822), .A(
        n17821), .ZN(n17827) );
  NOR2_X1 U21025 ( .A1(n18182), .A2(n18158), .ZN(n18167) );
  OAI21_X1 U21026 ( .B1(n17823), .B2(n18167), .A(n17874), .ZN(n17836) );
  OAI221_X1 U21027 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17840), 
        .C1(n18182), .C2(n17834), .A(n17824), .ZN(n17825) );
  XOR2_X1 U21028 ( .A(n18148), .B(n17825), .Z(n18171) );
  AOI22_X1 U21029 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17836), .B1(
        n17973), .B2(n18171), .ZN(n17826) );
  OAI211_X1 U21030 ( .C1(n17839), .C2(n18176), .A(n17827), .B(n17826), .ZN(
        P3_U2810) );
  AOI21_X1 U21031 ( .B1(n17907), .B2(n17829), .A(n18022), .ZN(n17852) );
  OAI21_X1 U21032 ( .B1(n17828), .B2(n18937), .A(n17852), .ZN(n17844) );
  NOR2_X1 U21033 ( .A1(n17910), .A2(n17829), .ZN(n17846) );
  OAI211_X1 U21034 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17846), .B(n17830), .ZN(n17831) );
  NAND2_X1 U21035 ( .A1(n18393), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18179) );
  OAI211_X1 U21036 ( .C1(n17911), .C2(n17832), .A(n17831), .B(n18179), .ZN(
        n17833) );
  AOI21_X1 U21037 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17844), .A(
        n17833), .ZN(n17838) );
  AOI21_X1 U21038 ( .B1(n17840), .B2(n17811), .A(n17834), .ZN(n17835) );
  XOR2_X1 U21039 ( .A(n18182), .B(n17835), .Z(n18178) );
  AOI22_X1 U21040 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17836), .B1(
        n17973), .B2(n18178), .ZN(n17837) );
  OAI211_X1 U21041 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17839), .A(
        n17838), .B(n17837), .ZN(P3_U2811) );
  AOI21_X1 U21042 ( .B1(n17955), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17840), .ZN(n17841) );
  XNOR2_X1 U21043 ( .A(n17811), .B(n17841), .ZN(n18199) );
  OAI22_X1 U21044 ( .A1(n9655), .A2(n18989), .B1(n17911), .B2(n17842), .ZN(
        n17843) );
  AOI221_X1 U21045 ( .B1(n17846), .B2(n17845), .C1(n17844), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17843), .ZN(n17849) );
  OAI21_X1 U21046 ( .B1(n18184), .B2(n17875), .A(n17874), .ZN(n17850) );
  NOR2_X1 U21047 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17847), .ZN(
        n18195) );
  AOI22_X1 U21048 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17850), .B1(
        n17858), .B2(n18195), .ZN(n17848) );
  OAI211_X1 U21049 ( .C1(n17991), .C2(n18199), .A(n17849), .B(n17848), .ZN(
        P3_U2812) );
  INV_X1 U21050 ( .A(n17850), .ZN(n17862) );
  AOI21_X1 U21051 ( .B1(n17851), .B2(n18798), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17853) );
  NAND2_X1 U21052 ( .A1(n18393), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18202) );
  OAI21_X1 U21053 ( .B1(n17853), .B2(n17852), .A(n18202), .ZN(n17854) );
  AOI21_X1 U21054 ( .B1(n17855), .B2(n18071), .A(n17854), .ZN(n17860) );
  OAI21_X1 U21055 ( .B1(n17857), .B2(n17861), .A(n17856), .ZN(n18201) );
  NOR2_X1 U21056 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18212), .ZN(
        n18200) );
  AOI22_X1 U21057 ( .A1(n17973), .A2(n18201), .B1(n17858), .B2(n18200), .ZN(
        n17859) );
  OAI211_X1 U21058 ( .C1(n17862), .C2(n17861), .A(n17860), .B(n17859), .ZN(
        P3_U2813) );
  NAND2_X1 U21059 ( .A1(n17955), .A2(n17904), .ZN(n17965) );
  INV_X1 U21060 ( .A(n17863), .ZN(n18193) );
  OAI22_X1 U21061 ( .A1(n17955), .A2(n17864), .B1(n17965), .B2(n18193), .ZN(
        n17865) );
  XOR2_X1 U21062 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17865), .Z(
        n18214) );
  AOI21_X1 U21063 ( .B1(n17907), .B2(n17867), .A(n18022), .ZN(n17893) );
  OAI21_X1 U21064 ( .B1(n17866), .B2(n18937), .A(n17893), .ZN(n17882) );
  AOI22_X1 U21065 ( .A1(n18393), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17882), .ZN(n17870) );
  NOR2_X1 U21066 ( .A1(n17910), .A2(n17867), .ZN(n17884) );
  OAI211_X1 U21067 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17884), .B(n17868), .ZN(n17869) );
  OAI211_X1 U21068 ( .C1(n17911), .C2(n17871), .A(n17870), .B(n17869), .ZN(
        n17872) );
  AOI21_X1 U21069 ( .B1(n17973), .B2(n18214), .A(n17872), .ZN(n17873) );
  OAI221_X1 U21070 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17875), 
        .C1(n18212), .C2(n17874), .A(n17873), .ZN(P3_U2814) );
  AOI21_X1 U21071 ( .B1(n17877), .B2(n17917), .A(n17876), .ZN(n17878) );
  AOI221_X1 U21072 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18269), 
        .C1(n17978), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17878), .ZN(
        n17879) );
  XOR2_X1 U21073 ( .A(n12657), .B(n17879), .Z(n18223) );
  OAI22_X1 U21074 ( .A1(n9655), .A2(n18983), .B1(n17911), .B2(n17880), .ZN(
        n17881) );
  AOI221_X1 U21075 ( .B1(n17884), .B2(n17883), .C1(n17882), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17881), .ZN(n17889) );
  AOI21_X1 U21076 ( .B1(n17890), .B2(n12657), .A(n17885), .ZN(n18226) );
  NOR2_X1 U21077 ( .A1(n17886), .A2(n17986), .ZN(n17887) );
  OAI21_X1 U21078 ( .B1(n18218), .B2(n18276), .A(n12657), .ZN(n18221) );
  AOI22_X1 U21079 ( .A1(n18069), .A2(n18226), .B1(n17887), .B2(n18221), .ZN(
        n17888) );
  OAI211_X1 U21080 ( .C1(n17991), .C2(n18223), .A(n17889), .B(n17888), .ZN(
        P3_U2815) );
  NOR3_X1 U21081 ( .A1(n18269), .A2(n18263), .A3(n18229), .ZN(n17898) );
  OAI221_X1 U21082 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17898), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17903), .A(n17890), .ZN(
        n18240) );
  NOR2_X1 U21083 ( .A1(n17891), .A2(n18444), .ZN(n17942) );
  AOI21_X1 U21084 ( .B1(n17914), .B2(n17942), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17892) );
  OAI22_X1 U21085 ( .A1(n17893), .A2(n17892), .B1(n9655), .B2(n18982), .ZN(
        n17900) );
  INV_X1 U21086 ( .A(n17898), .ZN(n18236) );
  OAI21_X1 U21087 ( .B1(n17965), .B2(n18236), .A(n17894), .ZN(n17895) );
  XOR2_X1 U21088 ( .A(n17895), .B(n12656), .Z(n18242) );
  NAND2_X1 U21089 ( .A1(n17896), .A2(n17904), .ZN(n17897) );
  OAI221_X1 U21090 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17904), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17898), .A(n17897), .ZN(
        n18241) );
  OAI22_X1 U21091 ( .A1(n18242), .A2(n17991), .B1(n17986), .B2(n18241), .ZN(
        n17899) );
  AOI211_X1 U21092 ( .C1(n17901), .C2(n18071), .A(n17900), .B(n17899), .ZN(
        n17902) );
  OAI21_X1 U21093 ( .B1(n18080), .B2(n18240), .A(n17902), .ZN(P3_U2816) );
  NOR2_X1 U21094 ( .A1(n18269), .A2(n18263), .ZN(n18231) );
  NAND2_X1 U21095 ( .A1(n17903), .A2(n18231), .ZN(n18247) );
  NAND2_X1 U21096 ( .A1(n17904), .A2(n18231), .ZN(n18252) );
  AOI22_X1 U21097 ( .A1(n18069), .A2(n18247), .B1(n17945), .B2(n18252), .ZN(
        n17934) );
  INV_X1 U21098 ( .A(n18937), .ZN(n17905) );
  AOI21_X1 U21099 ( .B1(n17907), .B2(n17906), .A(n17905), .ZN(n17908) );
  INV_X1 U21100 ( .A(n17907), .ZN(n18048) );
  OAI21_X1 U21101 ( .B1(n18048), .B2(n17939), .A(n9676), .ZN(n17997) );
  INV_X1 U21102 ( .A(n17997), .ZN(n17983) );
  OAI21_X1 U21103 ( .B1(n17909), .B2(n17908), .A(n17983), .ZN(n17928) );
  NOR2_X1 U21104 ( .A1(n9655), .A2(n18979), .ZN(n17916) );
  INV_X1 U21105 ( .A(n17910), .ZN(n17924) );
  OAI211_X1 U21106 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17925), .B(n17924), .ZN(n17913) );
  OAI22_X1 U21107 ( .A1(n17914), .A2(n17913), .B1(n17912), .B2(n17911), .ZN(
        n17915) );
  AOI211_X1 U21108 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17928), .A(
        n17916), .B(n17915), .ZN(n17921) );
  AOI22_X1 U21109 ( .A1(n18231), .A2(n17917), .B1(n18269), .B2(n17978), .ZN(
        n17918) );
  AOI21_X1 U21110 ( .B1(n17978), .B2(n17922), .A(n17918), .ZN(n17919) );
  XNOR2_X1 U21111 ( .A(n18229), .B(n17919), .ZN(n18257) );
  INV_X1 U21112 ( .A(n18231), .ZN(n18260) );
  NOR2_X1 U21113 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18260), .ZN(
        n18256) );
  AOI22_X1 U21114 ( .A1(n17973), .A2(n18257), .B1(n18256), .B2(n17944), .ZN(
        n17920) );
  OAI211_X1 U21115 ( .C1(n17934), .C2(n18229), .A(n17921), .B(n17920), .ZN(
        P3_U2817) );
  OAI21_X1 U21116 ( .B1(n18263), .B2(n17965), .A(n17922), .ZN(n17923) );
  XOR2_X1 U21117 ( .A(n17923), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18266) );
  INV_X1 U21118 ( .A(n17944), .ZN(n17976) );
  NOR3_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17976), .A3(
        n18263), .ZN(n17932) );
  NAND2_X1 U21120 ( .A1(n17925), .A2(n17924), .ZN(n17930) );
  AOI22_X1 U21121 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17928), .B1(
        n17927), .B2(n17926), .ZN(n17929) );
  NAND2_X1 U21122 ( .A1(n18393), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18267) );
  OAI211_X1 U21123 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17930), .A(
        n17929), .B(n18267), .ZN(n17931) );
  AOI211_X1 U21124 ( .C1(n17973), .C2(n18266), .A(n17932), .B(n17931), .ZN(
        n17933) );
  OAI21_X1 U21125 ( .B1(n17934), .B2(n18269), .A(n17933), .ZN(P3_U2818) );
  INV_X1 U21126 ( .A(n18281), .ZN(n17937) );
  NOR2_X1 U21127 ( .A1(n17937), .A2(n17965), .ZN(n17958) );
  NOR2_X1 U21128 ( .A1(n17958), .A2(n17935), .ZN(n17936) );
  XOR2_X1 U21129 ( .A(n17936), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18287) );
  NOR2_X1 U21130 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17937), .ZN(
        n18272) );
  NOR2_X1 U21131 ( .A1(n9655), .A2(n18975), .ZN(n18270) );
  INV_X1 U21132 ( .A(n18012), .ZN(n18072) );
  NAND4_X1 U21133 ( .A1(n17939), .A2(n17938), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(n18798), .ZN(n17967) );
  NOR2_X1 U21134 ( .A1(n17950), .A2(n17967), .ZN(n17949) );
  AOI21_X1 U21135 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18072), .A(
        n17949), .ZN(n17941) );
  OAI22_X1 U21136 ( .A1(n17942), .A2(n17941), .B1(n18062), .B2(n17940), .ZN(
        n17943) );
  AOI211_X1 U21137 ( .C1(n18272), .C2(n17944), .A(n18270), .B(n17943), .ZN(
        n17948) );
  NOR2_X1 U21138 ( .A1(n18281), .A2(n17976), .ZN(n17961) );
  AOI22_X1 U21139 ( .A1(n18276), .A2(n17945), .B1(n18069), .B2(n18274), .ZN(
        n17975) );
  INV_X1 U21140 ( .A(n17975), .ZN(n17946) );
  OAI21_X1 U21141 ( .B1(n17961), .B2(n17946), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17947) );
  OAI211_X1 U21142 ( .C1(n18287), .C2(n17991), .A(n17948), .B(n17947), .ZN(
        P3_U2819) );
  AOI211_X1 U21143 ( .C1(n17967), .C2(n17950), .A(n18012), .B(n17949), .ZN(
        n17952) );
  INV_X1 U21144 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18973) );
  NOR2_X1 U21145 ( .A1(n9655), .A2(n18973), .ZN(n17951) );
  AOI211_X1 U21146 ( .C1(n17953), .C2(n18071), .A(n17952), .B(n17951), .ZN(
        n17963) );
  NOR3_X1 U21147 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17955), .A3(
        n17954), .ZN(n17959) );
  OAI221_X1 U21148 ( .B1(n12654), .B2(n17965), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17964), .A(n12653), .ZN(
        n17956) );
  INV_X1 U21149 ( .A(n17956), .ZN(n17957) );
  AOI211_X1 U21150 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17959), .A(
        n17958), .B(n17957), .ZN(n18288) );
  AOI22_X1 U21151 ( .A1(n17973), .A2(n18288), .B1(n17961), .B2(n17960), .ZN(
        n17962) );
  OAI211_X1 U21152 ( .C1(n17975), .C2(n12653), .A(n17963), .B(n17962), .ZN(
        P3_U2820) );
  NAND2_X1 U21153 ( .A1(n17965), .A2(n17964), .ZN(n17966) );
  XOR2_X1 U21154 ( .A(n17966), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18298) );
  NOR2_X1 U21155 ( .A1(n9655), .A2(n18971), .ZN(n18297) );
  INV_X1 U21156 ( .A(n17967), .ZN(n17971) );
  NOR3_X1 U21157 ( .A1(n17994), .A2(n17979), .A3(n18444), .ZN(n17968) );
  AOI21_X1 U21158 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18072), .A(
        n17968), .ZN(n17970) );
  OAI22_X1 U21159 ( .A1(n17971), .A2(n17970), .B1(n18062), .B2(n17969), .ZN(
        n17972) );
  AOI211_X1 U21160 ( .C1(n17973), .C2(n18298), .A(n18297), .B(n17972), .ZN(
        n17974) );
  OAI221_X1 U21161 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17976), .C1(
        n12654), .C2(n17975), .A(n17974), .ZN(P3_U2821) );
  AOI21_X1 U21162 ( .B1(n17978), .B2(n18311), .A(n17977), .ZN(n18313) );
  NAND2_X1 U21163 ( .A1(n18393), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18309) );
  OAI211_X1 U21164 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17980), .A(
        n18798), .B(n17979), .ZN(n17981) );
  OAI211_X1 U21165 ( .C1(n17983), .C2(n17982), .A(n18309), .B(n17981), .ZN(
        n17988) );
  OAI21_X1 U21166 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17985), .A(
        n17984), .ZN(n18318) );
  OAI22_X1 U21167 ( .A1(n18080), .A2(n18318), .B1(n17986), .B2(n18311), .ZN(
        n17987) );
  AOI211_X1 U21168 ( .C1(n17989), .C2(n18071), .A(n17988), .B(n17987), .ZN(
        n17990) );
  OAI21_X1 U21169 ( .B1(n18313), .B2(n17991), .A(n17990), .ZN(P3_U2822) );
  OAI21_X1 U21170 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17993), .A(
        n17992), .ZN(n18321) );
  NOR2_X1 U21171 ( .A1(n17994), .A2(n18444), .ZN(n17996) );
  NOR2_X1 U21172 ( .A1(n9655), .A2(n18967), .ZN(n18325) );
  AOI221_X1 U21173 ( .B1(n17997), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17996), .C2(n17995), .A(n18325), .ZN(n18004) );
  AOI21_X1 U21174 ( .B1(n18000), .B2(n17999), .A(n17998), .ZN(n18001) );
  XOR2_X1 U21175 ( .A(n18001), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18319) );
  AOI22_X1 U21176 ( .A1(n18069), .A2(n18319), .B1(n18002), .B2(n18071), .ZN(
        n18003) );
  OAI211_X1 U21177 ( .C1(n18079), .C2(n18321), .A(n18004), .B(n18003), .ZN(
        P3_U2823) );
  OAI21_X1 U21178 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18006), .A(
        n18005), .ZN(n18330) );
  NAND2_X1 U21179 ( .A1(n18013), .A2(n18798), .ZN(n18010) );
  OAI21_X1 U21180 ( .B1(n18009), .B2(n9666), .A(n18007), .ZN(n18329) );
  OAI22_X1 U21181 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18010), .B1(
        n18079), .B2(n18329), .ZN(n18011) );
  AOI21_X1 U21182 ( .B1(n18393), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18011), .ZN(
        n18016) );
  AOI21_X1 U21183 ( .B1(n18798), .B2(n18013), .A(n18012), .ZN(n18028) );
  AOI22_X1 U21184 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18028), .B1(
        n18014), .B2(n18071), .ZN(n18015) );
  OAI211_X1 U21185 ( .C1(n18080), .C2(n18330), .A(n18016), .B(n18015), .ZN(
        P3_U2824) );
  OAI21_X1 U21186 ( .B1(n18019), .B2(n18018), .A(n18017), .ZN(n18342) );
  OAI21_X1 U21187 ( .B1(n18022), .B2(n18021), .A(n18020), .ZN(n18027) );
  OAI21_X1 U21188 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18024), .A(
        n9667), .ZN(n18338) );
  OAI22_X1 U21189 ( .A1(n18062), .A2(n18025), .B1(n18079), .B2(n18338), .ZN(
        n18026) );
  AOI21_X1 U21190 ( .B1(n18028), .B2(n18027), .A(n18026), .ZN(n18029) );
  NAND2_X1 U21191 ( .A1(n18393), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18337) );
  OAI211_X1 U21192 ( .C1(n18080), .C2(n18342), .A(n18029), .B(n18337), .ZN(
        P3_U2825) );
  OAI21_X1 U21193 ( .B1(n18032), .B2(n18031), .A(n18030), .ZN(n18346) );
  OAI21_X1 U21194 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18034), .A(
        n18033), .ZN(n18352) );
  OAI22_X1 U21195 ( .A1(n18080), .A2(n18352), .B1(n18444), .B2(n18035), .ZN(
        n18036) );
  AOI21_X1 U21196 ( .B1(n18393), .B2(P3_REIP_REG_4__SCAN_IN), .A(n18036), .ZN(
        n18039) );
  OAI21_X1 U21197 ( .B1(n18047), .B2(n18048), .A(n9676), .ZN(n18052) );
  AOI22_X1 U21198 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18052), .B1(
        n18037), .B2(n18071), .ZN(n18038) );
  OAI211_X1 U21199 ( .C1(n18079), .C2(n18346), .A(n18039), .B(n18038), .ZN(
        P3_U2826) );
  OAI21_X1 U21200 ( .B1(n18042), .B2(n18041), .A(n9668), .ZN(n18043) );
  XOR2_X1 U21201 ( .A(n18043), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18356) );
  INV_X1 U21202 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18959) );
  OAI22_X1 U21203 ( .A1(n18079), .A2(n18356), .B1(n9655), .B2(n18959), .ZN(
        n18051) );
  OAI21_X1 U21204 ( .B1(n18046), .B2(n18045), .A(n18044), .ZN(n18361) );
  OR2_X1 U21205 ( .A1(n18048), .A2(n18047), .ZN(n18049) );
  NAND2_X1 U21206 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n9676), .ZN(
        n18064) );
  OAI22_X1 U21207 ( .A1(n18080), .A2(n18361), .B1(n18049), .B2(n18064), .ZN(
        n18050) );
  AOI211_X1 U21208 ( .C1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n18052), .A(
        n18051), .B(n18050), .ZN(n18053) );
  OAI21_X1 U21209 ( .B1(n18062), .B2(n18054), .A(n18053), .ZN(P3_U2827) );
  OAI21_X1 U21210 ( .B1(n18057), .B2(n18056), .A(n18055), .ZN(n18372) );
  OAI21_X1 U21211 ( .B1(n18060), .B2(n18059), .A(n18058), .ZN(n18373) );
  OAI22_X1 U21212 ( .A1(n18062), .A2(n18061), .B1(n18080), .B2(n18373), .ZN(
        n18063) );
  AOI221_X1 U21213 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18064), .C1(
        n18798), .C2(n18064), .A(n18063), .ZN(n18065) );
  NAND2_X1 U21214 ( .A1(n18393), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18378) );
  OAI211_X1 U21215 ( .C1(n18079), .C2(n18372), .A(n18065), .B(n18378), .ZN(
        P3_U2828) );
  OAI21_X1 U21216 ( .B1(n18067), .B2(n18075), .A(n18066), .ZN(n18392) );
  NAND2_X1 U21217 ( .A1(n18385), .A2(n12815), .ZN(n18068) );
  XNOR2_X1 U21218 ( .A(n18068), .B(n18067), .ZN(n18388) );
  AOI22_X1 U21219 ( .A1(n18069), .A2(n18388), .B1(n18393), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U21220 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18072), .B1(
        n18071), .B2(n18070), .ZN(n18073) );
  OAI211_X1 U21221 ( .C1(n18079), .C2(n18392), .A(n18074), .B(n18073), .ZN(
        P3_U2829) );
  AOI21_X1 U21222 ( .B1(n12815), .B2(n18385), .A(n18075), .ZN(n18397) );
  INV_X1 U21223 ( .A(n18397), .ZN(n18395) );
  NAND3_X1 U21224 ( .A1(n19049), .A2(n18937), .A3(n9676), .ZN(n18077) );
  AOI22_X1 U21225 ( .A1(n18393), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18077), .ZN(n18078) );
  OAI221_X1 U21226 ( .B1(n18397), .B2(n18080), .C1(n18395), .C2(n18079), .A(
        n18078), .ZN(P3_U2830) );
  INV_X1 U21227 ( .A(n18081), .ZN(n18082) );
  AOI221_X1 U21228 ( .B1(n18152), .B2(n9991), .C1(n18082), .C2(n9991), .A(
        n18399), .ZN(n18092) );
  NAND2_X1 U21229 ( .A1(n18864), .A2(n18385), .ZN(n18366) );
  NAND2_X1 U21230 ( .A1(n18143), .A2(n18366), .ZN(n18185) );
  NOR2_X1 U21231 ( .A1(n18135), .A2(n18185), .ZN(n18122) );
  NOR2_X1 U21232 ( .A1(n18897), .A2(n18864), .ZN(n18365) );
  AOI21_X1 U21233 ( .B1(n18106), .B2(n18122), .A(n18365), .ZN(n18102) );
  AOI22_X1 U21234 ( .A1(n18897), .A2(n18107), .B1(n18864), .B2(n18083), .ZN(
        n18084) );
  INV_X1 U21235 ( .A(n18084), .ZN(n18085) );
  AOI211_X1 U21236 ( .C1(n18087), .C2(n18852), .A(n18086), .B(n18085), .ZN(
        n18088) );
  INV_X1 U21237 ( .A(n18088), .ZN(n18089) );
  AOI211_X1 U21238 ( .C1(n18277), .C2(n18090), .A(n18102), .B(n18089), .ZN(
        n18096) );
  OAI211_X1 U21239 ( .C1(n18872), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18096), .ZN(n18091) );
  AOI22_X1 U21240 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18359), .B1(
        n18092), .B2(n18091), .ZN(n18094) );
  NAND2_X1 U21241 ( .A1(n18393), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18093) );
  OAI211_X1 U21242 ( .C1(n18095), .C2(n18312), .A(n18094), .B(n18093), .ZN(
        P3_U2835) );
  AOI21_X1 U21243 ( .B1(n18382), .B2(n18096), .A(n9990), .ZN(n18099) );
  NOR3_X1 U21244 ( .A1(n18135), .A2(n18156), .A3(n18097), .ZN(n18098) );
  AOI221_X1 U21245 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n18393), .C1(n18099), 
        .C2(n9655), .A(n18098), .ZN(n18100) );
  OAI21_X1 U21246 ( .B1(n18101), .B2(n18312), .A(n18100), .ZN(P3_U2836) );
  OAI21_X1 U21247 ( .B1(n18105), .B2(n18363), .A(n18183), .ZN(n18124) );
  AOI211_X1 U21248 ( .C1(n18881), .C2(n18103), .A(n18102), .B(n18124), .ZN(
        n18109) );
  NAND3_X1 U21249 ( .A1(n18106), .A2(n18105), .A3(n18104), .ZN(n18108) );
  AOI221_X1 U21250 ( .B1(n18109), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n18108), .C2(n18107), .A(n18399), .ZN(n18110) );
  AOI21_X1 U21251 ( .B1(n18359), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18110), .ZN(n18112) );
  OAI211_X1 U21252 ( .C1(n18113), .C2(n18312), .A(n18112), .B(n18111), .ZN(
        n18114) );
  AOI21_X1 U21253 ( .B1(n18116), .B2(n18115), .A(n18114), .ZN(n18117) );
  OAI21_X1 U21254 ( .B1(n18374), .B2(n18118), .A(n18117), .ZN(P3_U2837) );
  NOR2_X1 U21255 ( .A1(n18135), .A2(n18156), .ZN(n18131) );
  AOI22_X1 U21256 ( .A1(n18852), .A2(n18120), .B1(n18277), .B2(n18119), .ZN(
        n18121) );
  OAI211_X1 U21257 ( .C1(n18365), .C2(n18122), .A(n18121), .B(n18383), .ZN(
        n18123) );
  INV_X1 U21258 ( .A(n18123), .ZN(n18128) );
  INV_X1 U21259 ( .A(n18124), .ZN(n18125) );
  NAND3_X1 U21260 ( .A1(n18125), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n18128), .ZN(n18126) );
  NAND2_X1 U21261 ( .A1(n9655), .A2(n18126), .ZN(n18140) );
  AOI211_X1 U21262 ( .C1(n18345), .C2(n18128), .A(n18127), .B(n18140), .ZN(
        n18129) );
  AOI211_X1 U21263 ( .C1(n18132), .C2(n18131), .A(n18130), .B(n18129), .ZN(
        n18133) );
  OAI21_X1 U21264 ( .B1(n18134), .B2(n18312), .A(n18133), .ZN(P3_U2838) );
  OR3_X1 U21265 ( .A1(n18135), .A2(n18359), .A3(n18152), .ZN(n18138) );
  AOI22_X1 U21266 ( .A1(n18393), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18299), 
        .B2(n18136), .ZN(n18137) );
  OAI221_X1 U21267 ( .B1(n18140), .B2(n18139), .C1(n18140), .C2(n18138), .A(
        n18137), .ZN(P3_U2839) );
  OAI21_X1 U21268 ( .B1(n18150), .B2(n18207), .A(n18864), .ZN(n18141) );
  NOR2_X1 U21269 ( .A1(n18852), .A2(n18277), .ZN(n18280) );
  AOI22_X1 U21270 ( .A1(n18852), .A2(n18142), .B1(n18277), .B2(n18217), .ZN(
        n18187) );
  OAI221_X1 U21271 ( .B1(n18872), .B2(n18143), .C1(n18872), .C2(n18167), .A(
        n18187), .ZN(n18144) );
  AOI221_X1 U21272 ( .B1(n18145), .B2(n18881), .C1(n18158), .C2(n18881), .A(
        n18144), .ZN(n18165) );
  OAI21_X1 U21273 ( .B1(n18146), .B2(n18280), .A(n18165), .ZN(n18147) );
  AOI21_X1 U21274 ( .B1(n18897), .B2(n18148), .A(n18147), .ZN(n18159) );
  NAND2_X1 U21275 ( .A1(n18393), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18153) );
  OAI211_X1 U21276 ( .C1(n18155), .C2(n18312), .A(n18154), .B(n18153), .ZN(
        P3_U2840) );
  NOR2_X1 U21277 ( .A1(n18156), .A2(n18158), .ZN(n18177) );
  INV_X1 U21278 ( .A(n18177), .ZN(n18175) );
  AOI22_X1 U21279 ( .A1(n18393), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18299), 
        .B2(n18157), .ZN(n18163) );
  NAND2_X1 U21280 ( .A1(n18363), .A2(n18894), .ZN(n18381) );
  INV_X1 U21281 ( .A(n18381), .ZN(n18170) );
  AOI221_X1 U21282 ( .B1(n18207), .B2(n18864), .C1(n18158), .C2(n18864), .A(
        n18399), .ZN(n18166) );
  OAI211_X1 U21283 ( .C1(n18160), .C2(n18170), .A(n18166), .B(n18159), .ZN(
        n18161) );
  NAND3_X1 U21284 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n9655), .A3(
        n18161), .ZN(n18162) );
  OAI211_X1 U21285 ( .C1(n18164), .C2(n18175), .A(n18163), .B(n18162), .ZN(
        P3_U2841) );
  NAND2_X1 U21286 ( .A1(n18182), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18169) );
  OAI211_X1 U21287 ( .C1(n18167), .C2(n18280), .A(n18166), .B(n18165), .ZN(
        n18168) );
  NAND2_X1 U21288 ( .A1(n9655), .A2(n18168), .ZN(n18181) );
  OAI21_X1 U21289 ( .B1(n18170), .B2(n18169), .A(n18181), .ZN(n18172) );
  AOI22_X1 U21290 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18172), .B1(
        n18299), .B2(n18171), .ZN(n18174) );
  NAND2_X1 U21291 ( .A1(n18393), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18173) );
  OAI211_X1 U21292 ( .C1(n18176), .C2(n18175), .A(n18174), .B(n18173), .ZN(
        P3_U2842) );
  AOI22_X1 U21293 ( .A1(n18299), .A2(n18178), .B1(n18177), .B2(n18182), .ZN(
        n18180) );
  OAI211_X1 U21294 ( .C1(n18182), .C2(n18181), .A(n18180), .B(n18179), .ZN(
        P3_U2843) );
  AOI22_X1 U21295 ( .A1(n18184), .A2(n18183), .B1(n18280), .B2(n18363), .ZN(
        n18189) );
  INV_X1 U21296 ( .A(n18185), .ZN(n18186) );
  AOI21_X1 U21297 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18186), .A(
        n18365), .ZN(n18188) );
  NAND2_X1 U21298 ( .A1(n18382), .A2(n18187), .ZN(n18211) );
  NOR3_X1 U21299 ( .A1(n18189), .A2(n18188), .A3(n18211), .ZN(n18205) );
  AOI221_X1 U21300 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18205), 
        .C1(n18365), .C2(n18205), .A(n18393), .ZN(n18196) );
  NOR2_X1 U21301 ( .A1(n18380), .A2(n19036), .ZN(n18303) );
  AOI22_X1 U21302 ( .A1(n18881), .A2(n18362), .B1(n18303), .B2(n18190), .ZN(
        n18355) );
  NOR2_X1 U21303 ( .A1(n18355), .A2(n18191), .ZN(n18320) );
  NAND2_X1 U21304 ( .A1(n18192), .A2(n18320), .ZN(n18237) );
  AOI211_X1 U21305 ( .C1(n18194), .C2(n18237), .A(n18193), .B(n18399), .ZN(
        n18213) );
  AOI22_X1 U21306 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18196), .B1(
        n18195), .B2(n18213), .ZN(n18198) );
  NAND2_X1 U21307 ( .A1(n18393), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18197) );
  OAI211_X1 U21308 ( .C1(n18199), .C2(n18312), .A(n18198), .B(n18197), .ZN(
        P3_U2844) );
  NAND2_X1 U21309 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n9655), .ZN(
        n18204) );
  AOI22_X1 U21310 ( .A1(n18299), .A2(n18201), .B1(n18213), .B2(n18200), .ZN(
        n18203) );
  OAI211_X1 U21311 ( .C1(n18205), .C2(n18204), .A(n18203), .B(n18202), .ZN(
        P3_U2845) );
  INV_X1 U21312 ( .A(n18248), .ZN(n18290) );
  NOR2_X1 U21313 ( .A1(n18872), .A2(n18206), .ZN(n18296) );
  NOR2_X1 U21314 ( .A1(n18232), .A2(n18363), .ZN(n18273) );
  NOR3_X1 U21315 ( .A1(n18296), .A2(n18273), .A3(n18218), .ZN(n18209) );
  OAI21_X1 U21316 ( .B1(n12657), .B2(n18864), .A(n18207), .ZN(n18208) );
  OAI21_X1 U21317 ( .B1(n18290), .B2(n18209), .A(n18208), .ZN(n18220) );
  OAI221_X1 U21318 ( .B1(n18211), .B2(n18210), .C1(n18211), .C2(n18220), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U21319 ( .A1(n18299), .A2(n18214), .B1(n18213), .B2(n18212), .ZN(
        n18215) );
  OAI221_X1 U21320 ( .B1(n18393), .B2(n18216), .C1(n9655), .C2(n18985), .A(
        n18215), .ZN(P3_U2846) );
  AND2_X1 U21321 ( .A1(n18217), .A2(n18277), .ZN(n18222) );
  OAI21_X1 U21322 ( .B1(n18218), .B2(n18237), .A(n12657), .ZN(n18219) );
  AOI22_X1 U21323 ( .A1(n18222), .A2(n18221), .B1(n18220), .B2(n18219), .ZN(
        n18224) );
  OAI22_X1 U21324 ( .A1(n18224), .A2(n18399), .B1(n18312), .B2(n18223), .ZN(
        n18225) );
  AOI21_X1 U21325 ( .B1(n18396), .B2(n18226), .A(n18225), .ZN(n18228) );
  NAND2_X1 U21326 ( .A1(n18393), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18227) );
  OAI211_X1 U21327 ( .C1(n18383), .C2(n12657), .A(n18228), .B(n18227), .ZN(
        P3_U2847) );
  AOI22_X1 U21328 ( .A1(n18897), .A2(n18236), .B1(n18229), .B2(n18381), .ZN(
        n18235) );
  AOI21_X1 U21329 ( .B1(n18230), .B2(n18231), .A(n18894), .ZN(n18254) );
  AOI21_X1 U21330 ( .B1(n18232), .B2(n18231), .A(n18363), .ZN(n18233) );
  NOR4_X1 U21331 ( .A1(n18254), .A2(n18296), .A3(n18233), .A4(n12656), .ZN(
        n18234) );
  AOI21_X1 U21332 ( .B1(n18235), .B2(n18234), .A(n18399), .ZN(n18239) );
  NOR2_X1 U21333 ( .A1(n18237), .A2(n18236), .ZN(n18238) );
  AOI222_X1 U21334 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18239), 
        .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18359), .C1(n18239), 
        .C2(n18238), .ZN(n18246) );
  INV_X1 U21335 ( .A(n18240), .ZN(n18244) );
  OAI22_X1 U21336 ( .A1(n18242), .A2(n18312), .B1(n18310), .B2(n18241), .ZN(
        n18243) );
  AOI21_X1 U21337 ( .B1(n18396), .B2(n18244), .A(n18243), .ZN(n18245) );
  OAI211_X1 U21338 ( .C1(n9655), .C2(n18982), .A(n18246), .B(n18245), .ZN(
        P3_U2848) );
  INV_X1 U21339 ( .A(n18247), .ZN(n18250) );
  OAI21_X1 U21340 ( .B1(n18296), .B2(n18263), .A(n18248), .ZN(n18283) );
  OAI21_X1 U21341 ( .B1(n18250), .B2(n18249), .A(n18283), .ZN(n18251) );
  AOI211_X1 U21342 ( .C1(n18277), .C2(n18252), .A(n18273), .B(n18251), .ZN(
        n18261) );
  OAI211_X1 U21343 ( .C1(n18290), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18261), .B(n18383), .ZN(n18253) );
  OAI21_X1 U21344 ( .B1(n18254), .B2(n18253), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18259) );
  NAND2_X1 U21345 ( .A1(n18382), .A2(n18320), .ZN(n18334) );
  OAI222_X1 U21346 ( .A1(n18310), .A2(n18276), .B1(n18374), .B2(n18274), .C1(
        n18255), .C2(n18334), .ZN(n18271) );
  AOI22_X1 U21347 ( .A1(n18299), .A2(n18257), .B1(n18256), .B2(n18271), .ZN(
        n18258) );
  OAI221_X1 U21348 ( .B1(n18393), .B2(n18259), .C1(n9655), .C2(n18979), .A(
        n18258), .ZN(P3_U2849) );
  NOR2_X1 U21349 ( .A1(n18275), .A2(n18260), .ZN(n18262) );
  OAI211_X1 U21350 ( .C1(n18262), .C2(n18894), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18261), .ZN(n18265) );
  INV_X1 U21351 ( .A(n18271), .ZN(n18302) );
  OAI22_X1 U21352 ( .A1(n18302), .A2(n18263), .B1(n18269), .B2(n18399), .ZN(
        n18264) );
  AOI22_X1 U21353 ( .A1(n18299), .A2(n18266), .B1(n18265), .B2(n18264), .ZN(
        n18268) );
  OAI211_X1 U21354 ( .C1(n18383), .C2(n18269), .A(n18268), .B(n18267), .ZN(
        P3_U2850) );
  AOI21_X1 U21355 ( .B1(n18272), .B2(n18271), .A(n18270), .ZN(n18286) );
  AOI211_X1 U21356 ( .C1(n18274), .C2(n18852), .A(n18273), .B(n18399), .ZN(
        n18279) );
  AOI22_X1 U21357 ( .A1(n18277), .A2(n18276), .B1(n18864), .B2(n18275), .ZN(
        n18278) );
  NAND2_X1 U21358 ( .A1(n18279), .A2(n18278), .ZN(n18295) );
  OAI22_X1 U21359 ( .A1(n18894), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n18281), .B2(n18280), .ZN(n18282) );
  NOR2_X1 U21360 ( .A1(n18295), .A2(n18282), .ZN(n18289) );
  OAI211_X1 U21361 ( .C1(n18894), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18289), .B(n18283), .ZN(n18284) );
  NAND3_X1 U21362 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n9655), .A3(
        n18284), .ZN(n18285) );
  OAI211_X1 U21363 ( .C1(n18287), .C2(n18312), .A(n18286), .B(n18285), .ZN(
        P3_U2851) );
  NAND2_X1 U21364 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n12653), .ZN(
        n18294) );
  AOI22_X1 U21365 ( .A1(n18393), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18299), 
        .B2(n18288), .ZN(n18293) );
  OAI21_X1 U21366 ( .B1(n18290), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18289), .ZN(n18291) );
  OAI211_X1 U21367 ( .C1(n18296), .C2(n18291), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n9655), .ZN(n18292) );
  OAI211_X1 U21368 ( .C1(n18302), .C2(n18294), .A(n18293), .B(n18292), .ZN(
        P3_U2852) );
  OAI21_X1 U21369 ( .B1(n18296), .B2(n18295), .A(n9655), .ZN(n18301) );
  AOI21_X1 U21370 ( .B1(n18299), .B2(n18298), .A(n18297), .ZN(n18300) );
  OAI221_X1 U21371 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18302), .C1(
        n12654), .C2(n18301), .A(n18300), .ZN(P3_U2853) );
  NOR3_X1 U21372 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18307), .A3(
        n18334), .ZN(n18316) );
  AOI21_X1 U21373 ( .B1(n18303), .B2(n18366), .A(n18365), .ZN(n18344) );
  AOI21_X1 U21374 ( .B1(n18881), .B2(n18304), .A(n18344), .ZN(n18305) );
  AOI221_X1 U21375 ( .B1(n18306), .B2(n18305), .C1(n18365), .C2(n18305), .A(
        n18399), .ZN(n18328) );
  AOI21_X1 U21376 ( .B1(n18308), .B2(n18307), .A(n18328), .ZN(n18323) );
  OAI221_X1 U21377 ( .B1(n9664), .B2(n18323), .C1(n9664), .C2(n18383), .A(
        n18309), .ZN(n18315) );
  OAI22_X1 U21378 ( .A1(n18313), .A2(n18312), .B1(n18311), .B2(n18310), .ZN(
        n18314) );
  NOR3_X1 U21379 ( .A1(n18316), .A2(n18315), .A3(n18314), .ZN(n18317) );
  OAI21_X1 U21380 ( .B1(n18374), .B2(n18318), .A(n18317), .ZN(P3_U2854) );
  INV_X1 U21381 ( .A(n18319), .ZN(n18327) );
  AOI21_X1 U21382 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18320), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18322) );
  OAI22_X1 U21383 ( .A1(n18323), .A2(n18322), .B1(n18391), .B2(n18321), .ZN(
        n18324) );
  AOI211_X1 U21384 ( .C1(n18359), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18325), .B(n18324), .ZN(n18326) );
  OAI21_X1 U21385 ( .B1(n18374), .B2(n18327), .A(n18326), .ZN(P3_U2855) );
  OR2_X1 U21386 ( .A1(n18359), .A2(n18328), .ZN(n18340) );
  NOR2_X1 U21387 ( .A1(n9655), .A2(n18965), .ZN(n18332) );
  OAI22_X1 U21388 ( .A1(n18374), .A2(n18330), .B1(n18391), .B2(n18329), .ZN(
        n18331) );
  AOI211_X1 U21389 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18340), .A(
        n18332), .B(n18331), .ZN(n18333) );
  OAI21_X1 U21390 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18334), .A(
        n18333), .ZN(P3_U2856) );
  NOR3_X1 U21391 ( .A1(n18355), .A2(n18399), .A3(n18354), .ZN(n18350) );
  INV_X1 U21392 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18335) );
  NAND3_X1 U21393 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18350), .A3(
        n18335), .ZN(n18336) );
  OAI211_X1 U21394 ( .C1(n18338), .C2(n18391), .A(n18337), .B(n18336), .ZN(
        n18339) );
  AOI21_X1 U21395 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18340), .A(
        n18339), .ZN(n18341) );
  OAI21_X1 U21396 ( .B1(n18374), .B2(n18342), .A(n18341), .ZN(P3_U2857) );
  INV_X1 U21397 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18349) );
  OAI21_X1 U21398 ( .B1(n18363), .B2(n18362), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18343) );
  OAI21_X1 U21399 ( .B1(n18344), .B2(n18343), .A(n18382), .ZN(n18353) );
  OAI21_X1 U21400 ( .B1(n18345), .B2(n18353), .A(n18383), .ZN(n18348) );
  OAI22_X1 U21401 ( .A1(n9655), .A2(n18961), .B1(n18391), .B2(n18346), .ZN(
        n18347) );
  AOI221_X1 U21402 ( .B1(n18350), .B2(n18349), .C1(n18348), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18347), .ZN(n18351) );
  OAI21_X1 U21403 ( .B1(n18374), .B2(n18352), .A(n18351), .ZN(P3_U2858) );
  AOI21_X1 U21404 ( .B1(n18355), .B2(n18354), .A(n18353), .ZN(n18358) );
  OAI22_X1 U21405 ( .A1(n9655), .A2(n18959), .B1(n18391), .B2(n18356), .ZN(
        n18357) );
  AOI211_X1 U21406 ( .C1(n18359), .C2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n18358), .B(n18357), .ZN(n18360) );
  OAI21_X1 U21407 ( .B1(n18374), .B2(n18361), .A(n18360), .ZN(P3_U2859) );
  NOR2_X1 U21408 ( .A1(n18363), .A2(n18362), .ZN(n18377) );
  NOR2_X1 U21409 ( .A1(n19036), .A2(n18364), .ZN(n18371) );
  NOR2_X1 U21410 ( .A1(n18385), .A2(n19036), .ZN(n18368) );
  AOI21_X1 U21411 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18366), .A(
        n18365), .ZN(n18367) );
  AOI21_X1 U21412 ( .B1(n18368), .B2(n18881), .A(n18367), .ZN(n18369) );
  INV_X1 U21413 ( .A(n18369), .ZN(n18370) );
  MUX2_X1 U21414 ( .A(n18371), .B(n18370), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18376) );
  OAI22_X1 U21415 ( .A1(n18374), .A2(n18373), .B1(n18391), .B2(n18372), .ZN(
        n18375) );
  AOI221_X1 U21416 ( .B1(n18377), .B2(n18382), .C1(n18376), .C2(n18382), .A(
        n18375), .ZN(n18379) );
  OAI211_X1 U21417 ( .C1(n18383), .C2(n18380), .A(n18379), .B(n18378), .ZN(
        P3_U2860) );
  NAND3_X1 U21418 ( .A1(n18382), .A2(n18385), .A3(n18381), .ZN(n18401) );
  AOI21_X1 U21419 ( .B1(n18383), .B2(n18401), .A(n19036), .ZN(n18387) );
  AOI211_X1 U21420 ( .C1(n18872), .C2(n18385), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18384), .ZN(n18386) );
  AOI211_X1 U21421 ( .C1(n18396), .C2(n18388), .A(n18387), .B(n18386), .ZN(
        n18390) );
  NAND2_X1 U21422 ( .A1(n18393), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18389) );
  OAI211_X1 U21423 ( .C1(n18392), .C2(n18391), .A(n18390), .B(n18389), .ZN(
        P3_U2861) );
  AND2_X1 U21424 ( .A1(n18393), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18394) );
  AOI221_X1 U21425 ( .B1(n18398), .B2(n18397), .C1(n18396), .C2(n18395), .A(
        n18394), .ZN(n18402) );
  OAI211_X1 U21426 ( .C1(n18897), .C2(n18399), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n9655), .ZN(n18400) );
  NAND3_X1 U21427 ( .A1(n18402), .A2(n18401), .A3(n18400), .ZN(P3_U2862) );
  INV_X1 U21428 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18411) );
  AOI211_X1 U21429 ( .C1(n18404), .C2(n18403), .A(n19086), .B(n19049), .ZN(
        n18919) );
  OAI21_X1 U21430 ( .B1(n18919), .B2(n18452), .A(n18409), .ZN(n18405) );
  OAI221_X1 U21431 ( .B1(n18411), .B2(n19068), .C1(n18411), .C2(n18409), .A(
        n18405), .ZN(P3_U2863) );
  INV_X1 U21432 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18907) );
  NOR2_X1 U21433 ( .A1(n18906), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18585) );
  INV_X1 U21434 ( .A(n18585), .ZN(n18539) );
  NOR2_X1 U21435 ( .A1(n18907), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18680) );
  NAND2_X1 U21436 ( .A1(n18758), .A2(n18680), .ZN(n18702) );
  AND2_X1 U21437 ( .A1(n18539), .A2(n18702), .ZN(n18407) );
  OAI22_X1 U21438 ( .A1(n18408), .A2(n18907), .B1(n18407), .B2(n18406), .ZN(
        P3_U2866) );
  NOR2_X1 U21439 ( .A1(n18908), .A2(n18409), .ZN(P3_U2867) );
  NAND2_X1 U21440 ( .A1(n18798), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18763) );
  NAND2_X1 U21441 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18412) );
  INV_X1 U21442 ( .A(n18412), .ZN(n18410) );
  NOR2_X1 U21443 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18679), .ZN(
        n18653) );
  NAND2_X1 U21444 ( .A1(n18410), .A2(n18653), .ZN(n18774) );
  INV_X1 U21445 ( .A(n18453), .ZN(n18705) );
  AND2_X1 U21446 ( .A1(n18705), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18793) );
  INV_X1 U21447 ( .A(n18792), .ZN(n18927) );
  NOR2_X1 U21448 ( .A1(n18679), .A2(n18411), .ZN(n18898) );
  NAND2_X1 U21449 ( .A1(n18898), .A2(n18410), .ZN(n18816) );
  NOR2_X1 U21450 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18899) );
  NOR2_X1 U21451 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18492) );
  NAND2_X1 U21452 ( .A1(n18899), .A2(n18492), .ZN(n18507) );
  NAND2_X1 U21453 ( .A1(n18816), .A2(n18507), .ZN(n18413) );
  INV_X1 U21454 ( .A(n18413), .ZN(n18472) );
  NOR2_X1 U21455 ( .A1(n18927), .A2(n18472), .ZN(n18446) );
  NOR2_X1 U21456 ( .A1(n18412), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18797) );
  NAND2_X1 U21457 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18797), .ZN(
        n18736) );
  INV_X1 U21458 ( .A(n18736), .ZN(n18844) );
  NOR2_X2 U21459 ( .A1(n15491), .A2(n18444), .ZN(n18799) );
  AOI22_X1 U21460 ( .A1(n18793), .A2(n18446), .B1(n18844), .B2(n18799), .ZN(
        n18418) );
  NOR2_X1 U21461 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18411), .ZN(
        n18628) );
  NOR2_X1 U21462 ( .A1(n18653), .A2(n18628), .ZN(n18703) );
  NOR2_X1 U21463 ( .A1(n18703), .A2(n18412), .ZN(n18759) );
  AOI21_X1 U21464 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18453), .ZN(n18756) );
  AOI22_X1 U21465 ( .A1(n18798), .A2(n18759), .B1(n18756), .B2(n18413), .ZN(
        n18449) );
  INV_X1 U21466 ( .A(n18507), .ZN(n18511) );
  NAND2_X1 U21467 ( .A1(n18415), .A2(n18414), .ZN(n18447) );
  NOR2_X1 U21468 ( .A1(n18416), .A2(n18447), .ZN(n18760) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n18760), .ZN(n18417) );
  OAI211_X1 U21470 ( .C1(n18763), .C2(n18774), .A(n18418), .B(n18417), .ZN(
        P3_U2868) );
  NAND2_X1 U21471 ( .A1(n18798), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18767) );
  AND2_X1 U21472 ( .A1(n18705), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18803) );
  NAND2_X1 U21473 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18798), .ZN(n18808) );
  INV_X1 U21474 ( .A(n18808), .ZN(n18764) );
  AOI22_X1 U21475 ( .A1(n18446), .A2(n18803), .B1(n18844), .B2(n18764), .ZN(
        n18420) );
  NOR2_X2 U21476 ( .A1(n19074), .A2(n18447), .ZN(n18805) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n18805), .ZN(n18419) );
  OAI211_X1 U21478 ( .C1(n18774), .C2(n18767), .A(n18420), .B(n18419), .ZN(
        P3_U2869) );
  NOR2_X1 U21479 ( .A1(n18421), .A2(n18444), .ZN(n18811) );
  INV_X1 U21480 ( .A(n18811), .ZN(n18742) );
  INV_X1 U21481 ( .A(n18774), .ZN(n18787) );
  AND2_X1 U21482 ( .A1(n18798), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18812) );
  NOR2_X2 U21483 ( .A1(n18453), .A2(n18422), .ZN(n18809) );
  AOI22_X1 U21484 ( .A1(n18787), .A2(n18812), .B1(n18446), .B2(n18809), .ZN(
        n18425) );
  NOR2_X1 U21485 ( .A1(n18423), .A2(n18447), .ZN(n18739) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n18739), .ZN(n18424) );
  OAI211_X1 U21487 ( .C1(n18736), .C2(n18742), .A(n18425), .B(n18424), .ZN(
        P3_U2870) );
  NOR2_X1 U21488 ( .A1(n18444), .A2(n15523), .ZN(n18818) );
  INV_X1 U21489 ( .A(n18818), .ZN(n18714) );
  NOR2_X2 U21490 ( .A1(n18453), .A2(n18426), .ZN(n18817) );
  NAND2_X1 U21491 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18798), .ZN(n18822) );
  INV_X1 U21492 ( .A(n18822), .ZN(n18770) );
  AOI22_X1 U21493 ( .A1(n18446), .A2(n18817), .B1(n18844), .B2(n18770), .ZN(
        n18429) );
  NOR2_X2 U21494 ( .A1(n18427), .A2(n18447), .ZN(n18819) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n18819), .ZN(n18428) );
  OAI211_X1 U21496 ( .C1(n18774), .C2(n18714), .A(n18429), .B(n18428), .ZN(
        P3_U2871) );
  INV_X1 U21497 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18430) );
  NOR2_X1 U21498 ( .A1(n18444), .A2(n18430), .ZN(n18824) );
  INV_X1 U21499 ( .A(n18824), .ZN(n18718) );
  NOR2_X2 U21500 ( .A1(n18453), .A2(n18431), .ZN(n18823) );
  NAND2_X1 U21501 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18798), .ZN(n18828) );
  INV_X1 U21502 ( .A(n18828), .ZN(n18715) );
  AOI22_X1 U21503 ( .A1(n18446), .A2(n18823), .B1(n18844), .B2(n18715), .ZN(
        n18434) );
  NOR2_X2 U21504 ( .A1(n18432), .A2(n18447), .ZN(n18825) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n18825), .ZN(n18433) );
  OAI211_X1 U21506 ( .C1(n18774), .C2(n18718), .A(n18434), .B(n18433), .ZN(
        P3_U2872) );
  NOR2_X1 U21507 ( .A1(n18444), .A2(n19483), .ZN(n18830) );
  INV_X1 U21508 ( .A(n18830), .ZN(n18780) );
  NOR2_X2 U21509 ( .A1(n18453), .A2(n18435), .ZN(n18829) );
  NAND2_X1 U21510 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18798), .ZN(n18834) );
  INV_X1 U21511 ( .A(n18834), .ZN(n18777) );
  AOI22_X1 U21512 ( .A1(n18446), .A2(n18829), .B1(n18844), .B2(n18777), .ZN(
        n18438) );
  NOR2_X2 U21513 ( .A1(n18436), .A2(n18447), .ZN(n18831) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n18831), .ZN(n18437) );
  OAI211_X1 U21515 ( .C1(n18774), .C2(n18780), .A(n18438), .B(n18437), .ZN(
        P3_U2873) );
  INV_X1 U21516 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18439) );
  NOR2_X1 U21517 ( .A1(n18444), .A2(n18439), .ZN(n18836) );
  INV_X1 U21518 ( .A(n18836), .ZN(n18725) );
  NOR2_X2 U21519 ( .A1(n18453), .A2(n18440), .ZN(n18835) );
  NAND2_X1 U21520 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18798), .ZN(n18840) );
  INV_X1 U21521 ( .A(n18840), .ZN(n18722) );
  AOI22_X1 U21522 ( .A1(n18446), .A2(n18835), .B1(n18844), .B2(n18722), .ZN(
        n18443) );
  NOR2_X2 U21523 ( .A1(n18441), .A2(n18447), .ZN(n18837) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n18837), .ZN(n18442) );
  OAI211_X1 U21525 ( .C1(n18774), .C2(n18725), .A(n18443), .B(n18442), .ZN(
        P3_U2874) );
  NOR2_X1 U21526 ( .A1(n18444), .A2(n19495), .ZN(n18786) );
  INV_X1 U21527 ( .A(n18786), .ZN(n18851) );
  NAND2_X1 U21528 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18798), .ZN(n18791) );
  INV_X1 U21529 ( .A(n18791), .ZN(n18843) );
  NOR2_X2 U21530 ( .A1(n18445), .A2(n18453), .ZN(n18842) );
  AOI22_X1 U21531 ( .A1(n18787), .A2(n18843), .B1(n18446), .B2(n18842), .ZN(
        n18451) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18449), .B1(
        n18511), .B2(n9636), .ZN(n18450) );
  OAI211_X1 U21533 ( .C1(n18736), .C2(n18851), .A(n18451), .B(n18450), .ZN(
        P3_U2875) );
  INV_X1 U21534 ( .A(n18492), .ZN(n18540) );
  NAND2_X1 U21535 ( .A1(n18679), .A2(n18792), .ZN(n18629) );
  NOR2_X1 U21536 ( .A1(n18540), .A2(n18629), .ZN(n18468) );
  AOI22_X1 U21537 ( .A1(n18787), .A2(n18799), .B1(n18793), .B2(n18468), .ZN(
        n18455) );
  NOR2_X1 U21538 ( .A1(n18907), .A2(n18630), .ZN(n18795) );
  NOR2_X1 U21539 ( .A1(n18453), .A2(n18452), .ZN(n18796) );
  INV_X1 U21540 ( .A(n18796), .ZN(n18583) );
  NOR2_X1 U21541 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18583), .ZN(
        n18541) );
  AOI22_X1 U21542 ( .A1(n18798), .A2(n18795), .B1(n18492), .B2(n18541), .ZN(
        n18469) );
  NAND2_X1 U21543 ( .A1(n18492), .A2(n18628), .ZN(n18528) );
  INV_X1 U21544 ( .A(n18528), .ZN(n18534) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18469), .B1(
        n18760), .B2(n18534), .ZN(n18454) );
  OAI211_X1 U21546 ( .C1(n18763), .C2(n18816), .A(n18455), .B(n18454), .ZN(
        P3_U2876) );
  INV_X1 U21547 ( .A(n18816), .ZN(n18846) );
  INV_X1 U21548 ( .A(n18767), .ZN(n18804) );
  AOI22_X1 U21549 ( .A1(n18846), .A2(n18804), .B1(n18803), .B2(n18468), .ZN(
        n18457) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18469), .B1(
        n18805), .B2(n18534), .ZN(n18456) );
  OAI211_X1 U21551 ( .C1(n18774), .C2(n18808), .A(n18457), .B(n18456), .ZN(
        P3_U2877) );
  AOI22_X1 U21552 ( .A1(n18846), .A2(n18812), .B1(n18809), .B2(n18468), .ZN(
        n18459) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18469), .B1(
        n18739), .B2(n18534), .ZN(n18458) );
  OAI211_X1 U21554 ( .C1(n18774), .C2(n18742), .A(n18459), .B(n18458), .ZN(
        P3_U2878) );
  AOI22_X1 U21555 ( .A1(n18787), .A2(n18770), .B1(n18817), .B2(n18468), .ZN(
        n18461) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18469), .B1(
        n18819), .B2(n18534), .ZN(n18460) );
  OAI211_X1 U21557 ( .C1(n18816), .C2(n18714), .A(n18461), .B(n18460), .ZN(
        P3_U2879) );
  AOI22_X1 U21558 ( .A1(n18846), .A2(n18824), .B1(n18823), .B2(n18468), .ZN(
        n18463) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18469), .B1(
        n18825), .B2(n18534), .ZN(n18462) );
  OAI211_X1 U21560 ( .C1(n18774), .C2(n18828), .A(n18463), .B(n18462), .ZN(
        P3_U2880) );
  AOI22_X1 U21561 ( .A1(n18846), .A2(n18830), .B1(n18829), .B2(n18468), .ZN(
        n18465) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18469), .B1(
        n18831), .B2(n18534), .ZN(n18464) );
  OAI211_X1 U21563 ( .C1(n18774), .C2(n18834), .A(n18465), .B(n18464), .ZN(
        P3_U2881) );
  AOI22_X1 U21564 ( .A1(n18787), .A2(n18722), .B1(n18835), .B2(n18468), .ZN(
        n18467) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18469), .B1(
        n18837), .B2(n18534), .ZN(n18466) );
  OAI211_X1 U21566 ( .C1(n18816), .C2(n18725), .A(n18467), .B(n18466), .ZN(
        P3_U2882) );
  AOI22_X1 U21567 ( .A1(n18846), .A2(n18843), .B1(n18842), .B2(n18468), .ZN(
        n18471) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18469), .B1(
        n9636), .B2(n18534), .ZN(n18470) );
  OAI211_X1 U21569 ( .C1(n18774), .C2(n18851), .A(n18471), .B(n18470), .ZN(
        P3_U2883) );
  INV_X1 U21570 ( .A(n18760), .ZN(n18802) );
  NAND2_X1 U21571 ( .A1(n18653), .A2(n18492), .ZN(n18538) );
  INV_X1 U21572 ( .A(n18763), .ZN(n18794) );
  INV_X1 U21573 ( .A(n18538), .ZN(n18558) );
  NOR2_X1 U21574 ( .A1(n18534), .A2(n18558), .ZN(n18516) );
  NOR2_X1 U21575 ( .A1(n18927), .A2(n18516), .ZN(n18488) );
  AOI22_X1 U21576 ( .A1(n18794), .A2(n18511), .B1(n18793), .B2(n18488), .ZN(
        n18475) );
  OAI21_X1 U21577 ( .B1(n18472), .B2(n18654), .A(n18516), .ZN(n18473) );
  OAI211_X1 U21578 ( .C1(n18558), .C2(n19028), .A(n18705), .B(n18473), .ZN(
        n18489) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18489), .B1(
        n18846), .B2(n18799), .ZN(n18474) );
  OAI211_X1 U21580 ( .C1(n18802), .C2(n18538), .A(n18475), .B(n18474), .ZN(
        P3_U2884) );
  AOI22_X1 U21581 ( .A1(n18511), .A2(n18804), .B1(n18803), .B2(n18488), .ZN(
        n18477) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18489), .B1(
        n18805), .B2(n18558), .ZN(n18476) );
  OAI211_X1 U21583 ( .C1(n18816), .C2(n18808), .A(n18477), .B(n18476), .ZN(
        P3_U2885) );
  INV_X1 U21584 ( .A(n18739), .ZN(n18815) );
  AOI22_X1 U21585 ( .A1(n18846), .A2(n18811), .B1(n18809), .B2(n18488), .ZN(
        n18479) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18489), .B1(
        n18511), .B2(n18812), .ZN(n18478) );
  OAI211_X1 U21587 ( .C1(n18815), .C2(n18538), .A(n18479), .B(n18478), .ZN(
        P3_U2886) );
  AOI22_X1 U21588 ( .A1(n18846), .A2(n18770), .B1(n18817), .B2(n18488), .ZN(
        n18481) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18489), .B1(
        n18819), .B2(n18558), .ZN(n18480) );
  OAI211_X1 U21590 ( .C1(n18507), .C2(n18714), .A(n18481), .B(n18480), .ZN(
        P3_U2887) );
  AOI22_X1 U21591 ( .A1(n18511), .A2(n18824), .B1(n18823), .B2(n18488), .ZN(
        n18483) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18489), .B1(
        n18825), .B2(n18558), .ZN(n18482) );
  OAI211_X1 U21593 ( .C1(n18816), .C2(n18828), .A(n18483), .B(n18482), .ZN(
        P3_U2888) );
  AOI22_X1 U21594 ( .A1(n18511), .A2(n18830), .B1(n18829), .B2(n18488), .ZN(
        n18485) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18489), .B1(
        n18831), .B2(n18558), .ZN(n18484) );
  OAI211_X1 U21596 ( .C1(n18816), .C2(n18834), .A(n18485), .B(n18484), .ZN(
        P3_U2889) );
  AOI22_X1 U21597 ( .A1(n18846), .A2(n18722), .B1(n18835), .B2(n18488), .ZN(
        n18487) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18489), .B1(
        n18837), .B2(n18558), .ZN(n18486) );
  OAI211_X1 U21599 ( .C1(n18507), .C2(n18725), .A(n18487), .B(n18486), .ZN(
        P3_U2890) );
  AOI22_X1 U21600 ( .A1(n18846), .A2(n18786), .B1(n18842), .B2(n18488), .ZN(
        n18491) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18489), .B1(
        n9636), .B2(n18558), .ZN(n18490) );
  OAI211_X1 U21602 ( .C1(n18507), .C2(n18791), .A(n18491), .B(n18490), .ZN(
        P3_U2891) );
  OAI211_X1 U21603 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18758), .A(
        n18492), .B(n18796), .ZN(n18512) );
  INV_X1 U21604 ( .A(n18512), .ZN(n18496) );
  AOI22_X1 U21605 ( .A1(n18511), .A2(n18799), .B1(n18793), .B2(n18510), .ZN(
        n18494) );
  NAND2_X1 U21606 ( .A1(n18898), .A2(n18492), .ZN(n18577) );
  INV_X1 U21607 ( .A(n18577), .ZN(n18579) );
  AOI22_X1 U21608 ( .A1(n18794), .A2(n18534), .B1(n18760), .B2(n18579), .ZN(
        n18493) );
  OAI211_X1 U21609 ( .C1(n18496), .C2(n18495), .A(n18494), .B(n18493), .ZN(
        P3_U2892) );
  AOI22_X1 U21610 ( .A1(n18511), .A2(n18764), .B1(n18803), .B2(n18510), .ZN(
        n18498) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18512), .B1(
        n18805), .B2(n18579), .ZN(n18497) );
  OAI211_X1 U21612 ( .C1(n18767), .C2(n18528), .A(n18498), .B(n18497), .ZN(
        P3_U2893) );
  AOI22_X1 U21613 ( .A1(n18812), .A2(n18534), .B1(n18809), .B2(n18510), .ZN(
        n18500) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18512), .B1(
        n18739), .B2(n18579), .ZN(n18499) );
  OAI211_X1 U21615 ( .C1(n18507), .C2(n18742), .A(n18500), .B(n18499), .ZN(
        P3_U2894) );
  AOI22_X1 U21616 ( .A1(n18511), .A2(n18770), .B1(n18817), .B2(n18510), .ZN(
        n18502) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18512), .B1(
        n18819), .B2(n18579), .ZN(n18501) );
  OAI211_X1 U21618 ( .C1(n18714), .C2(n18528), .A(n18502), .B(n18501), .ZN(
        P3_U2895) );
  AOI22_X1 U21619 ( .A1(n18511), .A2(n18715), .B1(n18823), .B2(n18510), .ZN(
        n18504) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18512), .B1(
        n18825), .B2(n18579), .ZN(n18503) );
  OAI211_X1 U21621 ( .C1(n18718), .C2(n18528), .A(n18504), .B(n18503), .ZN(
        P3_U2896) );
  AOI22_X1 U21622 ( .A1(n18830), .A2(n18534), .B1(n18829), .B2(n18510), .ZN(
        n18506) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18512), .B1(
        n18831), .B2(n18579), .ZN(n18505) );
  OAI211_X1 U21624 ( .C1(n18507), .C2(n18834), .A(n18506), .B(n18505), .ZN(
        P3_U2897) );
  AOI22_X1 U21625 ( .A1(n18511), .A2(n18722), .B1(n18835), .B2(n18510), .ZN(
        n18509) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18512), .B1(
        n18837), .B2(n18579), .ZN(n18508) );
  OAI211_X1 U21627 ( .C1(n18725), .C2(n18528), .A(n18509), .B(n18508), .ZN(
        P3_U2898) );
  AOI22_X1 U21628 ( .A1(n18511), .A2(n18786), .B1(n18842), .B2(n18510), .ZN(
        n18514) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18512), .B1(
        n9636), .B2(n18579), .ZN(n18513) );
  OAI211_X1 U21630 ( .C1(n18791), .C2(n18528), .A(n18514), .B(n18513), .ZN(
        P3_U2899) );
  NAND2_X1 U21631 ( .A1(n18899), .A2(n18585), .ZN(n18605) );
  NAND2_X1 U21632 ( .A1(n18577), .A2(n18605), .ZN(n18562) );
  INV_X1 U21633 ( .A(n18562), .ZN(n18515) );
  NOR2_X1 U21634 ( .A1(n18927), .A2(n18515), .ZN(n18533) );
  AOI22_X1 U21635 ( .A1(n18793), .A2(n18533), .B1(n18799), .B2(n18534), .ZN(
        n18519) );
  INV_X1 U21636 ( .A(n18605), .ZN(n18598) );
  OAI21_X1 U21637 ( .B1(n18516), .B2(n18654), .A(n18515), .ZN(n18517) );
  OAI211_X1 U21638 ( .C1(n18598), .C2(n19028), .A(n18705), .B(n18517), .ZN(
        n18535) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18535), .B1(
        n18760), .B2(n18598), .ZN(n18518) );
  OAI211_X1 U21640 ( .C1(n18763), .C2(n18538), .A(n18519), .B(n18518), .ZN(
        P3_U2900) );
  AOI22_X1 U21641 ( .A1(n18764), .A2(n18534), .B1(n18803), .B2(n18533), .ZN(
        n18521) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18535), .B1(
        n18805), .B2(n18598), .ZN(n18520) );
  OAI211_X1 U21643 ( .C1(n18767), .C2(n18538), .A(n18521), .B(n18520), .ZN(
        P3_U2901) );
  AOI22_X1 U21644 ( .A1(n18811), .A2(n18534), .B1(n18809), .B2(n18533), .ZN(
        n18523) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18535), .B1(
        n18812), .B2(n18558), .ZN(n18522) );
  OAI211_X1 U21646 ( .C1(n18815), .C2(n18605), .A(n18523), .B(n18522), .ZN(
        P3_U2902) );
  AOI22_X1 U21647 ( .A1(n18770), .A2(n18534), .B1(n18817), .B2(n18533), .ZN(
        n18525) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18535), .B1(
        n18819), .B2(n18598), .ZN(n18524) );
  OAI211_X1 U21649 ( .C1(n18714), .C2(n18538), .A(n18525), .B(n18524), .ZN(
        P3_U2903) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18535), .B1(
        n18823), .B2(n18533), .ZN(n18527) );
  AOI22_X1 U21651 ( .A1(n18824), .A2(n18558), .B1(n18825), .B2(n18598), .ZN(
        n18526) );
  OAI211_X1 U21652 ( .C1(n18828), .C2(n18528), .A(n18527), .B(n18526), .ZN(
        P3_U2904) );
  AOI22_X1 U21653 ( .A1(n18777), .A2(n18534), .B1(n18829), .B2(n18533), .ZN(
        n18530) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18535), .B1(
        n18831), .B2(n18598), .ZN(n18529) );
  OAI211_X1 U21655 ( .C1(n18780), .C2(n18538), .A(n18530), .B(n18529), .ZN(
        P3_U2905) );
  AOI22_X1 U21656 ( .A1(n18722), .A2(n18534), .B1(n18835), .B2(n18533), .ZN(
        n18532) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18535), .B1(
        n18837), .B2(n18598), .ZN(n18531) );
  OAI211_X1 U21658 ( .C1(n18725), .C2(n18538), .A(n18532), .B(n18531), .ZN(
        P3_U2906) );
  AOI22_X1 U21659 ( .A1(n18786), .A2(n18534), .B1(n18842), .B2(n18533), .ZN(
        n18537) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18535), .B1(
        n9636), .B2(n18598), .ZN(n18536) );
  OAI211_X1 U21661 ( .C1(n18791), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P3_U2907) );
  NAND2_X1 U21662 ( .A1(n18628), .A2(n18585), .ZN(n18622) );
  NOR2_X1 U21663 ( .A1(n18629), .A2(n18539), .ZN(n18557) );
  AOI22_X1 U21664 ( .A1(n18794), .A2(n18579), .B1(n18793), .B2(n18557), .ZN(
        n18544) );
  NOR2_X1 U21665 ( .A1(n18679), .A2(n18540), .ZN(n18542) );
  AOI22_X1 U21666 ( .A1(n18798), .A2(n18542), .B1(n18541), .B2(n18585), .ZN(
        n18559) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18559), .B1(
        n18799), .B2(n18558), .ZN(n18543) );
  OAI211_X1 U21668 ( .C1(n18802), .C2(n18622), .A(n18544), .B(n18543), .ZN(
        P3_U2908) );
  INV_X1 U21669 ( .A(n18805), .ZN(n18661) );
  AOI22_X1 U21670 ( .A1(n18764), .A2(n18558), .B1(n18803), .B2(n18557), .ZN(
        n18546) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18559), .B1(
        n18804), .B2(n18579), .ZN(n18545) );
  OAI211_X1 U21672 ( .C1(n18661), .C2(n18622), .A(n18546), .B(n18545), .ZN(
        P3_U2909) );
  AOI22_X1 U21673 ( .A1(n18812), .A2(n18579), .B1(n18809), .B2(n18557), .ZN(
        n18548) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18559), .B1(
        n18811), .B2(n18558), .ZN(n18547) );
  OAI211_X1 U21675 ( .C1(n18815), .C2(n18622), .A(n18548), .B(n18547), .ZN(
        P3_U2910) );
  AOI22_X1 U21676 ( .A1(n18770), .A2(n18558), .B1(n18817), .B2(n18557), .ZN(
        n18550) );
  INV_X1 U21677 ( .A(n18622), .ZN(n18625) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18559), .B1(
        n18819), .B2(n18625), .ZN(n18549) );
  OAI211_X1 U21679 ( .C1(n18714), .C2(n18577), .A(n18550), .B(n18549), .ZN(
        P3_U2911) );
  AOI22_X1 U21680 ( .A1(n18715), .A2(n18558), .B1(n18823), .B2(n18557), .ZN(
        n18552) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18559), .B1(
        n18825), .B2(n18625), .ZN(n18551) );
  OAI211_X1 U21682 ( .C1(n18718), .C2(n18577), .A(n18552), .B(n18551), .ZN(
        P3_U2912) );
  AOI22_X1 U21683 ( .A1(n18777), .A2(n18558), .B1(n18829), .B2(n18557), .ZN(
        n18554) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18559), .B1(
        n18831), .B2(n18625), .ZN(n18553) );
  OAI211_X1 U21685 ( .C1(n18780), .C2(n18577), .A(n18554), .B(n18553), .ZN(
        P3_U2913) );
  AOI22_X1 U21686 ( .A1(n18722), .A2(n18558), .B1(n18835), .B2(n18557), .ZN(
        n18556) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18559), .B1(
        n18837), .B2(n18625), .ZN(n18555) );
  OAI211_X1 U21688 ( .C1(n18725), .C2(n18577), .A(n18556), .B(n18555), .ZN(
        P3_U2914) );
  AOI22_X1 U21689 ( .A1(n18786), .A2(n18558), .B1(n18842), .B2(n18557), .ZN(
        n18561) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18559), .B1(
        n9636), .B2(n18625), .ZN(n18560) );
  OAI211_X1 U21691 ( .C1(n18791), .C2(n18577), .A(n18561), .B(n18560), .ZN(
        P3_U2915) );
  NAND2_X1 U21692 ( .A1(n18653), .A2(n18585), .ZN(n18652) );
  NAND2_X1 U21693 ( .A1(n18622), .A2(n18652), .ZN(n18606) );
  OAI221_X1 U21694 ( .B1(n18606), .B2(n18758), .C1(n18606), .C2(n18562), .A(
        n18756), .ZN(n18580) );
  AND2_X1 U21695 ( .A1(n18792), .A2(n18606), .ZN(n18578) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18580), .B1(
        n18793), .B2(n18578), .ZN(n18564) );
  AOI22_X1 U21697 ( .A1(n18794), .A2(n18598), .B1(n18799), .B2(n18579), .ZN(
        n18563) );
  OAI211_X1 U21698 ( .C1(n18802), .C2(n18652), .A(n18564), .B(n18563), .ZN(
        P3_U2916) );
  AOI22_X1 U21699 ( .A1(n18764), .A2(n18579), .B1(n18803), .B2(n18578), .ZN(
        n18566) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18580), .B1(
        n18804), .B2(n18598), .ZN(n18565) );
  OAI211_X1 U21701 ( .C1(n18661), .C2(n18652), .A(n18566), .B(n18565), .ZN(
        P3_U2917) );
  AOI22_X1 U21702 ( .A1(n18811), .A2(n18579), .B1(n18809), .B2(n18578), .ZN(
        n18568) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18580), .B1(
        n18812), .B2(n18598), .ZN(n18567) );
  OAI211_X1 U21704 ( .C1(n18815), .C2(n18652), .A(n18568), .B(n18567), .ZN(
        P3_U2918) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18580), .B1(
        n18817), .B2(n18578), .ZN(n18570) );
  INV_X1 U21706 ( .A(n18652), .ZN(n18643) );
  AOI22_X1 U21707 ( .A1(n18819), .A2(n18643), .B1(n18770), .B2(n18579), .ZN(
        n18569) );
  OAI211_X1 U21708 ( .C1(n18714), .C2(n18605), .A(n18570), .B(n18569), .ZN(
        P3_U2919) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18580), .B1(
        n18823), .B2(n18578), .ZN(n18572) );
  AOI22_X1 U21710 ( .A1(n18824), .A2(n18598), .B1(n18825), .B2(n18643), .ZN(
        n18571) );
  OAI211_X1 U21711 ( .C1(n18828), .C2(n18577), .A(n18572), .B(n18571), .ZN(
        P3_U2920) );
  AOI22_X1 U21712 ( .A1(n18830), .A2(n18598), .B1(n18829), .B2(n18578), .ZN(
        n18574) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18580), .B1(
        n18831), .B2(n18643), .ZN(n18573) );
  OAI211_X1 U21714 ( .C1(n18834), .C2(n18577), .A(n18574), .B(n18573), .ZN(
        P3_U2921) );
  AOI22_X1 U21715 ( .A1(n18836), .A2(n18598), .B1(n18835), .B2(n18578), .ZN(
        n18576) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18580), .B1(
        n18837), .B2(n18643), .ZN(n18575) );
  OAI211_X1 U21717 ( .C1(n18840), .C2(n18577), .A(n18576), .B(n18575), .ZN(
        P3_U2922) );
  AOI22_X1 U21718 ( .A1(n18786), .A2(n18579), .B1(n18842), .B2(n18578), .ZN(
        n18582) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18580), .B1(
        n9636), .B2(n18643), .ZN(n18581) );
  OAI211_X1 U21720 ( .C1(n18791), .C2(n18605), .A(n18582), .B(n18581), .ZN(
        P3_U2923) );
  AOI22_X1 U21721 ( .A1(n18793), .A2(n18601), .B1(n18799), .B2(n18598), .ZN(
        n18587) );
  AOI21_X1 U21722 ( .B1(n18679), .B2(n18654), .A(n18583), .ZN(n18584) );
  NAND2_X1 U21723 ( .A1(n18584), .A2(n18585), .ZN(n18602) );
  NAND2_X1 U21724 ( .A1(n18898), .A2(n18585), .ZN(n18670) );
  INV_X1 U21725 ( .A(n18670), .ZN(n18674) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18602), .B1(
        n18760), .B2(n18674), .ZN(n18586) );
  OAI211_X1 U21727 ( .C1(n18763), .C2(n18622), .A(n18587), .B(n18586), .ZN(
        P3_U2924) );
  AOI22_X1 U21728 ( .A1(n18804), .A2(n18625), .B1(n18803), .B2(n18601), .ZN(
        n18589) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18602), .B1(
        n18805), .B2(n18674), .ZN(n18588) );
  OAI211_X1 U21730 ( .C1(n18808), .C2(n18605), .A(n18589), .B(n18588), .ZN(
        P3_U2925) );
  AOI22_X1 U21731 ( .A1(n18812), .A2(n18625), .B1(n18809), .B2(n18601), .ZN(
        n18591) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18602), .B1(
        n18739), .B2(n18674), .ZN(n18590) );
  OAI211_X1 U21733 ( .C1(n18742), .C2(n18605), .A(n18591), .B(n18590), .ZN(
        P3_U2926) );
  AOI22_X1 U21734 ( .A1(n18818), .A2(n18625), .B1(n18817), .B2(n18601), .ZN(
        n18593) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18602), .B1(
        n18819), .B2(n18674), .ZN(n18592) );
  OAI211_X1 U21736 ( .C1(n18822), .C2(n18605), .A(n18593), .B(n18592), .ZN(
        P3_U2927) );
  AOI22_X1 U21737 ( .A1(n18824), .A2(n18625), .B1(n18823), .B2(n18601), .ZN(
        n18595) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18602), .B1(
        n18825), .B2(n18674), .ZN(n18594) );
  OAI211_X1 U21739 ( .C1(n18828), .C2(n18605), .A(n18595), .B(n18594), .ZN(
        P3_U2928) );
  AOI22_X1 U21740 ( .A1(n18777), .A2(n18598), .B1(n18829), .B2(n18601), .ZN(
        n18597) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18602), .B1(
        n18831), .B2(n18674), .ZN(n18596) );
  OAI211_X1 U21742 ( .C1(n18780), .C2(n18622), .A(n18597), .B(n18596), .ZN(
        P3_U2929) );
  AOI22_X1 U21743 ( .A1(n18722), .A2(n18598), .B1(n18835), .B2(n18601), .ZN(
        n18600) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18602), .B1(
        n18837), .B2(n18674), .ZN(n18599) );
  OAI211_X1 U21745 ( .C1(n18725), .C2(n18622), .A(n18600), .B(n18599), .ZN(
        P3_U2930) );
  AOI22_X1 U21746 ( .A1(n18843), .A2(n18625), .B1(n18842), .B2(n18601), .ZN(
        n18604) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18602), .B1(
        n9636), .B2(n18674), .ZN(n18603) );
  OAI211_X1 U21748 ( .C1(n18851), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2931) );
  NAND2_X1 U21749 ( .A1(n18899), .A2(n18680), .ZN(n18695) );
  NAND2_X1 U21750 ( .A1(n18670), .A2(n18695), .ZN(n18607) );
  INV_X1 U21751 ( .A(n18607), .ZN(n18655) );
  NOR2_X1 U21752 ( .A1(n18927), .A2(n18655), .ZN(n18623) );
  AOI22_X1 U21753 ( .A1(n18793), .A2(n18623), .B1(n18799), .B2(n18625), .ZN(
        n18609) );
  OAI221_X1 U21754 ( .B1(n18607), .B2(n18758), .C1(n18607), .C2(n18606), .A(
        n18756), .ZN(n18624) );
  INV_X1 U21755 ( .A(n18695), .ZN(n18697) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18624), .B1(
        n18760), .B2(n18697), .ZN(n18608) );
  OAI211_X1 U21757 ( .C1(n18763), .C2(n18652), .A(n18609), .B(n18608), .ZN(
        P3_U2932) );
  AOI22_X1 U21758 ( .A1(n18804), .A2(n18643), .B1(n18803), .B2(n18623), .ZN(
        n18611) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18624), .B1(
        n18805), .B2(n18697), .ZN(n18610) );
  OAI211_X1 U21760 ( .C1(n18808), .C2(n18622), .A(n18611), .B(n18610), .ZN(
        P3_U2933) );
  AOI22_X1 U21761 ( .A1(n18812), .A2(n18643), .B1(n18809), .B2(n18623), .ZN(
        n18613) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18624), .B1(
        n18739), .B2(n18697), .ZN(n18612) );
  OAI211_X1 U21763 ( .C1(n18742), .C2(n18622), .A(n18613), .B(n18612), .ZN(
        P3_U2934) );
  AOI22_X1 U21764 ( .A1(n18770), .A2(n18625), .B1(n18817), .B2(n18623), .ZN(
        n18615) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18624), .B1(
        n18819), .B2(n18697), .ZN(n18614) );
  OAI211_X1 U21766 ( .C1(n18714), .C2(n18652), .A(n18615), .B(n18614), .ZN(
        P3_U2935) );
  AOI22_X1 U21767 ( .A1(n18824), .A2(n18643), .B1(n18823), .B2(n18623), .ZN(
        n18617) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18624), .B1(
        n18825), .B2(n18697), .ZN(n18616) );
  OAI211_X1 U21769 ( .C1(n18828), .C2(n18622), .A(n18617), .B(n18616), .ZN(
        P3_U2936) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18624), .B1(
        n18829), .B2(n18623), .ZN(n18619) );
  AOI22_X1 U21771 ( .A1(n18830), .A2(n18643), .B1(n18831), .B2(n18697), .ZN(
        n18618) );
  OAI211_X1 U21772 ( .C1(n18834), .C2(n18622), .A(n18619), .B(n18618), .ZN(
        P3_U2937) );
  AOI22_X1 U21773 ( .A1(n18836), .A2(n18643), .B1(n18835), .B2(n18623), .ZN(
        n18621) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18624), .B1(
        n18837), .B2(n18697), .ZN(n18620) );
  OAI211_X1 U21775 ( .C1(n18840), .C2(n18622), .A(n18621), .B(n18620), .ZN(
        P3_U2938) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18624), .B1(
        n18842), .B2(n18623), .ZN(n18627) );
  AOI22_X1 U21777 ( .A1(n18786), .A2(n18625), .B1(n9636), .B2(n18697), .ZN(
        n18626) );
  OAI211_X1 U21778 ( .C1(n18791), .C2(n18652), .A(n18627), .B(n18626), .ZN(
        P3_U2939) );
  NAND2_X1 U21779 ( .A1(n18628), .A2(n18680), .ZN(n18721) );
  INV_X1 U21780 ( .A(n18680), .ZN(n18678) );
  NOR2_X1 U21781 ( .A1(n18629), .A2(n18678), .ZN(n18648) );
  AOI22_X1 U21782 ( .A1(n18793), .A2(n18648), .B1(n18799), .B2(n18643), .ZN(
        n18634) );
  NOR2_X1 U21783 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18630), .ZN(
        n18632) );
  NOR2_X1 U21784 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18678), .ZN(
        n18631) );
  AOI22_X1 U21785 ( .A1(n18798), .A2(n18632), .B1(n18796), .B2(n18631), .ZN(
        n18649) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18649), .B1(
        n18794), .B2(n18674), .ZN(n18633) );
  OAI211_X1 U21787 ( .C1(n18802), .C2(n18721), .A(n18634), .B(n18633), .ZN(
        P3_U2940) );
  AOI22_X1 U21788 ( .A1(n18764), .A2(n18643), .B1(n18803), .B2(n18648), .ZN(
        n18636) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18649), .B1(
        n18804), .B2(n18674), .ZN(n18635) );
  OAI211_X1 U21790 ( .C1(n18661), .C2(n18721), .A(n18636), .B(n18635), .ZN(
        P3_U2941) );
  AOI22_X1 U21791 ( .A1(n18812), .A2(n18674), .B1(n18809), .B2(n18648), .ZN(
        n18638) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18649), .B1(
        n18811), .B2(n18643), .ZN(n18637) );
  OAI211_X1 U21793 ( .C1(n18815), .C2(n18721), .A(n18638), .B(n18637), .ZN(
        P3_U2942) );
  INV_X1 U21794 ( .A(n18819), .ZN(n18773) );
  AOI22_X1 U21795 ( .A1(n18770), .A2(n18643), .B1(n18817), .B2(n18648), .ZN(
        n18640) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18649), .B1(
        n18818), .B2(n18674), .ZN(n18639) );
  OAI211_X1 U21797 ( .C1(n18773), .C2(n18721), .A(n18640), .B(n18639), .ZN(
        P3_U2943) );
  AOI22_X1 U21798 ( .A1(n18824), .A2(n18674), .B1(n18823), .B2(n18648), .ZN(
        n18642) );
  INV_X1 U21799 ( .A(n18721), .ZN(n18727) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18649), .B1(
        n18825), .B2(n18727), .ZN(n18641) );
  OAI211_X1 U21801 ( .C1(n18828), .C2(n18652), .A(n18642), .B(n18641), .ZN(
        P3_U2944) );
  AOI22_X1 U21802 ( .A1(n18777), .A2(n18643), .B1(n18829), .B2(n18648), .ZN(
        n18645) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18649), .B1(
        n18831), .B2(n18727), .ZN(n18644) );
  OAI211_X1 U21804 ( .C1(n18780), .C2(n18670), .A(n18645), .B(n18644), .ZN(
        P3_U2945) );
  AOI22_X1 U21805 ( .A1(n18836), .A2(n18674), .B1(n18835), .B2(n18648), .ZN(
        n18647) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18649), .B1(
        n18837), .B2(n18727), .ZN(n18646) );
  OAI211_X1 U21807 ( .C1(n18840), .C2(n18652), .A(n18647), .B(n18646), .ZN(
        P3_U2946) );
  AOI22_X1 U21808 ( .A1(n18843), .A2(n18674), .B1(n18842), .B2(n18648), .ZN(
        n18651) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18649), .B1(
        n9636), .B2(n18727), .ZN(n18650) );
  OAI211_X1 U21810 ( .C1(n18851), .C2(n18652), .A(n18651), .B(n18650), .ZN(
        P3_U2947) );
  NAND2_X1 U21811 ( .A1(n18653), .A2(n18680), .ZN(n18755) );
  AOI21_X1 U21812 ( .B1(n18721), .B2(n18755), .A(n18927), .ZN(n18673) );
  AOI22_X1 U21813 ( .A1(n18793), .A2(n18673), .B1(n18799), .B2(n18674), .ZN(
        n18658) );
  INV_X1 U21814 ( .A(n18755), .ZN(n18733) );
  OAI211_X1 U21815 ( .C1(n18655), .C2(n18654), .A(n18721), .B(n18755), .ZN(
        n18656) );
  OAI211_X1 U21816 ( .C1(n18733), .C2(n19028), .A(n18705), .B(n18656), .ZN(
        n18675) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18675), .B1(
        n18794), .B2(n18697), .ZN(n18657) );
  OAI211_X1 U21818 ( .C1(n18802), .C2(n18755), .A(n18658), .B(n18657), .ZN(
        P3_U2948) );
  AOI22_X1 U21819 ( .A1(n18764), .A2(n18674), .B1(n18803), .B2(n18673), .ZN(
        n18660) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18675), .B1(
        n18804), .B2(n18697), .ZN(n18659) );
  OAI211_X1 U21821 ( .C1(n18661), .C2(n18755), .A(n18660), .B(n18659), .ZN(
        P3_U2949) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18675), .B1(
        n18809), .B2(n18673), .ZN(n18663) );
  AOI22_X1 U21823 ( .A1(n18739), .A2(n18733), .B1(n18812), .B2(n18697), .ZN(
        n18662) );
  OAI211_X1 U21824 ( .C1(n18742), .C2(n18670), .A(n18663), .B(n18662), .ZN(
        P3_U2950) );
  AOI22_X1 U21825 ( .A1(n18770), .A2(n18674), .B1(n18817), .B2(n18673), .ZN(
        n18665) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18675), .B1(
        n18818), .B2(n18697), .ZN(n18664) );
  OAI211_X1 U21827 ( .C1(n18773), .C2(n18755), .A(n18665), .B(n18664), .ZN(
        P3_U2951) );
  AOI22_X1 U21828 ( .A1(n18715), .A2(n18674), .B1(n18823), .B2(n18673), .ZN(
        n18667) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18675), .B1(
        n18825), .B2(n18733), .ZN(n18666) );
  OAI211_X1 U21830 ( .C1(n18718), .C2(n18695), .A(n18667), .B(n18666), .ZN(
        P3_U2952) );
  AOI22_X1 U21831 ( .A1(n18830), .A2(n18697), .B1(n18829), .B2(n18673), .ZN(
        n18669) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18675), .B1(
        n18831), .B2(n18733), .ZN(n18668) );
  OAI211_X1 U21833 ( .C1(n18834), .C2(n18670), .A(n18669), .B(n18668), .ZN(
        P3_U2953) );
  AOI22_X1 U21834 ( .A1(n18722), .A2(n18674), .B1(n18835), .B2(n18673), .ZN(
        n18672) );
  AOI22_X1 U21835 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18675), .B1(
        n18837), .B2(n18733), .ZN(n18671) );
  OAI211_X1 U21836 ( .C1(n18725), .C2(n18695), .A(n18672), .B(n18671), .ZN(
        P3_U2954) );
  AOI22_X1 U21837 ( .A1(n18786), .A2(n18674), .B1(n18842), .B2(n18673), .ZN(
        n18677) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18675), .B1(
        n9636), .B2(n18733), .ZN(n18676) );
  OAI211_X1 U21839 ( .C1(n18791), .C2(n18695), .A(n18677), .B(n18676), .ZN(
        P3_U2955) );
  NOR2_X1 U21840 ( .A1(n18679), .A2(n18678), .ZN(n18732) );
  AND2_X1 U21841 ( .A1(n18792), .A2(n18732), .ZN(n18696) );
  AOI22_X1 U21842 ( .A1(n18793), .A2(n18696), .B1(n18799), .B2(n18697), .ZN(
        n18682) );
  OAI211_X1 U21843 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18798), .A(
        n18796), .B(n18680), .ZN(n18698) );
  NAND2_X1 U21844 ( .A1(n18898), .A2(n18680), .ZN(n18783) );
  INV_X1 U21845 ( .A(n18783), .ZN(n18785) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18698), .B1(
        n18760), .B2(n18785), .ZN(n18681) );
  OAI211_X1 U21847 ( .C1(n18763), .C2(n18721), .A(n18682), .B(n18681), .ZN(
        P3_U2956) );
  AOI22_X1 U21848 ( .A1(n18804), .A2(n18727), .B1(n18803), .B2(n18696), .ZN(
        n18684) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18698), .B1(
        n18805), .B2(n18785), .ZN(n18683) );
  OAI211_X1 U21850 ( .C1(n18808), .C2(n18695), .A(n18684), .B(n18683), .ZN(
        P3_U2957) );
  AOI22_X1 U21851 ( .A1(n18812), .A2(n18727), .B1(n18809), .B2(n18696), .ZN(
        n18686) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18698), .B1(
        n18739), .B2(n18785), .ZN(n18685) );
  OAI211_X1 U21853 ( .C1(n18742), .C2(n18695), .A(n18686), .B(n18685), .ZN(
        P3_U2958) );
  AOI22_X1 U21854 ( .A1(n18818), .A2(n18727), .B1(n18817), .B2(n18696), .ZN(
        n18688) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18698), .B1(
        n18819), .B2(n18785), .ZN(n18687) );
  OAI211_X1 U21856 ( .C1(n18822), .C2(n18695), .A(n18688), .B(n18687), .ZN(
        P3_U2959) );
  AOI22_X1 U21857 ( .A1(n18715), .A2(n18697), .B1(n18823), .B2(n18696), .ZN(
        n18690) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18698), .B1(
        n18825), .B2(n18785), .ZN(n18689) );
  OAI211_X1 U21859 ( .C1(n18718), .C2(n18721), .A(n18690), .B(n18689), .ZN(
        P3_U2960) );
  AOI22_X1 U21860 ( .A1(n18777), .A2(n18697), .B1(n18829), .B2(n18696), .ZN(
        n18692) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18698), .B1(
        n18831), .B2(n18785), .ZN(n18691) );
  OAI211_X1 U21862 ( .C1(n18780), .C2(n18721), .A(n18692), .B(n18691), .ZN(
        P3_U2961) );
  AOI22_X1 U21863 ( .A1(n18836), .A2(n18727), .B1(n18835), .B2(n18696), .ZN(
        n18694) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18698), .B1(
        n18837), .B2(n18785), .ZN(n18693) );
  OAI211_X1 U21865 ( .C1(n18840), .C2(n18695), .A(n18694), .B(n18693), .ZN(
        P3_U2962) );
  AOI22_X1 U21866 ( .A1(n18786), .A2(n18697), .B1(n18842), .B2(n18696), .ZN(
        n18700) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18698), .B1(
        n9636), .B2(n18785), .ZN(n18699) );
  OAI211_X1 U21868 ( .C1(n18791), .C2(n18721), .A(n18700), .B(n18699), .ZN(
        P3_U2963) );
  INV_X1 U21869 ( .A(n18797), .ZN(n18731) );
  NOR2_X2 U21870 ( .A1(n18731), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18810) );
  INV_X1 U21871 ( .A(n18810), .ZN(n18850) );
  NAND2_X1 U21872 ( .A1(n18783), .A2(n18850), .ZN(n18757) );
  INV_X1 U21873 ( .A(n18757), .ZN(n18701) );
  NOR2_X1 U21874 ( .A1(n18927), .A2(n18701), .ZN(n18726) );
  AOI22_X1 U21875 ( .A1(n18794), .A2(n18733), .B1(n18793), .B2(n18726), .ZN(
        n18707) );
  OAI21_X1 U21876 ( .B1(n18703), .B2(n18702), .A(n18701), .ZN(n18704) );
  OAI211_X1 U21877 ( .C1(n18810), .C2(n19028), .A(n18705), .B(n18704), .ZN(
        n18728) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18728), .B1(
        n18799), .B2(n18727), .ZN(n18706) );
  OAI211_X1 U21879 ( .C1(n18802), .C2(n18850), .A(n18707), .B(n18706), .ZN(
        P3_U2964) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18728), .B1(
        n18803), .B2(n18726), .ZN(n18709) );
  AOI22_X1 U21881 ( .A1(n18805), .A2(n18810), .B1(n18764), .B2(n18727), .ZN(
        n18708) );
  OAI211_X1 U21882 ( .C1(n18767), .C2(n18755), .A(n18709), .B(n18708), .ZN(
        P3_U2965) );
  AOI22_X1 U21883 ( .A1(n18811), .A2(n18727), .B1(n18809), .B2(n18726), .ZN(
        n18711) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18728), .B1(
        n18812), .B2(n18733), .ZN(n18710) );
  OAI211_X1 U21885 ( .C1(n18815), .C2(n18850), .A(n18711), .B(n18710), .ZN(
        P3_U2966) );
  AOI22_X1 U21886 ( .A1(n18770), .A2(n18727), .B1(n18817), .B2(n18726), .ZN(
        n18713) );
  AOI22_X1 U21887 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18728), .B1(
        n18819), .B2(n18810), .ZN(n18712) );
  OAI211_X1 U21888 ( .C1(n18714), .C2(n18755), .A(n18713), .B(n18712), .ZN(
        P3_U2967) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18728), .B1(
        n18823), .B2(n18726), .ZN(n18717) );
  AOI22_X1 U21890 ( .A1(n18825), .A2(n18810), .B1(n18715), .B2(n18727), .ZN(
        n18716) );
  OAI211_X1 U21891 ( .C1(n18718), .C2(n18755), .A(n18717), .B(n18716), .ZN(
        P3_U2968) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18728), .B1(
        n18829), .B2(n18726), .ZN(n18720) );
  AOI22_X1 U21893 ( .A1(n18830), .A2(n18733), .B1(n18831), .B2(n18810), .ZN(
        n18719) );
  OAI211_X1 U21894 ( .C1(n18834), .C2(n18721), .A(n18720), .B(n18719), .ZN(
        P3_U2969) );
  AOI22_X1 U21895 ( .A1(n18722), .A2(n18727), .B1(n18835), .B2(n18726), .ZN(
        n18724) );
  AOI22_X1 U21896 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18728), .B1(
        n18837), .B2(n18810), .ZN(n18723) );
  OAI211_X1 U21897 ( .C1(n18725), .C2(n18755), .A(n18724), .B(n18723), .ZN(
        P3_U2970) );
  AOI22_X1 U21898 ( .A1(n18786), .A2(n18727), .B1(n18842), .B2(n18726), .ZN(
        n18730) );
  AOI22_X1 U21899 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18728), .B1(
        n9636), .B2(n18810), .ZN(n18729) );
  OAI211_X1 U21900 ( .C1(n18791), .C2(n18755), .A(n18730), .B(n18729), .ZN(
        P3_U2971) );
  NOR2_X1 U21901 ( .A1(n18927), .A2(n18731), .ZN(n18751) );
  AOI22_X1 U21902 ( .A1(n18794), .A2(n18785), .B1(n18793), .B2(n18751), .ZN(
        n18735) );
  AOI22_X1 U21903 ( .A1(n18798), .A2(n18732), .B1(n18797), .B2(n18796), .ZN(
        n18752) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18752), .B1(
        n18799), .B2(n18733), .ZN(n18734) );
  OAI211_X1 U21905 ( .C1(n18802), .C2(n18736), .A(n18735), .B(n18734), .ZN(
        P3_U2972) );
  AOI22_X1 U21906 ( .A1(n18804), .A2(n18785), .B1(n18803), .B2(n18751), .ZN(
        n18738) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18752), .B1(
        n18844), .B2(n18805), .ZN(n18737) );
  OAI211_X1 U21908 ( .C1(n18808), .C2(n18755), .A(n18738), .B(n18737), .ZN(
        P3_U2973) );
  AOI22_X1 U21909 ( .A1(n18812), .A2(n18785), .B1(n18809), .B2(n18751), .ZN(
        n18741) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18752), .B1(
        n18844), .B2(n18739), .ZN(n18740) );
  OAI211_X1 U21911 ( .C1(n18742), .C2(n18755), .A(n18741), .B(n18740), .ZN(
        P3_U2974) );
  AOI22_X1 U21912 ( .A1(n18818), .A2(n18785), .B1(n18817), .B2(n18751), .ZN(
        n18744) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18752), .B1(
        n18844), .B2(n18819), .ZN(n18743) );
  OAI211_X1 U21914 ( .C1(n18822), .C2(n18755), .A(n18744), .B(n18743), .ZN(
        P3_U2975) );
  AOI22_X1 U21915 ( .A1(n18824), .A2(n18785), .B1(n18823), .B2(n18751), .ZN(
        n18746) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18752), .B1(
        n18844), .B2(n18825), .ZN(n18745) );
  OAI211_X1 U21917 ( .C1(n18828), .C2(n18755), .A(n18746), .B(n18745), .ZN(
        P3_U2976) );
  AOI22_X1 U21918 ( .A1(n18830), .A2(n18785), .B1(n18829), .B2(n18751), .ZN(
        n18748) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18752), .B1(
        n18844), .B2(n18831), .ZN(n18747) );
  OAI211_X1 U21920 ( .C1(n18834), .C2(n18755), .A(n18748), .B(n18747), .ZN(
        P3_U2977) );
  AOI22_X1 U21921 ( .A1(n18836), .A2(n18785), .B1(n18835), .B2(n18751), .ZN(
        n18750) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18752), .B1(
        n18844), .B2(n18837), .ZN(n18749) );
  OAI211_X1 U21923 ( .C1(n18840), .C2(n18755), .A(n18750), .B(n18749), .ZN(
        P3_U2978) );
  AOI22_X1 U21924 ( .A1(n18843), .A2(n18785), .B1(n18842), .B2(n18751), .ZN(
        n18754) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18752), .B1(
        n18844), .B2(n9636), .ZN(n18753) );
  OAI211_X1 U21926 ( .C1(n18851), .C2(n18755), .A(n18754), .B(n18753), .ZN(
        P3_U2979) );
  AND2_X1 U21927 ( .A1(n18792), .A2(n18759), .ZN(n18784) );
  AOI22_X1 U21928 ( .A1(n18793), .A2(n18784), .B1(n18799), .B2(n18785), .ZN(
        n18762) );
  OAI221_X1 U21929 ( .B1(n18759), .B2(n18758), .C1(n18759), .C2(n18757), .A(
        n18756), .ZN(n18788) );
  AOI22_X1 U21930 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18788), .B1(
        n18787), .B2(n18760), .ZN(n18761) );
  OAI211_X1 U21931 ( .C1(n18763), .C2(n18850), .A(n18762), .B(n18761), .ZN(
        P3_U2980) );
  AOI22_X1 U21932 ( .A1(n18764), .A2(n18785), .B1(n18803), .B2(n18784), .ZN(
        n18766) );
  AOI22_X1 U21933 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18788), .B1(
        n18787), .B2(n18805), .ZN(n18765) );
  OAI211_X1 U21934 ( .C1(n18767), .C2(n18850), .A(n18766), .B(n18765), .ZN(
        P3_U2981) );
  AOI22_X1 U21935 ( .A1(n18811), .A2(n18785), .B1(n18809), .B2(n18784), .ZN(
        n18769) );
  AOI22_X1 U21936 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18788), .B1(
        n18812), .B2(n18810), .ZN(n18768) );
  OAI211_X1 U21937 ( .C1(n18774), .C2(n18815), .A(n18769), .B(n18768), .ZN(
        P3_U2982) );
  AOI22_X1 U21938 ( .A1(n18818), .A2(n18810), .B1(n18817), .B2(n18784), .ZN(
        n18772) );
  AOI22_X1 U21939 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18788), .B1(
        n18770), .B2(n18785), .ZN(n18771) );
  OAI211_X1 U21940 ( .C1(n18774), .C2(n18773), .A(n18772), .B(n18771), .ZN(
        P3_U2983) );
  AOI22_X1 U21941 ( .A1(n18824), .A2(n18810), .B1(n18823), .B2(n18784), .ZN(
        n18776) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18788), .B1(
        n18787), .B2(n18825), .ZN(n18775) );
  OAI211_X1 U21943 ( .C1(n18828), .C2(n18783), .A(n18776), .B(n18775), .ZN(
        P3_U2984) );
  AOI22_X1 U21944 ( .A1(n18777), .A2(n18785), .B1(n18829), .B2(n18784), .ZN(
        n18779) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18788), .B1(
        n18787), .B2(n18831), .ZN(n18778) );
  OAI211_X1 U21946 ( .C1(n18780), .C2(n18850), .A(n18779), .B(n18778), .ZN(
        P3_U2985) );
  AOI22_X1 U21947 ( .A1(n18836), .A2(n18810), .B1(n18835), .B2(n18784), .ZN(
        n18782) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18788), .B1(
        n18787), .B2(n18837), .ZN(n18781) );
  OAI211_X1 U21949 ( .C1(n18840), .C2(n18783), .A(n18782), .B(n18781), .ZN(
        P3_U2986) );
  AOI22_X1 U21950 ( .A1(n18786), .A2(n18785), .B1(n18842), .B2(n18784), .ZN(
        n18790) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18788), .B1(
        n18787), .B2(n9636), .ZN(n18789) );
  OAI211_X1 U21952 ( .C1(n18791), .C2(n18850), .A(n18790), .B(n18789), .ZN(
        P3_U2987) );
  AND2_X1 U21953 ( .A1(n18792), .A2(n18795), .ZN(n18841) );
  AOI22_X1 U21954 ( .A1(n18794), .A2(n18844), .B1(n18793), .B2(n18841), .ZN(
        n18801) );
  AOI22_X1 U21955 ( .A1(n18798), .A2(n18797), .B1(n18796), .B2(n18795), .ZN(
        n18847) );
  AOI22_X1 U21956 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18847), .B1(
        n18799), .B2(n18810), .ZN(n18800) );
  OAI211_X1 U21957 ( .C1(n18816), .C2(n18802), .A(n18801), .B(n18800), .ZN(
        P3_U2988) );
  AOI22_X1 U21958 ( .A1(n18844), .A2(n18804), .B1(n18803), .B2(n18841), .ZN(
        n18807) );
  AOI22_X1 U21959 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18847), .B1(
        n18846), .B2(n18805), .ZN(n18806) );
  OAI211_X1 U21960 ( .C1(n18808), .C2(n18850), .A(n18807), .B(n18806), .ZN(
        P3_U2989) );
  AOI22_X1 U21961 ( .A1(n18811), .A2(n18810), .B1(n18809), .B2(n18841), .ZN(
        n18814) );
  AOI22_X1 U21962 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18847), .B1(
        n18844), .B2(n18812), .ZN(n18813) );
  OAI211_X1 U21963 ( .C1(n18816), .C2(n18815), .A(n18814), .B(n18813), .ZN(
        P3_U2990) );
  AOI22_X1 U21964 ( .A1(n18844), .A2(n18818), .B1(n18817), .B2(n18841), .ZN(
        n18821) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18847), .B1(
        n18846), .B2(n18819), .ZN(n18820) );
  OAI211_X1 U21966 ( .C1(n18822), .C2(n18850), .A(n18821), .B(n18820), .ZN(
        P3_U2991) );
  AOI22_X1 U21967 ( .A1(n18844), .A2(n18824), .B1(n18823), .B2(n18841), .ZN(
        n18827) );
  AOI22_X1 U21968 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18847), .B1(
        n18846), .B2(n18825), .ZN(n18826) );
  OAI211_X1 U21969 ( .C1(n18828), .C2(n18850), .A(n18827), .B(n18826), .ZN(
        P3_U2992) );
  AOI22_X1 U21970 ( .A1(n18844), .A2(n18830), .B1(n18829), .B2(n18841), .ZN(
        n18833) );
  AOI22_X1 U21971 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18847), .B1(
        n18846), .B2(n18831), .ZN(n18832) );
  OAI211_X1 U21972 ( .C1(n18834), .C2(n18850), .A(n18833), .B(n18832), .ZN(
        P3_U2993) );
  AOI22_X1 U21973 ( .A1(n18844), .A2(n18836), .B1(n18835), .B2(n18841), .ZN(
        n18839) );
  AOI22_X1 U21974 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18847), .B1(
        n18846), .B2(n18837), .ZN(n18838) );
  OAI211_X1 U21975 ( .C1(n18840), .C2(n18850), .A(n18839), .B(n18838), .ZN(
        P3_U2994) );
  AOI22_X1 U21976 ( .A1(n18844), .A2(n18843), .B1(n18842), .B2(n18841), .ZN(
        n18849) );
  AOI22_X1 U21977 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18847), .B1(
        n18846), .B2(n9636), .ZN(n18848) );
  OAI211_X1 U21978 ( .C1(n18851), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        P3_U2995) );
  NOR2_X1 U21979 ( .A1(n18881), .A2(n18852), .ZN(n18854) );
  OAI222_X1 U21980 ( .A1(n18858), .A2(n18857), .B1(n18856), .B2(n18855), .C1(
        n18854), .C2(n18853), .ZN(n19066) );
  OAI21_X1 U21981 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18859), .ZN(n18860) );
  OAI211_X1 U21982 ( .C1(n18862), .C2(n18900), .A(n18861), .B(n18860), .ZN(
        n18914) );
  AOI21_X1 U21983 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18864), .A(
        n18863), .ZN(n18889) );
  NAND2_X1 U21984 ( .A1(n18889), .A2(n18865), .ZN(n18895) );
  AOI22_X1 U21985 ( .A1(n18873), .A2(n18895), .B1(n18881), .B2(n18866), .ZN(
        n18867) );
  NOR2_X1 U21986 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18867), .ZN(
        n19030) );
  AOI21_X1 U21987 ( .B1(n18870), .B2(n18869), .A(n18868), .ZN(n18878) );
  OAI22_X1 U21988 ( .A1(n18873), .A2(n18872), .B1(n18871), .B2(n18878), .ZN(
        n18874) );
  AOI21_X1 U21989 ( .B1(n12678), .B2(n18875), .A(n18874), .ZN(n19031) );
  AOI21_X1 U21990 ( .B1(n19031), .B2(n18900), .A(n12533), .ZN(n18876) );
  AOI21_X1 U21991 ( .B1(n18900), .B2(n19030), .A(n18876), .ZN(n18912) );
  INV_X1 U21992 ( .A(n18900), .ZN(n18891) );
  INV_X1 U21993 ( .A(n18877), .ZN(n18883) );
  OAI21_X1 U21994 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18879), .A(
        n18878), .ZN(n18882) );
  AOI22_X1 U21995 ( .A1(n18883), .A2(n18882), .B1(n18881), .B2(n18880), .ZN(
        n18887) );
  NAND3_X1 U21996 ( .A1(n18885), .A2(n18884), .A3(n12540), .ZN(n18886) );
  OAI211_X1 U21997 ( .C1(n18889), .C2(n18888), .A(n18887), .B(n18886), .ZN(
        n19039) );
  AOI22_X1 U21998 ( .A1(n18891), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19039), .B2(n18900), .ZN(n18903) );
  INV_X1 U21999 ( .A(n18892), .ZN(n19045) );
  NAND2_X1 U22000 ( .A1(n18894), .A2(n18893), .ZN(n18896) );
  AOI22_X1 U22001 ( .A1(n19045), .A2(n18896), .B1(n19048), .B2(n18895), .ZN(
        n19041) );
  AOI22_X1 U22002 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18897), .B1(
        n18896), .B2(n12679), .ZN(n19050) );
  AOI222_X1 U22003 ( .A1(n19041), .A2(n19050), .B1(n19041), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n19050), .C2(n18898), .ZN(
        n18901) );
  AOI21_X1 U22004 ( .B1(n18901), .B2(n18900), .A(n18899), .ZN(n18902) );
  AOI21_X1 U22005 ( .B1(n18903), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n18902), .ZN(n18904) );
  INV_X1 U22006 ( .A(n18903), .ZN(n18905) );
  AOI221_X1 U22007 ( .B1(n18904), .B2(n18908), .C1(n18907), .C2(n18908), .A(
        n18905), .ZN(n18911) );
  AOI21_X1 U22008 ( .B1(n18906), .B2(n18905), .A(n18904), .ZN(n18910) );
  NAND2_X1 U22009 ( .A1(n18908), .A2(n18907), .ZN(n18909) );
  OAI22_X1 U22010 ( .A1(n18912), .A2(n18911), .B1(n18910), .B2(n18909), .ZN(
        n18913) );
  NOR4_X1 U22011 ( .A1(n18915), .A2(n19066), .A3(n18914), .A4(n18913), .ZN(
        n18925) );
  AOI22_X1 U22012 ( .A1(n19053), .A2(n19078), .B1(n18943), .B2(n19071), .ZN(
        n18916) );
  INV_X1 U22013 ( .A(n18916), .ZN(n18921) );
  OAI211_X1 U22014 ( .C1(n18918), .C2(n18917), .A(n19069), .B(n18925), .ZN(
        n19027) );
  OAI21_X1 U22015 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19075), .A(n19027), 
        .ZN(n18928) );
  NOR2_X1 U22016 ( .A1(n18919), .A2(n18928), .ZN(n18920) );
  MUX2_X1 U22017 ( .A(n18921), .B(n18920), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18923) );
  OAI211_X1 U22018 ( .C1(n18925), .C2(n18924), .A(n18923), .B(n18922), .ZN(
        P3_U2996) );
  NAND2_X1 U22019 ( .A1(n18943), .A2(n19071), .ZN(n18932) );
  NOR4_X1 U22020 ( .A1(n18926), .A2(n19049), .A3(n19075), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18935) );
  INV_X1 U22021 ( .A(n18935), .ZN(n18931) );
  OR3_X1 U22022 ( .A1(n18929), .A2(n18928), .A3(n18927), .ZN(n18930) );
  NAND4_X1 U22023 ( .A1(n18933), .A2(n18932), .A3(n18931), .A4(n18930), .ZN(
        P3_U2997) );
  OAI21_X1 U22024 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18934), .ZN(n18936) );
  AOI21_X1 U22025 ( .B1(n18937), .B2(n18936), .A(n18935), .ZN(P3_U2998) );
  INV_X1 U22026 ( .A(n19025), .ZN(n18938) );
  AND2_X1 U22027 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18938), .ZN(
        P3_U2999) );
  AND2_X1 U22028 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18938), .ZN(
        P3_U3000) );
  AND2_X1 U22029 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18938), .ZN(
        P3_U3001) );
  AND2_X1 U22030 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18938), .ZN(
        P3_U3002) );
  AND2_X1 U22031 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18938), .ZN(
        P3_U3003) );
  AND2_X1 U22032 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18938), .ZN(
        P3_U3004) );
  AND2_X1 U22033 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18938), .ZN(
        P3_U3005) );
  AND2_X1 U22034 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18938), .ZN(
        P3_U3006) );
  AND2_X1 U22035 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18938), .ZN(
        P3_U3007) );
  AND2_X1 U22036 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18938), .ZN(
        P3_U3008) );
  AND2_X1 U22037 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18938), .ZN(
        P3_U3009) );
  AND2_X1 U22038 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18938), .ZN(
        P3_U3010) );
  AND2_X1 U22039 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18938), .ZN(
        P3_U3011) );
  AND2_X1 U22040 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18938), .ZN(
        P3_U3012) );
  AND2_X1 U22041 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18938), .ZN(
        P3_U3013) );
  AND2_X1 U22042 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18938), .ZN(
        P3_U3014) );
  AND2_X1 U22043 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18938), .ZN(
        P3_U3015) );
  AND2_X1 U22044 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18938), .ZN(
        P3_U3016) );
  AND2_X1 U22045 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18938), .ZN(
        P3_U3017) );
  AND2_X1 U22046 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18938), .ZN(
        P3_U3018) );
  AND2_X1 U22047 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18938), .ZN(
        P3_U3019) );
  AND2_X1 U22048 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18938), .ZN(
        P3_U3020) );
  AND2_X1 U22049 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18938), .ZN(P3_U3021) );
  AND2_X1 U22050 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18938), .ZN(P3_U3022) );
  AND2_X1 U22051 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18938), .ZN(P3_U3023) );
  AND2_X1 U22052 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18938), .ZN(P3_U3024) );
  AND2_X1 U22053 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18938), .ZN(P3_U3025) );
  AND2_X1 U22054 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18938), .ZN(P3_U3026) );
  AND2_X1 U22055 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18938), .ZN(P3_U3027) );
  AND2_X1 U22056 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18938), .ZN(P3_U3028) );
  OAI21_X1 U22057 ( .B1(n18939), .B2(n21071), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18940) );
  AOI22_X1 U22058 ( .A1(n18952), .A2(n18954), .B1(n19084), .B2(n18940), .ZN(
        n18942) );
  INV_X1 U22059 ( .A(NA), .ZN(n21000) );
  OR3_X1 U22060 ( .A1(n21000), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18941) );
  OAI211_X1 U22061 ( .C1(n19075), .C2(n18946), .A(n18942), .B(n18941), .ZN(
        P3_U3029) );
  NOR2_X1 U22062 ( .A1(n18954), .A2(n21071), .ZN(n18950) );
  NOR2_X1 U22063 ( .A1(n18952), .A2(n18950), .ZN(n18944) );
  NAND2_X1 U22064 ( .A1(n18943), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18948) );
  INV_X1 U22065 ( .A(n18948), .ZN(n18947) );
  AOI21_X1 U22066 ( .B1(n18944), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n18947), .ZN(n18945) );
  OAI211_X1 U22067 ( .C1(n21071), .C2(n18946), .A(n18945), .B(n19072), .ZN(
        P3_U3030) );
  AOI221_X1 U22068 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18952), .C1(n21000), 
        .C2(n18952), .A(n18947), .ZN(n18953) );
  OAI22_X1 U22069 ( .A1(NA), .A2(n18948), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18949) );
  OAI22_X1 U22070 ( .A1(n18950), .A2(n18949), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18951) );
  OAI22_X1 U22071 ( .A1(n18953), .A2(n18954), .B1(n18952), .B2(n18951), .ZN(
        P3_U3031) );
  OAI222_X1 U22072 ( .A1(n18956), .A2(n19017), .B1(n18955), .B2(n19083), .C1(
        n18957), .C2(n19013), .ZN(P3_U3032) );
  OAI222_X1 U22073 ( .A1(n19013), .A2(n18959), .B1(n18958), .B2(n19083), .C1(
        n18957), .C2(n19017), .ZN(P3_U3033) );
  OAI222_X1 U22074 ( .A1(n19013), .A2(n18961), .B1(n18960), .B2(n19083), .C1(
        n18959), .C2(n19017), .ZN(P3_U3034) );
  OAI222_X1 U22075 ( .A1(n19013), .A2(n18964), .B1(n18962), .B2(n19083), .C1(
        n18961), .C2(n19017), .ZN(P3_U3035) );
  OAI222_X1 U22076 ( .A1(n18964), .A2(n19017), .B1(n18963), .B2(n19083), .C1(
        n18965), .C2(n19013), .ZN(P3_U3036) );
  OAI222_X1 U22077 ( .A1(n19013), .A2(n18967), .B1(n18966), .B2(n19083), .C1(
        n18965), .C2(n19017), .ZN(P3_U3037) );
  INV_X1 U22078 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18970) );
  OAI222_X1 U22079 ( .A1(n19013), .A2(n18970), .B1(n18968), .B2(n19083), .C1(
        n18967), .C2(n19017), .ZN(P3_U3038) );
  OAI222_X1 U22080 ( .A1(n18970), .A2(n19017), .B1(n18969), .B2(n19083), .C1(
        n18971), .C2(n19013), .ZN(P3_U3039) );
  OAI222_X1 U22081 ( .A1(n19013), .A2(n18973), .B1(n18972), .B2(n19083), .C1(
        n18971), .C2(n19017), .ZN(P3_U3040) );
  OAI222_X1 U22082 ( .A1(n19013), .A2(n18975), .B1(n18974), .B2(n19083), .C1(
        n18973), .C2(n19017), .ZN(P3_U3041) );
  INV_X1 U22083 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18977) );
  OAI222_X1 U22084 ( .A1(n19013), .A2(n18977), .B1(n18976), .B2(n19083), .C1(
        n18975), .C2(n19017), .ZN(P3_U3042) );
  OAI222_X1 U22085 ( .A1(n19013), .A2(n18979), .B1(n18978), .B2(n19083), .C1(
        n18977), .C2(n19017), .ZN(P3_U3043) );
  OAI222_X1 U22086 ( .A1(n19013), .A2(n18982), .B1(n18980), .B2(n19083), .C1(
        n18979), .C2(n19017), .ZN(P3_U3044) );
  OAI222_X1 U22087 ( .A1(n18982), .A2(n19017), .B1(n18981), .B2(n19083), .C1(
        n18983), .C2(n19013), .ZN(P3_U3045) );
  OAI222_X1 U22088 ( .A1(n19013), .A2(n18985), .B1(n18984), .B2(n19083), .C1(
        n18983), .C2(n19017), .ZN(P3_U3046) );
  OAI222_X1 U22089 ( .A1(n19013), .A2(n18988), .B1(n18986), .B2(n19083), .C1(
        n18985), .C2(n19017), .ZN(P3_U3047) );
  OAI222_X1 U22090 ( .A1(n18988), .A2(n19017), .B1(n18987), .B2(n19083), .C1(
        n18989), .C2(n19013), .ZN(P3_U3048) );
  INV_X1 U22091 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18991) );
  OAI222_X1 U22092 ( .A1(n19013), .A2(n18991), .B1(n18990), .B2(n19083), .C1(
        n18989), .C2(n19017), .ZN(P3_U3049) );
  OAI222_X1 U22093 ( .A1(n19013), .A2(n18993), .B1(n18992), .B2(n19083), .C1(
        n18991), .C2(n19017), .ZN(P3_U3050) );
  OAI222_X1 U22094 ( .A1(n19013), .A2(n18996), .B1(n18994), .B2(n19083), .C1(
        n18993), .C2(n19017), .ZN(P3_U3051) );
  OAI222_X1 U22095 ( .A1(n18996), .A2(n19017), .B1(n18995), .B2(n19083), .C1(
        n18997), .C2(n19013), .ZN(P3_U3052) );
  OAI222_X1 U22096 ( .A1(n19013), .A2(n19000), .B1(n18998), .B2(n19083), .C1(
        n18997), .C2(n19017), .ZN(P3_U3053) );
  OAI222_X1 U22097 ( .A1(n19000), .A2(n19017), .B1(n18999), .B2(n19083), .C1(
        n19001), .C2(n19013), .ZN(P3_U3054) );
  INV_X1 U22098 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19003) );
  OAI222_X1 U22099 ( .A1(n19013), .A2(n19003), .B1(n19002), .B2(n19083), .C1(
        n19001), .C2(n19017), .ZN(P3_U3055) );
  INV_X1 U22100 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19005) );
  OAI222_X1 U22101 ( .A1(n19013), .A2(n19005), .B1(n19004), .B2(n19083), .C1(
        n19003), .C2(n19017), .ZN(P3_U3056) );
  OAI222_X1 U22102 ( .A1(n19013), .A2(n19007), .B1(n19006), .B2(n19083), .C1(
        n19005), .C2(n19017), .ZN(P3_U3057) );
  OAI222_X1 U22103 ( .A1(n19013), .A2(n19010), .B1(n19008), .B2(n19083), .C1(
        n19007), .C2(n19017), .ZN(P3_U3058) );
  OAI222_X1 U22104 ( .A1(n19010), .A2(n19017), .B1(n19009), .B2(n19083), .C1(
        n19011), .C2(n19013), .ZN(P3_U3059) );
  OAI222_X1 U22105 ( .A1(n19013), .A2(n19016), .B1(n19012), .B2(n19083), .C1(
        n19011), .C2(n19017), .ZN(P3_U3060) );
  INV_X1 U22106 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19015) );
  OAI222_X1 U22107 ( .A1(n19017), .A2(n19016), .B1(n19015), .B2(n19083), .C1(
        n19014), .C2(n19013), .ZN(P3_U3061) );
  OAI22_X1 U22108 ( .A1(n19084), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19083), .ZN(n19018) );
  INV_X1 U22109 ( .A(n19018), .ZN(P3_U3274) );
  OAI22_X1 U22110 ( .A1(n19084), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19083), .ZN(n19019) );
  INV_X1 U22111 ( .A(n19019), .ZN(P3_U3275) );
  OAI22_X1 U22112 ( .A1(n19084), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19083), .ZN(n19020) );
  INV_X1 U22113 ( .A(n19020), .ZN(P3_U3276) );
  OAI22_X1 U22114 ( .A1(n19084), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19083), .ZN(n19021) );
  INV_X1 U22115 ( .A(n19021), .ZN(P3_U3277) );
  OAI21_X1 U22116 ( .B1(n19025), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19023), 
        .ZN(n19022) );
  INV_X1 U22117 ( .A(n19022), .ZN(P3_U3280) );
  OAI21_X1 U22118 ( .B1(n19025), .B2(n19024), .A(n19023), .ZN(P3_U3281) );
  OAI221_X1 U22119 ( .B1(n19028), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19028), 
        .C2(n19027), .A(n19026), .ZN(P3_U3282) );
  AOI22_X1 U22120 ( .A1(n19087), .A2(n19030), .B1(n19053), .B2(n19029), .ZN(
        n19035) );
  OAI21_X1 U22121 ( .B1(n19032), .B2(n19031), .A(n19054), .ZN(n19033) );
  INV_X1 U22122 ( .A(n19033), .ZN(n19034) );
  OAI22_X1 U22123 ( .A1(n19056), .A2(n19035), .B1(n19034), .B2(n12533), .ZN(
        P3_U3285) );
  OAI22_X1 U22124 ( .A1(n19037), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19036), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19042) );
  NAND2_X1 U22125 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19052) );
  INV_X1 U22126 ( .A(n19052), .ZN(n19043) );
  AOI222_X1 U22127 ( .A1(n19039), .A2(n19087), .B1(n19042), .B2(n19043), .C1(
        n19053), .C2(n19038), .ZN(n19040) );
  AOI22_X1 U22128 ( .A1(n19056), .A2(n12678), .B1(n19040), .B2(n19054), .ZN(
        P3_U3288) );
  INV_X1 U22129 ( .A(n19041), .ZN(n19046) );
  INV_X1 U22130 ( .A(n19042), .ZN(n19044) );
  AOI222_X1 U22131 ( .A1(n19046), .A2(n19087), .B1(n19053), .B2(n19045), .C1(
        n19044), .C2(n19043), .ZN(n19047) );
  AOI22_X1 U22132 ( .A1(n19056), .A2(n19048), .B1(n19047), .B2(n19054), .ZN(
        P3_U3289) );
  OAI21_X1 U22133 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19050), .A(n19049), 
        .ZN(n19051) );
  AOI22_X1 U22134 ( .A1(n19053), .A2(n12679), .B1(n19052), .B2(n19051), .ZN(
        n19055) );
  AOI22_X1 U22135 ( .A1(n19056), .A2(n12679), .B1(n19055), .B2(n19054), .ZN(
        P3_U3290) );
  AOI211_X1 U22136 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19057) );
  AOI21_X1 U22137 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19057), .ZN(n19059) );
  INV_X1 U22138 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19058) );
  AOI22_X1 U22139 ( .A1(n19063), .A2(n19059), .B1(n19058), .B2(n19060), .ZN(
        P3_U3292) );
  NOR2_X1 U22140 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19062) );
  INV_X1 U22141 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19061) );
  AOI22_X1 U22142 ( .A1(n19063), .A2(n19062), .B1(n19061), .B2(n19060), .ZN(
        P3_U3293) );
  INV_X1 U22143 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19090) );
  OAI22_X1 U22144 ( .A1(n19084), .A2(n19090), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n19083), .ZN(n19064) );
  INV_X1 U22145 ( .A(n19064), .ZN(P3_U3294) );
  MUX2_X1 U22146 ( .A(P3_MORE_REG_SCAN_IN), .B(n19066), .S(n19065), .Z(
        P3_U3295) );
  OAI21_X1 U22147 ( .B1(n19069), .B2(n19068), .A(n19067), .ZN(n19070) );
  AOI21_X1 U22148 ( .B1(n19071), .B2(n19075), .A(n19070), .ZN(n19082) );
  AOI21_X1 U22149 ( .B1(n19074), .B2(n19073), .A(n19072), .ZN(n19076) );
  OAI211_X1 U22150 ( .C1(n19077), .C2(n19076), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19075), .ZN(n19079) );
  AOI21_X1 U22151 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19079), .A(n19078), 
        .ZN(n19081) );
  NAND2_X1 U22152 ( .A1(n19082), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19080) );
  OAI21_X1 U22153 ( .B1(n19082), .B2(n19081), .A(n19080), .ZN(P3_U3296) );
  OAI22_X1 U22154 ( .A1(n19084), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19083), .ZN(n19085) );
  INV_X1 U22155 ( .A(n19085), .ZN(P3_U3297) );
  AOI21_X1 U22156 ( .B1(n19087), .B2(n19086), .A(n19089), .ZN(n19093) );
  AOI22_X1 U22157 ( .A1(n19093), .A2(n19090), .B1(n19089), .B2(n19088), .ZN(
        P3_U3298) );
  INV_X1 U22158 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19092) );
  AOI21_X1 U22159 ( .B1(n19093), .B2(n19092), .A(n19091), .ZN(P3_U3299) );
  INV_X1 U22160 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20046) );
  NAND2_X1 U22161 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20046), .ZN(n20037) );
  NOR2_X1 U22162 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20033) );
  INV_X1 U22163 ( .A(n20033), .ZN(n19094) );
  OAI21_X1 U22164 ( .B1(n20043), .B2(n20037), .A(n19094), .ZN(n20096) );
  AOI21_X1 U22165 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20096), .ZN(n19095) );
  INV_X1 U22166 ( .A(n19095), .ZN(P2_U2815) );
  INV_X1 U22167 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19099) );
  OAI22_X1 U22168 ( .A1(n19098), .A2(n19099), .B1(n19097), .B2(n19096), .ZN(
        P2_U2816) );
  INV_X1 U22169 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n19101) );
  AOI21_X1 U22170 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n19099), .A(n20040), 
        .ZN(n19100) );
  OAI22_X1 U22171 ( .A1(n20159), .A2(n19101), .B1(P2_STATE_REG_0__SCAN_IN), 
        .B2(n19100), .ZN(P2_U2817) );
  OAI21_X1 U22172 ( .B1(n20040), .B2(BS16), .A(n20096), .ZN(n20094) );
  OAI21_X1 U22173 ( .B1(n20096), .B2(n20098), .A(n20094), .ZN(P2_U2818) );
  NOR4_X1 U22174 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19105) );
  NOR4_X1 U22175 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19104) );
  NOR4_X1 U22176 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19103) );
  NOR4_X1 U22177 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19102) );
  NAND4_X1 U22178 ( .A1(n19105), .A2(n19104), .A3(n19103), .A4(n19102), .ZN(
        n19111) );
  NOR4_X1 U22179 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19109) );
  AOI211_X1 U22180 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19108) );
  NOR4_X1 U22181 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19107) );
  NOR4_X1 U22182 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19106) );
  NAND4_X1 U22183 ( .A1(n19109), .A2(n19108), .A3(n19107), .A4(n19106), .ZN(
        n19110) );
  NOR2_X1 U22184 ( .A1(n19111), .A2(n19110), .ZN(n19122) );
  INV_X1 U22185 ( .A(n19122), .ZN(n19120) );
  NOR2_X1 U22186 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19120), .ZN(n19114) );
  INV_X1 U22187 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19112) );
  AOI22_X1 U22188 ( .A1(n19114), .A2(n19115), .B1(n19120), .B2(n19112), .ZN(
        P2_U2820) );
  OR3_X1 U22189 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19119) );
  INV_X1 U22190 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19113) );
  AOI22_X1 U22191 ( .A1(n19114), .A2(n19119), .B1(n19120), .B2(n19113), .ZN(
        P2_U2821) );
  INV_X1 U22192 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20095) );
  NAND2_X1 U22193 ( .A1(n19114), .A2(n20095), .ZN(n19118) );
  OAI21_X1 U22194 ( .B1(n19115), .B2(n13256), .A(n19122), .ZN(n19116) );
  OAI21_X1 U22195 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19122), .A(n19116), 
        .ZN(n19117) );
  OAI221_X1 U22196 ( .B1(n19118), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19118), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19117), .ZN(P2_U2822) );
  INV_X1 U22197 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19121) );
  OAI221_X1 U22198 ( .B1(n19122), .B2(n19121), .C1(n19120), .C2(n19119), .A(
        n19118), .ZN(P2_U2823) );
  NAND2_X1 U22199 ( .A1(n19123), .A2(n19125), .ZN(n19137) );
  AOI211_X1 U22200 ( .C1(n19257), .C2(n19125), .A(n19124), .B(n19289), .ZN(
        n19127) );
  OAI22_X1 U22201 ( .A1(n10783), .A2(n19180), .B1(n20070), .B2(n19262), .ZN(
        n19126) );
  AOI211_X1 U22202 ( .C1(n19323), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n19127), .B(n19126), .ZN(n19135) );
  INV_X1 U22203 ( .A(n19128), .ZN(n19131) );
  INV_X1 U22204 ( .A(n19129), .ZN(n19130) );
  OAI22_X1 U22205 ( .A1(n19131), .A2(n19320), .B1(n19130), .B2(n19302), .ZN(
        n19132) );
  AOI21_X1 U22206 ( .B1(n19133), .B2(n19305), .A(n19132), .ZN(n19134) );
  OAI211_X1 U22207 ( .C1(n19136), .C2(n19137), .A(n19135), .B(n19134), .ZN(
        P2_U2834) );
  INV_X1 U22208 ( .A(n19137), .ZN(n19138) );
  OAI21_X1 U22209 ( .B1(n19143), .B2(n19139), .A(n19138), .ZN(n19140) );
  INV_X1 U22210 ( .A(n19140), .ZN(n19141) );
  AOI21_X1 U22211 ( .B1(n19317), .B2(n19142), .A(n19141), .ZN(n19150) );
  NAND2_X1 U22212 ( .A1(n19311), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n19146) );
  OAI22_X1 U22213 ( .A1(n20068), .A2(n19262), .B1(n19143), .B2(n19310), .ZN(
        n19144) );
  AOI21_X1 U22214 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19323), .A(
        n19144), .ZN(n19145) );
  NAND2_X1 U22215 ( .A1(n19146), .A2(n19145), .ZN(n19147) );
  AOI21_X1 U22216 ( .B1(n19148), .B2(n19285), .A(n19147), .ZN(n19149) );
  OAI211_X1 U22217 ( .C1(n19151), .C2(n19315), .A(n19150), .B(n19149), .ZN(
        P2_U2835) );
  NAND2_X1 U22218 ( .A1(n19257), .A2(n19152), .ZN(n19153) );
  XOR2_X1 U22219 ( .A(n19154), .B(n19153), .Z(n19163) );
  AOI22_X1 U22220 ( .A1(n19311), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19323), .ZN(n19155) );
  OAI21_X1 U22221 ( .B1(n19156), .B2(n19302), .A(n19155), .ZN(n19157) );
  AOI211_X1 U22222 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19312), .A(n19420), 
        .B(n19157), .ZN(n19162) );
  OAI22_X1 U22223 ( .A1(n19159), .A2(n19320), .B1(n19158), .B2(n19315), .ZN(
        n19160) );
  INV_X1 U22224 ( .A(n19160), .ZN(n19161) );
  OAI211_X1 U22225 ( .C1(n19289), .C2(n19163), .A(n19162), .B(n19161), .ZN(
        P2_U2836) );
  OAI21_X1 U22226 ( .B1(n19164), .B2(n19180), .A(n19178), .ZN(n19167) );
  OAI22_X1 U22227 ( .A1(n19165), .A2(n19302), .B1(n20065), .B2(n19262), .ZN(
        n19166) );
  AOI211_X1 U22228 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19323), .A(
        n19167), .B(n19166), .ZN(n19173) );
  NOR2_X1 U22229 ( .A1(n19288), .A2(n19175), .ZN(n19169) );
  XNOR2_X1 U22230 ( .A(n19169), .B(n19168), .ZN(n19171) );
  AOI22_X1 U22231 ( .A1(n19171), .A2(n19306), .B1(n19170), .B2(n19285), .ZN(
        n19172) );
  OAI211_X1 U22232 ( .C1(n19174), .C2(n19315), .A(n19173), .B(n19172), .ZN(
        P2_U2837) );
  INV_X1 U22233 ( .A(n19176), .ZN(n19190) );
  AOI211_X1 U22234 ( .C1(n19177), .C2(n19176), .A(n19329), .B(n19175), .ZN(
        n19182) );
  AOI22_X1 U22235 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19323), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19312), .ZN(n19179) );
  OAI211_X1 U22236 ( .C1(n19180), .C2(n10752), .A(n19179), .B(n19178), .ZN(
        n19181) );
  AOI211_X1 U22237 ( .C1(n19183), .C2(n19317), .A(n19182), .B(n19181), .ZN(
        n19189) );
  OR2_X1 U22238 ( .A1(n19184), .A2(n19320), .ZN(n19187) );
  NAND2_X1 U22239 ( .A1(n19185), .A2(n19305), .ZN(n19186) );
  AND2_X1 U22240 ( .A1(n19187), .A2(n19186), .ZN(n19188) );
  OAI211_X1 U22241 ( .C1(n19190), .C2(n19310), .A(n19189), .B(n19188), .ZN(
        P2_U2838) );
  OAI21_X1 U22242 ( .B1(n20062), .B2(n19262), .A(n19178), .ZN(n19194) );
  INV_X1 U22243 ( .A(n19191), .ZN(n19192) );
  OAI22_X1 U22244 ( .A1(n19192), .A2(n19302), .B1(n19297), .B2(n10035), .ZN(
        n19193) );
  AOI211_X1 U22245 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19311), .A(n19194), .B(
        n19193), .ZN(n19201) );
  NOR2_X1 U22246 ( .A1(n19288), .A2(n19195), .ZN(n19197) );
  XNOR2_X1 U22247 ( .A(n19197), .B(n19196), .ZN(n19199) );
  AOI22_X1 U22248 ( .A1(n19199), .A2(n19306), .B1(n19285), .B2(n19198), .ZN(
        n19200) );
  OAI211_X1 U22249 ( .C1(n19202), .C2(n19315), .A(n19201), .B(n19200), .ZN(
        P2_U2839) );
  AOI22_X1 U22250 ( .A1(n19311), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19323), .ZN(n19203) );
  OAI21_X1 U22251 ( .B1(n19204), .B2(n19302), .A(n19203), .ZN(n19205) );
  AOI211_X1 U22252 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19312), .A(n19420), 
        .B(n19205), .ZN(n19212) );
  NOR2_X1 U22253 ( .A1(n19288), .A2(n19206), .ZN(n19208) );
  XNOR2_X1 U22254 ( .A(n19208), .B(n19207), .ZN(n19210) );
  AOI22_X1 U22255 ( .A1(n19210), .A2(n19306), .B1(n19285), .B2(n19209), .ZN(
        n19211) );
  OAI211_X1 U22256 ( .C1(n19344), .C2(n19315), .A(n19212), .B(n19211), .ZN(
        P2_U2841) );
  NAND2_X1 U22257 ( .A1(n19257), .A2(n19213), .ZN(n19214) );
  XOR2_X1 U22258 ( .A(n19215), .B(n19214), .Z(n19223) );
  AOI22_X1 U22259 ( .A1(n19216), .A2(n19317), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19323), .ZN(n19217) );
  OAI211_X1 U22260 ( .C1(n11095), .C2(n19262), .A(n19217), .B(n19178), .ZN(
        n19218) );
  AOI21_X1 U22261 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n19311), .A(n19218), .ZN(
        n19222) );
  AOI22_X1 U22262 ( .A1(n19220), .A2(n19285), .B1(n19305), .B2(n19219), .ZN(
        n19221) );
  OAI211_X1 U22263 ( .C1(n19289), .C2(n19223), .A(n19222), .B(n19221), .ZN(
        P2_U2842) );
  AOI22_X1 U22264 ( .A1(n19311), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19323), .ZN(n19224) );
  OAI21_X1 U22265 ( .B1(n19225), .B2(n19302), .A(n19224), .ZN(n19226) );
  AOI211_X1 U22266 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19312), .A(n19420), 
        .B(n19226), .ZN(n19233) );
  NOR2_X1 U22267 ( .A1(n19288), .A2(n19227), .ZN(n19229) );
  XNOR2_X1 U22268 ( .A(n19229), .B(n19228), .ZN(n19231) );
  AOI22_X1 U22269 ( .A1(n19231), .A2(n19306), .B1(n19285), .B2(n19230), .ZN(
        n19232) );
  OAI211_X1 U22270 ( .C1(n19234), .C2(n19315), .A(n19233), .B(n19232), .ZN(
        P2_U2843) );
  AOI22_X1 U22271 ( .A1(n19311), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19323), .ZN(n19235) );
  OAI21_X1 U22272 ( .B1(n19236), .B2(n19302), .A(n19235), .ZN(n19237) );
  AOI211_X1 U22273 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19312), .A(n19420), 
        .B(n19237), .ZN(n19243) );
  NOR2_X1 U22274 ( .A1(n19288), .A2(n19238), .ZN(n19240) );
  XNOR2_X1 U22275 ( .A(n19240), .B(n19239), .ZN(n19241) );
  AOI22_X1 U22276 ( .A1(n19241), .A2(n19306), .B1(n19285), .B2(n9761), .ZN(
        n19242) );
  OAI211_X1 U22277 ( .C1(n19244), .C2(n19315), .A(n19243), .B(n19242), .ZN(
        P2_U2845) );
  AOI22_X1 U22278 ( .A1(n19245), .A2(n19317), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19323), .ZN(n19246) );
  OAI211_X1 U22279 ( .C1(n11030), .C2(n19262), .A(n19246), .B(n19178), .ZN(
        n19247) );
  AOI21_X1 U22280 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19311), .A(n19247), .ZN(
        n19254) );
  NOR2_X1 U22281 ( .A1(n19288), .A2(n19248), .ZN(n19250) );
  XNOR2_X1 U22282 ( .A(n19250), .B(n19249), .ZN(n19252) );
  AOI22_X1 U22283 ( .A1(n19252), .A2(n19306), .B1(n19285), .B2(n19251), .ZN(
        n19253) );
  OAI211_X1 U22284 ( .C1(n19315), .C2(n19255), .A(n19254), .B(n19253), .ZN(
        P2_U2847) );
  NAND2_X1 U22285 ( .A1(n19257), .A2(n19256), .ZN(n19259) );
  XOR2_X1 U22286 ( .A(n19259), .B(n19258), .Z(n19269) );
  AOI22_X1 U22287 ( .A1(n19260), .A2(n19317), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19311), .ZN(n19261) );
  OAI211_X1 U22288 ( .C1(n11012), .C2(n19262), .A(n19261), .B(n19178), .ZN(
        n19267) );
  INV_X1 U22289 ( .A(n19263), .ZN(n19265) );
  OAI22_X1 U22290 ( .A1(n19265), .A2(n19320), .B1(n19315), .B2(n19264), .ZN(
        n19266) );
  AOI211_X1 U22291 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19323), .A(
        n19267), .B(n19266), .ZN(n19268) );
  OAI21_X1 U22292 ( .B1(n19269), .B2(n19289), .A(n19268), .ZN(P2_U2848) );
  NOR2_X1 U22293 ( .A1(n19288), .A2(n19270), .ZN(n19272) );
  XOR2_X1 U22294 ( .A(n19272), .B(n19271), .Z(n19280) );
  AOI22_X1 U22295 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19323), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19312), .ZN(n19273) );
  OAI21_X1 U22296 ( .B1(n19274), .B2(n19302), .A(n19273), .ZN(n19275) );
  AOI211_X1 U22297 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19311), .A(n19420), .B(
        n19275), .ZN(n19279) );
  OAI22_X1 U22298 ( .A1(n19276), .A2(n19320), .B1(n19315), .B2(n19350), .ZN(
        n19277) );
  INV_X1 U22299 ( .A(n19277), .ZN(n19278) );
  OAI211_X1 U22300 ( .C1(n19289), .C2(n19280), .A(n19279), .B(n19278), .ZN(
        P2_U2849) );
  AOI22_X1 U22301 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19323), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19312), .ZN(n19296) );
  INV_X1 U22302 ( .A(n19281), .ZN(n19282) );
  OAI22_X1 U22303 ( .A1(n19302), .A2(n19283), .B1(n19315), .B2(n19282), .ZN(
        n19284) );
  AOI211_X1 U22304 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n19311), .A(n19420), .B(
        n19284), .ZN(n19295) );
  INV_X1 U22305 ( .A(n19357), .ZN(n19286) );
  AOI22_X1 U22306 ( .A1(n19286), .A2(n19327), .B1(n19285), .B2(n19427), .ZN(
        n19294) );
  INV_X1 U22307 ( .A(n19431), .ZN(n19292) );
  NOR2_X1 U22308 ( .A1(n19288), .A2(n19287), .ZN(n19291) );
  AOI21_X1 U22309 ( .B1(n19292), .B2(n19291), .A(n19289), .ZN(n19290) );
  OAI21_X1 U22310 ( .B1(n19292), .B2(n19291), .A(n19290), .ZN(n19293) );
  NAND4_X1 U22311 ( .A1(n19296), .A2(n19295), .A3(n19294), .A4(n19293), .ZN(
        P2_U2851) );
  NOR2_X1 U22312 ( .A1(n19297), .A2(n13261), .ZN(n19298) );
  AOI21_X1 U22313 ( .B1(n19311), .B2(P2_EBX_REG_1__SCAN_IN), .A(n19298), .ZN(
        n19300) );
  NAND2_X1 U22314 ( .A1(n19312), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19299) );
  OAI211_X1 U22315 ( .C1(n19302), .C2(n19301), .A(n19300), .B(n19299), .ZN(
        n19304) );
  NOR2_X1 U22316 ( .A1(n13277), .A2(n19320), .ZN(n19303) );
  AOI211_X1 U22317 ( .C1(n19305), .C2(n20123), .A(n19304), .B(n19303), .ZN(
        n19309) );
  AOI22_X1 U22318 ( .A1(n19307), .A2(n19306), .B1(n19327), .B2(n20121), .ZN(
        n19308) );
  OAI211_X1 U22319 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19310), .A(
        n19309), .B(n19308), .ZN(P2_U2854) );
  AOI22_X1 U22320 ( .A1(n19312), .A2(P2_REIP_REG_0__SCAN_IN), .B1(
        P2_EBX_REG_0__SCAN_IN), .B2(n19311), .ZN(n19313) );
  OAI21_X1 U22321 ( .B1(n19315), .B2(n19314), .A(n19313), .ZN(n19316) );
  AOI21_X1 U22322 ( .B1(n19318), .B2(n19317), .A(n19316), .ZN(n19319) );
  OAI21_X1 U22323 ( .B1(n19321), .B2(n19320), .A(n19319), .ZN(n19326) );
  OAI21_X1 U22324 ( .B1(n19323), .B2(n19322), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19324) );
  INV_X1 U22325 ( .A(n19324), .ZN(n19325) );
  AOI211_X1 U22326 ( .C1(n19327), .C2(n19713), .A(n19326), .B(n19325), .ZN(
        n19328) );
  OAI21_X1 U22327 ( .B1(n19330), .B2(n19329), .A(n19328), .ZN(P2_U2855) );
  AOI22_X1 U22328 ( .A1(n19332), .A2(n19380), .B1(n19331), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19335) );
  AOI22_X1 U22329 ( .A1(n19333), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19379), .ZN(n19334) );
  NAND2_X1 U22330 ( .A1(n19335), .A2(n19334), .ZN(P2_U2888) );
  OAI22_X1 U22331 ( .A1(n19351), .A2(n19337), .B1(n19349), .B2(n19336), .ZN(
        n19338) );
  INV_X1 U22332 ( .A(n19338), .ZN(n19339) );
  OAI21_X1 U22333 ( .B1(n19386), .B2(n19340), .A(n19339), .ZN(P2_U2904) );
  AOI22_X1 U22334 ( .A1(n19342), .A2(n19341), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19379), .ZN(n19343) );
  OAI21_X1 U22335 ( .B1(n19351), .B2(n19344), .A(n19343), .ZN(P2_U2905) );
  INV_X1 U22336 ( .A(n19351), .ZN(n19355) );
  AOI22_X1 U22337 ( .A1(n19355), .A2(n19345), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n19379), .ZN(n19346) );
  OAI21_X1 U22338 ( .B1(n19347), .B2(n19386), .A(n19346), .ZN(P2_U2908) );
  OAI22_X1 U22339 ( .A1(n19351), .A2(n19350), .B1(n19349), .B2(n19348), .ZN(
        n19352) );
  INV_X1 U22340 ( .A(n19352), .ZN(n19353) );
  OAI21_X1 U22341 ( .B1(n19489), .B2(n19386), .A(n19353), .ZN(P2_U2913) );
  AOI22_X1 U22342 ( .A1(n19355), .A2(n19354), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19379), .ZN(n19360) );
  OR3_X1 U22343 ( .A1(n19358), .A2(n19357), .A3(n19356), .ZN(n19359) );
  OAI211_X1 U22344 ( .C1(n19486), .C2(n19386), .A(n19360), .B(n19359), .ZN(
        P2_U2914) );
  AOI22_X1 U22345 ( .A1(n19380), .A2(n19361), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19379), .ZN(n19367) );
  OAI21_X1 U22346 ( .B1(n19364), .B2(n19363), .A(n19362), .ZN(n19365) );
  NAND2_X1 U22347 ( .A1(n19365), .A2(n19381), .ZN(n19366) );
  OAI211_X1 U22348 ( .C1(n19475), .C2(n19386), .A(n19367), .B(n19366), .ZN(
        P2_U2916) );
  AOI22_X1 U22349 ( .A1(n19380), .A2(n20110), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19379), .ZN(n19373) );
  OAI21_X1 U22350 ( .B1(n19370), .B2(n19369), .A(n19368), .ZN(n19371) );
  NAND2_X1 U22351 ( .A1(n19371), .A2(n19381), .ZN(n19372) );
  OAI211_X1 U22352 ( .C1(n19471), .C2(n19386), .A(n19373), .B(n19372), .ZN(
        P2_U2917) );
  AOI22_X1 U22353 ( .A1(n19380), .A2(n20123), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19379), .ZN(n19378) );
  OAI21_X1 U22354 ( .B1(n19375), .B2(n19382), .A(n19374), .ZN(n19376) );
  NAND2_X1 U22355 ( .A1(n19376), .A2(n19381), .ZN(n19377) );
  OAI211_X1 U22356 ( .C1(n19467), .C2(n19386), .A(n19378), .B(n19377), .ZN(
        P2_U2918) );
  AOI22_X1 U22357 ( .A1(n19380), .A2(n19383), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19379), .ZN(n19385) );
  OAI211_X1 U22358 ( .C1(n19713), .C2(n19383), .A(n19382), .B(n19381), .ZN(
        n19384) );
  OAI211_X1 U22359 ( .C1(n19459), .C2(n19386), .A(n19385), .B(n19384), .ZN(
        P2_U2919) );
  AND2_X1 U22360 ( .A1(n19387), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22361 ( .A1(n19417), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19389) );
  OAI21_X1 U22362 ( .B1(n19336), .B2(n19419), .A(n19389), .ZN(P2_U2936) );
  AOI22_X1 U22363 ( .A1(n20146), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19390) );
  OAI21_X1 U22364 ( .B1(n19391), .B2(n19419), .A(n19390), .ZN(P2_U2937) );
  AOI22_X1 U22365 ( .A1(n20146), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19392) );
  OAI21_X1 U22366 ( .B1(n19393), .B2(n19419), .A(n19392), .ZN(P2_U2938) );
  AOI22_X1 U22367 ( .A1(n20146), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19394) );
  OAI21_X1 U22368 ( .B1(n19395), .B2(n19419), .A(n19394), .ZN(P2_U2939) );
  AOI22_X1 U22369 ( .A1(n20146), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19396) );
  OAI21_X1 U22370 ( .B1(n13188), .B2(n19419), .A(n19396), .ZN(P2_U2940) );
  AOI22_X1 U22371 ( .A1(n20146), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19397) );
  OAI21_X1 U22372 ( .B1(n19398), .B2(n19419), .A(n19397), .ZN(P2_U2941) );
  AOI22_X1 U22373 ( .A1(n20146), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19399) );
  OAI21_X1 U22374 ( .B1(n19400), .B2(n19419), .A(n19399), .ZN(P2_U2942) );
  AOI22_X1 U22375 ( .A1(n20146), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19401) );
  OAI21_X1 U22376 ( .B1(n19402), .B2(n19419), .A(n19401), .ZN(P2_U2943) );
  AOI22_X1 U22377 ( .A1(n19417), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19403) );
  OAI21_X1 U22378 ( .B1(n19404), .B2(n19419), .A(n19403), .ZN(P2_U2944) );
  AOI22_X1 U22379 ( .A1(n19417), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19405) );
  OAI21_X1 U22380 ( .B1(n19348), .B2(n19419), .A(n19405), .ZN(P2_U2945) );
  INV_X1 U22381 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19407) );
  AOI22_X1 U22382 ( .A1(n19417), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19406) );
  OAI21_X1 U22383 ( .B1(n19407), .B2(n19419), .A(n19406), .ZN(P2_U2946) );
  INV_X1 U22384 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19409) );
  AOI22_X1 U22385 ( .A1(n19417), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19408) );
  OAI21_X1 U22386 ( .B1(n19409), .B2(n19419), .A(n19408), .ZN(P2_U2947) );
  INV_X1 U22387 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19411) );
  AOI22_X1 U22388 ( .A1(n19417), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19410) );
  OAI21_X1 U22389 ( .B1(n19411), .B2(n19419), .A(n19410), .ZN(P2_U2948) );
  INV_X1 U22390 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19413) );
  AOI22_X1 U22391 ( .A1(n19417), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19412) );
  OAI21_X1 U22392 ( .B1(n19413), .B2(n19419), .A(n19412), .ZN(P2_U2949) );
  INV_X1 U22393 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19415) );
  AOI22_X1 U22394 ( .A1(n19417), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19414) );
  OAI21_X1 U22395 ( .B1(n19415), .B2(n19419), .A(n19414), .ZN(P2_U2950) );
  AOI22_X1 U22396 ( .A1(n19417), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19416), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19418) );
  OAI21_X1 U22397 ( .B1(n13182), .B2(n19419), .A(n19418), .ZN(P2_U2951) );
  AOI22_X1 U22398 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19421), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19420), .ZN(n19430) );
  OAI22_X1 U22399 ( .A1(n19425), .A2(n19424), .B1(n19423), .B2(n19422), .ZN(
        n19426) );
  AOI21_X1 U22400 ( .B1(n19428), .B2(n19427), .A(n19426), .ZN(n19429) );
  OAI211_X1 U22401 ( .C1(n19432), .C2(n19431), .A(n19430), .B(n19429), .ZN(
        P2_U3010) );
  OAI211_X1 U22402 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19434), .B(n19433), .ZN(n19446) );
  INV_X1 U22403 ( .A(n19435), .ZN(n19437) );
  AOI22_X1 U22404 ( .A1(n19438), .A2(n19437), .B1(n19436), .B2(n20123), .ZN(
        n19445) );
  NAND2_X1 U22405 ( .A1(n19440), .A2(n19439), .ZN(n19444) );
  OR2_X1 U22406 ( .A1(n19442), .A2(n19441), .ZN(n19443) );
  AND4_X1 U22407 ( .A1(n19446), .A2(n19445), .A3(n19444), .A4(n19443), .ZN(
        n19448) );
  OAI211_X1 U22408 ( .C1(n19450), .C2(n19449), .A(n19448), .B(n19447), .ZN(
        P2_U3045) );
  AOI22_X1 U22409 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19492), .ZN(n19933) );
  NAND2_X1 U22410 ( .A1(n19895), .A2(n19920), .ZN(n20026) );
  AOI22_X1 U22411 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19492), .ZN(n19898) );
  NOR2_X2 U22412 ( .A1(n20152), .A2(n19498), .ZN(n19971) );
  NOR3_X2 U22413 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19535), .ZN(n19500) );
  AOI22_X1 U22414 ( .A1(n20005), .A2(n19974), .B1(n19971), .B2(n19500), .ZN(
        n19466) );
  AOI21_X1 U22415 ( .B1(n19454), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19458) );
  AOI21_X1 U22416 ( .B1(n20026), .B2(n19530), .A(n20098), .ZN(n19455) );
  NOR2_X1 U22417 ( .A1(n19455), .A2(n19969), .ZN(n19460) );
  NOR2_X1 U22418 ( .A1(n19456), .A2(n20109), .ZN(n20017) );
  NOR2_X1 U22419 ( .A1(n20017), .A2(n19500), .ZN(n19463) );
  NAND2_X1 U22420 ( .A1(n19460), .A2(n19463), .ZN(n19457) );
  OAI211_X1 U22421 ( .C1(n19500), .C2(n19458), .A(n19457), .B(n19964), .ZN(
        n19503) );
  NOR2_X2 U22422 ( .A1(n19459), .A2(n19889), .ZN(n19972) );
  INV_X1 U22423 ( .A(n19460), .ZN(n19464) );
  OAI21_X1 U22424 ( .B1(n19461), .B2(n19500), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19462) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19503), .B1(
        n19972), .B2(n19502), .ZN(n19465) );
  OAI211_X1 U22426 ( .C1(n19933), .C2(n19530), .A(n19466), .B(n19465), .ZN(
        P2_U3048) );
  AOI22_X1 U22427 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19492), .ZN(n19937) );
  AOI22_X1 U22428 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19492), .ZN(n19983) );
  INV_X1 U22429 ( .A(n19983), .ZN(n19934) );
  NOR2_X2 U22430 ( .A1(n10458), .A2(n19498), .ZN(n19978) );
  AOI22_X1 U22431 ( .A1(n20005), .A2(n19934), .B1(n19978), .B2(n19500), .ZN(
        n19469) );
  NOR2_X2 U22432 ( .A1(n19467), .A2(n19889), .ZN(n19979) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19503), .B1(
        n19979), .B2(n19502), .ZN(n19468) );
  OAI211_X1 U22434 ( .C1(n19937), .C2(n19530), .A(n19469), .B(n19468), .ZN(
        P2_U3049) );
  AOI22_X1 U22435 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19492), .ZN(n19868) );
  AOI22_X1 U22436 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19492), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19493), .ZN(n19989) );
  NOR2_X2 U22437 ( .A1(n19470), .A2(n19498), .ZN(n19984) );
  AOI22_X1 U22438 ( .A1(n20005), .A2(n19865), .B1(n19500), .B2(n19984), .ZN(
        n19473) );
  NOR2_X2 U22439 ( .A1(n19471), .A2(n19889), .ZN(n19985) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19503), .B1(
        n19985), .B2(n19502), .ZN(n19472) );
  OAI211_X1 U22441 ( .C1(n19868), .C2(n19530), .A(n19473), .B(n19472), .ZN(
        P2_U3050) );
  AOI22_X1 U22442 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19492), .ZN(n19995) );
  AOI22_X1 U22443 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19492), .ZN(n19906) );
  NOR2_X2 U22444 ( .A1(n19474), .A2(n19498), .ZN(n19990) );
  AOI22_X1 U22445 ( .A1(n20005), .A2(n19992), .B1(n19990), .B2(n19500), .ZN(
        n19477) );
  NOR2_X2 U22446 ( .A1(n19475), .A2(n19889), .ZN(n19991) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19503), .B1(
        n19991), .B2(n19502), .ZN(n19476) );
  OAI211_X1 U22448 ( .C1(n19995), .C2(n19530), .A(n19477), .B(n19476), .ZN(
        P2_U3051) );
  AOI22_X1 U22449 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19492), .ZN(n19945) );
  OAI22_X2 U22450 ( .A1(n19479), .A2(n19496), .B1(n19478), .B2(n19494), .ZN(
        n19942) );
  NOR2_X2 U22451 ( .A1(n10321), .A2(n19498), .ZN(n19996) );
  AOI22_X1 U22452 ( .A1(n19942), .A2(n20005), .B1(n19996), .B2(n19500), .ZN(
        n19482) );
  NOR2_X2 U22453 ( .A1(n19480), .A2(n19889), .ZN(n19997) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19503), .B1(
        n19997), .B2(n19502), .ZN(n19481) );
  OAI211_X1 U22455 ( .C1(n19945), .C2(n19530), .A(n19482), .B(n19481), .ZN(
        P2_U3052) );
  INV_X1 U22456 ( .A(n20004), .ZN(n19875) );
  AOI22_X1 U22457 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19492), .ZN(n19948) );
  AOI22_X1 U22458 ( .A1(n20005), .A2(n20006), .B1(n19500), .B2(n19485), .ZN(
        n19488) );
  NOR2_X2 U22459 ( .A1(n19486), .A2(n19889), .ZN(n20003) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19503), .B1(
        n20003), .B2(n19502), .ZN(n19487) );
  OAI211_X1 U22461 ( .C1(n19875), .C2(n19530), .A(n19488), .B(n19487), .ZN(
        P2_U3053) );
  AOI22_X2 U22462 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19492), .ZN(n20016) );
  AOI22_X1 U22463 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19492), .ZN(n19914) );
  NOR2_X2 U22464 ( .A1(n13269), .A2(n19498), .ZN(n20011) );
  AOI22_X1 U22465 ( .A1(n20005), .A2(n20013), .B1(n20011), .B2(n19500), .ZN(
        n19491) );
  NOR2_X2 U22466 ( .A1(n19489), .A2(n19889), .ZN(n20012) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19503), .B1(
        n20012), .B2(n19502), .ZN(n19490) );
  OAI211_X1 U22468 ( .C1(n20016), .C2(n19530), .A(n19491), .B(n19490), .ZN(
        P2_U3054) );
  AOI22_X1 U22469 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19493), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19492), .ZN(n20027) );
  OAI22_X2 U22470 ( .A1(n19497), .A2(n19496), .B1(n19495), .B2(n19494), .ZN(
        n20021) );
  NOR2_X2 U22471 ( .A1(n19499), .A2(n19498), .ZN(n20018) );
  AOI22_X1 U22472 ( .A1(n20021), .A2(n20005), .B1(n20018), .B2(n19500), .ZN(
        n19505) );
  NOR2_X2 U22473 ( .A1(n19889), .A2(n19501), .ZN(n20019) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19503), .B1(
        n20019), .B2(n19502), .ZN(n19504) );
  OAI211_X1 U22475 ( .C1(n20027), .C2(n19530), .A(n19505), .B(n19504), .ZN(
        P2_U3055) );
  NOR2_X1 U22476 ( .A1(n19535), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19510) );
  INV_X1 U22477 ( .A(n19510), .ZN(n19506) );
  NOR2_X1 U22478 ( .A1(n19745), .A2(n19535), .ZN(n19525) );
  NOR3_X1 U22479 ( .A1(n10589), .A2(n19525), .A3(n19884), .ZN(n19507) );
  AOI211_X2 U22480 ( .C1(n19506), .C2(n19884), .A(n19686), .B(n19507), .ZN(
        n19526) );
  AOI22_X1 U22481 ( .A1(n19526), .A2(n19972), .B1(n19971), .B2(n19525), .ZN(
        n19512) );
  INV_X1 U22482 ( .A(n19525), .ZN(n19508) );
  AOI211_X1 U22483 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19508), .A(n19889), 
        .B(n19507), .ZN(n19509) );
  OAI221_X1 U22484 ( .B1(n19510), .B2(n19755), .C1(n19510), .C2(n19687), .A(
        n19509), .ZN(n19527) );
  INV_X1 U22485 ( .A(n19933), .ZN(n19973) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n19973), .ZN(n19511) );
  OAI211_X1 U22487 ( .C1(n19898), .C2(n19530), .A(n19512), .B(n19511), .ZN(
        P2_U3056) );
  AOI22_X1 U22488 ( .A1(n19526), .A2(n19979), .B1(n19978), .B2(n19525), .ZN(
        n19514) );
  INV_X1 U22489 ( .A(n19937), .ZN(n19980) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n19980), .ZN(n19513) );
  OAI211_X1 U22491 ( .C1(n19983), .C2(n19530), .A(n19514), .B(n19513), .ZN(
        P2_U3057) );
  AOI22_X1 U22492 ( .A1(n19526), .A2(n19985), .B1(n19984), .B2(n19525), .ZN(
        n19516) );
  INV_X1 U22493 ( .A(n19868), .ZN(n19986) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n19986), .ZN(n19515) );
  OAI211_X1 U22495 ( .C1(n19989), .C2(n19530), .A(n19516), .B(n19515), .ZN(
        P2_U3058) );
  AOI22_X1 U22496 ( .A1(n19526), .A2(n19991), .B1(n19990), .B2(n19525), .ZN(
        n19518) );
  INV_X1 U22497 ( .A(n19995), .ZN(n19903) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n19903), .ZN(n19517) );
  OAI211_X1 U22499 ( .C1(n19906), .C2(n19530), .A(n19518), .B(n19517), .ZN(
        P2_U3059) );
  INV_X1 U22500 ( .A(n19942), .ZN(n20002) );
  AOI22_X1 U22501 ( .A1(n19526), .A2(n19997), .B1(n19996), .B2(n19525), .ZN(
        n19520) );
  INV_X1 U22502 ( .A(n19945), .ZN(n19998) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n19998), .ZN(n19519) );
  OAI211_X1 U22504 ( .C1(n20002), .C2(n19530), .A(n19520), .B(n19519), .ZN(
        P2_U3060) );
  AOI22_X1 U22505 ( .A1(n19526), .A2(n20003), .B1(n19485), .B2(n19525), .ZN(
        n19522) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n20004), .ZN(n19521) );
  OAI211_X1 U22507 ( .C1(n19948), .C2(n19530), .A(n19522), .B(n19521), .ZN(
        P2_U3061) );
  AOI22_X1 U22508 ( .A1(n19526), .A2(n20012), .B1(n20011), .B2(n19525), .ZN(
        n19524) );
  INV_X1 U22509 ( .A(n20016), .ZN(n19911) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n19911), .ZN(n19523) );
  OAI211_X1 U22511 ( .C1(n19914), .C2(n19530), .A(n19524), .B(n19523), .ZN(
        P2_U3062) );
  AOI22_X1 U22512 ( .A1(n19526), .A2(n20019), .B1(n20018), .B2(n19525), .ZN(
        n19529) );
  INV_X1 U22513 ( .A(n20027), .ZN(n19953) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19527), .B1(
        n19554), .B2(n19953), .ZN(n19528) );
  OAI211_X1 U22515 ( .C1(n19959), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U3063) );
  INV_X1 U22516 ( .A(n19531), .ZN(n19785) );
  NOR2_X1 U22517 ( .A1(n19782), .A2(n19535), .ZN(n19552) );
  OAI21_X1 U22518 ( .B1(n19532), .B2(n19552), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19533) );
  OAI21_X1 U22519 ( .B1(n19535), .B2(n19785), .A(n19533), .ZN(n19553) );
  AOI22_X1 U22520 ( .A1(n19553), .A2(n19972), .B1(n19971), .B2(n19552), .ZN(
        n19539) );
  AOI21_X1 U22521 ( .B1(n10581), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19537) );
  INV_X1 U22522 ( .A(n19593), .ZN(n19663) );
  OAI21_X1 U22523 ( .B1(n19554), .B2(n19583), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19534) );
  OAI21_X1 U22524 ( .B1(n19663), .B2(n19535), .A(n19534), .ZN(n19536) );
  OAI211_X1 U22525 ( .C1(n19552), .C2(n19537), .A(n19536), .B(n19964), .ZN(
        n19555) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19974), .ZN(n19538) );
  OAI211_X1 U22527 ( .C1(n19933), .C2(n19591), .A(n19539), .B(n19538), .ZN(
        P2_U3064) );
  AOI22_X1 U22528 ( .A1(n19553), .A2(n19979), .B1(n19978), .B2(n19552), .ZN(
        n19541) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19934), .ZN(n19540) );
  OAI211_X1 U22530 ( .C1(n19937), .C2(n19591), .A(n19541), .B(n19540), .ZN(
        P2_U3065) );
  AOI22_X1 U22531 ( .A1(n19553), .A2(n19985), .B1(n19984), .B2(n19552), .ZN(
        n19543) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19865), .ZN(n19542) );
  OAI211_X1 U22533 ( .C1(n19868), .C2(n19591), .A(n19543), .B(n19542), .ZN(
        P2_U3066) );
  AOI22_X1 U22534 ( .A1(n19553), .A2(n19991), .B1(n19990), .B2(n19552), .ZN(
        n19545) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19992), .ZN(n19544) );
  OAI211_X1 U22536 ( .C1(n19995), .C2(n19591), .A(n19545), .B(n19544), .ZN(
        P2_U3067) );
  AOI22_X1 U22537 ( .A1(n19553), .A2(n19997), .B1(n19996), .B2(n19552), .ZN(
        n19547) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19942), .ZN(n19546) );
  OAI211_X1 U22539 ( .C1(n19945), .C2(n19591), .A(n19547), .B(n19546), .ZN(
        P2_U3068) );
  AOI22_X1 U22540 ( .A1(n19553), .A2(n20003), .B1(n19485), .B2(n19552), .ZN(
        n19549) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n20006), .ZN(n19548) );
  OAI211_X1 U22542 ( .C1(n19875), .C2(n19591), .A(n19549), .B(n19548), .ZN(
        P2_U3069) );
  AOI22_X1 U22543 ( .A1(n19553), .A2(n20012), .B1(n20011), .B2(n19552), .ZN(
        n19551) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n20013), .ZN(n19550) );
  OAI211_X1 U22545 ( .C1(n20016), .C2(n19591), .A(n19551), .B(n19550), .ZN(
        P2_U3070) );
  AOI22_X1 U22546 ( .A1(n19553), .A2(n20019), .B1(n20018), .B2(n19552), .ZN(
        n19557) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n20021), .ZN(n19556) );
  OAI211_X1 U22548 ( .C1(n20027), .C2(n19591), .A(n19557), .B(n19556), .ZN(
        P2_U3071) );
  NAND2_X1 U22549 ( .A1(n19687), .A2(n19822), .ZN(n19565) );
  NAND2_X1 U22550 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19558), .ZN(
        n19563) );
  NAND2_X1 U22551 ( .A1(n19565), .A2(n19563), .ZN(n19562) );
  OAI21_X1 U22552 ( .B1(n19566), .B2(n19884), .A(n19854), .ZN(n19560) );
  AND2_X1 U22553 ( .A1(n19812), .A2(n19558), .ZN(n19586) );
  INV_X1 U22554 ( .A(n19586), .ZN(n19559) );
  AOI21_X1 U22555 ( .B1(n19560), .B2(n19559), .A(n19889), .ZN(n19561) );
  INV_X1 U22556 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19571) );
  AOI22_X1 U22557 ( .A1(n19973), .A2(n19619), .B1(n19586), .B2(n19971), .ZN(
        n19570) );
  INV_X1 U22558 ( .A(n19563), .ZN(n19564) );
  NAND3_X1 U22559 ( .A1(n19565), .A2(n20107), .A3(n19564), .ZN(n19568) );
  OAI21_X1 U22560 ( .B1(n19566), .B2(n19586), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19567) );
  NAND2_X1 U22561 ( .A1(n19568), .A2(n19567), .ZN(n19587) );
  AOI22_X1 U22562 ( .A1(n19972), .A2(n19587), .B1(n19583), .B2(n19974), .ZN(
        n19569) );
  OAI211_X1 U22563 ( .C1(n19572), .C2(n19571), .A(n19570), .B(n19569), .ZN(
        P2_U3072) );
  AOI22_X1 U22564 ( .A1(n19980), .A2(n19619), .B1(n19586), .B2(n19978), .ZN(
        n19574) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19588), .B1(
        n19979), .B2(n19587), .ZN(n19573) );
  OAI211_X1 U22566 ( .C1(n19983), .C2(n19591), .A(n19574), .B(n19573), .ZN(
        P2_U3073) );
  AOI22_X1 U22567 ( .A1(n19865), .A2(n19583), .B1(n19586), .B2(n19984), .ZN(
        n19576) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19588), .B1(
        n19985), .B2(n19587), .ZN(n19575) );
  OAI211_X1 U22569 ( .C1(n19868), .C2(n19607), .A(n19576), .B(n19575), .ZN(
        P2_U3074) );
  AOI22_X1 U22570 ( .A1(n19903), .A2(n19619), .B1(n19586), .B2(n19990), .ZN(
        n19578) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19588), .B1(
        n19991), .B2(n19587), .ZN(n19577) );
  OAI211_X1 U22572 ( .C1(n19906), .C2(n19591), .A(n19578), .B(n19577), .ZN(
        P2_U3075) );
  AOI22_X1 U22573 ( .A1(n19942), .A2(n19583), .B1(n19586), .B2(n19996), .ZN(
        n19580) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19588), .B1(
        n19997), .B2(n19587), .ZN(n19579) );
  OAI211_X1 U22575 ( .C1(n19945), .C2(n19607), .A(n19580), .B(n19579), .ZN(
        P2_U3076) );
  AOI22_X1 U22576 ( .A1(n20006), .A2(n19583), .B1(n19586), .B2(n19485), .ZN(
        n19582) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19588), .B1(
        n20003), .B2(n19587), .ZN(n19581) );
  OAI211_X1 U22578 ( .C1(n19875), .C2(n19607), .A(n19582), .B(n19581), .ZN(
        P2_U3077) );
  AOI22_X1 U22579 ( .A1(n20013), .A2(n19583), .B1(n19586), .B2(n20011), .ZN(
        n19585) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19588), .B1(
        n20012), .B2(n19587), .ZN(n19584) );
  OAI211_X1 U22581 ( .C1(n20016), .C2(n19607), .A(n19585), .B(n19584), .ZN(
        P2_U3078) );
  AOI22_X1 U22582 ( .A1(n19953), .A2(n19619), .B1(n19586), .B2(n20018), .ZN(
        n19590) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19588), .B1(
        n20019), .B2(n19587), .ZN(n19589) );
  OAI211_X1 U22584 ( .C1(n19959), .C2(n19591), .A(n19590), .B(n19589), .ZN(
        P2_U3079) );
  INV_X1 U22585 ( .A(n19625), .ZN(n19662) );
  NOR3_X2 U22586 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19662), .ZN(n19618) );
  AOI22_X1 U22587 ( .A1(n19973), .A2(n19650), .B1(n19971), .B2(n19618), .ZN(
        n19604) );
  OAI21_X1 U22588 ( .B1(n19650), .B2(n19619), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19592) );
  NAND2_X1 U22589 ( .A1(n19592), .A2(n20107), .ZN(n19602) );
  OR2_X1 U22590 ( .A1(n19594), .A2(n19593), .ZN(n19853) );
  NOR2_X1 U22591 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19853), .ZN(
        n19598) );
  INV_X1 U22592 ( .A(n19599), .ZN(n19596) );
  INV_X1 U22593 ( .A(n19618), .ZN(n19595) );
  OAI211_X1 U22594 ( .C1(n19596), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19595), 
        .B(n19969), .ZN(n19597) );
  OAI211_X1 U22595 ( .C1(n19602), .C2(n19598), .A(n19964), .B(n19597), .ZN(
        n19621) );
  INV_X1 U22596 ( .A(n19598), .ZN(n19601) );
  OAI21_X1 U22597 ( .B1(n19599), .B2(n19618), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19600) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19621), .B1(
        n19972), .B2(n19620), .ZN(n19603) );
  OAI211_X1 U22599 ( .C1(n19898), .C2(n19607), .A(n19604), .B(n19603), .ZN(
        P2_U3080) );
  AOI22_X1 U22600 ( .A1(n19980), .A2(n19650), .B1(n19978), .B2(n19618), .ZN(
        n19606) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19621), .B1(
        n19979), .B2(n19620), .ZN(n19605) );
  OAI211_X1 U22602 ( .C1(n19983), .C2(n19607), .A(n19606), .B(n19605), .ZN(
        P2_U3081) );
  AOI22_X1 U22603 ( .A1(n19865), .A2(n19619), .B1(n19984), .B2(n19618), .ZN(
        n19609) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19621), .B1(
        n19985), .B2(n19620), .ZN(n19608) );
  OAI211_X1 U22605 ( .C1(n19868), .C2(n19638), .A(n19609), .B(n19608), .ZN(
        P2_U3082) );
  AOI22_X1 U22606 ( .A1(n19992), .A2(n19619), .B1(n19990), .B2(n19618), .ZN(
        n19611) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19621), .B1(
        n19991), .B2(n19620), .ZN(n19610) );
  OAI211_X1 U22608 ( .C1(n19995), .C2(n19638), .A(n19611), .B(n19610), .ZN(
        P2_U3083) );
  AOI22_X1 U22609 ( .A1(n19942), .A2(n19619), .B1(n19996), .B2(n19618), .ZN(
        n19613) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19621), .B1(
        n19997), .B2(n19620), .ZN(n19612) );
  OAI211_X1 U22611 ( .C1(n19945), .C2(n19638), .A(n19613), .B(n19612), .ZN(
        P2_U3084) );
  AOI22_X1 U22612 ( .A1(n20006), .A2(n19619), .B1(n19485), .B2(n19618), .ZN(
        n19615) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19621), .B1(
        n20003), .B2(n19620), .ZN(n19614) );
  OAI211_X1 U22614 ( .C1(n19875), .C2(n19638), .A(n19615), .B(n19614), .ZN(
        P2_U3085) );
  AOI22_X1 U22615 ( .A1(n19619), .A2(n20013), .B1(n20011), .B2(n19618), .ZN(
        n19617) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19621), .B1(
        n20012), .B2(n19620), .ZN(n19616) );
  OAI211_X1 U22617 ( .C1(n20016), .C2(n19638), .A(n19617), .B(n19616), .ZN(
        P2_U3086) );
  AOI22_X1 U22618 ( .A1(n20021), .A2(n19619), .B1(n20018), .B2(n19618), .ZN(
        n19623) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19621), .B1(
        n20019), .B2(n19620), .ZN(n19622) );
  OAI211_X1 U22620 ( .C1(n20027), .C2(n19638), .A(n19623), .B(n19622), .ZN(
        P2_U3087) );
  NOR2_X1 U22621 ( .A1(n19662), .A2(n19745), .ZN(n19649) );
  AOI22_X1 U22622 ( .A1(n19650), .A2(n19974), .B1(n19971), .B2(n19649), .ZN(
        n19635) );
  AOI21_X1 U22623 ( .B1(n19624), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19627) );
  NAND2_X1 U22624 ( .A1(n20125), .A2(n19625), .ZN(n19628) );
  NAND2_X1 U22625 ( .A1(n19687), .A2(n19894), .ZN(n19630) );
  NAND2_X1 U22626 ( .A1(n19628), .A2(n19630), .ZN(n19626) );
  OAI211_X1 U22627 ( .C1(n19649), .C2(n19627), .A(n19626), .B(n19964), .ZN(
        n19652) );
  INV_X1 U22628 ( .A(n19628), .ZN(n19629) );
  NAND3_X1 U22629 ( .A1(n19630), .A2(n20107), .A3(n19629), .ZN(n19633) );
  OAI21_X1 U22630 ( .B1(n19631), .B2(n19649), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19632) );
  NAND2_X1 U22631 ( .A1(n19633), .A2(n19632), .ZN(n19651) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19652), .B1(
        n19972), .B2(n19651), .ZN(n19634) );
  OAI211_X1 U22633 ( .C1(n19933), .C2(n19655), .A(n19635), .B(n19634), .ZN(
        P2_U3088) );
  AOI22_X1 U22634 ( .A1(n19980), .A2(n19682), .B1(n19978), .B2(n19649), .ZN(
        n19637) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19652), .B1(
        n19979), .B2(n19651), .ZN(n19636) );
  OAI211_X1 U22636 ( .C1(n19983), .C2(n19638), .A(n19637), .B(n19636), .ZN(
        P2_U3089) );
  AOI22_X1 U22637 ( .A1(n19865), .A2(n19650), .B1(n19984), .B2(n19649), .ZN(
        n19640) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19652), .B1(
        n19985), .B2(n19651), .ZN(n19639) );
  OAI211_X1 U22639 ( .C1(n19868), .C2(n19655), .A(n19640), .B(n19639), .ZN(
        P2_U3090) );
  AOI22_X1 U22640 ( .A1(n19650), .A2(n19992), .B1(n19990), .B2(n19649), .ZN(
        n19642) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19652), .B1(
        n19991), .B2(n19651), .ZN(n19641) );
  OAI211_X1 U22642 ( .C1(n19995), .C2(n19655), .A(n19642), .B(n19641), .ZN(
        P2_U3091) );
  AOI22_X1 U22643 ( .A1(n19942), .A2(n19650), .B1(n19996), .B2(n19649), .ZN(
        n19644) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19652), .B1(
        n19997), .B2(n19651), .ZN(n19643) );
  OAI211_X1 U22645 ( .C1(n19945), .C2(n19655), .A(n19644), .B(n19643), .ZN(
        P2_U3092) );
  AOI22_X1 U22646 ( .A1(n19650), .A2(n20006), .B1(n19485), .B2(n19649), .ZN(
        n19646) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19652), .B1(
        n20003), .B2(n19651), .ZN(n19645) );
  OAI211_X1 U22648 ( .C1(n19875), .C2(n19655), .A(n19646), .B(n19645), .ZN(
        P2_U3093) );
  AOI22_X1 U22649 ( .A1(n19650), .A2(n20013), .B1(n20011), .B2(n19649), .ZN(
        n19648) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19652), .B1(
        n20012), .B2(n19651), .ZN(n19647) );
  OAI211_X1 U22651 ( .C1(n20016), .C2(n19655), .A(n19648), .B(n19647), .ZN(
        P2_U3094) );
  AOI22_X1 U22652 ( .A1(n20021), .A2(n19650), .B1(n20018), .B2(n19649), .ZN(
        n19654) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19652), .B1(
        n20019), .B2(n19651), .ZN(n19653) );
  OAI211_X1 U22654 ( .C1(n20027), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U3095) );
  NOR2_X1 U22655 ( .A1(n19662), .A2(n19782), .ZN(n19680) );
  OAI21_X1 U22656 ( .B1(n10596), .B2(n19680), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19657) );
  OAI21_X1 U22657 ( .B1(n19785), .B2(n19662), .A(n19657), .ZN(n19681) );
  AOI22_X1 U22658 ( .A1(n19681), .A2(n19972), .B1(n19971), .B2(n19680), .ZN(
        n19667) );
  INV_X1 U22659 ( .A(n19680), .ZN(n19658) );
  OAI211_X1 U22660 ( .C1(n19659), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19658), 
        .B(n19969), .ZN(n19665) );
  INV_X1 U22661 ( .A(n19712), .ZN(n19660) );
  OAI21_X1 U22662 ( .B1(n19682), .B2(n19660), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19661) );
  OAI21_X1 U22663 ( .B1(n19663), .B2(n19662), .A(n19661), .ZN(n19664) );
  NAND3_X1 U22664 ( .A1(n19665), .A2(n19964), .A3(n19664), .ZN(n19683) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19974), .ZN(n19666) );
  OAI211_X1 U22666 ( .C1(n19933), .C2(n19712), .A(n19667), .B(n19666), .ZN(
        P2_U3096) );
  AOI22_X1 U22667 ( .A1(n19681), .A2(n19979), .B1(n19978), .B2(n19680), .ZN(
        n19669) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19934), .ZN(n19668) );
  OAI211_X1 U22669 ( .C1(n19937), .C2(n19712), .A(n19669), .B(n19668), .ZN(
        P2_U3097) );
  AOI22_X1 U22670 ( .A1(n19681), .A2(n19985), .B1(n19984), .B2(n19680), .ZN(
        n19671) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19865), .ZN(n19670) );
  OAI211_X1 U22672 ( .C1(n19868), .C2(n19712), .A(n19671), .B(n19670), .ZN(
        P2_U3098) );
  AOI22_X1 U22673 ( .A1(n19681), .A2(n19991), .B1(n19990), .B2(n19680), .ZN(
        n19673) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19992), .ZN(n19672) );
  OAI211_X1 U22675 ( .C1(n19995), .C2(n19712), .A(n19673), .B(n19672), .ZN(
        P2_U3099) );
  AOI22_X1 U22676 ( .A1(n19681), .A2(n19997), .B1(n19996), .B2(n19680), .ZN(
        n19675) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n19942), .ZN(n19674) );
  OAI211_X1 U22678 ( .C1(n19945), .C2(n19712), .A(n19675), .B(n19674), .ZN(
        P2_U3100) );
  AOI22_X1 U22679 ( .A1(n19681), .A2(n20003), .B1(n19485), .B2(n19680), .ZN(
        n19677) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n20006), .ZN(n19676) );
  OAI211_X1 U22681 ( .C1(n19875), .C2(n19712), .A(n19677), .B(n19676), .ZN(
        P2_U3101) );
  AOI22_X1 U22682 ( .A1(n19681), .A2(n20012), .B1(n20011), .B2(n19680), .ZN(
        n19679) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n20013), .ZN(n19678) );
  OAI211_X1 U22684 ( .C1(n20016), .C2(n19712), .A(n19679), .B(n19678), .ZN(
        P2_U3102) );
  AOI22_X1 U22685 ( .A1(n19681), .A2(n20019), .B1(n20018), .B2(n19680), .ZN(
        n19685) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19683), .B1(
        n19682), .B2(n20021), .ZN(n19684) );
  OAI211_X1 U22687 ( .C1(n20027), .C2(n19712), .A(n19685), .B(n19684), .ZN(
        P2_U3103) );
  NAND3_X1 U22688 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20109), .ZN(n19690) );
  NOR3_X1 U22689 ( .A1(n10591), .A2(n19719), .A3(n19884), .ZN(n19689) );
  AOI211_X2 U22690 ( .C1(n19690), .C2(n19884), .A(n19686), .B(n19689), .ZN(
        n19708) );
  AOI22_X1 U22691 ( .A1(n19708), .A2(n19972), .B1(n19719), .B2(n19971), .ZN(
        n19695) );
  INV_X1 U22692 ( .A(n19687), .ZN(n19688) );
  INV_X1 U22693 ( .A(n19920), .ZN(n19960) );
  NOR2_X1 U22694 ( .A1(n19688), .A2(n19960), .ZN(n20106) );
  INV_X1 U22695 ( .A(n20106), .ZN(n19691) );
  AOI211_X1 U22696 ( .C1(n19691), .C2(n19690), .A(n19889), .B(n19689), .ZN(
        n19692) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n19973), .ZN(n19694) );
  OAI211_X1 U22698 ( .C1(n19898), .C2(n19712), .A(n19695), .B(n19694), .ZN(
        P2_U3104) );
  AOI22_X1 U22699 ( .A1(n19708), .A2(n19979), .B1(n19719), .B2(n19978), .ZN(
        n19697) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n19980), .ZN(n19696) );
  OAI211_X1 U22701 ( .C1(n19983), .C2(n19712), .A(n19697), .B(n19696), .ZN(
        P2_U3105) );
  AOI22_X1 U22702 ( .A1(n19708), .A2(n19985), .B1(n19719), .B2(n19984), .ZN(
        n19699) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n19986), .ZN(n19698) );
  OAI211_X1 U22704 ( .C1(n19989), .C2(n19712), .A(n19699), .B(n19698), .ZN(
        P2_U3106) );
  AOI22_X1 U22705 ( .A1(n19708), .A2(n19991), .B1(n19719), .B2(n19990), .ZN(
        n19701) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n19903), .ZN(n19700) );
  OAI211_X1 U22707 ( .C1(n19906), .C2(n19712), .A(n19701), .B(n19700), .ZN(
        P2_U3107) );
  AOI22_X1 U22708 ( .A1(n19708), .A2(n19997), .B1(n19719), .B2(n19996), .ZN(
        n19703) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n19998), .ZN(n19702) );
  OAI211_X1 U22710 ( .C1(n20002), .C2(n19712), .A(n19703), .B(n19702), .ZN(
        P2_U3108) );
  AOI22_X1 U22711 ( .A1(n19708), .A2(n20003), .B1(n19719), .B2(n19485), .ZN(
        n19705) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n20004), .ZN(n19704) );
  OAI211_X1 U22713 ( .C1(n19948), .C2(n19712), .A(n19705), .B(n19704), .ZN(
        P2_U3109) );
  AOI22_X1 U22714 ( .A1(n19708), .A2(n20012), .B1(n19719), .B2(n20011), .ZN(
        n19707) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n19911), .ZN(n19706) );
  OAI211_X1 U22716 ( .C1(n19914), .C2(n19712), .A(n19707), .B(n19706), .ZN(
        P2_U3110) );
  AOI22_X1 U22717 ( .A1(n19708), .A2(n20019), .B1(n19719), .B2(n20018), .ZN(
        n19711) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19709), .B1(
        n19733), .B2(n19953), .ZN(n19710) );
  OAI211_X1 U22719 ( .C1(n19959), .C2(n19712), .A(n19711), .B(n19710), .ZN(
        P2_U3111) );
  NAND2_X1 U22720 ( .A1(n19921), .A2(n19755), .ZN(n19773) );
  NAND2_X1 U22721 ( .A1(n20116), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19786) );
  INV_X1 U22722 ( .A(n19786), .ZN(n19811) );
  NAND2_X1 U22723 ( .A1(n19811), .A2(n20125), .ZN(n19751) );
  NOR2_X1 U22724 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19751), .ZN(
        n19738) );
  AOI22_X1 U22725 ( .A1(n19733), .A2(n19974), .B1(n19738), .B2(n19971), .ZN(
        n19724) );
  AOI21_X1 U22726 ( .B1(n19773), .B2(n19743), .A(n20098), .ZN(n19714) );
  NOR2_X1 U22727 ( .A1(n19714), .A2(n19969), .ZN(n19718) );
  OAI21_X1 U22728 ( .B1(n19720), .B2(n19884), .A(n19854), .ZN(n19715) );
  AOI21_X1 U22729 ( .B1(n19718), .B2(n19716), .A(n19715), .ZN(n19717) );
  OAI21_X1 U22730 ( .B1(n19738), .B2(n19717), .A(n19964), .ZN(n19740) );
  OAI21_X1 U22731 ( .B1(n19719), .B2(n19738), .A(n19718), .ZN(n19722) );
  OAI21_X1 U22732 ( .B1(n19720), .B2(n19738), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19721) );
  NAND2_X1 U22733 ( .A1(n19722), .A2(n19721), .ZN(n19739) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19740), .B1(
        n19972), .B2(n19739), .ZN(n19723) );
  OAI211_X1 U22735 ( .C1(n19933), .C2(n19773), .A(n19724), .B(n19723), .ZN(
        P2_U3112) );
  AOI22_X1 U22736 ( .A1(n19934), .A2(n19733), .B1(n19738), .B2(n19978), .ZN(
        n19726) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19979), .ZN(n19725) );
  OAI211_X1 U22738 ( .C1(n19937), .C2(n19773), .A(n19726), .B(n19725), .ZN(
        P2_U3113) );
  AOI22_X1 U22739 ( .A1(n19865), .A2(n19733), .B1(n19738), .B2(n19984), .ZN(
        n19728) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19985), .ZN(n19727) );
  OAI211_X1 U22741 ( .C1(n19868), .C2(n19773), .A(n19728), .B(n19727), .ZN(
        P2_U3114) );
  AOI22_X1 U22742 ( .A1(n19903), .A2(n19776), .B1(n19738), .B2(n19990), .ZN(
        n19730) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19991), .ZN(n19729) );
  OAI211_X1 U22744 ( .C1(n19906), .C2(n19743), .A(n19730), .B(n19729), .ZN(
        P2_U3115) );
  AOI22_X1 U22745 ( .A1(n19998), .A2(n19776), .B1(n19738), .B2(n19996), .ZN(
        n19732) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19997), .ZN(n19731) );
  OAI211_X1 U22747 ( .C1(n20002), .C2(n19743), .A(n19732), .B(n19731), .ZN(
        P2_U3116) );
  AOI22_X1 U22748 ( .A1(n20006), .A2(n19733), .B1(n19738), .B2(n19485), .ZN(
        n19735) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n20003), .ZN(n19734) );
  OAI211_X1 U22750 ( .C1(n19875), .C2(n19773), .A(n19735), .B(n19734), .ZN(
        P2_U3117) );
  AOI22_X1 U22751 ( .A1(n19911), .A2(n19776), .B1(n19738), .B2(n20011), .ZN(
        n19737) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n20012), .ZN(n19736) );
  OAI211_X1 U22753 ( .C1(n19914), .C2(n19743), .A(n19737), .B(n19736), .ZN(
        P2_U3118) );
  AOI22_X1 U22754 ( .A1(n19776), .A2(n19953), .B1(n19738), .B2(n20018), .ZN(
        n19742) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n20019), .ZN(n19741) );
  OAI211_X1 U22756 ( .C1(n19959), .C2(n19743), .A(n19742), .B(n19741), .ZN(
        P2_U3119) );
  OR2_X1 U22757 ( .A1(n20103), .A2(n20098), .ZN(n19961) );
  INV_X1 U22758 ( .A(n19961), .ZN(n19892) );
  NAND2_X1 U22759 ( .A1(n19892), .A2(n19755), .ZN(n19744) );
  NAND2_X1 U22760 ( .A1(n19744), .A2(n19751), .ZN(n19749) );
  NAND2_X1 U22761 ( .A1(n10588), .A2(n19854), .ZN(n19747) );
  NOR2_X1 U22762 ( .A1(n19745), .A2(n19786), .ZN(n19787) );
  INV_X1 U22763 ( .A(n19787), .ZN(n19746) );
  NAND2_X1 U22764 ( .A1(n19747), .A2(n19746), .ZN(n19748) );
  MUX2_X1 U22765 ( .A(n19749), .B(n19748), .S(n19969), .Z(n19750) );
  NAND2_X1 U22766 ( .A1(n19750), .A2(n19964), .ZN(n19778) );
  INV_X1 U22767 ( .A(n19778), .ZN(n19764) );
  INV_X1 U22768 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U22769 ( .A1(n19776), .A2(n19974), .B1(n19971), .B2(n19787), .ZN(
        n19759) );
  INV_X1 U22770 ( .A(n19751), .ZN(n19752) );
  NAND2_X1 U22771 ( .A1(n19752), .A2(n20107), .ZN(n19754) );
  OAI21_X1 U22772 ( .B1(n10588), .B2(n19787), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19753) );
  NAND2_X1 U22773 ( .A1(n19754), .A2(n19753), .ZN(n19777) );
  INV_X1 U22774 ( .A(n19755), .ZN(n19756) );
  AOI22_X1 U22775 ( .A1(n19972), .A2(n19777), .B1(n19807), .B2(n19973), .ZN(
        n19758) );
  OAI211_X1 U22776 ( .C1(n19764), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P2_U3120) );
  INV_X1 U22777 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U22778 ( .A1(n19776), .A2(n19934), .B1(n19787), .B2(n19978), .ZN(
        n19762) );
  AOI22_X1 U22779 ( .A1(n19979), .A2(n19777), .B1(n19807), .B2(n19980), .ZN(
        n19761) );
  OAI211_X1 U22780 ( .C1(n19764), .C2(n19763), .A(n19762), .B(n19761), .ZN(
        P2_U3121) );
  AOI22_X1 U22781 ( .A1(n19986), .A2(n19807), .B1(n19787), .B2(n19984), .ZN(
        n19766) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19778), .B1(
        n19985), .B2(n19777), .ZN(n19765) );
  OAI211_X1 U22783 ( .C1(n19989), .C2(n19773), .A(n19766), .B(n19765), .ZN(
        P2_U3122) );
  INV_X1 U22784 ( .A(n19807), .ZN(n19781) );
  AOI22_X1 U22785 ( .A1(n19776), .A2(n19992), .B1(n19990), .B2(n19787), .ZN(
        n19768) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19778), .B1(
        n19991), .B2(n19777), .ZN(n19767) );
  OAI211_X1 U22787 ( .C1(n19995), .C2(n19781), .A(n19768), .B(n19767), .ZN(
        P2_U3123) );
  AOI22_X1 U22788 ( .A1(n19942), .A2(n19776), .B1(n19996), .B2(n19787), .ZN(
        n19770) );
  AOI22_X1 U22789 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19778), .B1(
        n19997), .B2(n19777), .ZN(n19769) );
  OAI211_X1 U22790 ( .C1(n19945), .C2(n19781), .A(n19770), .B(n19769), .ZN(
        P2_U3124) );
  AOI22_X1 U22791 ( .A1(n20004), .A2(n19807), .B1(n19787), .B2(n19485), .ZN(
        n19772) );
  AOI22_X1 U22792 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19778), .B1(
        n20003), .B2(n19777), .ZN(n19771) );
  OAI211_X1 U22793 ( .C1(n19948), .C2(n19773), .A(n19772), .B(n19771), .ZN(
        P2_U3125) );
  AOI22_X1 U22794 ( .A1(n19776), .A2(n20013), .B1(n20011), .B2(n19787), .ZN(
        n19775) );
  AOI22_X1 U22795 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19778), .B1(
        n20012), .B2(n19777), .ZN(n19774) );
  OAI211_X1 U22796 ( .C1(n20016), .C2(n19781), .A(n19775), .B(n19774), .ZN(
        P2_U3126) );
  AOI22_X1 U22797 ( .A1(n20021), .A2(n19776), .B1(n20018), .B2(n19787), .ZN(
        n19780) );
  AOI22_X1 U22798 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19778), .B1(
        n20019), .B2(n19777), .ZN(n19779) );
  OAI211_X1 U22799 ( .C1(n20027), .C2(n19781), .A(n19780), .B(n19779), .ZN(
        P2_U3127) );
  NOR2_X1 U22800 ( .A1(n19782), .A2(n19786), .ZN(n19805) );
  OAI21_X1 U22801 ( .B1(n19783), .B2(n19805), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19784) );
  OAI21_X1 U22802 ( .B1(n19786), .B2(n19785), .A(n19784), .ZN(n19806) );
  AOI22_X1 U22803 ( .A1(n19806), .A2(n19972), .B1(n19971), .B2(n19805), .ZN(
        n19792) );
  AOI221_X1 U22804 ( .B1(n19844), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19807), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19787), .ZN(n19788) );
  AOI211_X1 U22805 ( .C1(n19789), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19788), .ZN(n19790) );
  OAI21_X1 U22806 ( .B1(n19790), .B2(n19805), .A(n19964), .ZN(n19808) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n19974), .ZN(n19791) );
  OAI211_X1 U22808 ( .C1(n19933), .C2(n19835), .A(n19792), .B(n19791), .ZN(
        P2_U3128) );
  AOI22_X1 U22809 ( .A1(n19806), .A2(n19979), .B1(n19978), .B2(n19805), .ZN(
        n19794) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n19934), .ZN(n19793) );
  OAI211_X1 U22811 ( .C1(n19937), .C2(n19835), .A(n19794), .B(n19793), .ZN(
        P2_U3129) );
  AOI22_X1 U22812 ( .A1(n19806), .A2(n19985), .B1(n19984), .B2(n19805), .ZN(
        n19796) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n19865), .ZN(n19795) );
  OAI211_X1 U22814 ( .C1(n19868), .C2(n19835), .A(n19796), .B(n19795), .ZN(
        P2_U3130) );
  AOI22_X1 U22815 ( .A1(n19806), .A2(n19991), .B1(n19990), .B2(n19805), .ZN(
        n19798) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n19992), .ZN(n19797) );
  OAI211_X1 U22817 ( .C1(n19995), .C2(n19835), .A(n19798), .B(n19797), .ZN(
        P2_U3131) );
  AOI22_X1 U22818 ( .A1(n19806), .A2(n19997), .B1(n19996), .B2(n19805), .ZN(
        n19800) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n19942), .ZN(n19799) );
  OAI211_X1 U22820 ( .C1(n19945), .C2(n19835), .A(n19800), .B(n19799), .ZN(
        P2_U3132) );
  AOI22_X1 U22821 ( .A1(n19806), .A2(n20003), .B1(n19485), .B2(n19805), .ZN(
        n19802) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n20006), .ZN(n19801) );
  OAI211_X1 U22823 ( .C1(n19875), .C2(n19835), .A(n19802), .B(n19801), .ZN(
        P2_U3133) );
  AOI22_X1 U22824 ( .A1(n19806), .A2(n20012), .B1(n20011), .B2(n19805), .ZN(
        n19804) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n20013), .ZN(n19803) );
  OAI211_X1 U22826 ( .C1(n20016), .C2(n19835), .A(n19804), .B(n19803), .ZN(
        P2_U3134) );
  AOI22_X1 U22827 ( .A1(n19806), .A2(n20019), .B1(n20018), .B2(n19805), .ZN(
        n19810) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19808), .B1(
        n19807), .B2(n20021), .ZN(n19809) );
  OAI211_X1 U22829 ( .C1(n20027), .C2(n19835), .A(n19810), .B(n19809), .ZN(
        P2_U3135) );
  INV_X1 U22830 ( .A(n19822), .ZN(n20097) );
  NAND2_X1 U22831 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19811), .ZN(
        n19819) );
  OAI21_X1 U22832 ( .B1(n19961), .B2(n20097), .A(n19819), .ZN(n19818) );
  NAND2_X1 U22833 ( .A1(n19812), .A2(n19811), .ZN(n19813) );
  INV_X1 U22834 ( .A(n19813), .ZN(n19842) );
  AND2_X1 U22835 ( .A1(n19813), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19814) );
  NAND2_X1 U22836 ( .A1(n19815), .A2(n19814), .ZN(n19821) );
  OAI211_X1 U22837 ( .C1(n19842), .C2(n19854), .A(n19821), .B(n19964), .ZN(
        n19816) );
  INV_X1 U22838 ( .A(n19816), .ZN(n19817) );
  INV_X1 U22839 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n19825) );
  OAI21_X1 U22840 ( .B1(n19819), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19884), 
        .ZN(n19820) );
  AND2_X1 U22841 ( .A1(n19821), .A2(n19820), .ZN(n19843) );
  AOI22_X1 U22842 ( .A1(n19843), .A2(n19972), .B1(n19971), .B2(n19842), .ZN(
        n19824) );
  NAND2_X1 U22843 ( .A1(n19895), .A2(n19822), .ZN(n19852) );
  AOI22_X1 U22844 ( .A1(n19844), .A2(n19974), .B1(n19880), .B2(n19973), .ZN(
        n19823) );
  OAI211_X1 U22845 ( .C1(n19848), .C2(n19825), .A(n19824), .B(n19823), .ZN(
        P2_U3136) );
  AOI22_X1 U22846 ( .A1(n19843), .A2(n19979), .B1(n19978), .B2(n19842), .ZN(
        n19827) );
  INV_X1 U22847 ( .A(n19848), .ZN(n19839) );
  AOI22_X1 U22848 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19839), .B1(
        n19880), .B2(n19980), .ZN(n19826) );
  OAI211_X1 U22849 ( .C1(n19983), .C2(n19835), .A(n19827), .B(n19826), .ZN(
        P2_U3137) );
  AOI22_X1 U22850 ( .A1(n19843), .A2(n19985), .B1(n19984), .B2(n19842), .ZN(
        n19829) );
  AOI22_X1 U22851 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19839), .B1(
        n19844), .B2(n19865), .ZN(n19828) );
  OAI211_X1 U22852 ( .C1(n19868), .C2(n19852), .A(n19829), .B(n19828), .ZN(
        P2_U3138) );
  AOI22_X1 U22853 ( .A1(n19843), .A2(n19991), .B1(n19990), .B2(n19842), .ZN(
        n19831) );
  AOI22_X1 U22854 ( .A1(n19880), .A2(n19903), .B1(n19844), .B2(n19992), .ZN(
        n19830) );
  OAI211_X1 U22855 ( .C1(n19848), .C2(n19832), .A(n19831), .B(n19830), .ZN(
        P2_U3139) );
  AOI22_X1 U22856 ( .A1(n19843), .A2(n19997), .B1(n19996), .B2(n19842), .ZN(
        n19834) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19839), .B1(
        n19880), .B2(n19998), .ZN(n19833) );
  OAI211_X1 U22858 ( .C1(n20002), .C2(n19835), .A(n19834), .B(n19833), .ZN(
        P2_U3140) );
  INV_X1 U22859 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n19838) );
  AOI22_X1 U22860 ( .A1(n19843), .A2(n20003), .B1(n19485), .B2(n19842), .ZN(
        n19837) );
  AOI22_X1 U22861 ( .A1(n19844), .A2(n20006), .B1(n19880), .B2(n20004), .ZN(
        n19836) );
  OAI211_X1 U22862 ( .C1(n19848), .C2(n19838), .A(n19837), .B(n19836), .ZN(
        P2_U3141) );
  AOI22_X1 U22863 ( .A1(n19843), .A2(n20012), .B1(n20011), .B2(n19842), .ZN(
        n19841) );
  AOI22_X1 U22864 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19839), .B1(
        n19844), .B2(n20013), .ZN(n19840) );
  OAI211_X1 U22865 ( .C1(n20016), .C2(n19852), .A(n19841), .B(n19840), .ZN(
        P2_U3142) );
  AOI22_X1 U22866 ( .A1(n19843), .A2(n20019), .B1(n20018), .B2(n19842), .ZN(
        n19846) );
  AOI22_X1 U22867 ( .A1(n19880), .A2(n19953), .B1(n19844), .B2(n20021), .ZN(
        n19845) );
  OAI211_X1 U22868 ( .C1(n19848), .C2(n19847), .A(n19846), .B(n19845), .ZN(
        P2_U3143) );
  INV_X1 U22869 ( .A(n19849), .ZN(n19851) );
  NAND3_X1 U22870 ( .A1(n20125), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19886) );
  NOR2_X1 U22871 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19886), .ZN(
        n19878) );
  OAI21_X1 U22872 ( .B1(n19855), .B2(n19878), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19850) );
  OAI21_X1 U22873 ( .B1(n19853), .B2(n19851), .A(n19850), .ZN(n19879) );
  AOI22_X1 U22874 ( .A1(n19879), .A2(n19972), .B1(n19971), .B2(n19878), .ZN(
        n19862) );
  AOI21_X1 U22875 ( .B1(n19852), .B2(n19919), .A(n20098), .ZN(n19860) );
  NOR2_X1 U22876 ( .A1(n20109), .A2(n19853), .ZN(n19859) );
  OAI21_X1 U22877 ( .B1(n19855), .B2(n19884), .A(n19854), .ZN(n19857) );
  INV_X1 U22878 ( .A(n19878), .ZN(n19856) );
  AOI21_X1 U22879 ( .B1(n19857), .B2(n19856), .A(n19889), .ZN(n19858) );
  AOI22_X1 U22880 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n19974), .ZN(n19861) );
  OAI211_X1 U22881 ( .C1(n19933), .C2(n19919), .A(n19862), .B(n19861), .ZN(
        P2_U3144) );
  AOI22_X1 U22882 ( .A1(n19879), .A2(n19979), .B1(n19978), .B2(n19878), .ZN(
        n19864) );
  AOI22_X1 U22883 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n19934), .ZN(n19863) );
  OAI211_X1 U22884 ( .C1(n19937), .C2(n19919), .A(n19864), .B(n19863), .ZN(
        P2_U3145) );
  AOI22_X1 U22885 ( .A1(n19879), .A2(n19985), .B1(n19984), .B2(n19878), .ZN(
        n19867) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n19865), .ZN(n19866) );
  OAI211_X1 U22887 ( .C1(n19868), .C2(n19919), .A(n19867), .B(n19866), .ZN(
        P2_U3146) );
  AOI22_X1 U22888 ( .A1(n19879), .A2(n19991), .B1(n19990), .B2(n19878), .ZN(
        n19870) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n19992), .ZN(n19869) );
  OAI211_X1 U22890 ( .C1(n19995), .C2(n19919), .A(n19870), .B(n19869), .ZN(
        P2_U3147) );
  AOI22_X1 U22891 ( .A1(n19879), .A2(n19997), .B1(n19996), .B2(n19878), .ZN(
        n19872) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n19942), .ZN(n19871) );
  OAI211_X1 U22893 ( .C1(n19945), .C2(n19919), .A(n19872), .B(n19871), .ZN(
        P2_U3148) );
  AOI22_X1 U22894 ( .A1(n19879), .A2(n20003), .B1(n19485), .B2(n19878), .ZN(
        n19874) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n20006), .ZN(n19873) );
  OAI211_X1 U22896 ( .C1(n19875), .C2(n19919), .A(n19874), .B(n19873), .ZN(
        P2_U3149) );
  AOI22_X1 U22897 ( .A1(n19879), .A2(n20012), .B1(n20011), .B2(n19878), .ZN(
        n19877) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n20013), .ZN(n19876) );
  OAI211_X1 U22899 ( .C1(n20016), .C2(n19919), .A(n19877), .B(n19876), .ZN(
        P2_U3150) );
  AOI22_X1 U22900 ( .A1(n19879), .A2(n20019), .B1(n20018), .B2(n19878), .ZN(
        n19883) );
  AOI22_X1 U22901 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19881), .B1(
        n19880), .B2(n20021), .ZN(n19882) );
  OAI211_X1 U22902 ( .C1(n20027), .C2(n19919), .A(n19883), .B(n19882), .ZN(
        P2_U3151) );
  NOR2_X1 U22903 ( .A1(n20135), .A2(n19886), .ZN(n19924) );
  NOR3_X1 U22904 ( .A1(n19885), .A2(n19924), .A3(n19884), .ZN(n19888) );
  INV_X1 U22905 ( .A(n19886), .ZN(n19893) );
  AOI21_X1 U22906 ( .B1(n19854), .B2(n19893), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19887) );
  NOR2_X1 U22907 ( .A1(n19888), .A2(n19887), .ZN(n19915) );
  AOI22_X1 U22908 ( .A1(n19915), .A2(n19972), .B1(n19971), .B2(n19924), .ZN(
        n19897) );
  INV_X1 U22909 ( .A(n19924), .ZN(n19890) );
  AOI211_X1 U22910 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19890), .A(n19889), 
        .B(n19888), .ZN(n19891) );
  OAI221_X1 U22911 ( .B1(n19893), .B2(n19894), .C1(n19893), .C2(n19892), .A(
        n19891), .ZN(n19916) );
  NAND2_X1 U22912 ( .A1(n19895), .A2(n19894), .ZN(n19958) );
  AOI22_X1 U22913 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n19973), .ZN(n19896) );
  OAI211_X1 U22914 ( .C1(n19898), .C2(n19919), .A(n19897), .B(n19896), .ZN(
        P2_U3152) );
  AOI22_X1 U22915 ( .A1(n19915), .A2(n19979), .B1(n19978), .B2(n19924), .ZN(
        n19900) );
  AOI22_X1 U22916 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n19980), .ZN(n19899) );
  OAI211_X1 U22917 ( .C1(n19983), .C2(n19919), .A(n19900), .B(n19899), .ZN(
        P2_U3153) );
  AOI22_X1 U22918 ( .A1(n19915), .A2(n19985), .B1(n19984), .B2(n19924), .ZN(
        n19902) );
  AOI22_X1 U22919 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n19986), .ZN(n19901) );
  OAI211_X1 U22920 ( .C1(n19989), .C2(n19919), .A(n19902), .B(n19901), .ZN(
        P2_U3154) );
  AOI22_X1 U22921 ( .A1(n19915), .A2(n19991), .B1(n19990), .B2(n19924), .ZN(
        n19905) );
  AOI22_X1 U22922 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n19903), .ZN(n19904) );
  OAI211_X1 U22923 ( .C1(n19906), .C2(n19919), .A(n19905), .B(n19904), .ZN(
        P2_U3155) );
  AOI22_X1 U22924 ( .A1(n19915), .A2(n19997), .B1(n19996), .B2(n19924), .ZN(
        n19908) );
  AOI22_X1 U22925 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n19998), .ZN(n19907) );
  OAI211_X1 U22926 ( .C1(n20002), .C2(n19919), .A(n19908), .B(n19907), .ZN(
        P2_U3156) );
  AOI22_X1 U22927 ( .A1(n19915), .A2(n20003), .B1(n19485), .B2(n19924), .ZN(
        n19910) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n20004), .ZN(n19909) );
  OAI211_X1 U22929 ( .C1(n19948), .C2(n19919), .A(n19910), .B(n19909), .ZN(
        P2_U3157) );
  AOI22_X1 U22930 ( .A1(n19915), .A2(n20012), .B1(n20011), .B2(n19924), .ZN(
        n19913) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n19911), .ZN(n19912) );
  OAI211_X1 U22932 ( .C1(n19914), .C2(n19919), .A(n19913), .B(n19912), .ZN(
        P2_U3158) );
  AOI22_X1 U22933 ( .A1(n19915), .A2(n20019), .B1(n20018), .B2(n19924), .ZN(
        n19918) );
  AOI22_X1 U22934 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19916), .B1(
        n19949), .B2(n19953), .ZN(n19917) );
  OAI211_X1 U22935 ( .C1(n19959), .C2(n19919), .A(n19918), .B(n19917), .ZN(
        P2_U3159) );
  NAND3_X1 U22936 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19970) );
  NOR2_X1 U22937 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19970), .ZN(
        n19952) );
  AOI22_X1 U22938 ( .A1(n19949), .A2(n19974), .B1(n19971), .B2(n19952), .ZN(
        n19932) );
  AOI21_X1 U22939 ( .B1(n19922), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19926) );
  AOI21_X1 U22940 ( .B1(n20001), .B2(n19958), .A(n20098), .ZN(n19923) );
  NOR2_X1 U22941 ( .A1(n19923), .A2(n19969), .ZN(n19927) );
  NOR2_X1 U22942 ( .A1(n19952), .A2(n19924), .ZN(n19929) );
  NAND2_X1 U22943 ( .A1(n19927), .A2(n19929), .ZN(n19925) );
  OAI211_X1 U22944 ( .C1(n19952), .C2(n19926), .A(n19925), .B(n19964), .ZN(
        n19955) );
  INV_X1 U22945 ( .A(n19927), .ZN(n19930) );
  OAI21_X1 U22946 ( .B1(n10590), .B2(n19952), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19928) );
  AOI22_X1 U22947 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19955), .B1(
        n19972), .B2(n19954), .ZN(n19931) );
  OAI211_X1 U22948 ( .C1(n19933), .C2(n20001), .A(n19932), .B(n19931), .ZN(
        P2_U3160) );
  AOI22_X1 U22949 ( .A1(n19949), .A2(n19934), .B1(n19978), .B2(n19952), .ZN(
        n19936) );
  AOI22_X1 U22950 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19955), .B1(
        n19979), .B2(n19954), .ZN(n19935) );
  OAI211_X1 U22951 ( .C1(n19937), .C2(n20001), .A(n19936), .B(n19935), .ZN(
        P2_U3161) );
  AOI22_X1 U22952 ( .A1(n19986), .A2(n20022), .B1(n19984), .B2(n19952), .ZN(
        n19939) );
  AOI22_X1 U22953 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19955), .B1(
        n19985), .B2(n19954), .ZN(n19938) );
  OAI211_X1 U22954 ( .C1(n19989), .C2(n19958), .A(n19939), .B(n19938), .ZN(
        P2_U3162) );
  AOI22_X1 U22955 ( .A1(n19949), .A2(n19992), .B1(n19990), .B2(n19952), .ZN(
        n19941) );
  AOI22_X1 U22956 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19955), .B1(
        n19991), .B2(n19954), .ZN(n19940) );
  OAI211_X1 U22957 ( .C1(n19995), .C2(n20001), .A(n19941), .B(n19940), .ZN(
        P2_U3163) );
  AOI22_X1 U22958 ( .A1(n19942), .A2(n19949), .B1(n19996), .B2(n19952), .ZN(
        n19944) );
  AOI22_X1 U22959 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19955), .B1(
        n19997), .B2(n19954), .ZN(n19943) );
  OAI211_X1 U22960 ( .C1(n19945), .C2(n20001), .A(n19944), .B(n19943), .ZN(
        P2_U3164) );
  AOI22_X1 U22961 ( .A1(n20004), .A2(n20022), .B1(n19485), .B2(n19952), .ZN(
        n19947) );
  AOI22_X1 U22962 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19955), .B1(
        n20003), .B2(n19954), .ZN(n19946) );
  OAI211_X1 U22963 ( .C1(n19948), .C2(n19958), .A(n19947), .B(n19946), .ZN(
        P2_U3165) );
  AOI22_X1 U22964 ( .A1(n19949), .A2(n20013), .B1(n20011), .B2(n19952), .ZN(
        n19951) );
  AOI22_X1 U22965 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19955), .B1(
        n20012), .B2(n19954), .ZN(n19950) );
  OAI211_X1 U22966 ( .C1(n20016), .C2(n20001), .A(n19951), .B(n19950), .ZN(
        P2_U3166) );
  AOI22_X1 U22967 ( .A1(n20022), .A2(n19953), .B1(n20018), .B2(n19952), .ZN(
        n19957) );
  AOI22_X1 U22968 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19955), .B1(
        n20019), .B2(n19954), .ZN(n19956) );
  OAI211_X1 U22969 ( .C1(n19959), .C2(n19958), .A(n19957), .B(n19956), .ZN(
        P2_U3167) );
  OAI21_X1 U22970 ( .B1(n19961), .B2(n19960), .A(n19970), .ZN(n19967) );
  INV_X1 U22971 ( .A(n20017), .ZN(n19962) );
  OAI211_X1 U22972 ( .C1(n19963), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19962), 
        .B(n19969), .ZN(n19965) );
  AND2_X1 U22973 ( .A1(n19965), .A2(n19964), .ZN(n19966) );
  AND2_X1 U22974 ( .A1(n19967), .A2(n19966), .ZN(n20010) );
  OAI21_X1 U22975 ( .B1(n10583), .B2(n20017), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19968) );
  OAI21_X1 U22976 ( .B1(n19970), .B2(n19969), .A(n19968), .ZN(n20020) );
  AOI22_X1 U22977 ( .A1(n20020), .A2(n19972), .B1(n19971), .B2(n20017), .ZN(
        n19976) );
  AOI22_X1 U22978 ( .A1(n20022), .A2(n19974), .B1(n20005), .B2(n19973), .ZN(
        n19975) );
  OAI211_X1 U22979 ( .C1(n20010), .C2(n19977), .A(n19976), .B(n19975), .ZN(
        P2_U3168) );
  AOI22_X1 U22980 ( .A1(n20020), .A2(n19979), .B1(n19978), .B2(n20017), .ZN(
        n19982) );
  INV_X1 U22981 ( .A(n20010), .ZN(n20023) );
  AOI22_X1 U22982 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20023), .B1(
        n20005), .B2(n19980), .ZN(n19981) );
  OAI211_X1 U22983 ( .C1(n19983), .C2(n20001), .A(n19982), .B(n19981), .ZN(
        P2_U3169) );
  AOI22_X1 U22984 ( .A1(n20020), .A2(n19985), .B1(n19984), .B2(n20017), .ZN(
        n19988) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20023), .B1(
        n20005), .B2(n19986), .ZN(n19987) );
  OAI211_X1 U22986 ( .C1(n19989), .C2(n20001), .A(n19988), .B(n19987), .ZN(
        P2_U3170) );
  AOI22_X1 U22987 ( .A1(n20020), .A2(n19991), .B1(n19990), .B2(n20017), .ZN(
        n19994) );
  AOI22_X1 U22988 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20023), .B1(
        n20022), .B2(n19992), .ZN(n19993) );
  OAI211_X1 U22989 ( .C1(n19995), .C2(n20026), .A(n19994), .B(n19993), .ZN(
        P2_U3171) );
  AOI22_X1 U22990 ( .A1(n20020), .A2(n19997), .B1(n19996), .B2(n20017), .ZN(
        n20000) );
  AOI22_X1 U22991 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20023), .B1(
        n20005), .B2(n19998), .ZN(n19999) );
  OAI211_X1 U22992 ( .C1(n20002), .C2(n20001), .A(n20000), .B(n19999), .ZN(
        P2_U3172) );
  INV_X1 U22993 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20009) );
  AOI22_X1 U22994 ( .A1(n20020), .A2(n20003), .B1(n19485), .B2(n20017), .ZN(
        n20008) );
  AOI22_X1 U22995 ( .A1(n20022), .A2(n20006), .B1(n20005), .B2(n20004), .ZN(
        n20007) );
  OAI211_X1 U22996 ( .C1(n20010), .C2(n20009), .A(n20008), .B(n20007), .ZN(
        P2_U3173) );
  AOI22_X1 U22997 ( .A1(n20020), .A2(n20012), .B1(n20011), .B2(n20017), .ZN(
        n20015) );
  AOI22_X1 U22998 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20023), .B1(
        n20022), .B2(n20013), .ZN(n20014) );
  OAI211_X1 U22999 ( .C1(n20016), .C2(n20026), .A(n20015), .B(n20014), .ZN(
        P2_U3174) );
  AOI22_X1 U23000 ( .A1(n20020), .A2(n20019), .B1(n20018), .B2(n20017), .ZN(
        n20025) );
  AOI22_X1 U23001 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20023), .B1(
        n20022), .B2(n20021), .ZN(n20024) );
  OAI211_X1 U23002 ( .C1(n20027), .C2(n20026), .A(n20025), .B(n20024), .ZN(
        P2_U3175) );
  INV_X1 U23003 ( .A(n20096), .ZN(n20028) );
  AND2_X1 U23004 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20028), .ZN(
        P2_U3179) );
  AND2_X1 U23005 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20028), .ZN(
        P2_U3180) );
  AND2_X1 U23006 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20028), .ZN(
        P2_U3181) );
  AND2_X1 U23007 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20028), .ZN(
        P2_U3182) );
  AND2_X1 U23008 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20028), .ZN(
        P2_U3183) );
  AND2_X1 U23009 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20028), .ZN(
        P2_U3184) );
  AND2_X1 U23010 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20028), .ZN(
        P2_U3185) );
  AND2_X1 U23011 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20028), .ZN(
        P2_U3186) );
  AND2_X1 U23012 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20028), .ZN(
        P2_U3187) );
  AND2_X1 U23013 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20028), .ZN(
        P2_U3188) );
  AND2_X1 U23014 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20028), .ZN(
        P2_U3189) );
  AND2_X1 U23015 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20028), .ZN(
        P2_U3190) );
  AND2_X1 U23016 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20028), .ZN(
        P2_U3191) );
  AND2_X1 U23017 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20028), .ZN(
        P2_U3192) );
  AND2_X1 U23018 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20028), .ZN(
        P2_U3193) );
  AND2_X1 U23019 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20028), .ZN(
        P2_U3194) );
  AND2_X1 U23020 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20028), .ZN(
        P2_U3195) );
  AND2_X1 U23021 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20028), .ZN(
        P2_U3196) );
  AND2_X1 U23022 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20028), .ZN(
        P2_U3197) );
  AND2_X1 U23023 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20028), .ZN(
        P2_U3198) );
  AND2_X1 U23024 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20028), .ZN(
        P2_U3199) );
  AND2_X1 U23025 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20028), .ZN(
        P2_U3200) );
  AND2_X1 U23026 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20028), .ZN(P2_U3201) );
  AND2_X1 U23027 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20028), .ZN(P2_U3202) );
  AND2_X1 U23028 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20028), .ZN(P2_U3203) );
  AND2_X1 U23029 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20028), .ZN(P2_U3204) );
  AND2_X1 U23030 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20028), .ZN(P2_U3205) );
  AND2_X1 U23031 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20028), .ZN(P2_U3206) );
  AND2_X1 U23032 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20028), .ZN(P2_U3207) );
  AND2_X1 U23033 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20028), .ZN(P2_U3208) );
  AND2_X1 U23034 ( .A1(n20029), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20039) );
  INV_X1 U23035 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20157) );
  NOR3_X1 U23036 ( .A1(n20039), .A2(n20157), .A3(n20043), .ZN(n20032) );
  OAI211_X1 U23037 ( .C1(HOLD), .C2(n20157), .A(n20160), .B(n20030), .ZN(
        n20031) );
  NAND2_X1 U23038 ( .A1(NA), .A2(n20033), .ZN(n20038) );
  OAI211_X1 U23039 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20032), .A(n20031), 
        .B(n20038), .ZN(P2_U3209) );
  OAI22_X1 U23040 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20033), .B1(HOLD), .B2(
        n20043), .ZN(n20034) );
  AOI21_X1 U23041 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n20034), .A(n20039), .ZN(n20036) );
  OAI211_X1 U23042 ( .C1(n21071), .C2(n20037), .A(n20036), .B(n20035), .ZN(
        P2_U3210) );
  INV_X1 U23043 ( .A(n20038), .ZN(n20045) );
  NOR3_X1 U23044 ( .A1(HOLD), .A2(n20039), .A3(n20043), .ZN(n20044) );
  NOR2_X1 U23045 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(HOLD), .ZN(n20042)
         );
  AOI22_X1 U23046 ( .A1(n20040), .A2(n20157), .B1(n20039), .B2(n21000), .ZN(
        n20041) );
  OAI33_X1 U23047 ( .A1(n20046), .A2(n20045), .A3(n20044), .B1(n20043), .B2(
        n20042), .B3(n20041), .ZN(P2_U3211) );
  OAI222_X1 U23048 ( .A1(n20089), .A2(n15371), .B1(n20047), .B2(n20159), .C1(
        n13256), .C2(n20086), .ZN(P2_U3212) );
  OAI222_X1 U23049 ( .A1(n20086), .A2(n15371), .B1(n20048), .B2(n20159), .C1(
        n13804), .C2(n20089), .ZN(P2_U3213) );
  OAI222_X1 U23050 ( .A1(n20086), .A2(n13804), .B1(n20049), .B2(n20159), .C1(
        n11000), .C2(n20089), .ZN(P2_U3214) );
  OAI222_X1 U23051 ( .A1(n20089), .A2(n13852), .B1(n20050), .B2(n20159), .C1(
        n11000), .C2(n20086), .ZN(P2_U3215) );
  OAI222_X1 U23052 ( .A1(n20089), .A2(n11007), .B1(n20051), .B2(n20159), .C1(
        n13852), .C2(n20086), .ZN(P2_U3216) );
  OAI222_X1 U23053 ( .A1(n20089), .A2(n11012), .B1(n20052), .B2(n20159), .C1(
        n11007), .C2(n20086), .ZN(P2_U3217) );
  OAI222_X1 U23054 ( .A1(n20089), .A2(n11030), .B1(n20053), .B2(n20159), .C1(
        n11012), .C2(n20086), .ZN(P2_U3218) );
  OAI222_X1 U23055 ( .A1(n20089), .A2(n11031), .B1(n20054), .B2(n20159), .C1(
        n11030), .C2(n20086), .ZN(P2_U3219) );
  OAI222_X1 U23056 ( .A1(n20089), .A2(n11063), .B1(n20055), .B2(n20159), .C1(
        n11031), .C2(n20086), .ZN(P2_U3220) );
  OAI222_X1 U23057 ( .A1(n20089), .A2(n11064), .B1(n20056), .B2(n20159), .C1(
        n11063), .C2(n20086), .ZN(P2_U3221) );
  OAI222_X1 U23058 ( .A1(n20089), .A2(n11094), .B1(n20057), .B2(n20159), .C1(
        n11064), .C2(n20086), .ZN(P2_U3222) );
  OAI222_X1 U23059 ( .A1(n20089), .A2(n11095), .B1(n20058), .B2(n20159), .C1(
        n11094), .C2(n20086), .ZN(P2_U3223) );
  OAI222_X1 U23060 ( .A1(n20089), .A2(n15845), .B1(n20059), .B2(n20159), .C1(
        n11095), .C2(n20086), .ZN(P2_U3224) );
  OAI222_X1 U23061 ( .A1(n20089), .A2(n11140), .B1(n20060), .B2(n20159), .C1(
        n15845), .C2(n20086), .ZN(P2_U3225) );
  OAI222_X1 U23062 ( .A1(n20089), .A2(n20062), .B1(n20061), .B2(n20159), .C1(
        n11140), .C2(n20086), .ZN(P2_U3226) );
  OAI222_X1 U23063 ( .A1(n20089), .A2(n10912), .B1(n20063), .B2(n20159), .C1(
        n20062), .C2(n20086), .ZN(P2_U3227) );
  OAI222_X1 U23064 ( .A1(n20089), .A2(n20065), .B1(n20064), .B2(n20159), .C1(
        n10912), .C2(n20086), .ZN(P2_U3228) );
  OAI222_X1 U23065 ( .A1(n20089), .A2(n11147), .B1(n20066), .B2(n20159), .C1(
        n20065), .C2(n20086), .ZN(P2_U3229) );
  OAI222_X1 U23066 ( .A1(n20089), .A2(n20068), .B1(n20067), .B2(n20159), .C1(
        n11147), .C2(n20086), .ZN(P2_U3230) );
  OAI222_X1 U23067 ( .A1(n20089), .A2(n20070), .B1(n20069), .B2(n20159), .C1(
        n20068), .C2(n20086), .ZN(P2_U3231) );
  OAI222_X1 U23068 ( .A1(n20089), .A2(n20072), .B1(n20071), .B2(n20159), .C1(
        n20070), .C2(n20086), .ZN(P2_U3232) );
  OAI222_X1 U23069 ( .A1(n20089), .A2(n20074), .B1(n20073), .B2(n20159), .C1(
        n20072), .C2(n20086), .ZN(P2_U3233) );
  OAI222_X1 U23070 ( .A1(n20089), .A2(n20076), .B1(n20075), .B2(n20159), .C1(
        n20074), .C2(n20086), .ZN(P2_U3234) );
  OAI222_X1 U23071 ( .A1(n20089), .A2(n11220), .B1(n20077), .B2(n20159), .C1(
        n20076), .C2(n20086), .ZN(P2_U3235) );
  OAI222_X1 U23072 ( .A1(n20089), .A2(n20079), .B1(n20078), .B2(n20159), .C1(
        n11220), .C2(n20086), .ZN(P2_U3236) );
  OAI222_X1 U23073 ( .A1(n20089), .A2(n20082), .B1(n20080), .B2(n20159), .C1(
        n20079), .C2(n20086), .ZN(P2_U3237) );
  OAI222_X1 U23074 ( .A1(n20086), .A2(n20082), .B1(n20081), .B2(n20159), .C1(
        n20083), .C2(n20089), .ZN(P2_U3238) );
  OAI222_X1 U23075 ( .A1(n20089), .A2(n16328), .B1(n20084), .B2(n20159), .C1(
        n20083), .C2(n20086), .ZN(P2_U3239) );
  OAI222_X1 U23076 ( .A1(n20089), .A2(n20087), .B1(n20085), .B2(n20159), .C1(
        n16328), .C2(n20086), .ZN(P2_U3240) );
  INV_X1 U23077 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20088) );
  OAI222_X1 U23078 ( .A1(n20089), .A2(n15271), .B1(n20088), .B2(n20159), .C1(
        n20087), .C2(n20086), .ZN(P2_U3241) );
  OAI22_X1 U23079 ( .A1(n20160), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20159), .ZN(n20090) );
  INV_X1 U23080 ( .A(n20090), .ZN(P2_U3585) );
  MUX2_X1 U23081 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20160), .Z(P2_U3586) );
  OAI22_X1 U23082 ( .A1(n20160), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20159), .ZN(n20091) );
  INV_X1 U23083 ( .A(n20091), .ZN(P2_U3587) );
  OAI22_X1 U23084 ( .A1(n20160), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20159), .ZN(n20092) );
  INV_X1 U23085 ( .A(n20092), .ZN(P2_U3588) );
  OAI21_X1 U23086 ( .B1(n20096), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20094), 
        .ZN(n20093) );
  INV_X1 U23087 ( .A(n20093), .ZN(P2_U3591) );
  OAI21_X1 U23088 ( .B1(n20096), .B2(n20095), .A(n20094), .ZN(P2_U3592) );
  NAND2_X1 U23089 ( .A1(n20107), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20120) );
  NOR2_X1 U23090 ( .A1(n20097), .A2(n20120), .ZN(n20113) );
  OAI21_X1 U23091 ( .B1(n20099), .B2(n20098), .A(n20107), .ZN(n20101) );
  NAND2_X1 U23092 ( .A1(n20101), .A2(n20100), .ZN(n20112) );
  NOR2_X1 U23093 ( .A1(n20113), .A2(n20112), .ZN(n20104) );
  OAI22_X1 U23094 ( .A1(n20104), .A2(n20103), .B1(n19854), .B2(n20102), .ZN(
        n20105) );
  AOI21_X1 U23095 ( .B1(n20107), .B2(n20106), .A(n20105), .ZN(n20108) );
  AOI22_X1 U23096 ( .A1(n20133), .A2(n20109), .B1(n20108), .B2(n20134), .ZN(
        P2_U3602) );
  AOI22_X1 U23097 ( .A1(n20112), .A2(n20111), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20110), .ZN(n20115) );
  NOR2_X1 U23098 ( .A1(n20133), .A2(n20113), .ZN(n20114) );
  AOI22_X1 U23099 ( .A1(n20116), .A2(n20133), .B1(n20115), .B2(n20114), .ZN(
        P2_U3603) );
  INV_X1 U23100 ( .A(n20117), .ZN(n20118) );
  NAND3_X1 U23101 ( .A1(n20121), .A2(n20126), .A3(n20118), .ZN(n20119) );
  OAI21_X1 U23102 ( .B1(n20121), .B2(n20120), .A(n20119), .ZN(n20122) );
  AOI21_X1 U23103 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20123), .A(n20122), 
        .ZN(n20124) );
  AOI22_X1 U23104 ( .A1(n20133), .A2(n20125), .B1(n20124), .B2(n20134), .ZN(
        P2_U3604) );
  INV_X1 U23105 ( .A(n20126), .ZN(n20129) );
  OAI22_X1 U23106 ( .A1(n20130), .A2(n20129), .B1(n20128), .B2(n20127), .ZN(
        n20131) );
  AOI21_X1 U23107 ( .B1(n20135), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20131), 
        .ZN(n20132) );
  OAI22_X1 U23108 ( .A1(n20135), .A2(n20134), .B1(n20133), .B2(n20132), .ZN(
        P2_U3605) );
  INV_X1 U23109 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20136) );
  AOI22_X1 U23110 ( .A1(n20159), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20136), 
        .B2(n20160), .ZN(P2_U3608) );
  AOI22_X1 U23111 ( .A1(n20140), .A2(n20139), .B1(n20138), .B2(n20137), .ZN(
        n20141) );
  NAND2_X1 U23112 ( .A1(n20142), .A2(n20141), .ZN(n20144) );
  MUX2_X1 U23113 ( .A(P2_MORE_REG_SCAN_IN), .B(n20144), .S(n20143), .Z(
        P2_U3609) );
  AOI22_X1 U23114 ( .A1(n20146), .A2(n20150), .B1(n19854), .B2(n20145), .ZN(
        n20147) );
  NAND2_X1 U23115 ( .A1(n20148), .A2(n20147), .ZN(n20158) );
  AOI21_X1 U23116 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20150), .A(n20149), 
        .ZN(n20155) );
  OAI21_X1 U23117 ( .B1(n20152), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20151), 
        .ZN(n20153) );
  AND3_X1 U23118 ( .A1(n13122), .A2(n20153), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20154) );
  OAI21_X1 U23119 ( .B1(n20155), .B2(n20154), .A(n20158), .ZN(n20156) );
  OAI21_X1 U23120 ( .B1(n20158), .B2(n20157), .A(n20156), .ZN(P2_U3610) );
  OAI22_X1 U23121 ( .A1(n20160), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20159), .ZN(n20161) );
  INV_X1 U23122 ( .A(n20161), .ZN(P2_U3611) );
  AOI21_X1 U23123 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20883), .A(n12994), 
        .ZN(n20879) );
  INV_X1 U23124 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21075) );
  NAND2_X1 U23125 ( .A1(n12994), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20916) );
  AOI21_X1 U23126 ( .B1(n20879), .B2(n21075), .A(n20962), .ZN(P1_U2802) );
  OAI21_X1 U23127 ( .B1(n20163), .B2(n20162), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20164) );
  OAI21_X1 U23128 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20165), .A(n20164), 
        .ZN(P1_U2803) );
  INV_X1 U23129 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20991) );
  NOR2_X1 U23130 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20882) );
  NOR2_X1 U23131 ( .A1(n20962), .A2(n20882), .ZN(n20166) );
  AOI22_X1 U23132 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20962), .B1(n20991), 
        .B2(n20166), .ZN(P1_U2804) );
  NOR2_X1 U23133 ( .A1(n20962), .A2(n20879), .ZN(n20934) );
  OAI21_X1 U23134 ( .B1(BS16), .B2(n20882), .A(n20934), .ZN(n20932) );
  OAI21_X1 U23135 ( .B1(n20934), .B2(n21022), .A(n20932), .ZN(P1_U2805) );
  OAI21_X1 U23136 ( .B1(n20169), .B2(n20168), .A(n20167), .ZN(P1_U2806) );
  NOR4_X1 U23137 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20173) );
  NOR4_X1 U23138 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20172) );
  NOR4_X1 U23139 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20171) );
  NOR4_X1 U23140 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20170) );
  NAND4_X1 U23141 ( .A1(n20173), .A2(n20172), .A3(n20171), .A4(n20170), .ZN(
        n20179) );
  NOR4_X1 U23142 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20177) );
  AOI211_X1 U23143 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20176) );
  NOR4_X1 U23144 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20175) );
  NOR4_X1 U23145 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20174) );
  NAND4_X1 U23146 ( .A1(n20177), .A2(n20176), .A3(n20175), .A4(n20174), .ZN(
        n20178) );
  NOR2_X1 U23147 ( .A1(n20179), .A2(n20178), .ZN(n20946) );
  INV_X1 U23148 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21081) );
  NOR3_X1 U23149 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20181) );
  OAI21_X1 U23150 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20181), .A(n20946), .ZN(
        n20180) );
  OAI21_X1 U23151 ( .B1(n20946), .B2(n21081), .A(n20180), .ZN(P1_U2807) );
  INV_X1 U23152 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20933) );
  AOI21_X1 U23153 ( .B1(n13825), .B2(n20933), .A(n20181), .ZN(n20183) );
  INV_X1 U23154 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20182) );
  INV_X1 U23155 ( .A(n20946), .ZN(n20944) );
  AOI22_X1 U23156 ( .A1(n20946), .A2(n20183), .B1(n20182), .B2(n20944), .ZN(
        P1_U2808) );
  NOR3_X1 U23157 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20220), .A3(n20184), .ZN(
        n20189) );
  AOI22_X1 U23158 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20215), .B1(
        n20185), .B2(n20229), .ZN(n20186) );
  OAI211_X1 U23159 ( .C1(n20243), .C2(n20187), .A(n20186), .B(n20351), .ZN(
        n20188) );
  AOI211_X1 U23160 ( .C1(n20250), .C2(P1_EBX_REG_8__SCAN_IN), .A(n20189), .B(
        n20188), .ZN(n20193) );
  AOI22_X1 U23161 ( .A1(n20191), .A2(n20210), .B1(P1_REIP_REG_8__SCAN_IN), 
        .B2(n20190), .ZN(n20192) );
  NAND2_X1 U23162 ( .A1(n20193), .A2(n20192), .ZN(P1_U2832) );
  NOR2_X1 U23163 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20220), .ZN(n20194) );
  AOI22_X1 U23164 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20250), .B1(n20202), .B2(
        n20194), .ZN(n20201) );
  OAI22_X1 U23165 ( .A1(n20196), .A2(n20245), .B1(n20195), .B2(n20244), .ZN(
        n20197) );
  AOI211_X1 U23166 ( .C1(n20257), .C2(n20260), .A(n20377), .B(n20197), .ZN(
        n20200) );
  OAI21_X1 U23167 ( .B1(n20220), .B2(n20202), .A(n20198), .ZN(n20209) );
  AOI22_X1 U23168 ( .A1(n20261), .A2(n20210), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20209), .ZN(n20199) );
  NAND3_X1 U23169 ( .A1(n20201), .A2(n20200), .A3(n20199), .ZN(P1_U2833) );
  OR2_X1 U23170 ( .A1(n20220), .A2(n20202), .ZN(n20214) );
  OAI21_X1 U23171 ( .B1(n20204), .B2(n20232), .A(n20203), .ZN(n20236) );
  NAND2_X1 U23172 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20236), .ZN(n20222) );
  AOI22_X1 U23173 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20250), .B1(n20257), .B2(
        n20205), .ZN(n20206) );
  OAI21_X1 U23174 ( .B1(n20207), .B2(n20244), .A(n20206), .ZN(n20208) );
  AOI211_X1 U23175 ( .C1(n20215), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20377), .B(n20208), .ZN(n20213) );
  AOI22_X1 U23176 ( .A1(n20211), .A2(n20210), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20209), .ZN(n20212) );
  OAI211_X1 U23177 ( .C1(n20214), .C2(n20222), .A(n20213), .B(n20212), .ZN(
        P1_U2834) );
  INV_X1 U23178 ( .A(n20264), .ZN(n20218) );
  AOI22_X1 U23179 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20215), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(n20250), .ZN(n20216) );
  INV_X1 U23180 ( .A(n20216), .ZN(n20217) );
  AOI211_X1 U23181 ( .C1(n20257), .C2(n20218), .A(n20377), .B(n20217), .ZN(
        n20225) );
  OAI21_X1 U23182 ( .B1(n20220), .B2(n20232), .A(n20219), .ZN(n20221) );
  AOI22_X1 U23183 ( .A1(n20223), .A2(n20247), .B1(n20222), .B2(n20221), .ZN(
        n20224) );
  OAI211_X1 U23184 ( .C1(n20226), .C2(n20244), .A(n20225), .B(n20224), .ZN(
        P1_U2835) );
  AOI22_X1 U23185 ( .A1(n20230), .A2(n20229), .B1(n20228), .B2(n20227), .ZN(
        n20242) );
  INV_X1 U23186 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20887) );
  NOR2_X1 U23187 ( .A1(n20887), .A2(n20231), .ZN(n20233) );
  NAND3_X1 U23188 ( .A1(n20233), .A2(n20248), .A3(n20232), .ZN(n20234) );
  OAI211_X1 U23189 ( .C1(n20245), .C2(n20235), .A(n20351), .B(n20234), .ZN(
        n20240) );
  OAI22_X1 U23190 ( .A1(n20238), .A2(n20237), .B1(n13957), .B2(n20236), .ZN(
        n20239) );
  AOI211_X1 U23191 ( .C1(P1_EBX_REG_4__SCAN_IN), .C2(n20250), .A(n20240), .B(
        n20239), .ZN(n20241) );
  OAI211_X1 U23192 ( .C1(n20243), .C2(n20353), .A(n20242), .B(n20241), .ZN(
        P1_U2836) );
  INV_X1 U23193 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20246) );
  OAI22_X1 U23194 ( .A1(n20246), .A2(n20245), .B1(n20337), .B2(n20244), .ZN(
        n20256) );
  NAND2_X1 U23195 ( .A1(n20334), .A2(n20247), .ZN(n20252) );
  AND4_X1 U23196 ( .A1(n20248), .A2(n20887), .A3(P1_REIP_REG_1__SCAN_IN), .A4(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20249) );
  AOI21_X1 U23197 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(n20250), .A(n20249), .ZN(
        n20251) );
  OAI211_X1 U23198 ( .C1(n20254), .C2(n20253), .A(n20252), .B(n20251), .ZN(
        n20255) );
  AOI211_X1 U23199 ( .C1(n20257), .C2(n20361), .A(n20256), .B(n20255), .ZN(
        n20258) );
  OAI21_X1 U23200 ( .B1(n20887), .B2(n20259), .A(n20258), .ZN(P1_U2837) );
  AOI22_X1 U23201 ( .A1(n20261), .A2(n12977), .B1(n12975), .B2(n20260), .ZN(
        n20262) );
  OAI21_X1 U23202 ( .B1(n20270), .B2(n20263), .A(n20262), .ZN(P1_U2865) );
  OAI22_X1 U23203 ( .A1(n20266), .A2(n14842), .B1(n20265), .B2(n20264), .ZN(
        n20267) );
  INV_X1 U23204 ( .A(n20267), .ZN(n20268) );
  OAI21_X1 U23205 ( .B1(n20270), .B2(n20269), .A(n20268), .ZN(P1_U2867) );
  AOI22_X1 U23206 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20274), .B1(n16031), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20271) );
  OAI21_X1 U23207 ( .B1(n20273), .B2(n20272), .A(n20271), .ZN(P1_U2921) );
  INV_X1 U23208 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20276) );
  AOI22_X1 U23209 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20275) );
  OAI21_X1 U23210 ( .B1(n20276), .B2(n20303), .A(n20275), .ZN(P1_U2922) );
  INV_X1 U23211 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20278) );
  AOI22_X1 U23212 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20277) );
  OAI21_X1 U23213 ( .B1(n20278), .B2(n20303), .A(n20277), .ZN(P1_U2923) );
  INV_X1 U23214 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20280) );
  AOI22_X1 U23215 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20279) );
  OAI21_X1 U23216 ( .B1(n20280), .B2(n20303), .A(n20279), .ZN(P1_U2924) );
  AOI22_X1 U23217 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20281) );
  OAI21_X1 U23218 ( .B1(n20282), .B2(n20303), .A(n20281), .ZN(P1_U2925) );
  INV_X1 U23219 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20284) );
  AOI22_X1 U23220 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20283) );
  OAI21_X1 U23221 ( .B1(n20284), .B2(n20303), .A(n20283), .ZN(P1_U2926) );
  INV_X1 U23222 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20286) );
  AOI22_X1 U23223 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20285) );
  OAI21_X1 U23224 ( .B1(n20286), .B2(n20303), .A(n20285), .ZN(P1_U2927) );
  INV_X1 U23225 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20288) );
  AOI22_X1 U23226 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20287) );
  OAI21_X1 U23227 ( .B1(n20288), .B2(n20303), .A(n20287), .ZN(P1_U2928) );
  AOI22_X1 U23228 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20289) );
  OAI21_X1 U23229 ( .B1(n11898), .B2(n20303), .A(n20289), .ZN(P1_U2929) );
  AOI22_X1 U23230 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20290) );
  OAI21_X1 U23231 ( .B1(n20291), .B2(n20303), .A(n20290), .ZN(P1_U2930) );
  AOI22_X1 U23232 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20292) );
  OAI21_X1 U23233 ( .B1(n11863), .B2(n20303), .A(n20292), .ZN(P1_U2931) );
  AOI22_X1 U23234 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20293) );
  OAI21_X1 U23235 ( .B1(n20294), .B2(n20303), .A(n20293), .ZN(P1_U2932) );
  AOI22_X1 U23236 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20295) );
  OAI21_X1 U23237 ( .B1(n20296), .B2(n20303), .A(n20295), .ZN(P1_U2933) );
  AOI22_X1 U23238 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20297) );
  OAI21_X1 U23239 ( .B1(n20298), .B2(n20303), .A(n20297), .ZN(P1_U2934) );
  AOI22_X1 U23240 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20299) );
  OAI21_X1 U23241 ( .B1(n20300), .B2(n20303), .A(n20299), .ZN(P1_U2935) );
  AOI22_X1 U23242 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20301), .B1(n16031), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20302) );
  OAI21_X1 U23243 ( .B1(n20304), .B2(n20303), .A(n20302), .ZN(P1_U2936) );
  AOI22_X1 U23244 ( .A1(n20327), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20326), .ZN(n20306) );
  NAND2_X1 U23245 ( .A1(n20314), .A2(n20305), .ZN(n20316) );
  NAND2_X1 U23246 ( .A1(n20306), .A2(n20316), .ZN(P1_U2945) );
  AOI22_X1 U23247 ( .A1(n20327), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20308) );
  NAND2_X1 U23248 ( .A1(n20314), .A2(n20307), .ZN(n20320) );
  NAND2_X1 U23249 ( .A1(n20308), .A2(n20320), .ZN(P1_U2947) );
  AOI22_X1 U23250 ( .A1(n20327), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20310) );
  NAND2_X1 U23251 ( .A1(n20314), .A2(n20309), .ZN(n20322) );
  NAND2_X1 U23252 ( .A1(n20310), .A2(n20322), .ZN(P1_U2949) );
  AOI22_X1 U23253 ( .A1(n20327), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20312) );
  NAND2_X1 U23254 ( .A1(n20314), .A2(n20311), .ZN(n20324) );
  NAND2_X1 U23255 ( .A1(n20312), .A2(n20324), .ZN(P1_U2950) );
  AOI22_X1 U23256 ( .A1(n20327), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20326), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20315) );
  NAND2_X1 U23257 ( .A1(n20314), .A2(n20313), .ZN(n20328) );
  NAND2_X1 U23258 ( .A1(n20315), .A2(n20328), .ZN(P1_U2951) );
  AOI22_X1 U23259 ( .A1(n20327), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20317) );
  NAND2_X1 U23260 ( .A1(n20317), .A2(n20316), .ZN(P1_U2960) );
  AOI22_X1 U23261 ( .A1(n20327), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20326), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20319) );
  NAND2_X1 U23262 ( .A1(n20319), .A2(n20318), .ZN(P1_U2961) );
  AOI22_X1 U23263 ( .A1(n20327), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20326), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20321) );
  NAND2_X1 U23264 ( .A1(n20321), .A2(n20320), .ZN(P1_U2962) );
  AOI22_X1 U23265 ( .A1(n20327), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20326), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20323) );
  NAND2_X1 U23266 ( .A1(n20323), .A2(n20322), .ZN(P1_U2964) );
  AOI22_X1 U23267 ( .A1(n20327), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20326), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20325) );
  NAND2_X1 U23268 ( .A1(n20325), .A2(n20324), .ZN(P1_U2965) );
  AOI22_X1 U23269 ( .A1(n20327), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20326), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20329) );
  NAND2_X1 U23270 ( .A1(n20329), .A2(n20328), .ZN(P1_U2966) );
  AOI22_X1 U23271 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n20336) );
  OAI21_X1 U23272 ( .B1(n20332), .B2(n20331), .A(n20330), .ZN(n20333) );
  INV_X1 U23273 ( .A(n20333), .ZN(n20360) );
  AOI22_X1 U23274 ( .A1(n20334), .A2(n20344), .B1(n20343), .B2(n20360), .ZN(
        n20335) );
  OAI211_X1 U23275 ( .C1(n20349), .C2(n20337), .A(n20336), .B(n20335), .ZN(
        P1_U2996) );
  AOI22_X1 U23276 ( .A1(n20338), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20377), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n20347) );
  OAI21_X1 U23277 ( .B1(n20341), .B2(n20340), .A(n20339), .ZN(n20342) );
  INV_X1 U23278 ( .A(n20342), .ZN(n20376) );
  AOI22_X1 U23279 ( .A1(n20345), .A2(n20344), .B1(n20343), .B2(n20376), .ZN(
        n20346) );
  OAI211_X1 U23280 ( .C1(n20349), .C2(n20348), .A(n20347), .B(n20346), .ZN(
        P1_U2997) );
  INV_X1 U23281 ( .A(n20350), .ZN(n20357) );
  OAI22_X1 U23282 ( .A1(n20353), .A2(n20352), .B1(n13957), .B2(n20351), .ZN(
        n20356) );
  AOI211_X1 U23283 ( .C1(n20359), .C2(n20364), .A(n20354), .B(n20365), .ZN(
        n20355) );
  AOI211_X1 U23284 ( .C1(n20357), .C2(n20375), .A(n20356), .B(n20355), .ZN(
        n20358) );
  OAI21_X1 U23285 ( .B1(n20363), .B2(n20359), .A(n20358), .ZN(P1_U3027) );
  AOI222_X1 U23286 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20377), .B1(n20372), 
        .B2(n20361), .C1(n20375), .C2(n20360), .ZN(n20362) );
  OAI221_X1 U23287 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20365), .C1(
        n20364), .C2(n20363), .A(n20362), .ZN(P1_U3028) );
  INV_X1 U23288 ( .A(n20366), .ZN(n20373) );
  NOR4_X1 U23289 ( .A1(n20369), .A2(n20368), .A3(n20367), .A4(n20380), .ZN(
        n20370) );
  AOI211_X1 U23290 ( .C1(n20373), .C2(n20372), .A(n20371), .B(n20370), .ZN(
        n20384) );
  AOI22_X1 U23291 ( .A1(n20376), .A2(n20375), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20374), .ZN(n20383) );
  NAND2_X1 U23292 ( .A1(n20377), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20382) );
  NAND4_X1 U23293 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20380), .A3(
        n20379), .A4(n20378), .ZN(n20381) );
  NAND4_X1 U23294 ( .A1(n20384), .A2(n20383), .A3(n20382), .A4(n20381), .ZN(
        P1_U3029) );
  NOR2_X1 U23295 ( .A1(n20386), .A2(n20385), .ZN(P1_U3032) );
  INV_X1 U23296 ( .A(n20804), .ZN(n20387) );
  OAI22_X1 U23297 ( .A1(n20863), .A2(n20657), .B1(n20400), .B2(n20387), .ZN(
        n20388) );
  INV_X1 U23298 ( .A(n20388), .ZN(n20390) );
  AOI22_X1 U23299 ( .A1(n20803), .A2(n20402), .B1(n20427), .B2(n20694), .ZN(
        n20389) );
  OAI211_X1 U23300 ( .C1(n20406), .C2(n20391), .A(n20390), .B(n20389), .ZN(
        P1_U3033) );
  INV_X1 U23301 ( .A(n20817), .ZN(n20443) );
  OAI22_X1 U23302 ( .A1(n20863), .A2(n20821), .B1(n20400), .B2(n20443), .ZN(
        n20392) );
  INV_X1 U23303 ( .A(n20392), .ZN(n20394) );
  AOI22_X1 U23304 ( .A1(n20816), .A2(n20402), .B1(n20427), .B2(n20818), .ZN(
        n20393) );
  OAI211_X1 U23305 ( .C1(n20406), .C2(n20395), .A(n20394), .B(n20393), .ZN(
        P1_U3034) );
  INV_X1 U23306 ( .A(n20840), .ZN(n20459) );
  OAI22_X1 U23307 ( .A1(n20863), .A2(n20847), .B1(n20400), .B2(n20459), .ZN(
        n20396) );
  INV_X1 U23308 ( .A(n20396), .ZN(n20398) );
  AOI22_X1 U23309 ( .A1(n20841), .A2(n20402), .B1(n20427), .B2(n20842), .ZN(
        n20397) );
  OAI211_X1 U23310 ( .C1(n20406), .C2(n20399), .A(n20398), .B(n20397), .ZN(
        P1_U3038) );
  INV_X1 U23311 ( .A(n20848), .ZN(n20463) );
  OAI22_X1 U23312 ( .A1(n20863), .A2(n9789), .B1(n20400), .B2(n20463), .ZN(
        n20401) );
  INV_X1 U23313 ( .A(n20401), .ZN(n20404) );
  AOI22_X1 U23314 ( .A1(n20849), .A2(n20402), .B1(n20427), .B2(n20715), .ZN(
        n20403) );
  OAI211_X1 U23315 ( .C1(n20406), .C2(n20405), .A(n20404), .B(n20403), .ZN(
        P1_U3039) );
  NOR2_X1 U23316 ( .A1(n20647), .A2(n20407), .ZN(n20425) );
  AOI21_X1 U23317 ( .B1(n20478), .B2(n20648), .A(n20425), .ZN(n20408) );
  OAI22_X1 U23318 ( .A1(n20408), .A2(n20802), .B1(n20407), .B2(n11760), .ZN(
        n20426) );
  AOI22_X1 U23319 ( .A1(n20426), .A2(n20803), .B1(n20804), .B2(n20425), .ZN(
        n20412) );
  OAI211_X1 U23320 ( .C1(n20485), .C2(n21022), .A(n20810), .B(n20408), .ZN(
        n20409) );
  OAI211_X1 U23321 ( .C1(n20677), .C2(n20410), .A(n20809), .B(n20409), .ZN(
        n20428) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20812), .ZN(n20411) );
  OAI211_X1 U23323 ( .C1(n20815), .C2(n20469), .A(n20412), .B(n20411), .ZN(
        P1_U3041) );
  AOI22_X1 U23324 ( .A1(n20426), .A2(n20816), .B1(n20817), .B2(n20425), .ZN(
        n20414) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20774), .ZN(n20413) );
  OAI211_X1 U23326 ( .C1(n20777), .C2(n20469), .A(n20414), .B(n20413), .ZN(
        P1_U3042) );
  INV_X1 U23327 ( .A(n20824), .ZN(n20781) );
  AOI22_X1 U23328 ( .A1(n20822), .A2(n20426), .B1(n20823), .B2(n20425), .ZN(
        n20416) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20778), .ZN(n20415) );
  OAI211_X1 U23330 ( .C1(n20781), .C2(n20469), .A(n20416), .B(n20415), .ZN(
        P1_U3043) );
  AOI22_X1 U23331 ( .A1(n20828), .A2(n20426), .B1(n20829), .B2(n20425), .ZN(
        n20418) );
  AOI22_X1 U23332 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n9792), .ZN(n20417) );
  OAI211_X1 U23333 ( .C1(n20833), .C2(n20469), .A(n20418), .B(n20417), .ZN(
        P1_U3044) );
  AOI22_X1 U23334 ( .A1(n20834), .A2(n20426), .B1(n20835), .B2(n20425), .ZN(
        n20420) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n9794), .ZN(n20419) );
  OAI211_X1 U23336 ( .C1(n20839), .C2(n20469), .A(n20420), .B(n20419), .ZN(
        P1_U3045) );
  INV_X1 U23337 ( .A(n20842), .ZN(n20789) );
  AOI22_X1 U23338 ( .A1(n20426), .A2(n20841), .B1(n20840), .B2(n20425), .ZN(
        n20422) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20786), .ZN(n20421) );
  OAI211_X1 U23340 ( .C1(n20789), .C2(n20469), .A(n20422), .B(n20421), .ZN(
        P1_U3046) );
  AOI22_X1 U23341 ( .A1(n20426), .A2(n20849), .B1(n20848), .B2(n20425), .ZN(
        n20424) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n9790), .ZN(n20423) );
  OAI211_X1 U23343 ( .C1(n20853), .C2(n20469), .A(n20424), .B(n20423), .ZN(
        P1_U3047) );
  AOI22_X1 U23344 ( .A1(n20855), .A2(n20426), .B1(n20857), .B2(n20425), .ZN(
        n20430) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20858), .ZN(n20429) );
  OAI211_X1 U23346 ( .C1(n20864), .C2(n20469), .A(n20430), .B(n20429), .ZN(
        P1_U3048) );
  NAND2_X1 U23347 ( .A1(n20469), .A2(n20677), .ZN(n20432) );
  NAND2_X1 U23348 ( .A1(n20810), .A2(n21022), .ZN(n20681) );
  OAI21_X1 U23349 ( .B1(n20501), .B2(n20432), .A(n20681), .ZN(n20435) );
  NOR2_X1 U23350 ( .A1(n20433), .A2(n20619), .ZN(n20438) );
  NOR3_X1 U23351 ( .A1(n20686), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20480) );
  NAND2_X1 U23352 ( .A1(n20647), .A2(n20480), .ZN(n20467) );
  INV_X1 U23353 ( .A(n20467), .ZN(n20434) );
  AOI22_X1 U23354 ( .A1(n20501), .A2(n20694), .B1(n20804), .B2(n20434), .ZN(
        n20442) );
  INV_X1 U23355 ( .A(n20435), .ZN(n20439) );
  NOR2_X1 U23356 ( .A1(n10195), .A2(n11760), .ZN(n20562) );
  AOI211_X1 U23357 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20467), .A(n20562), 
        .B(n20436), .ZN(n20437) );
  INV_X1 U23358 ( .A(n20469), .ZN(n20440) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20471), .B1(
        n20440), .B2(n20812), .ZN(n20441) );
  OAI211_X1 U23360 ( .C1(n20474), .C2(n20697), .A(n20442), .B(n20441), .ZN(
        P1_U3049) );
  OAI22_X1 U23361 ( .A1(n20469), .A2(n20821), .B1(n20443), .B2(n20467), .ZN(
        n20444) );
  INV_X1 U23362 ( .A(n20444), .ZN(n20446) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20471), .B1(
        n20501), .B2(n20818), .ZN(n20445) );
  OAI211_X1 U23364 ( .C1(n20474), .C2(n20700), .A(n20446), .B(n20445), .ZN(
        P1_U3050) );
  INV_X1 U23365 ( .A(n20822), .ZN(n20703) );
  OAI22_X1 U23366 ( .A1(n20469), .A2(n20827), .B1(n20447), .B2(n20467), .ZN(
        n20448) );
  INV_X1 U23367 ( .A(n20448), .ZN(n20450) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20471), .B1(
        n20501), .B2(n20824), .ZN(n20449) );
  OAI211_X1 U23369 ( .C1(n20474), .C2(n20703), .A(n20450), .B(n20449), .ZN(
        P1_U3051) );
  OAI22_X1 U23370 ( .A1(n20469), .A2(n9791), .B1(n20451), .B2(n20467), .ZN(
        n20452) );
  INV_X1 U23371 ( .A(n20452), .ZN(n20454) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20471), .B1(
        n20501), .B2(n20704), .ZN(n20453) );
  OAI211_X1 U23373 ( .C1(n20474), .C2(n20707), .A(n20454), .B(n20453), .ZN(
        P1_U3052) );
  OAI22_X1 U23374 ( .A1(n20469), .A2(n9793), .B1(n20455), .B2(n20467), .ZN(
        n20456) );
  INV_X1 U23375 ( .A(n20456), .ZN(n20458) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20471), .B1(
        n20501), .B2(n20708), .ZN(n20457) );
  OAI211_X1 U23377 ( .C1(n20474), .C2(n20711), .A(n20458), .B(n20457), .ZN(
        P1_U3053) );
  INV_X1 U23378 ( .A(n20841), .ZN(n20714) );
  OAI22_X1 U23379 ( .A1(n20469), .A2(n20847), .B1(n20459), .B2(n20467), .ZN(
        n20460) );
  INV_X1 U23380 ( .A(n20460), .ZN(n20462) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20471), .B1(
        n20501), .B2(n20842), .ZN(n20461) );
  OAI211_X1 U23382 ( .C1(n20474), .C2(n20714), .A(n20462), .B(n20461), .ZN(
        P1_U3054) );
  OAI22_X1 U23383 ( .A1(n20469), .A2(n9789), .B1(n20463), .B2(n20467), .ZN(
        n20464) );
  INV_X1 U23384 ( .A(n20464), .ZN(n20466) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20471), .B1(
        n20501), .B2(n20715), .ZN(n20465) );
  OAI211_X1 U23386 ( .C1(n20474), .C2(n20718), .A(n20466), .B(n20465), .ZN(
        P1_U3055) );
  OAI22_X1 U23387 ( .A1(n20469), .A2(n20676), .B1(n20468), .B2(n20467), .ZN(
        n20470) );
  INV_X1 U23388 ( .A(n20470), .ZN(n20473) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20471), .B1(
        n20501), .B2(n20721), .ZN(n20472) );
  OAI211_X1 U23390 ( .C1(n20474), .C2(n20725), .A(n20473), .B(n20472), .ZN(
        P1_U3056) );
  INV_X1 U23391 ( .A(n20485), .ZN(n20476) );
  INV_X1 U23392 ( .A(n20806), .ZN(n20475) );
  AOI21_X1 U23393 ( .B1(n20476), .B2(n20475), .A(n20802), .ZN(n20483) );
  AND2_X1 U23394 ( .A1(n20477), .A2(n11775), .ZN(n20799) );
  NOR2_X1 U23395 ( .A1(n20728), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20500) );
  AOI21_X1 U23396 ( .B1(n20478), .B2(n20799), .A(n20500), .ZN(n20482) );
  INV_X1 U23397 ( .A(n20482), .ZN(n20479) );
  AOI22_X1 U23398 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20480), .B1(n20483), 
        .B2(n20479), .ZN(n20505) );
  AOI22_X1 U23399 ( .A1(n20501), .A2(n20812), .B1(n20804), .B2(n20500), .ZN(
        n20487) );
  OAI21_X1 U23400 ( .B1(n20810), .B2(n20480), .A(n20809), .ZN(n20481) );
  AOI21_X1 U23401 ( .B1(n20483), .B2(n20482), .A(n20481), .ZN(n20484) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20502), .B1(
        n20529), .B2(n20694), .ZN(n20486) );
  OAI211_X1 U23403 ( .C1(n20505), .C2(n20697), .A(n20487), .B(n20486), .ZN(
        P1_U3057) );
  AOI22_X1 U23404 ( .A1(n20501), .A2(n20774), .B1(n20817), .B2(n20500), .ZN(
        n20489) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20502), .B1(
        n20529), .B2(n20818), .ZN(n20488) );
  OAI211_X1 U23406 ( .C1(n20505), .C2(n20700), .A(n20489), .B(n20488), .ZN(
        P1_U3058) );
  AOI22_X1 U23407 ( .A1(n20529), .A2(n20824), .B1(n20823), .B2(n20500), .ZN(
        n20491) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20778), .ZN(n20490) );
  OAI211_X1 U23409 ( .C1(n20505), .C2(n20703), .A(n20491), .B(n20490), .ZN(
        P1_U3059) );
  AOI22_X1 U23410 ( .A1(n20529), .A2(n20704), .B1(n20829), .B2(n20500), .ZN(
        n20493) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n9792), .ZN(n20492) );
  OAI211_X1 U23412 ( .C1(n20505), .C2(n20707), .A(n20493), .B(n20492), .ZN(
        P1_U3060) );
  AOI22_X1 U23413 ( .A1(n20501), .A2(n9794), .B1(n20835), .B2(n20500), .ZN(
        n20495) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20502), .B1(
        n20529), .B2(n20708), .ZN(n20494) );
  OAI211_X1 U23415 ( .C1(n20505), .C2(n20711), .A(n20495), .B(n20494), .ZN(
        P1_U3061) );
  AOI22_X1 U23416 ( .A1(n20529), .A2(n20842), .B1(n20840), .B2(n20500), .ZN(
        n20497) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n20786), .ZN(n20496) );
  OAI211_X1 U23418 ( .C1(n20505), .C2(n20714), .A(n20497), .B(n20496), .ZN(
        P1_U3062) );
  AOI22_X1 U23419 ( .A1(n20529), .A2(n20715), .B1(n20848), .B2(n20500), .ZN(
        n20499) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20502), .B1(
        n20501), .B2(n9790), .ZN(n20498) );
  OAI211_X1 U23421 ( .C1(n20505), .C2(n20718), .A(n20499), .B(n20498), .ZN(
        P1_U3063) );
  AOI22_X1 U23422 ( .A1(n20501), .A2(n20858), .B1(n20857), .B2(n20500), .ZN(
        n20504) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20502), .B1(
        n20529), .B2(n20721), .ZN(n20503) );
  OAI211_X1 U23424 ( .C1(n20505), .C2(n20725), .A(n20504), .B(n20503), .ZN(
        P1_U3064) );
  NOR3_X1 U23425 ( .A1(n12290), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20537) );
  INV_X1 U23426 ( .A(n20537), .ZN(n20533) );
  NOR2_X1 U23427 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20533), .ZN(
        n20528) );
  NAND3_X1 U23428 ( .A1(n20589), .A2(n20810), .A3(n20619), .ZN(n20507) );
  OAI21_X1 U23429 ( .B1(n20766), .B2(n20508), .A(n20507), .ZN(n20527) );
  AOI22_X1 U23430 ( .A1(n20804), .A2(n20528), .B1(n20803), .B2(n20527), .ZN(
        n20514) );
  INV_X1 U23431 ( .A(n20529), .ZN(n20509) );
  AOI21_X1 U23432 ( .B1(n20509), .B2(n20557), .A(n21022), .ZN(n20510) );
  AOI21_X1 U23433 ( .B1(n20589), .B2(n20619), .A(n20510), .ZN(n20511) );
  NOR2_X1 U23434 ( .A1(n20511), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20512) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20812), .ZN(n20513) );
  OAI211_X1 U23436 ( .C1(n20815), .C2(n20557), .A(n20514), .B(n20513), .ZN(
        P1_U3065) );
  AOI22_X1 U23437 ( .A1(n20817), .A2(n20528), .B1(n20816), .B2(n20527), .ZN(
        n20516) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20774), .ZN(n20515) );
  OAI211_X1 U23439 ( .C1(n20777), .C2(n20557), .A(n20516), .B(n20515), .ZN(
        P1_U3066) );
  AOI22_X1 U23440 ( .A1(n20823), .A2(n20528), .B1(n20822), .B2(n20527), .ZN(
        n20518) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20778), .ZN(n20517) );
  OAI211_X1 U23442 ( .C1(n20781), .C2(n20557), .A(n20518), .B(n20517), .ZN(
        P1_U3067) );
  AOI22_X1 U23443 ( .A1(n20829), .A2(n20528), .B1(n20828), .B2(n20527), .ZN(
        n20520) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n9792), .ZN(n20519) );
  OAI211_X1 U23445 ( .C1(n20833), .C2(n20557), .A(n20520), .B(n20519), .ZN(
        P1_U3068) );
  AOI22_X1 U23446 ( .A1(n20835), .A2(n20528), .B1(n20834), .B2(n20527), .ZN(
        n20522) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n9794), .ZN(n20521) );
  OAI211_X1 U23448 ( .C1(n20839), .C2(n20557), .A(n20522), .B(n20521), .ZN(
        P1_U3069) );
  AOI22_X1 U23449 ( .A1(n20841), .A2(n20527), .B1(n20840), .B2(n20528), .ZN(
        n20524) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20786), .ZN(n20523) );
  OAI211_X1 U23451 ( .C1(n20789), .C2(n20557), .A(n20524), .B(n20523), .ZN(
        P1_U3070) );
  AOI22_X1 U23452 ( .A1(n20849), .A2(n20527), .B1(n20848), .B2(n20528), .ZN(
        n20526) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n9790), .ZN(n20525) );
  OAI211_X1 U23454 ( .C1(n20853), .C2(n20557), .A(n20526), .B(n20525), .ZN(
        P1_U3071) );
  AOI22_X1 U23455 ( .A1(n20857), .A2(n20528), .B1(n20855), .B2(n20527), .ZN(
        n20532) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20530), .B1(
        n20529), .B2(n20858), .ZN(n20531) );
  OAI211_X1 U23457 ( .C1(n20864), .C2(n20557), .A(n20532), .B(n20531), .ZN(
        P1_U3072) );
  NOR2_X1 U23458 ( .A1(n20647), .A2(n20533), .ZN(n20553) );
  AOI21_X1 U23459 ( .B1(n20589), .B2(n20648), .A(n20553), .ZN(n20534) );
  OAI22_X1 U23460 ( .A1(n20534), .A2(n20802), .B1(n20533), .B2(n11760), .ZN(
        n20552) );
  AOI22_X1 U23461 ( .A1(n20804), .A2(n20553), .B1(n20552), .B2(n20803), .ZN(
        n20539) );
  INV_X1 U23462 ( .A(n20681), .ZN(n20535) );
  OAI21_X1 U23463 ( .B1(n20587), .B2(n20535), .A(n20534), .ZN(n20536) );
  OAI211_X1 U23464 ( .C1(n20677), .C2(n20537), .A(n20809), .B(n20536), .ZN(
        n20554) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20694), .ZN(n20538) );
  OAI211_X1 U23466 ( .C1(n20657), .C2(n20557), .A(n20539), .B(n20538), .ZN(
        P1_U3073) );
  AOI22_X1 U23467 ( .A1(n20817), .A2(n20553), .B1(n20552), .B2(n20816), .ZN(
        n20541) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20818), .ZN(n20540) );
  OAI211_X1 U23469 ( .C1(n20821), .C2(n20557), .A(n20541), .B(n20540), .ZN(
        P1_U3074) );
  AOI22_X1 U23470 ( .A1(n20823), .A2(n20553), .B1(n20822), .B2(n20552), .ZN(
        n20543) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20824), .ZN(n20542) );
  OAI211_X1 U23472 ( .C1(n20827), .C2(n20557), .A(n20543), .B(n20542), .ZN(
        P1_U3075) );
  AOI22_X1 U23473 ( .A1(n20829), .A2(n20553), .B1(n20828), .B2(n20552), .ZN(
        n20545) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20704), .ZN(n20544) );
  OAI211_X1 U23475 ( .C1(n9791), .C2(n20557), .A(n20545), .B(n20544), .ZN(
        P1_U3076) );
  AOI22_X1 U23476 ( .A1(n20835), .A2(n20553), .B1(n20834), .B2(n20552), .ZN(
        n20547) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20708), .ZN(n20546) );
  OAI211_X1 U23478 ( .C1(n9793), .C2(n20557), .A(n20547), .B(n20546), .ZN(
        P1_U3077) );
  AOI22_X1 U23479 ( .A1(n20841), .A2(n20552), .B1(n20840), .B2(n20553), .ZN(
        n20549) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20842), .ZN(n20548) );
  OAI211_X1 U23481 ( .C1(n20847), .C2(n20557), .A(n20549), .B(n20548), .ZN(
        P1_U3078) );
  AOI22_X1 U23482 ( .A1(n20849), .A2(n20552), .B1(n20848), .B2(n20553), .ZN(
        n20551) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20715), .ZN(n20550) );
  OAI211_X1 U23484 ( .C1(n9789), .C2(n20557), .A(n20551), .B(n20550), .ZN(
        P1_U3079) );
  AOI22_X1 U23485 ( .A1(n20857), .A2(n20553), .B1(n20855), .B2(n20552), .ZN(
        n20556) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20554), .B1(
        n20581), .B2(n20721), .ZN(n20555) );
  OAI211_X1 U23487 ( .C1(n20676), .C2(n20557), .A(n20556), .B(n20555), .ZN(
        P1_U3080) );
  INV_X1 U23488 ( .A(n20581), .ZN(n20558) );
  NAND2_X1 U23489 ( .A1(n20558), .A2(n20810), .ZN(n20559) );
  OAI21_X1 U23490 ( .B1(n20559), .B2(n20612), .A(n20681), .ZN(n20564) );
  AND2_X1 U23491 ( .A1(n20589), .A2(n11751), .ZN(n20561) );
  NOR2_X1 U23492 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20590), .ZN(
        n20580) );
  AOI22_X1 U23493 ( .A1(n20581), .A2(n20812), .B1(n20804), .B2(n20580), .ZN(
        n20567) );
  INV_X1 U23494 ( .A(n20561), .ZN(n20563) );
  AOI21_X1 U23495 ( .B1(n20564), .B2(n20563), .A(n20562), .ZN(n20565) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20582), .B1(
        n20612), .B2(n20694), .ZN(n20566) );
  OAI211_X1 U23497 ( .C1(n20585), .C2(n20697), .A(n20567), .B(n20566), .ZN(
        P1_U3081) );
  AOI22_X1 U23498 ( .A1(n20612), .A2(n20818), .B1(n20817), .B2(n20580), .ZN(
        n20569) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20774), .ZN(n20568) );
  OAI211_X1 U23500 ( .C1(n20585), .C2(n20700), .A(n20569), .B(n20568), .ZN(
        P1_U3082) );
  AOI22_X1 U23501 ( .A1(n20581), .A2(n20778), .B1(n20823), .B2(n20580), .ZN(
        n20571) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20582), .B1(
        n20612), .B2(n20824), .ZN(n20570) );
  OAI211_X1 U23503 ( .C1(n20585), .C2(n20703), .A(n20571), .B(n20570), .ZN(
        P1_U3083) );
  AOI22_X1 U23504 ( .A1(n20581), .A2(n9792), .B1(n20829), .B2(n20580), .ZN(
        n20573) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20582), .B1(
        n20612), .B2(n20704), .ZN(n20572) );
  OAI211_X1 U23506 ( .C1(n20585), .C2(n20707), .A(n20573), .B(n20572), .ZN(
        P1_U3084) );
  AOI22_X1 U23507 ( .A1(n20581), .A2(n9794), .B1(n20835), .B2(n20580), .ZN(
        n20575) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20582), .B1(
        n20612), .B2(n20708), .ZN(n20574) );
  OAI211_X1 U23509 ( .C1(n20585), .C2(n20711), .A(n20575), .B(n20574), .ZN(
        P1_U3085) );
  AOI22_X1 U23510 ( .A1(n20612), .A2(n20842), .B1(n20840), .B2(n20580), .ZN(
        n20577) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20786), .ZN(n20576) );
  OAI211_X1 U23512 ( .C1(n20585), .C2(n20714), .A(n20577), .B(n20576), .ZN(
        P1_U3086) );
  AOI22_X1 U23513 ( .A1(n20612), .A2(n20715), .B1(n20848), .B2(n20580), .ZN(
        n20579) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n9790), .ZN(n20578) );
  OAI211_X1 U23515 ( .C1(n20585), .C2(n20718), .A(n20579), .B(n20578), .ZN(
        P1_U3087) );
  AOI22_X1 U23516 ( .A1(n20581), .A2(n20858), .B1(n20857), .B2(n20580), .ZN(
        n20584) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20582), .B1(
        n20612), .B2(n20721), .ZN(n20583) );
  OAI211_X1 U23518 ( .C1(n20585), .C2(n20725), .A(n20584), .B(n20583), .ZN(
        P1_U3088) );
  INV_X1 U23519 ( .A(n20588), .ZN(n20611) );
  AOI21_X1 U23520 ( .B1(n20589), .B2(n20799), .A(n20611), .ZN(n20592) );
  OAI22_X1 U23521 ( .A1(n20592), .A2(n20802), .B1(n20590), .B2(n11760), .ZN(
        n20610) );
  AOI22_X1 U23522 ( .A1(n20804), .A2(n20611), .B1(n20610), .B2(n20803), .ZN(
        n20597) );
  INV_X1 U23523 ( .A(n20591), .ZN(n20593) );
  NAND2_X1 U23524 ( .A1(n20593), .A2(n20592), .ZN(n20594) );
  OAI221_X1 U23525 ( .B1(n20810), .B2(n20595), .C1(n20802), .C2(n20594), .A(
        n20809), .ZN(n20613) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20812), .ZN(n20596) );
  OAI211_X1 U23527 ( .C1(n20815), .C2(n20622), .A(n20597), .B(n20596), .ZN(
        P1_U3089) );
  AOI22_X1 U23528 ( .A1(n20817), .A2(n20611), .B1(n20610), .B2(n20816), .ZN(
        n20599) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20774), .ZN(n20598) );
  OAI211_X1 U23530 ( .C1(n20777), .C2(n20622), .A(n20599), .B(n20598), .ZN(
        P1_U3090) );
  AOI22_X1 U23531 ( .A1(n20823), .A2(n20611), .B1(n20822), .B2(n20610), .ZN(
        n20601) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20778), .ZN(n20600) );
  OAI211_X1 U23533 ( .C1(n20781), .C2(n20622), .A(n20601), .B(n20600), .ZN(
        P1_U3091) );
  AOI22_X1 U23534 ( .A1(n20829), .A2(n20611), .B1(n20828), .B2(n20610), .ZN(
        n20603) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n9792), .ZN(n20602) );
  OAI211_X1 U23536 ( .C1(n20833), .C2(n20622), .A(n20603), .B(n20602), .ZN(
        P1_U3092) );
  AOI22_X1 U23537 ( .A1(n20835), .A2(n20611), .B1(n20834), .B2(n20610), .ZN(
        n20605) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n9794), .ZN(n20604) );
  OAI211_X1 U23539 ( .C1(n20839), .C2(n20622), .A(n20605), .B(n20604), .ZN(
        P1_U3093) );
  AOI22_X1 U23540 ( .A1(n20841), .A2(n20610), .B1(n20840), .B2(n20611), .ZN(
        n20607) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20786), .ZN(n20606) );
  OAI211_X1 U23542 ( .C1(n20789), .C2(n20622), .A(n20607), .B(n20606), .ZN(
        P1_U3094) );
  AOI22_X1 U23543 ( .A1(n20849), .A2(n20610), .B1(n20848), .B2(n20611), .ZN(
        n20609) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n9790), .ZN(n20608) );
  OAI211_X1 U23545 ( .C1(n20853), .C2(n20622), .A(n20609), .B(n20608), .ZN(
        P1_U3095) );
  AOI22_X1 U23546 ( .A1(n20857), .A2(n20611), .B1(n20855), .B2(n20610), .ZN(
        n20615) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20613), .B1(
        n20612), .B2(n20858), .ZN(n20614) );
  OAI211_X1 U23548 ( .C1(n20864), .C2(n20622), .A(n20615), .B(n20614), .ZN(
        P1_U3096) );
  INV_X1 U23549 ( .A(n20616), .ZN(n20617) );
  AND2_X1 U23550 ( .A1(n20618), .A2(n9689), .ZN(n20729) );
  NOR3_X1 U23551 ( .A1(n20727), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20652) );
  INV_X1 U23552 ( .A(n20652), .ZN(n20649) );
  NOR2_X1 U23553 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20649), .ZN(
        n20642) );
  AOI21_X1 U23554 ( .B1(n20729), .B2(n20619), .A(n20642), .ZN(n20624) );
  OAI22_X1 U23555 ( .A1(n20624), .A2(n20802), .B1(n20621), .B2(n20620), .ZN(
        n20641) );
  AOI22_X1 U23556 ( .A1(n20641), .A2(n20803), .B1(n20804), .B2(n20642), .ZN(
        n20628) );
  INV_X1 U23557 ( .A(n20675), .ZN(n20623) );
  OAI21_X1 U23558 ( .B1(n20623), .B2(n20643), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20625) );
  NAND2_X1 U23559 ( .A1(n20625), .A2(n20624), .ZN(n20626) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20812), .ZN(n20627) );
  OAI211_X1 U23561 ( .C1(n20815), .C2(n20675), .A(n20628), .B(n20627), .ZN(
        P1_U3097) );
  AOI22_X1 U23562 ( .A1(n20641), .A2(n20816), .B1(n20817), .B2(n20642), .ZN(
        n20630) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20774), .ZN(n20629) );
  OAI211_X1 U23564 ( .C1(n20777), .C2(n20675), .A(n20630), .B(n20629), .ZN(
        P1_U3098) );
  AOI22_X1 U23565 ( .A1(n20823), .A2(n20642), .B1(n20641), .B2(n20822), .ZN(
        n20632) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20778), .ZN(n20631) );
  OAI211_X1 U23567 ( .C1(n20781), .C2(n20675), .A(n20632), .B(n20631), .ZN(
        P1_U3099) );
  AOI22_X1 U23568 ( .A1(n20829), .A2(n20642), .B1(n20641), .B2(n20828), .ZN(
        n20634) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n9792), .ZN(n20633) );
  OAI211_X1 U23570 ( .C1(n20833), .C2(n20675), .A(n20634), .B(n20633), .ZN(
        P1_U3100) );
  AOI22_X1 U23571 ( .A1(n20835), .A2(n20642), .B1(n20641), .B2(n20834), .ZN(
        n20636) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n9794), .ZN(n20635) );
  OAI211_X1 U23573 ( .C1(n20839), .C2(n20675), .A(n20636), .B(n20635), .ZN(
        P1_U3101) );
  AOI22_X1 U23574 ( .A1(n20641), .A2(n20841), .B1(n20840), .B2(n20642), .ZN(
        n20638) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20786), .ZN(n20637) );
  OAI211_X1 U23576 ( .C1(n20789), .C2(n20675), .A(n20638), .B(n20637), .ZN(
        P1_U3102) );
  AOI22_X1 U23577 ( .A1(n20641), .A2(n20849), .B1(n20848), .B2(n20642), .ZN(
        n20640) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n9790), .ZN(n20639) );
  OAI211_X1 U23579 ( .C1(n20853), .C2(n20675), .A(n20640), .B(n20639), .ZN(
        P1_U3103) );
  AOI22_X1 U23580 ( .A1(n20857), .A2(n20642), .B1(n20641), .B2(n20855), .ZN(
        n20646) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20644), .B1(
        n20643), .B2(n20858), .ZN(n20645) );
  OAI211_X1 U23582 ( .C1(n20864), .C2(n20675), .A(n20646), .B(n20645), .ZN(
        P1_U3104) );
  NOR2_X1 U23583 ( .A1(n20647), .A2(n20649), .ZN(n20671) );
  AOI21_X1 U23584 ( .B1(n20729), .B2(n20648), .A(n20671), .ZN(n20650) );
  OAI22_X1 U23585 ( .A1(n20650), .A2(n20802), .B1(n20649), .B2(n11760), .ZN(
        n20670) );
  AOI22_X1 U23586 ( .A1(n20670), .A2(n20803), .B1(n20804), .B2(n20671), .ZN(
        n20656) );
  INV_X1 U23587 ( .A(n20680), .ZN(n20732) );
  OAI211_X1 U23588 ( .C1(n20732), .C2(n21022), .A(n20810), .B(n20650), .ZN(
        n20651) );
  OAI211_X1 U23589 ( .C1(n20810), .C2(n20652), .A(n20809), .B(n20651), .ZN(
        n20672) );
  INV_X1 U23590 ( .A(n20653), .ZN(n20654) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20694), .ZN(n20655) );
  OAI211_X1 U23592 ( .C1(n20657), .C2(n20675), .A(n20656), .B(n20655), .ZN(
        P1_U3105) );
  AOI22_X1 U23593 ( .A1(n20670), .A2(n20816), .B1(n20817), .B2(n20671), .ZN(
        n20659) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20818), .ZN(n20658) );
  OAI211_X1 U23595 ( .C1(n20821), .C2(n20675), .A(n20659), .B(n20658), .ZN(
        P1_U3106) );
  AOI22_X1 U23596 ( .A1(n20823), .A2(n20671), .B1(n20670), .B2(n20822), .ZN(
        n20661) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20824), .ZN(n20660) );
  OAI211_X1 U23598 ( .C1(n20827), .C2(n20675), .A(n20661), .B(n20660), .ZN(
        P1_U3107) );
  AOI22_X1 U23599 ( .A1(n20829), .A2(n20671), .B1(n20670), .B2(n20828), .ZN(
        n20663) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20704), .ZN(n20662) );
  OAI211_X1 U23601 ( .C1(n9791), .C2(n20675), .A(n20663), .B(n20662), .ZN(
        P1_U3108) );
  AOI22_X1 U23602 ( .A1(n20835), .A2(n20671), .B1(n20670), .B2(n20834), .ZN(
        n20665) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20708), .ZN(n20664) );
  OAI211_X1 U23604 ( .C1(n9793), .C2(n20675), .A(n20665), .B(n20664), .ZN(
        P1_U3109) );
  AOI22_X1 U23605 ( .A1(n20670), .A2(n20841), .B1(n20840), .B2(n20671), .ZN(
        n20667) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20842), .ZN(n20666) );
  OAI211_X1 U23607 ( .C1(n20847), .C2(n20675), .A(n20667), .B(n20666), .ZN(
        P1_U3110) );
  AOI22_X1 U23608 ( .A1(n20670), .A2(n20849), .B1(n20848), .B2(n20671), .ZN(
        n20669) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20715), .ZN(n20668) );
  OAI211_X1 U23610 ( .C1(n9789), .C2(n20675), .A(n20669), .B(n20668), .ZN(
        P1_U3111) );
  AOI22_X1 U23611 ( .A1(n20857), .A2(n20671), .B1(n20670), .B2(n20855), .ZN(
        n20674) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20672), .B1(
        n20720), .B2(n20721), .ZN(n20673) );
  OAI211_X1 U23613 ( .C1(n20676), .C2(n20675), .A(n20674), .B(n20673), .ZN(
        P1_U3112) );
  INV_X1 U23614 ( .A(n20720), .ZN(n20678) );
  NAND2_X1 U23615 ( .A1(n20678), .A2(n20677), .ZN(n20682) );
  INV_X1 U23616 ( .A(n20764), .ZN(n20679) );
  OAI21_X1 U23617 ( .B1(n20682), .B2(n20751), .A(n20681), .ZN(n20692) );
  AND2_X1 U23618 ( .A1(n20729), .A2(n11751), .ZN(n20687) );
  OR2_X1 U23619 ( .A1(n20683), .A2(n20727), .ZN(n20765) );
  INV_X1 U23620 ( .A(n20765), .ZN(n20684) );
  NOR3_X1 U23621 ( .A1(n20727), .A2(n20686), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20734) );
  INV_X1 U23622 ( .A(n20734), .ZN(n20730) );
  NOR2_X1 U23623 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20730), .ZN(
        n20719) );
  AOI22_X1 U23624 ( .A1(n20720), .A2(n20812), .B1(n20804), .B2(n20719), .ZN(
        n20696) );
  INV_X1 U23625 ( .A(n20687), .ZN(n20691) );
  NAND2_X1 U23626 ( .A1(n20765), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20770) );
  OAI211_X1 U23627 ( .C1(n20689), .C2(n20719), .A(n20770), .B(n20688), .ZN(
        n20690) );
  AOI21_X1 U23628 ( .B1(n20692), .B2(n20691), .A(n20690), .ZN(n20693) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20722), .B1(
        n20751), .B2(n20694), .ZN(n20695) );
  OAI211_X1 U23630 ( .C1(n20726), .C2(n20697), .A(n20696), .B(n20695), .ZN(
        P1_U3113) );
  AOI22_X1 U23631 ( .A1(n20751), .A2(n20818), .B1(n20817), .B2(n20719), .ZN(
        n20699) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20722), .B1(
        n20720), .B2(n20774), .ZN(n20698) );
  OAI211_X1 U23633 ( .C1(n20726), .C2(n20700), .A(n20699), .B(n20698), .ZN(
        P1_U3114) );
  AOI22_X1 U23634 ( .A1(n20751), .A2(n20824), .B1(n20823), .B2(n20719), .ZN(
        n20702) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20722), .B1(
        n20720), .B2(n20778), .ZN(n20701) );
  OAI211_X1 U23636 ( .C1(n20726), .C2(n20703), .A(n20702), .B(n20701), .ZN(
        P1_U3115) );
  AOI22_X1 U23637 ( .A1(n20720), .A2(n9792), .B1(n20829), .B2(n20719), .ZN(
        n20706) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20722), .B1(
        n20751), .B2(n20704), .ZN(n20705) );
  OAI211_X1 U23639 ( .C1(n20726), .C2(n20707), .A(n20706), .B(n20705), .ZN(
        P1_U3116) );
  AOI22_X1 U23640 ( .A1(n20720), .A2(n9794), .B1(n20835), .B2(n20719), .ZN(
        n20710) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20722), .B1(
        n20751), .B2(n20708), .ZN(n20709) );
  OAI211_X1 U23642 ( .C1(n20726), .C2(n20711), .A(n20710), .B(n20709), .ZN(
        P1_U3117) );
  AOI22_X1 U23643 ( .A1(n20751), .A2(n20842), .B1(n20840), .B2(n20719), .ZN(
        n20713) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20722), .B1(
        n20720), .B2(n20786), .ZN(n20712) );
  OAI211_X1 U23645 ( .C1(n20726), .C2(n20714), .A(n20713), .B(n20712), .ZN(
        P1_U3118) );
  AOI22_X1 U23646 ( .A1(n20751), .A2(n20715), .B1(n20848), .B2(n20719), .ZN(
        n20717) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20722), .B1(
        n20720), .B2(n9790), .ZN(n20716) );
  OAI211_X1 U23648 ( .C1(n20726), .C2(n20718), .A(n20717), .B(n20716), .ZN(
        P1_U3119) );
  AOI22_X1 U23649 ( .A1(n20720), .A2(n20858), .B1(n20857), .B2(n20719), .ZN(
        n20724) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20722), .B1(
        n20751), .B2(n20721), .ZN(n20723) );
  OAI211_X1 U23651 ( .C1(n20726), .C2(n20725), .A(n20724), .B(n20723), .ZN(
        P1_U3120) );
  NOR2_X1 U23652 ( .A1(n20728), .A2(n20727), .ZN(n20750) );
  AOI21_X1 U23653 ( .B1(n20729), .B2(n20799), .A(n20750), .ZN(n20731) );
  OAI22_X1 U23654 ( .A1(n20731), .A2(n20802), .B1(n20730), .B2(n11760), .ZN(
        n20749) );
  AOI22_X1 U23655 ( .A1(n20749), .A2(n20803), .B1(n20804), .B2(n20750), .ZN(
        n20736) );
  OAI211_X1 U23656 ( .C1(n20732), .C2(n20806), .A(n20810), .B(n20731), .ZN(
        n20733) );
  OAI211_X1 U23657 ( .C1(n20810), .C2(n20734), .A(n20809), .B(n20733), .ZN(
        n20752) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20812), .ZN(n20735) );
  OAI211_X1 U23659 ( .C1(n20815), .C2(n20763), .A(n20736), .B(n20735), .ZN(
        P1_U3121) );
  AOI22_X1 U23660 ( .A1(n20749), .A2(n20816), .B1(n20817), .B2(n20750), .ZN(
        n20738) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20774), .ZN(n20737) );
  OAI211_X1 U23662 ( .C1(n20777), .C2(n20763), .A(n20738), .B(n20737), .ZN(
        P1_U3122) );
  AOI22_X1 U23663 ( .A1(n20823), .A2(n20750), .B1(n20749), .B2(n20822), .ZN(
        n20740) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20778), .ZN(n20739) );
  OAI211_X1 U23665 ( .C1(n20781), .C2(n20763), .A(n20740), .B(n20739), .ZN(
        P1_U3123) );
  AOI22_X1 U23666 ( .A1(n20829), .A2(n20750), .B1(n20749), .B2(n20828), .ZN(
        n20742) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n9792), .ZN(n20741) );
  OAI211_X1 U23668 ( .C1(n20833), .C2(n20763), .A(n20742), .B(n20741), .ZN(
        P1_U3124) );
  AOI22_X1 U23669 ( .A1(n20835), .A2(n20750), .B1(n20749), .B2(n20834), .ZN(
        n20744) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n9794), .ZN(n20743) );
  OAI211_X1 U23671 ( .C1(n20839), .C2(n20763), .A(n20744), .B(n20743), .ZN(
        P1_U3125) );
  AOI22_X1 U23672 ( .A1(n20749), .A2(n20841), .B1(n20840), .B2(n20750), .ZN(
        n20746) );
  AOI22_X1 U23673 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20786), .ZN(n20745) );
  OAI211_X1 U23674 ( .C1(n20789), .C2(n20763), .A(n20746), .B(n20745), .ZN(
        P1_U3126) );
  AOI22_X1 U23675 ( .A1(n20749), .A2(n20849), .B1(n20848), .B2(n20750), .ZN(
        n20748) );
  AOI22_X1 U23676 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n9790), .ZN(n20747) );
  OAI211_X1 U23677 ( .C1(n20853), .C2(n20763), .A(n20748), .B(n20747), .ZN(
        P1_U3127) );
  AOI22_X1 U23678 ( .A1(n20857), .A2(n20750), .B1(n20749), .B2(n20855), .ZN(
        n20754) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20752), .B1(
        n20751), .B2(n20858), .ZN(n20753) );
  OAI211_X1 U23680 ( .C1(n20864), .C2(n20763), .A(n20754), .B(n20753), .ZN(
        P1_U3128) );
  AOI22_X1 U23681 ( .A1(n20758), .A2(n20824), .B1(n20823), .B2(n20757), .ZN(
        n20756) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20760), .B1(
        n20822), .B2(n20759), .ZN(n20755) );
  OAI211_X1 U23683 ( .C1(n20827), .C2(n20763), .A(n20756), .B(n20755), .ZN(
        P1_U3131) );
  AOI22_X1 U23684 ( .A1(n20758), .A2(n20842), .B1(n20757), .B2(n20840), .ZN(
        n20762) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20760), .B1(
        n20841), .B2(n20759), .ZN(n20761) );
  OAI211_X1 U23686 ( .C1(n20847), .C2(n20763), .A(n20762), .B(n20761), .ZN(
        P1_U3134) );
  INV_X1 U23687 ( .A(n20811), .ZN(n20801) );
  NOR2_X1 U23688 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20801), .ZN(
        n20793) );
  NAND2_X1 U23689 ( .A1(n20800), .A2(n11751), .ZN(n20767) );
  OAI22_X1 U23690 ( .A1(n20767), .A2(n20802), .B1(n20766), .B2(n20765), .ZN(
        n20792) );
  AOI22_X1 U23691 ( .A1(n20804), .A2(n20793), .B1(n20803), .B2(n20792), .ZN(
        n20773) );
  OAI21_X1 U23692 ( .B1(n20859), .B2(n20794), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20768) );
  AOI21_X1 U23693 ( .B1(n20768), .B2(n20767), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20771) );
  AOI22_X1 U23694 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n20812), .B2(n20794), .ZN(n20772) );
  OAI211_X1 U23695 ( .C1(n20815), .C2(n20846), .A(n20773), .B(n20772), .ZN(
        P1_U3145) );
  AOI22_X1 U23696 ( .A1(n20817), .A2(n20793), .B1(n20816), .B2(n20792), .ZN(
        n20776) );
  AOI22_X1 U23697 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20774), .B2(n20794), .ZN(n20775) );
  OAI211_X1 U23698 ( .C1(n20777), .C2(n20846), .A(n20776), .B(n20775), .ZN(
        P1_U3146) );
  AOI22_X1 U23699 ( .A1(n20823), .A2(n20793), .B1(n20822), .B2(n20792), .ZN(
        n20780) );
  AOI22_X1 U23700 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20778), .B2(n20794), .ZN(n20779) );
  OAI211_X1 U23701 ( .C1(n20781), .C2(n20846), .A(n20780), .B(n20779), .ZN(
        P1_U3147) );
  AOI22_X1 U23702 ( .A1(n20829), .A2(n20793), .B1(n20828), .B2(n20792), .ZN(
        n20783) );
  AOI22_X1 U23703 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9792), .B2(n20794), .ZN(n20782) );
  OAI211_X1 U23704 ( .C1(n20833), .C2(n20846), .A(n20783), .B(n20782), .ZN(
        P1_U3148) );
  AOI22_X1 U23705 ( .A1(n20835), .A2(n20793), .B1(n20834), .B2(n20792), .ZN(
        n20785) );
  AOI22_X1 U23706 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9794), .B2(n20794), .ZN(n20784) );
  OAI211_X1 U23707 ( .C1(n20839), .C2(n20846), .A(n20785), .B(n20784), .ZN(
        P1_U3149) );
  AOI22_X1 U23708 ( .A1(n20841), .A2(n20792), .B1(n20840), .B2(n20793), .ZN(
        n20788) );
  AOI22_X1 U23709 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n20794), .B2(n20786), .ZN(n20787) );
  OAI211_X1 U23710 ( .C1(n20789), .C2(n20846), .A(n20788), .B(n20787), .ZN(
        P1_U3150) );
  AOI22_X1 U23711 ( .A1(n20849), .A2(n20792), .B1(n20848), .B2(n20793), .ZN(
        n20791) );
  AOI22_X1 U23712 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9790), .B2(n20794), .ZN(n20790) );
  OAI211_X1 U23713 ( .C1(n20853), .C2(n20846), .A(n20791), .B(n20790), .ZN(
        P1_U3151) );
  AOI22_X1 U23714 ( .A1(n20857), .A2(n20793), .B1(n20855), .B2(n20792), .ZN(
        n20797) );
  AOI22_X1 U23715 ( .A1(n20795), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20858), .B2(n20794), .ZN(n20796) );
  OAI211_X1 U23716 ( .C1(n20864), .C2(n20846), .A(n20797), .B(n20796), .ZN(
        P1_U3152) );
  INV_X1 U23717 ( .A(n20798), .ZN(n20856) );
  AOI21_X1 U23718 ( .B1(n20800), .B2(n20799), .A(n20856), .ZN(n20805) );
  OAI22_X1 U23719 ( .A1(n20805), .A2(n20802), .B1(n20801), .B2(n11760), .ZN(
        n20854) );
  AOI22_X1 U23720 ( .A1(n20804), .A2(n20856), .B1(n20854), .B2(n20803), .ZN(
        n20814) );
  OAI211_X1 U23721 ( .C1(n20807), .C2(n20806), .A(n20810), .B(n20805), .ZN(
        n20808) );
  OAI211_X1 U23722 ( .C1(n20811), .C2(n20810), .A(n20809), .B(n20808), .ZN(
        n20860) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20860), .B1(
        n20859), .B2(n20812), .ZN(n20813) );
  OAI211_X1 U23724 ( .C1(n20815), .C2(n20863), .A(n20814), .B(n20813), .ZN(
        P1_U3153) );
  AOI22_X1 U23725 ( .A1(n20817), .A2(n20856), .B1(n20854), .B2(n20816), .ZN(
        n20820) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20860), .B1(
        n20843), .B2(n20818), .ZN(n20819) );
  OAI211_X1 U23727 ( .C1(n20821), .C2(n20846), .A(n20820), .B(n20819), .ZN(
        P1_U3154) );
  AOI22_X1 U23728 ( .A1(n20823), .A2(n20856), .B1(n20822), .B2(n20854), .ZN(
        n20826) );
  AOI22_X1 U23729 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20860), .B1(
        n20843), .B2(n20824), .ZN(n20825) );
  OAI211_X1 U23730 ( .C1(n20827), .C2(n20846), .A(n20826), .B(n20825), .ZN(
        P1_U3155) );
  AOI22_X1 U23731 ( .A1(n20829), .A2(n20856), .B1(n20828), .B2(n20854), .ZN(
        n20832) );
  AOI22_X1 U23732 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20860), .B1(
        n20859), .B2(n9792), .ZN(n20831) );
  OAI211_X1 U23733 ( .C1(n20833), .C2(n20863), .A(n20832), .B(n20831), .ZN(
        P1_U3156) );
  AOI22_X1 U23734 ( .A1(n20835), .A2(n20856), .B1(n20834), .B2(n20854), .ZN(
        n20838) );
  AOI22_X1 U23735 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20860), .B1(
        n20859), .B2(n9794), .ZN(n20837) );
  OAI211_X1 U23736 ( .C1(n20839), .C2(n20863), .A(n20838), .B(n20837), .ZN(
        P1_U3157) );
  AOI22_X1 U23737 ( .A1(n20841), .A2(n20854), .B1(n20840), .B2(n20856), .ZN(
        n20845) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20860), .B1(
        n20843), .B2(n20842), .ZN(n20844) );
  OAI211_X1 U23739 ( .C1(n20847), .C2(n20846), .A(n20845), .B(n20844), .ZN(
        P1_U3158) );
  AOI22_X1 U23740 ( .A1(n20849), .A2(n20854), .B1(n20848), .B2(n20856), .ZN(
        n20852) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20860), .B1(
        n20859), .B2(n9790), .ZN(n20851) );
  OAI211_X1 U23742 ( .C1(n20853), .C2(n20863), .A(n20852), .B(n20851), .ZN(
        P1_U3159) );
  AOI22_X1 U23743 ( .A1(n20857), .A2(n20856), .B1(n20855), .B2(n20854), .ZN(
        n20862) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20860), .B1(
        n20859), .B2(n20858), .ZN(n20861) );
  OAI211_X1 U23745 ( .C1(n20864), .C2(n20863), .A(n20862), .B(n20861), .ZN(
        P1_U3160) );
  NOR2_X1 U23746 ( .A1(n20865), .A2(n13651), .ZN(n20867) );
  AOI22_X1 U23747 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20867), .B1(n20866), 
        .B2(n11760), .ZN(P1_U3163) );
  AND2_X1 U23748 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20868), .ZN(
        P1_U3164) );
  AND2_X1 U23749 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20868), .ZN(
        P1_U3165) );
  AND2_X1 U23750 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20868), .ZN(
        P1_U3166) );
  AND2_X1 U23751 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20868), .ZN(
        P1_U3167) );
  AND2_X1 U23752 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20868), .ZN(
        P1_U3168) );
  AND2_X1 U23753 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20868), .ZN(
        P1_U3169) );
  AND2_X1 U23754 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20868), .ZN(
        P1_U3170) );
  AND2_X1 U23755 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20868), .ZN(
        P1_U3171) );
  AND2_X1 U23756 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20868), .ZN(
        P1_U3172) );
  AND2_X1 U23757 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20868), .ZN(
        P1_U3173) );
  AND2_X1 U23758 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20868), .ZN(
        P1_U3174) );
  AND2_X1 U23759 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20868), .ZN(
        P1_U3175) );
  AND2_X1 U23760 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20868), .ZN(
        P1_U3176) );
  AND2_X1 U23761 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20868), .ZN(
        P1_U3177) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20868), .ZN(
        P1_U3178) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20868), .ZN(
        P1_U3179) );
  AND2_X1 U23764 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20868), .ZN(
        P1_U3180) );
  AND2_X1 U23765 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20868), .ZN(
        P1_U3181) );
  AND2_X1 U23766 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20868), .ZN(
        P1_U3182) );
  AND2_X1 U23767 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20868), .ZN(
        P1_U3183) );
  AND2_X1 U23768 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20868), .ZN(
        P1_U3184) );
  AND2_X1 U23769 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20868), .ZN(
        P1_U3185) );
  AND2_X1 U23770 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20868), .ZN(P1_U3186) );
  AND2_X1 U23771 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20868), .ZN(P1_U3187) );
  AND2_X1 U23772 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20868), .ZN(P1_U3188) );
  AND2_X1 U23773 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20868), .ZN(P1_U3189) );
  AND2_X1 U23774 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20868), .ZN(P1_U3190) );
  AND2_X1 U23775 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20868), .ZN(P1_U3191) );
  AND2_X1 U23776 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20868), .ZN(P1_U3192) );
  AND2_X1 U23777 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20868), .ZN(P1_U3193) );
  NAND2_X1 U23778 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20883), .ZN(n20873) );
  NOR2_X1 U23779 ( .A1(NA), .A2(n21122), .ZN(n20877) );
  NOR2_X1 U23780 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20869) );
  OAI22_X1 U23781 ( .A1(n20870), .A2(n20877), .B1(n20869), .B2(n21071), .ZN(
        n20871) );
  AOI21_X1 U23782 ( .B1(n20916), .B2(n20871), .A(n20882), .ZN(n20872) );
  OAI21_X1 U23783 ( .B1(n20953), .B2(n20873), .A(n20872), .ZN(P1_U3194) );
  NOR2_X1 U23784 ( .A1(n20874), .A2(n20953), .ZN(n20876) );
  AOI21_X1 U23785 ( .B1(NA), .B2(n20874), .A(P1_STATE_REG_0__SCAN_IN), .ZN(
        n20875) );
  OAI22_X1 U23786 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20877), .B1(n20876), 
        .B2(n20875), .ZN(n20881) );
  NOR3_X1 U23787 ( .A1(NA), .A2(n12994), .A3(n20953), .ZN(n20878) );
  OAI22_X1 U23788 ( .A1(n20879), .A2(n20878), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21122), .ZN(n20880) );
  OAI22_X1 U23789 ( .A1(n20882), .A2(n20881), .B1(n21071), .B2(n20880), .ZN(
        P1_U3196) );
  OR2_X1 U23790 ( .A1(n20929), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20911) );
  INV_X1 U23791 ( .A(n20962), .ZN(n20929) );
  OR2_X1 U23792 ( .A1(n20883), .A2(n20929), .ZN(n20909) );
  AOI222_X1 U23793 ( .A1(n20923), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20924), .ZN(n20884) );
  INV_X1 U23794 ( .A(n20884), .ZN(P1_U3197) );
  AOI222_X1 U23795 ( .A1(n20924), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20923), .ZN(n20885) );
  INV_X1 U23796 ( .A(n20885), .ZN(P1_U3198) );
  OAI222_X1 U23797 ( .A1(n20909), .A2(n20887), .B1(n20886), .B2(n20962), .C1(
        n13957), .C2(n20911), .ZN(P1_U3199) );
  AOI222_X1 U23798 ( .A1(n20924), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20923), .ZN(n20888) );
  INV_X1 U23799 ( .A(n20888), .ZN(P1_U3200) );
  AOI222_X1 U23800 ( .A1(n20924), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20923), .ZN(n20889) );
  INV_X1 U23801 ( .A(n20889), .ZN(P1_U3201) );
  AOI22_X1 U23802 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20923), .ZN(n20890) );
  OAI21_X1 U23803 ( .B1(n20891), .B2(n20909), .A(n20890), .ZN(P1_U3202) );
  AOI22_X1 U23804 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20924), .ZN(n20892) );
  OAI21_X1 U23805 ( .B1(n20894), .B2(n20911), .A(n20892), .ZN(P1_U3203) );
  AOI22_X1 U23806 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20923), .ZN(n20893) );
  OAI21_X1 U23807 ( .B1(n20894), .B2(n20909), .A(n20893), .ZN(P1_U3204) );
  AOI22_X1 U23808 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20924), .ZN(n20895) );
  OAI21_X1 U23809 ( .B1(n20896), .B2(n20911), .A(n20895), .ZN(P1_U3205) );
  AOI222_X1 U23810 ( .A1(n20923), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20924), .ZN(n20897) );
  INV_X1 U23811 ( .A(n20897), .ZN(P1_U3206) );
  AOI22_X1 U23812 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20923), .ZN(n20898) );
  OAI21_X1 U23813 ( .B1(n20899), .B2(n20909), .A(n20898), .ZN(P1_U3207) );
  AOI22_X1 U23814 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20924), .ZN(n20900) );
  OAI21_X1 U23815 ( .B1(n20901), .B2(n20911), .A(n20900), .ZN(P1_U3208) );
  AOI222_X1 U23816 ( .A1(n20924), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20923), .ZN(n20902) );
  INV_X1 U23817 ( .A(n20902), .ZN(P1_U3209) );
  AOI222_X1 U23818 ( .A1(n20924), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20923), .ZN(n20903) );
  INV_X1 U23819 ( .A(n20903), .ZN(P1_U3210) );
  AOI222_X1 U23820 ( .A1(n20923), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20924), .ZN(n20904) );
  INV_X1 U23821 ( .A(n20904), .ZN(P1_U3211) );
  AOI22_X1 U23822 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20923), .ZN(n20905) );
  OAI21_X1 U23823 ( .B1(n20906), .B2(n20909), .A(n20905), .ZN(P1_U3212) );
  AOI22_X1 U23824 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20924), .ZN(n20907) );
  OAI21_X1 U23825 ( .B1(n14761), .B2(n20911), .A(n20907), .ZN(P1_U3213) );
  AOI22_X1 U23826 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20923), .ZN(n20908) );
  OAI21_X1 U23827 ( .B1(n14761), .B2(n20909), .A(n20908), .ZN(P1_U3214) );
  AOI22_X1 U23828 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20929), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20924), .ZN(n20910) );
  OAI21_X1 U23829 ( .B1(n21123), .B2(n20911), .A(n20910), .ZN(P1_U3215) );
  AOI222_X1 U23830 ( .A1(n20924), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20923), .ZN(n20912) );
  INV_X1 U23831 ( .A(n20912), .ZN(P1_U3216) );
  AOI222_X1 U23832 ( .A1(n20924), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20923), .ZN(n20913) );
  INV_X1 U23833 ( .A(n20913), .ZN(P1_U3217) );
  AOI222_X1 U23834 ( .A1(n20924), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20923), .ZN(n20914) );
  INV_X1 U23835 ( .A(n20914), .ZN(P1_U3218) );
  AOI222_X1 U23836 ( .A1(n20923), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20924), .ZN(n20915) );
  INV_X1 U23837 ( .A(n20915), .ZN(P1_U3219) );
  AOI222_X1 U23838 ( .A1(n20924), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20923), .ZN(n20917) );
  INV_X1 U23839 ( .A(n20917), .ZN(P1_U3220) );
  AOI222_X1 U23840 ( .A1(n20924), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20923), .ZN(n20918) );
  INV_X1 U23841 ( .A(n20918), .ZN(P1_U3221) );
  AOI222_X1 U23842 ( .A1(n20923), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20924), .ZN(n20919) );
  INV_X1 U23843 ( .A(n20919), .ZN(P1_U3222) );
  AOI222_X1 U23844 ( .A1(n20923), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20924), .ZN(n20920) );
  INV_X1 U23845 ( .A(n20920), .ZN(P1_U3223) );
  AOI222_X1 U23846 ( .A1(n20923), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20924), .ZN(n20921) );
  INV_X1 U23847 ( .A(n20921), .ZN(P1_U3224) );
  AOI222_X1 U23848 ( .A1(n20923), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20924), .ZN(n20922) );
  INV_X1 U23849 ( .A(n20922), .ZN(P1_U3225) );
  AOI222_X1 U23850 ( .A1(n20924), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20923), .ZN(n20925) );
  INV_X1 U23851 ( .A(n20925), .ZN(P1_U3226) );
  OAI22_X1 U23852 ( .A1(n20916), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20962), .ZN(n20926) );
  INV_X1 U23853 ( .A(n20926), .ZN(P1_U3458) );
  OAI22_X1 U23854 ( .A1(n20916), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20962), .ZN(n20927) );
  INV_X1 U23855 ( .A(n20927), .ZN(P1_U3459) );
  OAI22_X1 U23856 ( .A1(n20929), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20962), .ZN(n20928) );
  INV_X1 U23857 ( .A(n20928), .ZN(P1_U3460) );
  OAI22_X1 U23858 ( .A1(n20929), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20962), .ZN(n20930) );
  INV_X1 U23859 ( .A(n20930), .ZN(P1_U3461) );
  OAI21_X1 U23860 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20934), .A(n20932), 
        .ZN(n20931) );
  INV_X1 U23861 ( .A(n20931), .ZN(P1_U3464) );
  OAI21_X1 U23862 ( .B1(n20934), .B2(n20933), .A(n20932), .ZN(P1_U3465) );
  AOI22_X1 U23863 ( .A1(n20938), .A2(n20937), .B1(n20936), .B2(n20935), .ZN(
        n20939) );
  INV_X1 U23864 ( .A(n20939), .ZN(n20941) );
  MUX2_X1 U23865 ( .A(n20941), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20940), .Z(P1_U3469) );
  AOI21_X1 U23866 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20942) );
  OAI22_X1 U23867 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n13825), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n20942), .ZN(n20943) );
  INV_X1 U23868 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20970) );
  AOI22_X1 U23869 ( .A1(n20946), .A2(n20943), .B1(n20970), .B2(n20944), .ZN(
        P1_U3481) );
  NOR2_X1 U23870 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20945) );
  INV_X1 U23871 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21062) );
  AOI22_X1 U23872 ( .A1(n20946), .A2(n20945), .B1(n21062), .B2(n20944), .ZN(
        P1_U3482) );
  AOI22_X1 U23873 ( .A1(n20962), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21068), 
        .B2(n20916), .ZN(P1_U3483) );
  NOR2_X1 U23874 ( .A1(n20948), .A2(n11760), .ZN(n20951) );
  AOI211_X1 U23875 ( .C1(n20952), .C2(n20951), .A(n20950), .B(n20949), .ZN(
        n20961) );
  AOI21_X1 U23876 ( .B1(n20954), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n11643), 
        .ZN(n20957) );
  OAI211_X1 U23877 ( .C1(n20955), .C2(n20954), .A(P1_STATE2_REG_2__SCAN_IN), 
        .B(n20953), .ZN(n20956) );
  OAI21_X1 U23878 ( .B1(n20957), .B2(n20956), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n20960) );
  NOR2_X1 U23879 ( .A1(n20961), .A2(n20958), .ZN(n20959) );
  AOI22_X1 U23880 ( .A1(n21122), .A2(n20961), .B1(n20960), .B2(n20959), .ZN(
        P1_U3485) );
  OAI22_X1 U23881 ( .A1(n20929), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20962), .ZN(n20963) );
  INV_X1 U23882 ( .A(n20963), .ZN(P1_U3486) );
  AOI22_X1 U23883 ( .A1(n16702), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16704), .ZN(n21162) );
  INV_X1 U23884 ( .A(READY1), .ZN(n20966) );
  AOI22_X1 U23885 ( .A1(n20966), .A2(keyinput_g36), .B1(keyinput_g8), .B2(
        n20965), .ZN(n20964) );
  OAI221_X1 U23886 ( .B1(n20966), .B2(keyinput_g36), .C1(n20965), .C2(
        keyinput_g8), .A(n20964), .ZN(n20977) );
  AOI22_X1 U23887 ( .A1(n20968), .A2(keyinput_g58), .B1(keyinput_g49), .B2(
        n21081), .ZN(n20967) );
  OAI221_X1 U23888 ( .B1(n20968), .B2(keyinput_g58), .C1(n21081), .C2(
        keyinput_g49), .A(n20967), .ZN(n20976) );
  AOI22_X1 U23889 ( .A1(n21122), .A2(keyinput_g43), .B1(keyinput_g50), .B2(
        n20970), .ZN(n20969) );
  OAI221_X1 U23890 ( .B1(n21122), .B2(keyinput_g43), .C1(n20970), .C2(
        keyinput_g50), .A(n20969), .ZN(n20975) );
  INV_X1 U23891 ( .A(DATAI_2_), .ZN(n20973) );
  AOI22_X1 U23892 ( .A1(n20973), .A2(keyinput_g30), .B1(n20972), .B2(
        keyinput_g12), .ZN(n20971) );
  OAI221_X1 U23893 ( .B1(n20973), .B2(keyinput_g30), .C1(n20972), .C2(
        keyinput_g12), .A(n20971), .ZN(n20974) );
  NOR4_X1 U23894 ( .A1(n20977), .A2(n20976), .A3(n20975), .A4(n20974), .ZN(
        n21013) );
  AOI22_X1 U23895 ( .A1(n13420), .A2(keyinput_g21), .B1(keyinput_g26), .B2(
        n13417), .ZN(n20978) );
  OAI221_X1 U23896 ( .B1(n13420), .B2(keyinput_g21), .C1(n13417), .C2(
        keyinput_g26), .A(n20978), .ZN(n20985) );
  AOI22_X1 U23897 ( .A1(DATAI_28_), .A2(keyinput_g4), .B1(DATAI_13_), .B2(
        keyinput_g19), .ZN(n20979) );
  OAI221_X1 U23898 ( .B1(DATAI_28_), .B2(keyinput_g4), .C1(DATAI_13_), .C2(
        keyinput_g19), .A(n20979), .ZN(n20984) );
  AOI22_X1 U23899 ( .A1(n21062), .A2(keyinput_g48), .B1(n21082), .B2(
        keyinput_g3), .ZN(n20980) );
  OAI221_X1 U23900 ( .B1(n21062), .B2(keyinput_g48), .C1(n21082), .C2(
        keyinput_g3), .A(n20980), .ZN(n20983) );
  INV_X1 U23901 ( .A(DATAI_1_), .ZN(n21118) );
  AOI22_X1 U23902 ( .A1(n21118), .A2(keyinput_g31), .B1(n21073), .B2(
        keyinput_g15), .ZN(n20981) );
  OAI221_X1 U23903 ( .B1(n21118), .B2(keyinput_g31), .C1(n21073), .C2(
        keyinput_g15), .A(n20981), .ZN(n20982) );
  NOR4_X1 U23904 ( .A1(n20985), .A2(n20984), .A3(n20983), .A4(n20982), .ZN(
        n21012) );
  INV_X1 U23905 ( .A(BS16), .ZN(n21136) );
  AOI22_X1 U23906 ( .A1(n21136), .A2(keyinput_g35), .B1(n13405), .B2(
        keyinput_g28), .ZN(n20986) );
  OAI221_X1 U23907 ( .B1(n21136), .B2(keyinput_g35), .C1(n13405), .C2(
        keyinput_g28), .A(n20986), .ZN(n20996) );
  AOI22_X1 U23908 ( .A1(n21074), .A2(keyinput_g20), .B1(n21084), .B2(
        keyinput_g2), .ZN(n20987) );
  OAI221_X1 U23909 ( .B1(n21074), .B2(keyinput_g20), .C1(n21084), .C2(
        keyinput_g2), .A(n20987), .ZN(n20995) );
  INV_X1 U23910 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21139) );
  AOI22_X1 U23911 ( .A1(n20989), .A2(keyinput_g62), .B1(keyinput_g45), .B2(
        n21139), .ZN(n20988) );
  OAI221_X1 U23912 ( .B1(n20989), .B2(keyinput_g62), .C1(n21139), .C2(
        keyinput_g45), .A(n20988), .ZN(n20994) );
  INV_X1 U23913 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20992) );
  AOI22_X1 U23914 ( .A1(n20992), .A2(keyinput_g38), .B1(keyinput_g42), .B2(
        n20991), .ZN(n20990) );
  OAI221_X1 U23915 ( .B1(n20992), .B2(keyinput_g38), .C1(n20991), .C2(
        keyinput_g42), .A(n20990), .ZN(n20993) );
  NOR4_X1 U23916 ( .A1(n20996), .A2(n20995), .A3(n20994), .A4(n20993), .ZN(
        n21011) );
  AOI22_X1 U23917 ( .A1(n13175), .A2(keyinput_g0), .B1(n20998), .B2(
        keyinput_g7), .ZN(n20997) );
  OAI221_X1 U23918 ( .B1(n13175), .B2(keyinput_g0), .C1(n20998), .C2(
        keyinput_g7), .A(n20997), .ZN(n21009) );
  AOI22_X1 U23919 ( .A1(n21125), .A2(keyinput_g18), .B1(keyinput_g34), .B2(
        n21000), .ZN(n20999) );
  OAI221_X1 U23920 ( .B1(n21125), .B2(keyinput_g18), .C1(n21000), .C2(
        keyinput_g34), .A(n20999), .ZN(n21008) );
  INV_X1 U23921 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21002) );
  AOI22_X1 U23922 ( .A1(n21002), .A2(keyinput_g40), .B1(keyinput_g33), .B2(
        n21071), .ZN(n21001) );
  OAI221_X1 U23923 ( .B1(n21002), .B2(keyinput_g40), .C1(n21071), .C2(
        keyinput_g33), .A(n21001), .ZN(n21007) );
  INV_X1 U23924 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21005) );
  AOI22_X1 U23925 ( .A1(n21005), .A2(keyinput_g53), .B1(n21004), .B2(
        keyinput_g52), .ZN(n21003) );
  OAI221_X1 U23926 ( .B1(n21005), .B2(keyinput_g53), .C1(n21004), .C2(
        keyinput_g52), .A(n21003), .ZN(n21006) );
  NOR4_X1 U23927 ( .A1(n21009), .A2(n21008), .A3(n21007), .A4(n21006), .ZN(
        n21010) );
  NAND4_X1 U23928 ( .A1(n21013), .A2(n21012), .A3(n21011), .A4(n21010), .ZN(
        n21160) );
  AOI22_X1 U23929 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g51), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .ZN(n21014) );
  OAI221_X1 U23930 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), 
        .C1(P1_REIP_REG_23__SCAN_IN), .C2(keyinput_g60), .A(n21014), .ZN(
        n21021) );
  AOI22_X1 U23931 ( .A1(DATAI_18_), .A2(keyinput_g14), .B1(DATAI_10_), .B2(
        keyinput_g22), .ZN(n21015) );
  OAI221_X1 U23932 ( .B1(DATAI_18_), .B2(keyinput_g14), .C1(DATAI_10_), .C2(
        keyinput_g22), .A(n21015), .ZN(n21020) );
  AOI22_X1 U23933 ( .A1(DATAI_0_), .A2(keyinput_g32), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n21016) );
  OAI221_X1 U23934 ( .B1(DATAI_0_), .B2(keyinput_g32), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n21016), .ZN(n21019)
         );
  AOI22_X1 U23935 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_g47), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .ZN(n21017) );
  OAI221_X1 U23936 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_g47), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_g61), .A(n21017), .ZN(n21018)
         );
  NOR4_X1 U23937 ( .A1(n21021), .A2(n21020), .A3(n21019), .A4(n21018), .ZN(
        n21050) );
  XOR2_X1 U23938 ( .A(n21022), .B(keyinput_g44), .Z(n21030) );
  AOI22_X1 U23939 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(n21024), .B2(
        keyinput_g6), .ZN(n21023) );
  OAI221_X1 U23940 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(n21024), .C2(
        keyinput_g6), .A(n21023), .ZN(n21029) );
  AOI22_X1 U23941 ( .A1(DATAI_7_), .A2(keyinput_g25), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .ZN(n21025) );
  OAI221_X1 U23942 ( .B1(DATAI_7_), .B2(keyinput_g25), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_g55), .A(n21025), .ZN(n21028)
         );
  AOI22_X1 U23943 ( .A1(DATAI_16_), .A2(keyinput_g16), .B1(DATAI_31_), .B2(
        keyinput_g1), .ZN(n21026) );
  OAI221_X1 U23944 ( .B1(DATAI_16_), .B2(keyinput_g16), .C1(DATAI_31_), .C2(
        keyinput_g1), .A(n21026), .ZN(n21027) );
  NOR4_X1 U23945 ( .A1(n21030), .A2(n21029), .A3(n21028), .A4(n21027), .ZN(
        n21049) );
  AOI22_X1 U23946 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(DATAI_27_), .B2(
        keyinput_g5), .ZN(n21031) );
  OAI221_X1 U23947 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(DATAI_27_), .C2(
        keyinput_g5), .A(n21031), .ZN(n21038) );
  AOI22_X1 U23948 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .ZN(n21032) );
  OAI221_X1 U23949 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_g57), .A(n21032), .ZN(n21037)
         );
  AOI22_X1 U23950 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_g46), .B1(READY2), 
        .B2(keyinput_g37), .ZN(n21033) );
  OAI221_X1 U23951 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .C1(READY2), 
        .C2(keyinput_g37), .A(n21033), .ZN(n21036) );
  AOI22_X1 U23952 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n21034) );
  OAI221_X1 U23953 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n21034), .ZN(n21035)
         );
  NOR4_X1 U23954 ( .A1(n21038), .A2(n21037), .A3(n21036), .A4(n21035), .ZN(
        n21048) );
  AOI22_X1 U23955 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .ZN(n21039) );
  OAI221_X1 U23956 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_g59), .A(n21039), .ZN(n21046)
         );
  AOI22_X1 U23957 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        DATAI_23_), .B2(keyinput_g9), .ZN(n21040) );
  OAI221_X1 U23958 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        DATAI_23_), .C2(keyinput_g9), .A(n21040), .ZN(n21045) );
  AOI22_X1 U23959 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_g39), .B1(DATAI_5_), .B2(keyinput_g27), .ZN(n21041) );
  OAI221_X1 U23960 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_5_), .C2(keyinput_g27), .A(n21041), .ZN(n21044) );
  AOI22_X1 U23961 ( .A1(DATAI_9_), .A2(keyinput_g23), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .ZN(n21042) );
  OAI221_X1 U23962 ( .B1(DATAI_9_), .B2(keyinput_g23), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_g63), .A(n21042), .ZN(n21043)
         );
  NOR4_X1 U23963 ( .A1(n21046), .A2(n21045), .A3(n21044), .A4(n21043), .ZN(
        n21047) );
  NAND4_X1 U23964 ( .A1(n21050), .A2(n21049), .A3(n21048), .A4(n21047), .ZN(
        n21159) );
  OAI22_X1 U23965 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_f58), .B1(
        DATAI_4_), .B2(keyinput_f28), .ZN(n21051) );
  AOI221_X1 U23966 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .C1(
        keyinput_f28), .C2(DATAI_4_), .A(n21051), .ZN(n21058) );
  OAI22_X1 U23967 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_f54), .B1(
        DATAI_23_), .B2(keyinput_f9), .ZN(n21052) );
  AOI221_X1 U23968 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_f54), .C1(
        keyinput_f9), .C2(DATAI_23_), .A(n21052), .ZN(n21057) );
  OAI22_X1 U23969 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_f62), .B1(
        keyinput_f10), .B2(DATAI_22_), .ZN(n21053) );
  AOI221_X1 U23970 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .C1(
        DATAI_22_), .C2(keyinput_f10), .A(n21053), .ZN(n21056) );
  OAI22_X1 U23971 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_f46), .B1(
        keyinput_f41), .B2(P1_M_IO_N_REG_SCAN_IN), .ZN(n21054) );
  AOI221_X1 U23972 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .C1(
        P1_M_IO_N_REG_SCAN_IN), .C2(keyinput_f41), .A(n21054), .ZN(n21055) );
  NAND4_X1 U23973 ( .A1(n21058), .A2(n21057), .A3(n21056), .A4(n21055), .ZN(
        n21152) );
  OAI22_X1 U23974 ( .A1(READY1), .A2(keyinput_f36), .B1(DATAI_20_), .B2(
        keyinput_f12), .ZN(n21059) );
  AOI221_X1 U23975 ( .B1(READY1), .B2(keyinput_f36), .C1(keyinput_f12), .C2(
        DATAI_20_), .A(n21059), .ZN(n21066) );
  OAI22_X1 U23976 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_f44), .B1(
        DATAI_11_), .B2(keyinput_f21), .ZN(n21060) );
  AOI221_X1 U23977 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .C1(
        keyinput_f21), .C2(DATAI_11_), .A(n21060), .ZN(n21065) );
  OAI22_X1 U23978 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(DATAI_2_), .B2(
        keyinput_f30), .ZN(n21061) );
  AOI221_X1 U23979 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(keyinput_f30), .C2(
        DATAI_2_), .A(n21061), .ZN(n21064) );
  XOR2_X1 U23980 ( .A(keyinput_f48), .B(n21062), .Z(n21063) );
  NAND4_X1 U23981 ( .A1(n21066), .A2(n21065), .A3(n21064), .A4(n21063), .ZN(
        n21151) );
  OAI22_X1 U23982 ( .A1(n21069), .A2(keyinput_f56), .B1(n21068), .B2(
        keyinput_f47), .ZN(n21067) );
  AOI221_X1 U23983 ( .B1(n21069), .B2(keyinput_f56), .C1(keyinput_f47), .C2(
        n21068), .A(n21067), .ZN(n21099) );
  OAI22_X1 U23984 ( .A1(keyinput_f33), .A2(n21071), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .ZN(n21070) );
  AOI221_X1 U23985 ( .B1(n21071), .B2(keyinput_f33), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_f40), .A(n21070), .ZN(n21098)
         );
  OAI22_X1 U23986 ( .A1(n21074), .A2(keyinput_f20), .B1(n21073), .B2(
        keyinput_f15), .ZN(n21072) );
  AOI221_X1 U23987 ( .B1(n21074), .B2(keyinput_f20), .C1(keyinput_f15), .C2(
        n21073), .A(n21072), .ZN(n21077) );
  XOR2_X1 U23988 ( .A(keyinput_f39), .B(n21075), .Z(n21076) );
  OAI211_X1 U23989 ( .C1(n21079), .C2(keyinput_f1), .A(n21077), .B(n21076), 
        .ZN(n21078) );
  AOI21_X1 U23990 ( .B1(n21079), .B2(keyinput_f1), .A(n21078), .ZN(n21097) );
  AOI22_X1 U23991 ( .A1(n21082), .A2(keyinput_f3), .B1(keyinput_f49), .B2(
        n21081), .ZN(n21080) );
  OAI221_X1 U23992 ( .B1(n21082), .B2(keyinput_f3), .C1(n21081), .C2(
        keyinput_f49), .A(n21080), .ZN(n21095) );
  AOI22_X1 U23993 ( .A1(n21085), .A2(keyinput_f5), .B1(n21084), .B2(
        keyinput_f2), .ZN(n21083) );
  OAI221_X1 U23994 ( .B1(n21085), .B2(keyinput_f5), .C1(n21084), .C2(
        keyinput_f2), .A(n21083), .ZN(n21094) );
  AOI22_X1 U23995 ( .A1(n21088), .A2(keyinput_f16), .B1(n21087), .B2(
        keyinput_f59), .ZN(n21086) );
  OAI221_X1 U23996 ( .B1(n21088), .B2(keyinput_f16), .C1(n21087), .C2(
        keyinput_f59), .A(n21086), .ZN(n21093) );
  AOI22_X1 U23997 ( .A1(n21091), .A2(keyinput_f19), .B1(keyinput_f4), .B2(
        n21090), .ZN(n21089) );
  OAI221_X1 U23998 ( .B1(n21091), .B2(keyinput_f19), .C1(n21090), .C2(
        keyinput_f4), .A(n21089), .ZN(n21092) );
  NOR4_X1 U23999 ( .A1(n21095), .A2(n21094), .A3(n21093), .A4(n21092), .ZN(
        n21096) );
  NAND4_X1 U24000 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21150) );
  AOI22_X1 U24001 ( .A1(keyinput_f50), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .ZN(n21100) );
  OAI221_X1 U24002 ( .B1(keyinput_f50), .B2(P1_BYTEENABLE_REG_2__SCAN_IN), 
        .C1(P1_REIP_REG_22__SCAN_IN), .C2(keyinput_f61), .A(n21100), .ZN(
        n21107) );
  AOI22_X1 U24003 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .ZN(n21101) );
  OAI221_X1 U24004 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_REIP_REG_31__SCAN_IN), .C2(keyinput_f52), .A(n21101), .ZN(n21106)
         );
  AOI22_X1 U24005 ( .A1(keyinput_f34), .A2(NA), .B1(DATAI_24_), .B2(
        keyinput_f8), .ZN(n21102) );
  OAI221_X1 U24006 ( .B1(keyinput_f34), .B2(NA), .C1(DATAI_24_), .C2(
        keyinput_f8), .A(n21102), .ZN(n21105) );
  AOI22_X1 U24007 ( .A1(DATAI_3_), .A2(keyinput_f29), .B1(DATAI_19_), .B2(
        keyinput_f13), .ZN(n21103) );
  OAI221_X1 U24008 ( .B1(DATAI_3_), .B2(keyinput_f29), .C1(DATAI_19_), .C2(
        keyinput_f13), .A(n21103), .ZN(n21104) );
  NOR4_X1 U24009 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        n21148) );
  AOI22_X1 U24010 ( .A1(keyinput_f42), .A2(P1_D_C_N_REG_SCAN_IN), .B1(DATAI_5_), .B2(keyinput_f27), .ZN(n21108) );
  OAI221_X1 U24011 ( .B1(keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .C1(
        DATAI_5_), .C2(keyinput_f27), .A(n21108), .ZN(n21115) );
  AOI22_X1 U24012 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f0), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .ZN(n21109) );
  OAI221_X1 U24013 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f0), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_f53), .A(n21109), .ZN(n21114)
         );
  AOI22_X1 U24014 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .ZN(n21110) );
  OAI221_X1 U24015 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n21110), .ZN(n21113)
         );
  AOI22_X1 U24016 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .ZN(n21111) );
  OAI221_X1 U24017 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_f38), .A(n21111), .ZN(
        n21112) );
  NOR4_X1 U24018 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21147) );
  AOI22_X1 U24019 ( .A1(n21118), .A2(keyinput_f31), .B1(n21117), .B2(
        keyinput_f23), .ZN(n21116) );
  OAI221_X1 U24020 ( .B1(n21118), .B2(keyinput_f31), .C1(n21117), .C2(
        keyinput_f23), .A(n21116), .ZN(n21129) );
  AOI22_X1 U24021 ( .A1(n21120), .A2(keyinput_f11), .B1(n13414), .B2(
        keyinput_f25), .ZN(n21119) );
  OAI221_X1 U24022 ( .B1(n21120), .B2(keyinput_f11), .C1(n13414), .C2(
        keyinput_f25), .A(n21119), .ZN(n21128) );
  AOI22_X1 U24023 ( .A1(n21123), .A2(keyinput_f63), .B1(keyinput_f43), .B2(
        n21122), .ZN(n21121) );
  OAI221_X1 U24024 ( .B1(n21123), .B2(keyinput_f63), .C1(n21122), .C2(
        keyinput_f43), .A(n21121), .ZN(n21127) );
  AOI22_X1 U24025 ( .A1(n13417), .A2(keyinput_f26), .B1(n21125), .B2(
        keyinput_f18), .ZN(n21124) );
  OAI221_X1 U24026 ( .B1(n13417), .B2(keyinput_f26), .C1(n21125), .C2(
        keyinput_f18), .A(n21124), .ZN(n21126) );
  NOR4_X1 U24027 ( .A1(n21129), .A2(n21128), .A3(n21127), .A4(n21126), .ZN(
        n21146) );
  INV_X1 U24028 ( .A(READY2), .ZN(n21131) );
  AOI22_X1 U24029 ( .A1(n21132), .A2(keyinput_f22), .B1(keyinput_f37), .B2(
        n21131), .ZN(n21130) );
  OAI221_X1 U24030 ( .B1(n21132), .B2(keyinput_f22), .C1(n21131), .C2(
        keyinput_f37), .A(n21130), .ZN(n21144) );
  AOI22_X1 U24031 ( .A1(n13298), .A2(keyinput_f17), .B1(n21134), .B2(
        keyinput_f55), .ZN(n21133) );
  OAI221_X1 U24032 ( .B1(n13298), .B2(keyinput_f17), .C1(n21134), .C2(
        keyinput_f55), .A(n21133), .ZN(n21143) );
  INV_X1 U24033 ( .A(DATAI_0_), .ZN(n21137) );
  AOI22_X1 U24034 ( .A1(n21137), .A2(keyinput_f32), .B1(keyinput_f35), .B2(
        n21136), .ZN(n21135) );
  OAI221_X1 U24035 ( .B1(n21137), .B2(keyinput_f32), .C1(n21136), .C2(
        keyinput_f35), .A(n21135), .ZN(n21142) );
  AOI22_X1 U24036 ( .A1(n21140), .A2(keyinput_f14), .B1(keyinput_f45), .B2(
        n21139), .ZN(n21138) );
  OAI221_X1 U24037 ( .B1(n21140), .B2(keyinput_f14), .C1(n21139), .C2(
        keyinput_f45), .A(n21138), .ZN(n21141) );
  NOR4_X1 U24038 ( .A1(n21144), .A2(n21143), .A3(n21142), .A4(n21141), .ZN(
        n21145) );
  NAND4_X1 U24039 ( .A1(n21148), .A2(n21147), .A3(n21146), .A4(n21145), .ZN(
        n21149) );
  NOR4_X1 U24040 ( .A1(n21152), .A2(n21151), .A3(n21150), .A4(n21149), .ZN(
        n21155) );
  INV_X1 U24041 ( .A(n21155), .ZN(n21153) );
  AOI211_X1 U24042 ( .C1(keyinput_f24), .C2(n21153), .A(DATAI_8_), .B(
        keyinput_g24), .ZN(n21154) );
  INV_X1 U24043 ( .A(n21154), .ZN(n21157) );
  OAI211_X1 U24044 ( .C1(n21155), .C2(keyinput_f24), .A(DATAI_8_), .B(
        keyinput_g24), .ZN(n21156) );
  NAND2_X1 U24045 ( .A1(n21157), .A2(n21156), .ZN(n21158) );
  OAI21_X1 U24046 ( .B1(n21160), .B2(n21159), .A(n21158), .ZN(n21161) );
  XOR2_X1 U24047 ( .A(n21162), .B(n21161), .Z(U355) );
  OAI211_X1 U13318 ( .C1(n10387), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        n10405) );
  AND2_X1 U13377 ( .A1(n14500), .A2(n10275), .ZN(n10632) );
  NAND2_X1 U13281 ( .A1(n19474), .A2(n19470), .ZN(n10342) );
  CLKBUF_X1 U11109 ( .A(n11545), .Z(n11868) );
  OR2_X1 U11111 ( .A1(n10569), .A2(n10568), .ZN(n10997) );
  CLKBUF_X1 U11169 ( .A(n10408), .Z(n13312) );
  CLKBUF_X1 U11187 ( .A(n12886), .Z(n12953) );
  CLKBUF_X1 U11188 ( .A(n15243), .Z(n19288) );
  INV_X1 U11428 ( .A(n17945), .ZN(n17986) );
  CLKBUF_X1 U11517 ( .A(n18076), .Z(n9676) );
  INV_X1 U11943 ( .A(n13895), .ZN(n14611) );
  CLKBUF_X1 U11946 ( .A(n19417), .Z(n20146) );
  CLKBUF_X1 U12242 ( .A(n10405), .Z(n10406) );
  CLKBUF_X1 U12294 ( .A(n13657), .Z(n9689) );
  OR2_X1 U12386 ( .A1(n18448), .A2(n18447), .ZN(n21163) );
  OR2_X1 U12558 ( .A1(n13281), .A2(n13280), .ZN(n21164) );
  CLKBUF_X1 U12833 ( .A(n17696), .Z(n17704) );
endmodule

