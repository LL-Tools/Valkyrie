

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259;

  AND4_X2 U2530 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n4141)
         );
  AND4_X1 U2531 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n4164)
         );
  OAI21_X1 U2532 ( .B1(n3388), .B2(n5085), .A(n4883), .ZN(n4042) );
  CLKBUF_X2 U2533 ( .A(n2828), .Z(n3650) );
  OAI211_X2 U2534 ( .C1(n2761), .C2(n2633), .A(n2851), .B(n2631), .ZN(n5003)
         );
  AND2_X1 U2535 ( .A1(n2496), .A2(n2766), .ZN(n2643) );
  INV_X1 U2536 ( .A(n3603), .ZN(n2800) );
  INV_X1 U2537 ( .A(n2864), .ZN(n2843) );
  INV_X1 U2538 ( .A(n2869), .ZN(n2496) );
  AOI22_X1 U2539 ( .A1(n4820), .A2(REG2_REG_1__SCAN_IN), .B1(n5024), .B2(n5003), .ZN(n4822) );
  INV_X1 U2540 ( .A(IR_REG_31__SCAN_IN), .ZN(n2761) );
  OR2_X1 U2541 ( .A1(n4344), .A2(n4343), .ZN(n5257) );
  XNOR2_X1 U2542 ( .A(n2780), .B(IR_REG_29__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U2543 ( .A1(n3143), .A2(n3127), .ZN(n2654) );
  NAND2_X2 U2544 ( .A1(n3113), .A2(n4769), .ZN(n2802) );
  NAND2_X1 U2545 ( .A1(n2802), .A2(n2790), .ZN(n2848) );
  OR2_X1 U2546 ( .A1(n4956), .A2(n2629), .ZN(n2628) );
  OR2_X1 U2547 ( .A1(n4068), .A2(n4069), .ZN(n4082) );
  OAI21_X1 U2548 ( .B1(n3769), .B2(n2707), .A(n2704), .ZN(n3023) );
  NAND2_X1 U2549 ( .A1(n4925), .A2(n2738), .ZN(n4048) );
  NAND2_X1 U2550 ( .A1(n4904), .A2(n2527), .ZN(n4045) );
  OR2_X2 U2551 ( .A1(n4344), .A2(n4342), .ZN(n5254) );
  NAND2_X1 U2552 ( .A1(n2791), .A2(n2790), .ZN(n2828) );
  NAND2_X1 U2553 ( .A1(n2744), .A2(n2822), .ZN(n5010) );
  NAND2_X1 U2554 ( .A1(n3093), .A2(n2763), .ZN(n2790) );
  INV_X2 U2555 ( .A(n2654), .ZN(n3603) );
  NAND2_X1 U2556 ( .A1(n4830), .A2(n4031), .ZN(n4032) );
  CLKBUF_X1 U2557 ( .A(n2830), .Z(n3826) );
  INV_X2 U2558 ( .A(n2830), .ZN(n3565) );
  OAI21_X1 U2559 ( .B1(n5049), .B2(n5027), .A(n4979), .ZN(n4030) );
  INV_X1 U2560 ( .A(n4766), .ZN(n2495) );
  XNOR2_X1 U2561 ( .A(n2799), .B(n4681), .ZN(n3127) );
  NAND2_X1 U2562 ( .A1(n2774), .A2(n4475), .ZN(n2777) );
  AND2_X1 U2563 ( .A1(n2980), .A2(n2746), .ZN(n2774) );
  INV_X1 U2564 ( .A(n5027), .ZN(n4975) );
  NAND2_X1 U2565 ( .A1(n2623), .A2(n2622), .ZN(n5027) );
  AND4_X1 U2566 ( .A1(n2757), .A2(n2508), .A3(n2756), .A4(n2755), .ZN(n2758)
         );
  AND2_X1 U2567 ( .A1(n2752), .A2(n2751), .ZN(n2757) );
  INV_X1 U2568 ( .A(n2709), .ZN(n2708) );
  INV_X1 U2569 ( .A(IR_REG_23__SCAN_IN), .ZN(n4480) );
  NOR2_X2 U2570 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2850)
         );
  AOI21_X1 U2571 ( .B1(IR_REG_31__SCAN_IN), .B2(IR_REG_18__SCAN_IN), .A(
        IR_REG_19__SCAN_IN), .ZN(n2709) );
  INV_X1 U2572 ( .A(IR_REG_20__SCAN_IN), .ZN(n4669) );
  INV_X1 U2573 ( .A(IR_REG_13__SCAN_IN), .ZN(n2982) );
  INV_X1 U2574 ( .A(IR_REG_4__SCAN_IN), .ZN(n2748) );
  NOR2_X1 U2575 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2752)
         );
  NOR2_X1 U2576 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2751)
         );
  NOR2_X1 U2577 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2749)
         );
  NOR2_X1 U2578 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2750)
         );
  AOI22_X1 U2579 ( .A1(n3992), .A2(n3665), .B1(n3063), .B2(n5004), .ZN(n2838)
         );
  AOI22_X1 U2580 ( .A1(n3601), .A2(n3889), .B1(n3672), .B2(n3981), .ZN(n3605)
         );
  NOR2_X2 U2581 ( .A1(n3356), .A2(n3357), .ZN(n3368) );
  INV_X1 U2582 ( .A(IR_REG_31__SCAN_IN), .ZN(n2497) );
  INV_X4 U2583 ( .A(n3063), .ZN(n2825) );
  INV_X2 U2584 ( .A(n3651), .ZN(n2855) );
  OR2_X2 U2585 ( .A1(n4141), .A2(n3644), .ZN(n3547) );
  AND4_X4 U2586 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n4105)
         );
  OAI22_X2 U2587 ( .A1(n3402), .A2(n3403), .B1(n2935), .B2(n2934), .ZN(n3448)
         );
  NAND2_X2 U2588 ( .A1(n2732), .A2(n2733), .ZN(n3402) );
  OAI22_X2 U2589 ( .A1(n4111), .A2(n3574), .B1(n4127), .B2(n3657), .ZN(n3601)
         );
  XNOR2_X2 U2590 ( .A(n2710), .B(n4669), .ZN(n3113) );
  OAI22_X2 U2591 ( .A1(n2553), .A2(n2549), .B1(n2675), .B2(n2678), .ZN(n4111)
         );
  INV_X1 U2592 ( .A(n2843), .ZN(n3195) );
  INV_X1 U2594 ( .A(n2667), .ZN(n2666) );
  INV_X1 U2595 ( .A(n4765), .ZN(n2784) );
  NOR2_X1 U2596 ( .A1(n2551), .A2(n3503), .ZN(n2550) );
  INV_X1 U2597 ( .A(n2554), .ZN(n2551) );
  INV_X1 U2598 ( .A(n2558), .ZN(n2557) );
  OAI22_X1 U2599 ( .A1(n3431), .A2(n2559), .B1(n3480), .B2(n3435), .ZN(n2558)
         );
  NAND2_X1 U2600 ( .A1(n2521), .A2(n3434), .ZN(n2559) );
  AOI21_X1 U2601 ( .B1(n2534), .B2(n2536), .A(n2519), .ZN(n2531) );
  OR2_X1 U2602 ( .A1(n3991), .A2(n3281), .ZN(n3929) );
  OR2_X1 U2603 ( .A1(n3237), .A2(n3236), .ZN(n5036) );
  NOR2_X1 U2604 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2755)
         );
  OAI21_X1 U2605 ( .B1(n2718), .B2(n2720), .A(n2717), .ZN(n2716) );
  NAND2_X1 U2606 ( .A1(n2720), .A2(n3662), .ZN(n2717) );
  NOR2_X1 U2607 ( .A1(n3686), .A2(n3661), .ZN(n2718) );
  NAND2_X1 U2608 ( .A1(n3748), .A2(n3751), .ZN(n3720) );
  AOI22_X1 U2609 ( .A1(n3237), .A2(n2855), .B1(n3665), .B2(n5014), .ZN(n2857)
         );
  OR2_X1 U2610 ( .A1(n2842), .A2(n4170), .ZN(n3181) );
  NAND2_X1 U2611 ( .A1(n4901), .A2(n2528), .ZN(n4012) );
  NAND2_X1 U2612 ( .A1(n4946), .A2(n4945), .ZN(n4944) );
  AND4_X1 U2613 ( .A1(n3573), .A2(n3572), .A3(n3571), .A4(n3570), .ZN(n4127)
         );
  OR2_X1 U2614 ( .A1(n2553), .A2(n2548), .ZN(n3505) );
  INV_X1 U2615 ( .A(n2550), .ZN(n2548) );
  OAI21_X1 U2616 ( .B1(n3288), .B2(n3286), .A(n2543), .ZN(n2545) );
  OR2_X1 U2617 ( .A1(n3150), .A2(D_REG_0__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U2618 ( .A1(n2653), .A2(n2652), .ZN(n5004) );
  NAND2_X1 U2619 ( .A1(n3143), .A2(n2498), .ZN(n2652) );
  NAND2_X1 U2620 ( .A1(n2654), .A2(DATAI_0_), .ZN(n2653) );
  AND4_X1 U2621 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(n3833)
         );
  NOR2_X1 U2622 ( .A1(n2511), .A2(n2590), .ZN(n2589) );
  INV_X1 U2623 ( .A(n2591), .ZN(n2590) );
  NOR2_X1 U2624 ( .A1(n3958), .A2(n2665), .ZN(n2664) );
  NOR2_X1 U2625 ( .A1(n2670), .A2(n2666), .ZN(n2665) );
  NOR2_X1 U2626 ( .A1(n3844), .A2(n2592), .ZN(n2591) );
  INV_X1 U2627 ( .A(n3846), .ZN(n2592) );
  INV_X1 U2628 ( .A(n3843), .ZN(n2640) );
  INV_X1 U2629 ( .A(n3310), .ZN(n2546) );
  NOR2_X1 U2630 ( .A1(n3532), .A2(n2668), .ZN(n2667) );
  INV_X1 U2631 ( .A(n3956), .ZN(n2668) );
  INV_X1 U2632 ( .A(n2950), .ZN(n2727) );
  NOR2_X1 U2633 ( .A1(n2517), .A2(n3454), .ZN(n2730) );
  AND2_X1 U2634 ( .A1(n2705), .A2(n3003), .ZN(n2704) );
  NAND2_X1 U2635 ( .A1(n3695), .A2(n2706), .ZN(n2705) );
  INV_X1 U2636 ( .A(n3695), .ZN(n2707) );
  NAND2_X1 U2637 ( .A1(n4840), .A2(n2621), .ZN(n4035) );
  NAND2_X1 U2638 ( .A1(n4027), .A2(REG2_REG_5__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U2639 ( .A1(n2514), .A2(n2676), .ZN(n2675) );
  NAND2_X1 U2640 ( .A1(n3563), .A2(n2677), .ZN(n2676) );
  INV_X1 U2641 ( .A(n3563), .ZN(n2680) );
  INV_X1 U2642 ( .A(n2664), .ZN(n2663) );
  AOI21_X1 U2643 ( .B1(n2664), .B2(n2666), .A(n2662), .ZN(n2661) );
  INV_X1 U2644 ( .A(n3849), .ZN(n2662) );
  NAND2_X1 U2645 ( .A1(n2594), .A2(n2670), .ZN(n2669) );
  NOR2_X1 U2646 ( .A1(n4179), .A2(n4166), .ZN(n2619) );
  OR2_X1 U2647 ( .A1(n4156), .A2(n4157), .ZN(n4159) );
  AND2_X1 U2648 ( .A1(n4205), .A2(n4179), .ZN(n4160) );
  AND2_X1 U2649 ( .A1(n2682), .A2(n3504), .ZN(n2681) );
  NOR2_X1 U2650 ( .A1(n3517), .A2(n2642), .ZN(n2641) );
  INV_X1 U2651 ( .A(n3872), .ZN(n2642) );
  NAND2_X1 U2652 ( .A1(n2688), .A2(n2687), .ZN(n3495) );
  AOI21_X1 U2653 ( .B1(n2689), .B2(n2690), .A(n4268), .ZN(n2687) );
  NAND2_X1 U2654 ( .A1(n2562), .A2(n4268), .ZN(n3496) );
  INV_X1 U2655 ( .A(n2571), .ZN(n2570) );
  OAI21_X1 U2656 ( .B1(n2573), .B2(n2572), .A(n4266), .ZN(n2571) );
  INV_X1 U2657 ( .A(n3944), .ZN(n2572) );
  NOR2_X1 U2658 ( .A1(n2574), .A2(n3512), .ZN(n2573) );
  INV_X1 U2659 ( .A(n3837), .ZN(n2574) );
  NOR2_X1 U2660 ( .A1(n5162), .A2(n3473), .ZN(n2617) );
  AND2_X1 U2661 ( .A1(n3913), .A2(n2579), .ZN(n2578) );
  NAND2_X1 U2662 ( .A1(n2580), .A2(n3916), .ZN(n2579) );
  INV_X1 U2663 ( .A(n3909), .ZN(n2580) );
  INV_X1 U2664 ( .A(n3916), .ZN(n2581) );
  OR2_X1 U2665 ( .A1(n5118), .A2(n3467), .ZN(n3916) );
  NAND2_X1 U2666 ( .A1(n2584), .A2(n2582), .ZN(n5125) );
  AOI21_X1 U2667 ( .B1(n2586), .B2(n2588), .A(n2583), .ZN(n2582) );
  INV_X1 U2668 ( .A(n3908), .ZN(n2583) );
  AND2_X1 U2669 ( .A1(n3411), .A2(n2539), .ZN(n2538) );
  NAND2_X1 U2670 ( .A1(n3385), .A2(n2540), .ZN(n2539) );
  NAND2_X1 U2671 ( .A1(n2595), .A2(n3876), .ZN(n3302) );
  NAND2_X1 U2672 ( .A1(n3282), .A2(n3928), .ZN(n2595) );
  OR2_X1 U2673 ( .A1(n2824), .A2(n5010), .ZN(n3923) );
  NAND2_X1 U2674 ( .A1(n5036), .A2(n3921), .ZN(n5012) );
  INV_X1 U2675 ( .A(IR_REG_26__SCAN_IN), .ZN(n2795) );
  NAND2_X1 U2676 ( .A1(n2770), .A2(n2771), .ZN(n2772) );
  INV_X1 U2677 ( .A(n2777), .ZN(n2770) );
  NAND2_X1 U2678 ( .A1(n2777), .A2(IR_REG_31__SCAN_IN), .ZN(n2613) );
  AOI21_X1 U2679 ( .B1(n2700), .B2(n3040), .A(n2699), .ZN(n2698) );
  INV_X1 U2680 ( .A(n3740), .ZN(n2700) );
  INV_X1 U2681 ( .A(n3793), .ZN(n2699) );
  AOI21_X1 U2682 ( .B1(n2698), .B2(n2701), .A(n2697), .ZN(n2696) );
  INV_X1 U2683 ( .A(n3040), .ZN(n2701) );
  INV_X1 U2684 ( .A(n3792), .ZN(n2697) );
  OR2_X1 U2685 ( .A1(n2825), .A2(n3239), .ZN(n2870) );
  OR2_X1 U2686 ( .A1(n3321), .A2(n3651), .ZN(n2835) );
  INV_X1 U2687 ( .A(n2829), .ZN(n2836) );
  AOI21_X1 U2688 ( .B1(n2696), .B2(n2603), .A(n2602), .ZN(n2601) );
  INV_X1 U2689 ( .A(n3713), .ZN(n2602) );
  INV_X1 U2690 ( .A(n2698), .ZN(n2603) );
  INV_X1 U2691 ( .A(n2696), .ZN(n2604) );
  AOI21_X1 U2692 ( .B1(n2609), .B2(n2973), .A(n2607), .ZN(n2606) );
  XNOR2_X1 U2693 ( .A(n2827), .B(n2958), .ZN(n2860) );
  AOI21_X1 U2694 ( .B1(n5010), .B2(n3665), .A(n2826), .ZN(n2827) );
  NOR2_X1 U2695 ( .A1(n2825), .A2(n2824), .ZN(n2826) );
  AOI22_X1 U2696 ( .A1(n2855), .A2(n5010), .B1(n3665), .B2(n5028), .ZN(n2861)
         );
  NOR2_X1 U2697 ( .A1(n2991), .A2(n3697), .ZN(n3007) );
  NAND2_X1 U2698 ( .A1(n3007), .A2(REG3_REG_15__SCAN_IN), .ZN(n3012) );
  OR2_X1 U2699 ( .A1(n2842), .A2(n3723), .ZN(n3206) );
  AND4_X1 U2700 ( .A1(n2979), .A2(n2978), .A3(n2977), .A4(n2976), .ZN(n3480)
         );
  INV_X1 U2701 ( .A(n3822), .ZN(n3030) );
  OR2_X1 U2702 ( .A1(n2842), .A2(REG3_REG_3__SCAN_IN), .ZN(n2866) );
  NAND4_X1 U2703 ( .A1(n2847), .A2(n2844), .A3(n2846), .A4(n2845), .ZN(n3237)
         );
  OR2_X1 U2704 ( .A1(n2842), .A2(n2841), .ZN(n2846) );
  NAND2_X1 U2705 ( .A1(n4976), .A2(n2509), .ZN(n4000) );
  NAND2_X1 U2706 ( .A1(n4831), .A2(REG2_REG_3__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U2707 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  XNOR2_X1 U2708 ( .A(n4035), .B(n4004), .ZN(n4850) );
  NAND2_X1 U2709 ( .A1(n4850), .A2(REG2_REG_6__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U2710 ( .A1(n4892), .A2(n4043), .ZN(n4906) );
  NAND2_X1 U2711 ( .A1(n4906), .A2(n4905), .ZN(n4904) );
  NAND2_X1 U2712 ( .A1(n4927), .A2(n4926), .ZN(n4925) );
  NAND2_X1 U2713 ( .A1(n4922), .A2(n2525), .ZN(n4017) );
  XNOR2_X1 U2714 ( .A(n4048), .B(n4016), .ZN(n4939) );
  XNOR2_X1 U2715 ( .A(n4072), .B(n4772), .ZN(n4051) );
  NAND2_X1 U2716 ( .A1(n4950), .A2(n4050), .ZN(n4072) );
  NAND2_X1 U2717 ( .A1(n4944), .A2(n4019), .ZN(n4064) );
  INV_X1 U2718 ( .A(n2630), .ZN(n2629) );
  AOI21_X1 U2719 ( .B1(n4770), .B2(REG1_REG_18__SCAN_IN), .A(n4083), .ZN(n2630) );
  NOR2_X1 U2720 ( .A1(n3606), .A2(n5217), .ZN(n3592) );
  NOR2_X2 U2721 ( .A1(n2620), .A2(n3726), .ZN(n4133) );
  NAND2_X1 U2722 ( .A1(n4162), .A2(n3558), .ZN(n4140) );
  NOR2_X1 U2723 ( .A1(n4175), .A2(n2682), .ZN(n4177) );
  NAND2_X1 U2724 ( .A1(n3505), .A2(n2681), .ZN(n4189) );
  NAND2_X1 U2725 ( .A1(n2555), .A2(n4224), .ZN(n2554) );
  INV_X1 U2726 ( .A(n5211), .ZN(n2555) );
  NOR2_X1 U2727 ( .A1(n4212), .A2(n3502), .ZN(n2553) );
  NAND2_X1 U2728 ( .A1(n3497), .A2(n3496), .ZN(n4227) );
  NAND2_X1 U2729 ( .A1(n3493), .A2(n3492), .ZN(n3494) );
  AND2_X1 U2730 ( .A1(n3902), .A2(n3841), .ZN(n4266) );
  NAND2_X1 U2731 ( .A1(n3679), .A2(n3341), .ZN(n2540) );
  AOI21_X1 U2732 ( .B1(n3873), .B2(n2685), .A(n2507), .ZN(n2683) );
  OAI21_X1 U2733 ( .B1(n3373), .B2(n3304), .A(n3935), .ZN(n3339) );
  AND2_X1 U2734 ( .A1(n3936), .A2(n3904), .ZN(n3874) );
  NAND2_X1 U2735 ( .A1(n3290), .A2(n3289), .ZN(n3311) );
  NAND2_X1 U2736 ( .A1(n2747), .A2(n2565), .ZN(n5033) );
  NAND2_X1 U2737 ( .A1(n2852), .A2(n2615), .ZN(n5014) );
  NAND2_X1 U2738 ( .A1(n3603), .A2(n4820), .ZN(n2852) );
  NAND2_X1 U2739 ( .A1(n3095), .A2(n4767), .ZN(n3150) );
  NAND2_X1 U2740 ( .A1(n2693), .A2(n4681), .ZN(n2692) );
  INV_X1 U2741 ( .A(n2694), .ZN(n2693) );
  NOR2_X1 U2742 ( .A1(n2797), .A2(IR_REG_27__SCAN_IN), .ZN(n2659) );
  NOR2_X1 U2743 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2658)
         );
  INV_X1 U2744 ( .A(IR_REG_1__SCAN_IN), .ZN(n2632) );
  NOR2_X1 U2745 ( .A1(n2714), .A2(n3815), .ZN(n2712) );
  AND2_X1 U2746 ( .A1(n2515), .A2(n2716), .ZN(n2714) );
  NAND2_X1 U2747 ( .A1(n2716), .A2(n2719), .ZN(n2715) );
  NAND2_X1 U2748 ( .A1(n3668), .A2(n3662), .ZN(n2719) );
  INV_X1 U2749 ( .A(n3720), .ZN(n3718) );
  NAND2_X1 U2750 ( .A1(n2734), .A2(n2737), .ZN(n2733) );
  NAND2_X1 U2751 ( .A1(n3676), .A2(n2506), .ZN(n2732) );
  INV_X1 U2752 ( .A(n2735), .ZN(n2734) );
  INV_X1 U2753 ( .A(n4230), .ZN(n3762) );
  AND4_X1 U2754 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n4178)
         );
  INV_X1 U2755 ( .A(n5034), .ZN(n3266) );
  AND4_X1 U2756 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n4182)
         );
  NAND4_X1 U2757 ( .A1(n2811), .A2(n2810), .A3(n2809), .A4(n2808), .ZN(n3990)
         );
  NAND4_X1 U2758 ( .A1(n2879), .A2(n2878), .A3(n2877), .A4(n2876), .ZN(n3991)
         );
  NAND2_X1 U2759 ( .A1(n4894), .A2(n4011), .ZN(n4903) );
  NAND2_X1 U2760 ( .A1(n4903), .A2(n4902), .ZN(n4901) );
  XNOR2_X1 U2761 ( .A(n4012), .B(n5143), .ZN(n4916) );
  NAND2_X1 U2762 ( .A1(n4924), .A2(n4923), .ZN(n4922) );
  NAND2_X1 U2763 ( .A1(n4951), .A2(n4952), .ZN(n4950) );
  XNOR2_X1 U2764 ( .A(n4064), .B(n4772), .ZN(n4020) );
  AOI21_X1 U2765 ( .B1(n4988), .B2(ADDR_REG_18__SCAN_IN), .A(n4961), .ZN(n2626) );
  AND2_X1 U2766 ( .A1(n2628), .A2(n4992), .ZN(n2627) );
  NAND2_X1 U2767 ( .A1(n3619), .A2(n5244), .ZN(n4304) );
  OAI21_X1 U2768 ( .B1(n2597), .B2(n5217), .A(n2634), .ZN(n3624) );
  INV_X1 U2769 ( .A(n3615), .ZN(n2634) );
  XNOR2_X1 U2770 ( .A(n3607), .B(n3891), .ZN(n2597) );
  XNOR2_X1 U2771 ( .A(n3605), .B(n3604), .ZN(n4306) );
  NAND2_X1 U2772 ( .A1(n4311), .A2(n3157), .ZN(n5224) );
  NOR2_X1 U2773 ( .A1(n2760), .A2(n2694), .ZN(n2798) );
  OR2_X1 U2774 ( .A1(n3553), .A2(n4120), .ZN(n3556) );
  INV_X1 U2775 ( .A(n2989), .ZN(n2706) );
  INV_X1 U2776 ( .A(n3507), .ZN(n2677) );
  INV_X1 U2777 ( .A(n2587), .ZN(n2586) );
  OAI21_X1 U2778 ( .B1(n3938), .B2(n2588), .A(n5096), .ZN(n2587) );
  INV_X1 U2779 ( .A(IR_REG_21__SCAN_IN), .ZN(n4475) );
  INV_X1 U2780 ( .A(IR_REG_14__SCAN_IN), .ZN(n4464) );
  NOR2_X1 U2781 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2756)
         );
  INV_X1 U2782 ( .A(n3767), .ZN(n2607) );
  NAND2_X1 U2783 ( .A1(n3565), .A2(REG2_REG_1__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U2784 ( .A1(n4861), .A2(n4037), .ZN(n4038) );
  NOR2_X1 U2785 ( .A1(n4099), .A2(n3672), .ZN(n3617) );
  NAND2_X1 U2786 ( .A1(n2593), .A2(n2660), .ZN(n4101) );
  AOI21_X1 U2787 ( .B1(n2512), .B2(n2661), .A(n3818), .ZN(n2660) );
  NAND2_X1 U2788 ( .A1(n3526), .A2(n2589), .ZN(n2593) );
  OR2_X1 U2789 ( .A1(n2842), .A2(n4116), .ZN(n3571) );
  OR2_X1 U2790 ( .A1(n3177), .A2(n4603), .ZN(n3196) );
  OR2_X1 U2791 ( .A1(n3885), .A2(n2674), .ZN(n2673) );
  NOR2_X1 U2792 ( .A1(n2639), .A2(n2638), .ZN(n2637) );
  INV_X1 U2793 ( .A(n3523), .ZN(n2638) );
  NOR2_X1 U2794 ( .A1(n2641), .A2(n2640), .ZN(n2639) );
  AND2_X1 U2795 ( .A1(REG3_REG_18__SCAN_IN), .A2(n3042), .ZN(n3055) );
  NOR2_X1 U2796 ( .A1(n5160), .A2(n4272), .ZN(n2690) );
  OR2_X1 U2797 ( .A1(n4247), .A2(n3514), .ZN(n2689) );
  NAND2_X1 U2798 ( .A1(n3423), .A2(n3916), .ZN(n3479) );
  AOI21_X1 U2799 ( .B1(n2538), .B2(n2535), .A(n2505), .ZN(n2534) );
  INV_X1 U2800 ( .A(n2540), .ZN(n2535) );
  INV_X1 U2801 ( .A(n3414), .ZN(n2691) );
  INV_X1 U2802 ( .A(n2538), .ZN(n2536) );
  INV_X1 U2803 ( .A(n3904), .ZN(n2649) );
  NOR2_X1 U2804 ( .A1(n3874), .A2(n2686), .ZN(n2685) );
  INV_X1 U2805 ( .A(n3315), .ZN(n2686) );
  AND2_X1 U2806 ( .A1(n3367), .A2(n3308), .ZN(n2616) );
  NOR2_X1 U2807 ( .A1(n2544), .A2(n2546), .ZN(n2543) );
  NOR2_X1 U2808 ( .A1(n3287), .A2(n3286), .ZN(n2544) );
  AND2_X1 U2809 ( .A1(n2542), .A2(n3312), .ZN(n2541) );
  OR2_X1 U2810 ( .A1(n2546), .A2(n3289), .ZN(n2542) );
  AND2_X1 U2811 ( .A1(n2892), .A2(REG3_REG_6__SCAN_IN), .ZN(n2906) );
  AOI21_X1 U2812 ( .B1(n3288), .B2(n3287), .A(n3286), .ZN(n3290) );
  INV_X1 U2813 ( .A(n3285), .ZN(n3239) );
  AND2_X1 U2814 ( .A1(n2669), .A2(n2667), .ZN(n3576) );
  OR2_X1 U2815 ( .A1(n2898), .A2(IR_REG_6__SCAN_IN), .ZN(n2929) );
  INV_X1 U2816 ( .A(n2730), .ZN(n2728) );
  NAND2_X1 U2817 ( .A1(n2727), .A2(n2731), .ZN(n2726) );
  NAND2_X1 U2818 ( .A1(n2517), .A2(n3454), .ZN(n2731) );
  INV_X1 U2819 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U2820 ( .A1(n3012), .A2(n4427), .ZN(n3028) );
  NOR2_X1 U2821 ( .A1(n3640), .A2(n2722), .ZN(n2721) );
  INV_X1 U2822 ( .A(n3638), .ZN(n2722) );
  NAND2_X1 U2823 ( .A1(n3706), .A2(n3638), .ZN(n2610) );
  XNOR2_X1 U2824 ( .A(n2884), .B(n2958), .ZN(n2885) );
  NAND2_X1 U2825 ( .A1(n2919), .A2(n2920), .ZN(n2737) );
  NOR2_X1 U2826 ( .A1(n3394), .A2(n2736), .ZN(n2735) );
  INV_X1 U2827 ( .A(n2917), .ZN(n2736) );
  OR2_X1 U2828 ( .A1(n2730), .A2(n3449), .ZN(n2729) );
  NAND2_X1 U2829 ( .A1(n2725), .A2(n3463), .ZN(n2609) );
  AND2_X1 U2830 ( .A1(n3126), .A2(n3157), .ZN(n3167) );
  NAND2_X1 U2831 ( .A1(n2703), .A2(n2702), .ZN(n5169) );
  AOI21_X1 U2832 ( .B1(n2704), .B2(n2707), .A(n2516), .ZN(n2702) );
  OR2_X1 U2833 ( .A1(n2842), .A2(n4134), .ZN(n3216) );
  XNOR2_X1 U2834 ( .A(n4030), .B(n4029), .ZN(n4831) );
  NAND2_X1 U2835 ( .A1(n4828), .A2(n4001), .ZN(n4002) );
  NAND2_X1 U2836 ( .A1(n4994), .A2(n4034), .ZN(n4842) );
  OAI21_X1 U2837 ( .B1(n5064), .B2(n5059), .A(n4837), .ZN(n4005) );
  NAND2_X1 U2838 ( .A1(n4849), .A2(n4036), .ZN(n4863) );
  NAND2_X1 U2839 ( .A1(n4863), .A2(n4862), .ZN(n4861) );
  XNOR2_X1 U2840 ( .A(n4038), .B(n4039), .ZN(n4875) );
  NAND2_X1 U2841 ( .A1(n4007), .A2(n4858), .ZN(n4008) );
  INV_X1 U2842 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4435) );
  XNOR2_X1 U2843 ( .A(n4042), .B(n4041), .ZN(n4893) );
  NAND2_X1 U2844 ( .A1(n4893), .A2(REG2_REG_10__SCAN_IN), .ZN(n4892) );
  OAI21_X1 U2845 ( .B1(n3996), .B2(n5085), .A(n4880), .ZN(n4010) );
  NAND2_X1 U2846 ( .A1(n4913), .A2(n4046), .ZN(n4927) );
  INV_X1 U2847 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U2848 ( .A1(n4935), .A2(n4018), .ZN(n4946) );
  NOR2_X1 U2849 ( .A1(n2680), .A2(n2679), .ZN(n2678) );
  INV_X1 U2850 ( .A(n2681), .ZN(n2679) );
  OR2_X1 U2851 ( .A1(n3588), .A2(n3819), .ZN(n4115) );
  OR2_X1 U2852 ( .A1(n4131), .A2(n4108), .ZN(n4099) );
  OAI21_X1 U2853 ( .B1(n3531), .B2(n2663), .A(n2661), .ZN(n4126) );
  NAND2_X1 U2854 ( .A1(n4133), .A2(n4132), .ZN(n4131) );
  AND2_X1 U2855 ( .A1(n3552), .A2(n3551), .ZN(n4120) );
  AND2_X1 U2856 ( .A1(n2619), .A2(n4149), .ZN(n2618) );
  NAND2_X1 U2857 ( .A1(n4189), .A2(n3507), .ZN(n3564) );
  NAND2_X1 U2858 ( .A1(n4200), .A2(n4191), .ZN(n4190) );
  NAND2_X1 U2859 ( .A1(n3128), .A2(REG3_REG_22__SCAN_IN), .ZN(n3177) );
  INV_X1 U2860 ( .A(n3129), .ZN(n3128) );
  NAND2_X1 U2861 ( .A1(n3081), .A2(REG3_REG_21__SCAN_IN), .ZN(n3129) );
  INV_X1 U2862 ( .A(n3082), .ZN(n3081) );
  NAND2_X1 U2863 ( .A1(n3526), .A2(n3846), .ZN(n4156) );
  AND2_X1 U2864 ( .A1(n4199), .A2(n3538), .ZN(n4200) );
  NAND2_X1 U2865 ( .A1(n3069), .A2(REG3_REG_20__SCAN_IN), .ZN(n3082) );
  INV_X1 U2866 ( .A(n3070), .ZN(n3069) );
  NOR2_X1 U2867 ( .A1(n5202), .A2(n4224), .ZN(n4199) );
  AND2_X1 U2868 ( .A1(n3842), .A2(n3522), .ZN(n4221) );
  NAND2_X1 U2869 ( .A1(n3055), .A2(REG3_REG_19__SCAN_IN), .ZN(n3070) );
  NAND2_X1 U2870 ( .A1(n3516), .A2(n2641), .ZN(n5207) );
  OR2_X1 U2871 ( .A1(n5205), .A2(n5215), .ZN(n5202) );
  INV_X1 U2872 ( .A(n3041), .ZN(n3042) );
  NAND2_X1 U2873 ( .A1(n3516), .A2(n3872), .ZN(n4229) );
  NAND2_X1 U2874 ( .A1(n4256), .A2(n4233), .ZN(n5205) );
  AOI21_X1 U2875 ( .B1(n2570), .B2(n2572), .A(n2567), .ZN(n2566) );
  NAND2_X1 U2876 ( .A1(n4286), .A2(n2570), .ZN(n2568) );
  INV_X1 U2877 ( .A(n3841), .ZN(n2567) );
  NAND2_X1 U2878 ( .A1(n2563), .A2(n2689), .ZN(n4252) );
  NAND2_X1 U2879 ( .A1(n3493), .A2(n2560), .ZN(n2563) );
  NOR2_X1 U2880 ( .A1(n2690), .A2(n2561), .ZN(n2560) );
  INV_X1 U2881 ( .A(n3492), .ZN(n2561) );
  NAND2_X1 U2882 ( .A1(n4285), .A2(n2502), .ZN(n4275) );
  NOR2_X1 U2883 ( .A1(n4275), .A2(n4253), .ZN(n4256) );
  NAND2_X1 U2884 ( .A1(n4286), .A2(n2573), .ZN(n2569) );
  NAND2_X1 U2885 ( .A1(n4285), .A2(n2617), .ZN(n4273) );
  INV_X1 U2886 ( .A(n5162), .ZN(n3511) );
  NAND2_X1 U2887 ( .A1(n4286), .A2(n3837), .ZN(n3513) );
  INV_X1 U2888 ( .A(n4293), .ZN(n3474) );
  AOI21_X1 U2889 ( .B1(n3420), .B2(n2578), .A(n2576), .ZN(n2575) );
  NAND2_X1 U2890 ( .A1(n2577), .A2(n3912), .ZN(n2576) );
  NAND2_X1 U2891 ( .A1(n2578), .A2(n2581), .ZN(n2577) );
  NAND2_X1 U2892 ( .A1(n3836), .A2(n4293), .ZN(n4286) );
  AND2_X1 U2893 ( .A1(n3837), .A2(n3946), .ZN(n4293) );
  NAND2_X1 U2894 ( .A1(n4285), .A2(n4290), .ZN(n4284) );
  INV_X1 U2895 ( .A(n5158), .ZN(n3775) );
  AND2_X1 U2896 ( .A1(n3436), .A2(n3435), .ZN(n4285) );
  AND2_X1 U2897 ( .A1(n2951), .A2(REG3_REG_11__SCAN_IN), .ZN(n2960) );
  NAND2_X1 U2898 ( .A1(n3420), .A2(n3909), .ZN(n3423) );
  NOR2_X1 U2899 ( .A1(n5112), .A2(n3433), .ZN(n3436) );
  OR2_X1 U2900 ( .A1(n5114), .A2(n5115), .ZN(n5112) );
  OR2_X1 U2901 ( .A1(n2921), .A2(n4435), .ZN(n2937) );
  INV_X1 U2902 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U2903 ( .A1(n2585), .A2(n3945), .ZN(n5095) );
  NAND2_X1 U2904 ( .A1(n3419), .A2(n3938), .ZN(n2585) );
  NAND2_X1 U2905 ( .A1(n2533), .A2(n2538), .ZN(n3415) );
  NAND2_X1 U2906 ( .A1(n3386), .A2(n2540), .ZN(n2533) );
  NAND2_X1 U2907 ( .A1(n2530), .A2(n2534), .ZN(n5097) );
  OR2_X1 U2908 ( .A1(n3386), .A2(n2536), .ZN(n2530) );
  NAND2_X1 U2909 ( .A1(n5093), .A2(n5092), .ZN(n5114) );
  NAND2_X1 U2910 ( .A1(n2644), .A2(n2645), .ZN(n3418) );
  AOI21_X1 U2911 ( .B1(n2648), .B2(n2647), .A(n2646), .ZN(n2645) );
  NAND2_X1 U2912 ( .A1(n3339), .A2(n2648), .ZN(n2644) );
  INV_X1 U2913 ( .A(n3936), .ZN(n2647) );
  AND3_X1 U2914 ( .A1(n2500), .A2(n3368), .A3(n3406), .ZN(n5093) );
  NAND2_X1 U2915 ( .A1(n2906), .A2(REG3_REG_7__SCAN_IN), .ZN(n2908) );
  OR2_X1 U2916 ( .A1(n2908), .A2(n4416), .ZN(n2921) );
  NAND2_X1 U2917 ( .A1(n2650), .A2(n3904), .ZN(n3381) );
  NAND2_X1 U2918 ( .A1(n2651), .A2(n3936), .ZN(n2650) );
  INV_X1 U2919 ( .A(n3339), .ZN(n2651) );
  NAND2_X1 U2920 ( .A1(n3368), .A2(n2616), .ZN(n3346) );
  INV_X1 U2921 ( .A(n3374), .ZN(n3367) );
  NAND2_X1 U2922 ( .A1(n3368), .A2(n3367), .ZN(n3366) );
  NAND2_X1 U2923 ( .A1(n3303), .A2(n3931), .ZN(n3373) );
  NOR2_X1 U2924 ( .A1(n2806), .A2(n4616), .ZN(n2892) );
  OR2_X1 U2925 ( .A1(n3296), .A2(n3309), .ZN(n3356) );
  OR2_X1 U2926 ( .A1(n2635), .A2(n2596), .ZN(n3282) );
  NOR2_X1 U2927 ( .A1(n3238), .A2(n2636), .ZN(n2596) );
  INV_X1 U2928 ( .A(n3923), .ZN(n2636) );
  INV_X1 U2929 ( .A(n5120), .ZN(n5212) );
  NAND2_X1 U2930 ( .A1(n3238), .A2(n5032), .ZN(n5039) );
  AND2_X1 U2931 ( .A1(n5011), .A2(n3240), .ZN(n2747) );
  AND2_X1 U2932 ( .A1(n4807), .A2(n3247), .ZN(n5120) );
  OR2_X1 U2933 ( .A1(n5014), .A2(n5004), .ZN(n5029) );
  INV_X1 U2934 ( .A(n5252), .ZN(n5204) );
  INV_X1 U2936 ( .A(n4767), .ZN(n3108) );
  INV_X1 U2937 ( .A(IR_REG_29__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U2938 ( .A1(n2513), .A2(n2759), .ZN(n2694) );
  INV_X1 U2939 ( .A(IR_REG_28__SCAN_IN), .ZN(n4681) );
  NAND2_X1 U2940 ( .A1(n2612), .A2(n2611), .ZN(n2773) );
  NAND2_X1 U2941 ( .A1(IR_REG_31__SCAN_IN), .A2(n2771), .ZN(n2611) );
  NAND2_X1 U2942 ( .A1(n2613), .A2(IR_REG_22__SCAN_IN), .ZN(n2612) );
  AND2_X1 U2943 ( .A1(n2643), .A2(n2695), .ZN(n2980) );
  INV_X1 U2944 ( .A(IR_REG_3__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U2945 ( .A1(n3694), .A2(n3695), .ZN(n3693) );
  NAND2_X1 U2946 ( .A1(n3769), .A2(n2989), .ZN(n3694) );
  INV_X1 U2947 ( .A(n3632), .ZN(n4166) );
  NOR2_X1 U2948 ( .A1(n3448), .A2(n3449), .ZN(n3447) );
  NAND2_X1 U2949 ( .A1(n3738), .A2(n2698), .ZN(n2600) );
  NAND2_X1 U2950 ( .A1(n3674), .A2(n2917), .ZN(n3393) );
  INV_X1 U2951 ( .A(n4253), .ZN(n3742) );
  OAI22_X1 U2952 ( .A1(n3651), .A2(n4164), .B1(n3650), .B2(n4149), .ZN(n3751)
         );
  INV_X1 U2953 ( .A(n5163), .ZN(n3743) );
  AOI21_X1 U2954 ( .B1(n2601), .B2(n2604), .A(n2520), .ZN(n2599) );
  OR2_X1 U2955 ( .A1(n2723), .A2(n2609), .ZN(n3771) );
  NOR2_X1 U2956 ( .A1(n3447), .A2(n2950), .ZN(n3456) );
  NAND2_X1 U2957 ( .A1(n2856), .A2(n2858), .ZN(n2859) );
  OR2_X1 U2958 ( .A1(n3135), .A2(n4807), .ZN(n3809) );
  OR2_X1 U2959 ( .A1(n2891), .A2(n2890), .ZN(n2605) );
  INV_X1 U2960 ( .A(n3809), .ZN(n5161) );
  INV_X1 U2961 ( .A(n5177), .ZN(n3796) );
  INV_X1 U2962 ( .A(n3810), .ZN(n5159) );
  OR2_X1 U2963 ( .A1(n3135), .A2(n3127), .ZN(n3810) );
  AND4_X1 U2964 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n4205)
         );
  AND4_X1 U2965 ( .A1(n3076), .A2(n3075), .A3(n3074), .A4(n3073), .ZN(n5211)
         );
  OR2_X1 U2966 ( .A1(n3009), .A2(n3008), .ZN(n4287) );
  OR2_X1 U2967 ( .A1(n2790), .A2(n2765), .ZN(n3984) );
  INV_X1 U2968 ( .A(n3480), .ZN(n4288) );
  NAND4_X1 U2969 ( .A1(n2944), .A2(n2943), .A3(n2942), .A4(n2941), .ZN(n5119)
         );
  NAND4_X1 U2970 ( .A1(n2868), .A2(n2867), .A3(n2866), .A4(n2865), .ZN(n5034)
         );
  OR2_X1 U2971 ( .A1(n2840), .A2(n5044), .ZN(n2822) );
  NAND2_X1 U2972 ( .A1(n4978), .A2(n4977), .ZN(n4976) );
  XNOR2_X1 U2973 ( .A(n4000), .B(n4029), .ZN(n4829) );
  NAND2_X1 U2974 ( .A1(n4829), .A2(REG1_REG_3__SCAN_IN), .ZN(n4828) );
  XNOR2_X1 U2975 ( .A(n4032), .B(n4033), .ZN(n4996) );
  NAND2_X1 U2976 ( .A1(n4915), .A2(n4013), .ZN(n4924) );
  NOR2_X1 U2977 ( .A1(n2742), .A2(n4015), .ZN(n4923) );
  XNOR2_X1 U2978 ( .A(n4017), .B(n4016), .ZN(n4936) );
  NAND2_X1 U2979 ( .A1(n4936), .A2(REG1_REG_14__SCAN_IN), .ZN(n4935) );
  INV_X1 U2980 ( .A(n4816), .ZN(n4992) );
  NAND2_X1 U2981 ( .A1(n4938), .A2(n4049), .ZN(n4951) );
  NOR2_X1 U2982 ( .A1(n4074), .A2(n4073), .ZN(n4078) );
  NOR2_X1 U2983 ( .A1(n4066), .A2(n4065), .ZN(n4068) );
  INV_X1 U2984 ( .A(n2628), .ZN(n4960) );
  AND2_X1 U2985 ( .A1(n3595), .A2(n2743), .ZN(n4314) );
  XNOR2_X1 U2986 ( .A(n3510), .B(n3509), .ZN(n4322) );
  NAND2_X1 U2987 ( .A1(n3508), .A2(n3548), .ZN(n3510) );
  AND2_X1 U2988 ( .A1(n4185), .A2(n4184), .ZN(n4329) );
  NAND2_X1 U2989 ( .A1(n3505), .A2(n3504), .ZN(n4187) );
  INV_X1 U2990 ( .A(n2553), .ZN(n2552) );
  NAND2_X1 U2991 ( .A1(n2672), .A2(n3498), .ZN(n5200) );
  NAND2_X1 U2992 ( .A1(n4227), .A2(n3885), .ZN(n2672) );
  INV_X1 U2993 ( .A(n3494), .ZN(n4264) );
  NAND2_X1 U2994 ( .A1(n2556), .A2(n3434), .ZN(n3472) );
  NAND2_X1 U2995 ( .A1(n3432), .A2(n3431), .ZN(n2556) );
  NAND2_X1 U2996 ( .A1(n2537), .A2(n2540), .ZN(n3412) );
  OR2_X1 U2997 ( .A1(n3386), .A2(n3385), .ZN(n2537) );
  NAND2_X1 U2998 ( .A1(n3364), .A2(n3315), .ZN(n3338) );
  NAND2_X1 U2999 ( .A1(n3311), .A2(n3310), .ZN(n3351) );
  NAND2_X1 U3000 ( .A1(n5140), .A2(n5227), .ZN(n4282) );
  INV_X1 U3001 ( .A(n5224), .ZN(n5135) );
  AND2_X1 U3002 ( .A1(n3970), .A2(n2504), .ZN(n5240) );
  OR2_X1 U3003 ( .A1(n3229), .A2(n4312), .ZN(n3230) );
  INV_X1 U3004 ( .A(n4278), .ZN(n4260) );
  OAI21_X1 U3005 ( .B1(n4306), .B2(n5144), .A(n2499), .ZN(n4345) );
  INV_X1 U3006 ( .A(n3624), .ZN(n4305) );
  INV_X2 U3007 ( .A(n5257), .ZN(n5259) );
  XNOR2_X1 U3008 ( .A(n2564), .B(IR_REG_30__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U3009 ( .A1(n4763), .A2(IR_REG_31__SCAN_IN), .ZN(n2564) );
  AND2_X1 U3010 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2656)
         );
  XNOR2_X1 U3011 ( .A(n2796), .B(IR_REG_26__SCAN_IN), .ZN(n4767) );
  XNOR2_X1 U3012 ( .A(n2762), .B(n2759), .ZN(n3140) );
  NAND2_X1 U3013 ( .A1(n2753), .A2(IR_REG_31__SCAN_IN), .ZN(n2754) );
  AND2_X1 U3014 ( .A1(n3158), .A2(STATE_REG_SCAN_IN), .ZN(n4777) );
  NOR2_X1 U3015 ( .A1(n2614), .A2(n2869), .ZN(n2945) );
  NAND2_X1 U3016 ( .A1(n2823), .A2(IR_REG_2__SCAN_IN), .ZN(n2623) );
  AOI21_X1 U3017 ( .B1(n2761), .B2(n4445), .A(n2496), .ZN(n2622) );
  NAND2_X1 U3018 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2633)
         );
  NAND2_X1 U3019 ( .A1(n2497), .A2(n2632), .ZN(n2631) );
  NAND2_X1 U3020 ( .A1(n2715), .A2(n5172), .ZN(n2713) );
  NAND2_X1 U3021 ( .A1(n4965), .A2(n2624), .ZN(U3258) );
  AOI21_X1 U3022 ( .B1(n2627), .B2(n4957), .A(n2625), .ZN(n2624) );
  OAI21_X1 U3023 ( .B1(n4958), .B2(n4959), .A(n2626), .ZN(n2625) );
  INV_X1 U3024 ( .A(n2958), .ZN(n3642) );
  AND2_X1 U3025 ( .A1(n3935), .A2(n3933), .ZN(n3873) );
  AND2_X1 U3026 ( .A1(n3127), .A2(IR_REG_0__SCAN_IN), .ZN(n2498) );
  AND2_X1 U3027 ( .A1(n4305), .A2(n4304), .ZN(n2499) );
  AND2_X1 U3028 ( .A1(n2616), .A2(n3341), .ZN(n2500) );
  NAND2_X1 U3029 ( .A1(n3738), .A2(n3740), .ZN(n3739) );
  INV_X2 U3030 ( .A(n2800), .ZN(n3828) );
  AND2_X1 U3031 ( .A1(n4200), .A2(n2619), .ZN(n2501) );
  NAND2_X1 U3032 ( .A1(n2568), .A2(n2566), .ZN(n4246) );
  AND2_X1 U3033 ( .A1(n2617), .A2(n3514), .ZN(n2502) );
  OAI21_X1 U3034 ( .B1(n3048), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2803) );
  AND2_X1 U3035 ( .A1(n2532), .A2(n2531), .ZN(n2503) );
  AND2_X1 U3036 ( .A1(n3233), .A2(n3886), .ZN(n2504) );
  OAI21_X1 U3037 ( .B1(n3516), .B2(n2640), .A(n2637), .ZN(n4213) );
  NAND2_X1 U3038 ( .A1(n2495), .A2(n4765), .ZN(n2830) );
  NAND2_X1 U3039 ( .A1(n2600), .A2(n2696), .ZN(n3712) );
  NAND2_X1 U3040 ( .A1(n2552), .A2(n2554), .ZN(n4198) );
  NAND2_X1 U3041 ( .A1(n3739), .A2(n3040), .ZN(n3791) );
  INV_X1 U3042 ( .A(n5028), .ZN(n2824) );
  OR2_X1 U3043 ( .A1(n5096), .A2(n2691), .ZN(n2505) );
  INV_X1 U3044 ( .A(IR_REG_30__SCAN_IN), .ZN(n4680) );
  AND2_X1 U3045 ( .A1(n3675), .A2(n2737), .ZN(n2506) );
  AND2_X1 U3046 ( .A1(n3988), .A2(n3681), .ZN(n2507) );
  AND4_X1 U3047 ( .A1(n4475), .A2(n4669), .A3(n4464), .A4(n4480), .ZN(n2508)
         );
  NAND2_X1 U3048 ( .A1(n3706), .A2(n2721), .ZN(n3748) );
  INV_X1 U3049 ( .A(IR_REG_2__SCAN_IN), .ZN(n4445) );
  OR2_X1 U3050 ( .A1(n5027), .A2(n3999), .ZN(n2509) );
  AND2_X1 U3051 ( .A1(n2905), .A2(n2904), .ZN(n2510) );
  NOR2_X1 U3052 ( .A1(n2649), .A2(n3380), .ZN(n2648) );
  NAND2_X1 U3053 ( .A1(n2661), .A2(n3850), .ZN(n2511) );
  AND2_X1 U3054 ( .A1(n2663), .A2(n3850), .ZN(n2512) );
  AND2_X1 U3055 ( .A1(n4487), .A2(n2795), .ZN(n2513) );
  INV_X1 U3056 ( .A(IR_REG_19__SCAN_IN), .ZN(n2804) );
  OR2_X1 U3057 ( .A1(n3562), .A2(n3561), .ZN(n2514) );
  INV_X1 U3058 ( .A(n2594), .ZN(n3531) );
  NAND2_X1 U3059 ( .A1(n3526), .A2(n2591), .ZN(n2594) );
  INV_X1 U3060 ( .A(n2725), .ZN(n2724) );
  NAND2_X1 U3061 ( .A1(n2728), .A2(n2726), .ZN(n2725) );
  INV_X1 U3062 ( .A(IR_REG_27__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U3063 ( .A1(n2720), .A2(n3686), .ZN(n2515) );
  XNOR2_X1 U3064 ( .A(n2754), .B(IR_REG_24__SCAN_IN), .ZN(n3093) );
  INV_X1 U3065 ( .A(IR_REG_5__SCAN_IN), .ZN(n4643) );
  NAND2_X1 U3066 ( .A1(n2695), .A2(n2496), .ZN(n2957) );
  OAI21_X1 U3067 ( .B1(n2957), .B2(n2767), .A(IR_REG_31__SCAN_IN), .ZN(n3010)
         );
  OAI21_X1 U3068 ( .B1(n3018), .B2(IR_REG_16__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n3035) );
  NAND2_X1 U3069 ( .A1(n2772), .A2(IR_REG_31__SCAN_IN), .ZN(n2764) );
  NAND2_X1 U3070 ( .A1(n2569), .A2(n3944), .ZN(n4265) );
  XOR2_X1 U3071 ( .A(n3011), .B(n2958), .Z(n2516) );
  XOR2_X1 U3072 ( .A(n2959), .B(n2958), .Z(n2517) );
  OAI21_X1 U3073 ( .B1(n3432), .B2(n2559), .A(n2557), .ZN(n4292) );
  AND2_X1 U3074 ( .A1(n3674), .A2(n2735), .ZN(n2518) );
  AND2_X1 U3075 ( .A1(n5119), .A2(n5102), .ZN(n2519) );
  INV_X1 U3076 ( .A(n3435), .ZN(n3777) );
  INV_X1 U3077 ( .A(n3473), .ZN(n4290) );
  NOR2_X1 U3078 ( .A1(n3067), .A2(n3066), .ZN(n2520) );
  NAND2_X1 U3079 ( .A1(n4200), .A2(n2618), .ZN(n2620) );
  INV_X1 U3080 ( .A(IR_REG_22__SCAN_IN), .ZN(n2771) );
  NOR2_X1 U3081 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2927)
         );
  INV_X1 U3082 ( .A(n4027), .ZN(n5059) );
  OR2_X1 U3083 ( .A1(n4288), .A2(n3777), .ZN(n2521) );
  AND2_X1 U3084 ( .A1(n5209), .A2(n2673), .ZN(n2522) );
  NOR2_X1 U3085 ( .A1(n2723), .A2(n2724), .ZN(n2523) );
  AND2_X1 U3086 ( .A1(n3528), .A2(n3506), .ZN(n4186) );
  INV_X1 U3087 ( .A(n4186), .ZN(n2682) );
  INV_X1 U3088 ( .A(n3413), .ZN(n3406) );
  INV_X1 U3089 ( .A(n3498), .ZN(n2674) );
  INV_X1 U3090 ( .A(n3815), .ZN(n5172) );
  AND2_X1 U3091 ( .A1(n2500), .A2(n3368), .ZN(n2524) );
  NAND4_X1 U3092 ( .A1(n2834), .A2(n2833), .A3(n2832), .A4(n2831), .ZN(n3992)
         );
  INV_X1 U3093 ( .A(n3945), .ZN(n2588) );
  OR2_X1 U3094 ( .A1(n4930), .A2(n4014), .ZN(n2525) );
  INV_X1 U3095 ( .A(n3519), .ZN(n4224) );
  NAND2_X1 U3096 ( .A1(n4231), .A2(n3742), .ZN(n2526) );
  OR2_X1 U3097 ( .A1(n3363), .A2(n3873), .ZN(n3364) );
  INV_X1 U3098 ( .A(n3939), .ZN(n2646) );
  NAND2_X1 U3099 ( .A1(n3676), .A2(n3675), .ZN(n3674) );
  OR2_X1 U3100 ( .A1(n4909), .A2(n5139), .ZN(n2527) );
  OR2_X1 U3101 ( .A1(n4909), .A2(n3994), .ZN(n2528) );
  AND2_X1 U3102 ( .A1(n3415), .A2(n3414), .ZN(n2529) );
  NAND2_X1 U3103 ( .A1(n2657), .A2(n2655), .ZN(n3143) );
  NAND2_X1 U3104 ( .A1(n3235), .A2(n3234), .ZN(n5008) );
  INV_X1 U3105 ( .A(n2565), .ZN(n5032) );
  NAND2_X1 U3106 ( .A1(n3925), .A2(n3923), .ZN(n2565) );
  NAND2_X1 U3107 ( .A1(n3386), .A2(n2534), .ZN(n2532) );
  NAND2_X1 U3108 ( .A1(n2545), .A2(n2541), .ZN(n3314) );
  INV_X1 U3109 ( .A(n2675), .ZN(n2547) );
  NAND2_X1 U3110 ( .A1(n2547), .A2(n2550), .ZN(n2549) );
  NAND2_X1 U3111 ( .A1(n3501), .A2(n3500), .ZN(n4212) );
  INV_X1 U3112 ( .A(n4292), .ZN(n3475) );
  INV_X1 U3113 ( .A(n4252), .ZN(n2562) );
  INV_X1 U3114 ( .A(n2575), .ZN(n3836) );
  NAND2_X1 U3115 ( .A1(n3419), .A2(n2586), .ZN(n2584) );
  NAND2_X2 U3116 ( .A1(n4766), .A2(n4765), .ZN(n2842) );
  NAND2_X1 U3117 ( .A1(n3738), .A2(n2601), .ZN(n2598) );
  NAND2_X1 U3118 ( .A1(n2598), .A2(n2599), .ZN(n3757) );
  AOI21_X2 U3119 ( .B1(n3331), .B2(n3330), .A(n2510), .ZN(n3676) );
  NAND2_X2 U3120 ( .A1(n3272), .A2(n2605), .ZN(n3331) );
  NAND2_X2 U3121 ( .A1(n3273), .A2(n3274), .ZN(n3272) );
  NAND2_X1 U3122 ( .A1(n2723), .A2(n2973), .ZN(n2608) );
  NAND2_X2 U3123 ( .A1(n2608), .A2(n2606), .ZN(n3769) );
  NAND3_X1 U3124 ( .A1(n3720), .A2(n3719), .A3(n3749), .ZN(n3803) );
  NAND2_X2 U3125 ( .A1(n2610), .A2(n3640), .ZN(n3749) );
  NOR2_X2 U3126 ( .A1(n2614), .A2(IR_REG_10__SCAN_IN), .ZN(n2695) );
  NAND4_X1 U3127 ( .A1(n2927), .A2(n2749), .A3(n2750), .A4(n2748), .ZN(n2614)
         );
  NAND2_X1 U3128 ( .A1(n2654), .A2(DATAI_1_), .ZN(n2615) );
  INV_X1 U3129 ( .A(n2620), .ZN(n4148) );
  XNOR2_X1 U3130 ( .A(n4010), .B(n4041), .ZN(n4895) );
  XNOR2_X1 U3131 ( .A(n4005), .B(n4004), .ZN(n4853) );
  XNOR2_X1 U3132 ( .A(n4045), .B(n5143), .ZN(n4914) );
  OAI21_X1 U3133 ( .B1(n5032), .B2(n2636), .A(n3875), .ZN(n2635) );
  NAND4_X1 U3134 ( .A1(n2643), .A2(n2758), .A3(n2759), .A4(n2695), .ZN(n2779)
         );
  NAND3_X1 U3135 ( .A1(n2643), .A2(n2758), .A3(n2695), .ZN(n2760) );
  NAND2_X1 U3136 ( .A1(n2797), .A2(n2656), .ZN(n2655) );
  NOR2_X1 U3137 ( .A1(n2659), .A2(n2658), .ZN(n2657) );
  NAND2_X1 U3138 ( .A1(n2669), .A2(n3956), .ZN(n4143) );
  INV_X1 U3139 ( .A(n3959), .ZN(n2670) );
  NAND2_X1 U3140 ( .A1(n2671), .A2(n2522), .ZN(n3501) );
  NAND3_X1 U3141 ( .A1(n3497), .A2(n3498), .A3(n3496), .ZN(n2671) );
  INV_X1 U3142 ( .A(n3237), .ZN(n3188) );
  NAND2_X1 U3143 ( .A1(n3363), .A2(n2685), .ZN(n2684) );
  NAND2_X1 U3144 ( .A1(n2684), .A2(n2683), .ZN(n3386) );
  NAND2_X1 U3145 ( .A1(n3494), .A2(n2689), .ZN(n2688) );
  NOR2_X1 U3146 ( .A1(n2760), .A2(n2692), .ZN(n2781) );
  NAND2_X1 U3147 ( .A1(n3769), .A2(n2704), .ZN(n2703) );
  OAI21_X2 U31480 ( .B1(n3048), .B2(n2708), .A(IR_REG_31__SCAN_IN), .ZN(n2710)
         );
  NAND2_X1 U31490 ( .A1(n3687), .A2(n2712), .ZN(n2711) );
  OAI211_X1 U3150 ( .C1(n3687), .C2(n2713), .A(n2711), .B(n3673), .ZN(U3217)
         );
  NAND2_X1 U3151 ( .A1(n3687), .A2(n3686), .ZN(n3685) );
  INV_X1 U3152 ( .A(n3668), .ZN(n2720) );
  NAND2_X2 U3153 ( .A1(n3703), .A2(n3635), .ZN(n3706) );
  NOR2_X2 U3154 ( .A1(n3448), .A2(n2729), .ZN(n2723) );
  OR2_X1 U3155 ( .A1(n2781), .A2(n2761), .ZN(n2780) );
  NAND2_X1 U3156 ( .A1(n2843), .A2(REG1_REG_1__SCAN_IN), .ZN(n2844) );
  NAND2_X1 U3157 ( .A1(n3564), .A2(n4163), .ZN(n4162) );
  INV_X1 U3158 ( .A(n2857), .ZN(n2858) );
  NAND2_X1 U3159 ( .A1(n5169), .A2(n5170), .ZN(n3730) );
  INV_X4 U3160 ( .A(n2828), .ZN(n3665) );
  OR2_X1 U3161 ( .A1(n2798), .A2(n2761), .ZN(n2799) );
  NAND2_X1 U3162 ( .A1(n2779), .A2(IR_REG_31__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U3163 ( .A1(n2838), .A2(n3642), .ZN(n2839) );
  NAND2_X1 U3164 ( .A1(n2784), .A2(n4766), .ZN(n2864) );
  NAND2_X1 U3165 ( .A1(n3230), .A2(n5224), .ZN(n4242) );
  INV_X1 U3166 ( .A(n5249), .ZN(n5140) );
  OR2_X1 U3167 ( .A1(n4930), .A2(n3438), .ZN(n2738) );
  AND2_X1 U3168 ( .A1(n2888), .A2(n2887), .ZN(n2739) );
  OR2_X1 U3169 ( .A1(n2957), .A2(n2996), .ZN(n2740) );
  INV_X1 U3170 ( .A(n4891), .ZN(n4041) );
  NAND2_X1 U3171 ( .A1(n3010), .A2(n2768), .ZN(n3018) );
  OR2_X1 U3172 ( .A1(n2790), .A2(n2837), .ZN(n2741) );
  AND2_X1 U3173 ( .A1(n4930), .A2(n4014), .ZN(n2742) );
  AND2_X1 U3174 ( .A1(n3594), .A2(n3593), .ZN(n2743) );
  AND3_X1 U3175 ( .A1(n2821), .A2(n2820), .A3(n2819), .ZN(n2744) );
  AND2_X1 U3176 ( .A1(n3895), .A2(n3929), .ZN(n2745) );
  AND4_X1 U3177 ( .A1(n2757), .A2(n2756), .A3(n4669), .A4(n4464), .ZN(n2746)
         );
  NAND2_X1 U3178 ( .A1(n3063), .A2(n5014), .ZN(n2853) );
  OR2_X1 U3179 ( .A1(n3560), .A2(n3559), .ZN(n3561) );
  OAI21_X1 U3180 ( .B1(n4104), .B2(n3588), .A(n3587), .ZN(n3606) );
  AND2_X1 U3181 ( .A1(n3884), .A2(n3575), .ZN(n3856) );
  INV_X1 U3182 ( .A(n4028), .ZN(n4029) );
  NOR2_X1 U3183 ( .A1(n4930), .A2(n4014), .ZN(n4015) );
  INV_X1 U3184 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4616) );
  INV_X1 U3185 ( .A(n3856), .ZN(n3958) );
  OR2_X1 U3186 ( .A1(n2996), .A2(IR_REG_14__SCAN_IN), .ZN(n2767) );
  INV_X1 U3187 ( .A(DATAI_1_), .ZN(n2849) );
  OR2_X1 U3188 ( .A1(n3212), .A2(n3211), .ZN(n3567) );
  NOR2_X1 U3189 ( .A1(n3108), .A2(n3140), .ZN(n2763) );
  NAND2_X1 U3190 ( .A1(n4895), .A2(REG1_REG_10__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U3191 ( .A1(n4914), .A2(REG2_REG_12__SCAN_IN), .ZN(n4913) );
  NOR2_X1 U3192 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  OR2_X1 U3193 ( .A1(n3196), .A2(n3752), .ZN(n3212) );
  AND2_X1 U3194 ( .A1(n2960), .A2(REG3_REG_12__SCAN_IN), .ZN(n2974) );
  INV_X1 U3195 ( .A(n5126), .ZN(n3416) );
  INV_X1 U3196 ( .A(n4240), .ZN(n4233) );
  OAI21_X1 U3197 ( .B1(n3718), .B2(n3653), .A(n3652), .ZN(n3656) );
  MUX2_X1 U3198 ( .A(DATAI_10_), .B(n4891), .S(n3828), .Z(n5102) );
  INV_X1 U3199 ( .A(n4287), .ZN(n4267) );
  NOR2_X1 U3200 ( .A1(n3263), .A2(n2739), .ZN(n3273) );
  NAND2_X1 U3201 ( .A1(n2974), .A2(REG3_REG_13__SCAN_IN), .ZN(n2991) );
  OR2_X1 U3202 ( .A1(n2842), .A2(n3669), .ZN(n3583) );
  INV_X1 U3203 ( .A(n4851), .ZN(n4004) );
  INV_X1 U3204 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4416) );
  OR2_X1 U3205 ( .A1(n3579), .A2(n4417), .ZN(n3620) );
  OR2_X1 U3206 ( .A1(n3550), .A2(n3549), .ZN(n4121) );
  AND2_X1 U3207 ( .A1(n3915), .A2(n3909), .ZN(n5126) );
  INV_X1 U3208 ( .A(n5210), .ZN(n5117) );
  INV_X1 U3209 ( .A(n3433), .ZN(n3467) );
  INV_X1 U32100 ( .A(n5240), .ZN(n5123) );
  INV_X1 U32110 ( .A(n5008), .ZN(n5217) );
  INV_X1 U32120 ( .A(n3657), .ZN(n4108) );
  INV_X1 U32130 ( .A(n5102), .ZN(n5092) );
  INV_X1 U32140 ( .A(n3663), .ZN(n3672) );
  INV_X1 U32150 ( .A(n4149), .ZN(n4147) );
  NAND2_X1 U32160 ( .A1(n3121), .A2(n5224), .ZN(n5163) );
  AND4_X1 U32170 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n4106)
         );
  OR2_X1 U32180 ( .A1(n2842), .A2(n4150), .ZN(n3200) );
  OR2_X1 U32190 ( .A1(n2830), .A2(n2862), .ZN(n2868) );
  OR2_X1 U32200 ( .A1(n3157), .A2(n3156), .ZN(n4022) );
  NAND2_X1 U32210 ( .A1(n4853), .A2(REG1_REG_6__SCAN_IN), .ZN(n4852) );
  INV_X1 U32220 ( .A(n4958), .ZN(n4990) );
  INV_X1 U32230 ( .A(n3891), .ZN(n3604) );
  NAND2_X1 U32240 ( .A1(n3586), .A2(n3889), .ZN(n3595) );
  AND2_X1 U32250 ( .A1(n5252), .A2(n3112), .ZN(n4311) );
  NAND2_X1 U32260 ( .A1(n3110), .A2(n3153), .ZN(n4342) );
  NAND2_X1 U32270 ( .A1(n3242), .A2(n2958), .ZN(n5144) );
  INV_X1 U32280 ( .A(n5144), .ZN(n5227) );
  OR3_X1 U32290 ( .A1(n4312), .A2(n4311), .A3(n4310), .ZN(n4344) );
  AND2_X1 U32300 ( .A1(n2790), .A2(n4777), .ZN(n3157) );
  NAND2_X1 U32310 ( .A1(n2778), .A2(n2777), .ZN(n3886) );
  AND2_X1 U32320 ( .A1(n2814), .A2(n2898), .ZN(n4027) );
  AND2_X1 U32330 ( .A1(n4022), .A2(n3160), .ZN(n4988) );
  INV_X1 U32340 ( .A(n5014), .ZN(n3236) );
  NAND2_X1 U32350 ( .A1(n3167), .A2(n3116), .ZN(n3815) );
  NAND2_X1 U32360 ( .A1(n3123), .A2(STATE_REG_SCAN_IN), .ZN(n5177) );
  OAI21_X1 U32370 ( .B1(n4257), .B2(n2842), .A(n3034), .ZN(n4231) );
  NAND2_X1 U32380 ( .A1(n4242), .A2(n5219), .ZN(n4278) );
  INV_X1 U32390 ( .A(n3886), .ZN(n4769) );
  NAND2_X2 U32400 ( .A1(n2850), .A2(n4445), .ZN(n2869) );
  NAND2_X1 U32410 ( .A1(n2764), .A2(n4480), .ZN(n2753) );
  INV_X1 U32420 ( .A(IR_REG_25__SCAN_IN), .ZN(n2759) );
  NAND2_X1 U32430 ( .A1(n2760), .A2(IR_REG_31__SCAN_IN), .ZN(n2762) );
  XNOR2_X1 U32440 ( .A(n2764), .B(n4480), .ZN(n3158) );
  INV_X1 U32450 ( .A(n4777), .ZN(n2765) );
  INV_X2 U32460 ( .A(n3984), .ZN(U4043) );
  NOR2_X1 U32470 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2766) );
  NAND2_X1 U32480 ( .A1(n2766), .A2(n2982), .ZN(n2996) );
  INV_X1 U32490 ( .A(IR_REG_15__SCAN_IN), .ZN(n2768) );
  NAND2_X1 U32500 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(
        n2769) );
  NAND2_X1 U32510 ( .A1(n3035), .A2(n2769), .ZN(n3048) );
  NAND2_X1 U32520 ( .A1(n2773), .A2(n2772), .ZN(n3233) );
  INV_X1 U32530 ( .A(n2774), .ZN(n2775) );
  NAND2_X1 U32540 ( .A1(n2775), .A2(IR_REG_31__SCAN_IN), .ZN(n2776) );
  MUX2_X1 U32550 ( .A(IR_REG_31__SCAN_IN), .B(n2776), .S(IR_REG_21__SCAN_IN), 
        .Z(n2778) );
  AND2_X1 U32560 ( .A1(n3113), .A2(n2504), .ZN(n3111) );
  OR2_X4 U32570 ( .A1(n3111), .A2(n2848), .ZN(n3651) );
  NAND2_X1 U32580 ( .A1(n2781), .A2(n4682), .ZN(n4763) );
  NAND2_X1 U32590 ( .A1(n2495), .A2(n2784), .ZN(n2840) );
  NAND2_X1 U32600 ( .A1(n3030), .A2(REG0_REG_8__SCAN_IN), .ZN(n2789) );
  INV_X1 U32610 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2782) );
  OR2_X1 U32620 ( .A1(n3826), .A2(n2782), .ZN(n2788) );
  INV_X1 U32630 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2783) );
  OR2_X1 U32640 ( .A1(n3195), .A2(n2783), .ZN(n2787) );
  NAND2_X1 U32650 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2806) );
  NAND2_X1 U32660 ( .A1(n2908), .A2(n4416), .ZN(n2785) );
  NAND2_X1 U32670 ( .A1(n2921), .A2(n2785), .ZN(n3395) );
  OR2_X1 U32680 ( .A1(n2842), .A2(n3395), .ZN(n2786) );
  NAND4_X1 U32690 ( .A1(n2789), .A2(n2788), .A3(n2787), .A4(n2786), .ZN(n3987)
         );
  INV_X1 U32700 ( .A(n2802), .ZN(n2791) );
  NAND2_X1 U32710 ( .A1(n2748), .A2(n2880), .ZN(n2792) );
  NOR2_X1 U32720 ( .A1(n2869), .A2(n2792), .ZN(n2812) );
  NAND2_X1 U32730 ( .A1(n2812), .A2(n4643), .ZN(n2898) );
  NAND2_X1 U32740 ( .A1(n2929), .A2(IR_REG_31__SCAN_IN), .ZN(n2913) );
  INV_X1 U32750 ( .A(IR_REG_7__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U32760 ( .A1(n2913), .A2(n4647), .ZN(n2793) );
  NAND2_X1 U32770 ( .A1(n2793), .A2(IR_REG_31__SCAN_IN), .ZN(n2794) );
  XNOR2_X1 U32780 ( .A(n2794), .B(IR_REG_8__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U32790 ( .A1(n2796), .A2(n2795), .ZN(n2797) );
  MUX2_X1 U32800 ( .A(DATAI_8_), .B(n4873), .S(n3828), .Z(n3398) );
  AOI22_X1 U32810 ( .A1(n2855), .A2(n3987), .B1(n3665), .B2(n3398), .ZN(n2920)
         );
  INV_X1 U32820 ( .A(n3987), .ZN(n3679) );
  INV_X2 U32830 ( .A(n2848), .ZN(n3063) );
  INV_X1 U32840 ( .A(n3398), .ZN(n3341) );
  OR2_X1 U32850 ( .A1(n2825), .A2(n3341), .ZN(n2801) );
  OAI21_X1 U32860 ( .B1(n3650), .B2(n3679), .A(n2801), .ZN(n2805) );
  XNOR2_X2 U32870 ( .A(n2803), .B(n2804), .ZN(n5219) );
  INV_X1 U32880 ( .A(n3233), .ZN(n4768) );
  NAND2_X1 U32890 ( .A1(n5219), .A2(n4768), .ZN(n3124) );
  NAND2_X4 U32900 ( .A1(n2802), .A2(n3124), .ZN(n2958) );
  XNOR2_X1 U32910 ( .A(n2805), .B(n2958), .ZN(n2918) );
  INV_X1 U32920 ( .A(n2918), .ZN(n2919) );
  NAND2_X1 U32930 ( .A1(n2843), .A2(REG1_REG_5__SCAN_IN), .ZN(n2811) );
  INV_X1 U32940 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3359) );
  OR2_X1 U32950 ( .A1(n3826), .A2(n3359), .ZN(n2810) );
  AND2_X1 U32960 ( .A1(n2806), .A2(n4616), .ZN(n2807) );
  OR2_X1 U32970 ( .A1(n2807), .A2(n2892), .ZN(n3358) );
  OR2_X1 U32980 ( .A1(n2842), .A2(n3358), .ZN(n2809) );
  INV_X1 U32990 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5065) );
  OR2_X1 U33000 ( .A1(n3822), .A2(n5065), .ZN(n2808) );
  OR2_X1 U33010 ( .A1(n2812), .A2(n2761), .ZN(n2813) );
  MUX2_X1 U33020 ( .A(IR_REG_31__SCAN_IN), .B(n2813), .S(IR_REG_5__SCAN_IN), 
        .Z(n2814) );
  MUX2_X1 U33030 ( .A(DATAI_5_), .B(n4027), .S(n3603), .Z(n3357) );
  AOI22_X1 U33040 ( .A1(n2855), .A2(n3990), .B1(n3665), .B2(n3357), .ZN(n2889)
         );
  INV_X1 U33050 ( .A(n2889), .ZN(n2891) );
  INV_X1 U33060 ( .A(n3990), .ZN(n2816) );
  INV_X1 U33070 ( .A(n3357), .ZN(n3903) );
  OR2_X1 U33080 ( .A1(n2825), .A2(n3903), .ZN(n2815) );
  OAI21_X1 U33090 ( .B1(n3650), .B2(n2816), .A(n2815), .ZN(n2817) );
  XNOR2_X1 U33100 ( .A(n2817), .B(n2958), .ZN(n2890) );
  INV_X1 U33110 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3999) );
  OR2_X1 U33120 ( .A1(n2864), .A2(n3999), .ZN(n2821) );
  INV_X1 U33130 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2818) );
  OR2_X1 U33140 ( .A1(n2842), .A2(n2818), .ZN(n2820) );
  NAND2_X1 U33150 ( .A1(n3565), .A2(REG2_REG_2__SCAN_IN), .ZN(n2819) );
  INV_X1 U33160 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5044) );
  NOR2_X1 U33170 ( .A1(n2850), .A2(n2761), .ZN(n2823) );
  MUX2_X1 U33180 ( .A(DATAI_2_), .B(n4975), .S(n3603), .Z(n5028) );
  INV_X1 U33190 ( .A(n5004), .ZN(n3328) );
  INV_X1 U33200 ( .A(IR_REG_0__SCAN_IN), .ZN(n4967) );
  OAI22_X1 U33210 ( .A1(n3328), .A2(n2828), .B1(n2790), .B2(n4967), .ZN(n2829)
         );
  INV_X1 U33220 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3324) );
  OR2_X1 U33230 ( .A1(n2842), .A2(n3324), .ZN(n2834) );
  INV_X1 U33240 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3325) );
  OR2_X1 U33250 ( .A1(n2830), .A2(n3325), .ZN(n2833) );
  INV_X1 U33260 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4737) );
  OR2_X1 U33270 ( .A1(n2840), .A2(n4737), .ZN(n2832) );
  NAND2_X1 U33280 ( .A1(n2843), .A2(REG1_REG_0__SCAN_IN), .ZN(n2831) );
  INV_X1 U33290 ( .A(n3992), .ZN(n3321) );
  NAND2_X1 U33300 ( .A1(n2836), .A2(n2835), .ZN(n3164) );
  INV_X1 U33310 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2837) );
  NAND2_X1 U33320 ( .A1(n2838), .A2(n2741), .ZN(n3165) );
  NAND2_X1 U33330 ( .A1(n3164), .A2(n3165), .ZN(n3163) );
  NAND2_X1 U33340 ( .A1(n3163), .A2(n2839), .ZN(n3172) );
  INV_X1 U33350 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5020) );
  OR2_X1 U33360 ( .A1(n2840), .A2(n5020), .ZN(n2847) );
  INV_X1 U33370 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2841) );
  INV_X1 U33380 ( .A(n2850), .ZN(n2851) );
  INV_X1 U33390 ( .A(n5003), .ZN(n4820) );
  OAI21_X1 U33400 ( .B1(n3188), .B2(n2828), .A(n2853), .ZN(n2854) );
  XNOR2_X1 U33410 ( .A(n2854), .B(n2958), .ZN(n2856) );
  XNOR2_X1 U33420 ( .A(n2856), .B(n2857), .ZN(n3170) );
  NAND2_X1 U33430 ( .A1(n3172), .A2(n3170), .ZN(n3171) );
  NAND2_X1 U33440 ( .A1(n3171), .A2(n2859), .ZN(n3186) );
  XNOR2_X1 U33450 ( .A(n2860), .B(n2861), .ZN(n3187) );
  NOR2_X1 U33460 ( .A1(n3186), .A2(n3187), .ZN(n3185) );
  AOI21_X1 U33470 ( .B1(n2861), .B2(n2860), .A(n3185), .ZN(n3220) );
  INV_X1 U33480 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2862) );
  INV_X1 U33490 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2863) );
  OR2_X1 U33500 ( .A1(n2864), .A2(n2863), .ZN(n2867) );
  INV_X1 U33510 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4741) );
  OR2_X1 U33520 ( .A1(n2840), .A2(n4741), .ZN(n2865) );
  NAND2_X1 U3353 ( .A1(n2869), .A2(IR_REG_31__SCAN_IN), .ZN(n2881) );
  XNOR2_X1 U33540 ( .A(n2881), .B(IR_REG_3__SCAN_IN), .ZN(n4028) );
  MUX2_X1 U3355 ( .A(DATAI_3_), .B(n4028), .S(n3603), .Z(n3285) );
  OAI21_X1 U3356 ( .B1(n3266), .B2(n3650), .A(n2870), .ZN(n2871) );
  XNOR2_X1 U3357 ( .A(n2871), .B(n2958), .ZN(n2874) );
  AOI22_X1 U3358 ( .A1(n2855), .A2(n5034), .B1(n3665), .B2(n3285), .ZN(n2872)
         );
  XOR2_X1 U3359 ( .A(n2874), .B(n2872), .Z(n3221) );
  INV_X1 U3360 ( .A(n2872), .ZN(n2873) );
  OAI22_X1 U3361 ( .A1(n3220), .A2(n3221), .B1(n2874), .B2(n2873), .ZN(n3264)
         );
  NAND2_X1 U3362 ( .A1(n3565), .A2(REG2_REG_4__SCAN_IN), .ZN(n2879) );
  INV_X1 U3363 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2875) );
  OR2_X1 U3364 ( .A1(n3195), .A2(n2875), .ZN(n2878) );
  XNOR2_X1 U3365 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3297) );
  OR2_X1 U3366 ( .A1(n2842), .A2(n3297), .ZN(n2877) );
  INV_X1 U3367 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4742) );
  OR2_X1 U3368 ( .A1(n3822), .A2(n4742), .ZN(n2876) );
  NAND2_X1 U3369 ( .A1(n2881), .A2(n2880), .ZN(n2882) );
  NAND2_X1 U3370 ( .A1(n2882), .A2(IR_REG_31__SCAN_IN), .ZN(n2883) );
  XNOR2_X1 U3371 ( .A(n2883), .B(IR_REG_4__SCAN_IN), .ZN(n4989) );
  MUX2_X1 U3372 ( .A(DATAI_4_), .B(n4989), .S(n3828), .Z(n3309) );
  AOI22_X1 U3373 ( .A1(n3665), .A2(n3991), .B1(n3063), .B2(n3309), .ZN(n2884)
         );
  AOI22_X1 U3374 ( .A1(n2855), .A2(n3991), .B1(n3665), .B2(n3309), .ZN(n2886)
         );
  XNOR2_X1 U3375 ( .A(n2885), .B(n2886), .ZN(n3265) );
  NOR2_X1 U3376 ( .A1(n3264), .A2(n3265), .ZN(n3263) );
  INV_X1 U3377 ( .A(n2885), .ZN(n2888) );
  INV_X1 U3378 ( .A(n2886), .ZN(n2887) );
  XNOR2_X1 U3379 ( .A(n2889), .B(n2890), .ZN(n3274) );
  NAND2_X1 U3380 ( .A1(n2843), .A2(REG1_REG_6__SCAN_IN), .ZN(n2897) );
  INV_X1 U3381 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5072) );
  OR2_X1 U3382 ( .A1(n3822), .A2(n5072), .ZN(n2896) );
  NOR2_X1 U3383 ( .A1(n2892), .A2(REG3_REG_6__SCAN_IN), .ZN(n2893) );
  OR2_X1 U3384 ( .A1(n2906), .A2(n2893), .ZN(n3369) );
  OR2_X1 U3385 ( .A1(n2842), .A2(n3369), .ZN(n2895) );
  INV_X1 U3386 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3370) );
  OR2_X1 U3387 ( .A1(n3826), .A2(n3370), .ZN(n2894) );
  NAND4_X1 U3388 ( .A1(n2897), .A2(n2896), .A3(n2895), .A4(n2894), .ZN(n3989)
         );
  NAND2_X1 U3389 ( .A1(n2898), .A2(IR_REG_31__SCAN_IN), .ZN(n2899) );
  XNOR2_X1 U3390 ( .A(n2899), .B(IR_REG_6__SCAN_IN), .ZN(n4851) );
  MUX2_X1 U3391 ( .A(DATAI_6_), .B(n4851), .S(n3828), .Z(n3374) );
  AOI22_X1 U3392 ( .A1(n2855), .A2(n3989), .B1(n3665), .B2(n3374), .ZN(n2904)
         );
  INV_X1 U3393 ( .A(n3989), .ZN(n2901) );
  OR2_X1 U3394 ( .A1(n2825), .A2(n3367), .ZN(n2900) );
  OAI21_X1 U3395 ( .B1(n3650), .B2(n2901), .A(n2900), .ZN(n2902) );
  XNOR2_X1 U3396 ( .A(n2902), .B(n2958), .ZN(n2903) );
  XNOR2_X1 U3397 ( .A(n2904), .B(n2903), .ZN(n3330) );
  INV_X1 U3398 ( .A(n2903), .ZN(n2905) );
  NAND2_X1 U3399 ( .A1(n3565), .A2(REG2_REG_7__SCAN_IN), .ZN(n2912) );
  OR2_X1 U3400 ( .A1(n3195), .A2(n5077), .ZN(n2911) );
  OR2_X1 U3401 ( .A1(n2906), .A2(REG3_REG_7__SCAN_IN), .ZN(n2907) );
  NAND2_X1 U3402 ( .A1(n2908), .A2(n2907), .ZN(n3677) );
  OR2_X1 U3403 ( .A1(n2842), .A2(n3677), .ZN(n2910) );
  INV_X1 U3404 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5078) );
  OR2_X1 U3405 ( .A1(n3822), .A2(n5078), .ZN(n2909) );
  NAND4_X1 U3406 ( .A1(n2912), .A2(n2911), .A3(n2910), .A4(n2909), .ZN(n3988)
         );
  XNOR2_X1 U3407 ( .A(n2913), .B(IR_REG_7__SCAN_IN), .ZN(n4776) );
  MUX2_X1 U3408 ( .A(DATAI_7_), .B(n4776), .S(n3828), .Z(n3681) );
  AOI22_X1 U3409 ( .A1(n2855), .A2(n3988), .B1(n3665), .B2(n3681), .ZN(n2915)
         );
  AOI22_X1 U3410 ( .A1(n3665), .A2(n3988), .B1(n3063), .B2(n3681), .ZN(n2914)
         );
  XNOR2_X1 U3411 ( .A(n2914), .B(n2958), .ZN(n2916) );
  XOR2_X1 U3412 ( .A(n2915), .B(n2916), .Z(n3675) );
  OR2_X1 U3413 ( .A1(n2916), .A2(n2915), .ZN(n2917) );
  XOR2_X1 U3414 ( .A(n2918), .B(n2920), .Z(n3394) );
  NAND2_X1 U3415 ( .A1(n3030), .A2(REG0_REG_9__SCAN_IN), .ZN(n2926) );
  INV_X1 U3416 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3388) );
  OR2_X1 U3417 ( .A1(n3826), .A2(n3388), .ZN(n2925) );
  INV_X1 U3418 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3996) );
  OR2_X1 U3419 ( .A1(n3195), .A2(n3996), .ZN(n2924) );
  NAND2_X1 U3420 ( .A1(n2921), .A2(n4435), .ZN(n2922) );
  NAND2_X1 U3421 ( .A1(n2937), .A2(n2922), .ZN(n3404) );
  OR2_X1 U3422 ( .A1(n2842), .A2(n3404), .ZN(n2923) );
  NAND4_X1 U3423 ( .A1(n2926), .A2(n2925), .A3(n2924), .A4(n2923), .ZN(n3986)
         );
  INV_X1 U3424 ( .A(n3986), .ZN(n5100) );
  INV_X1 U3425 ( .A(n2927), .ZN(n2928) );
  OAI21_X1 U3426 ( .B1(n2929), .B2(n2928), .A(IR_REG_31__SCAN_IN), .ZN(n2930)
         );
  XNOR2_X1 U3427 ( .A(n2930), .B(IR_REG_9__SCAN_IN), .ZN(n4025) );
  MUX2_X1 U3428 ( .A(DATAI_9_), .B(n4025), .S(n3828), .Z(n3413) );
  OR2_X1 U3429 ( .A1(n2825), .A2(n3406), .ZN(n2931) );
  OAI21_X1 U3430 ( .B1(n3650), .B2(n5100), .A(n2931), .ZN(n2932) );
  XNOR2_X1 U3431 ( .A(n2932), .B(n2958), .ZN(n2935) );
  AOI22_X1 U3432 ( .A1(n2855), .A2(n3986), .B1(n3665), .B2(n3413), .ZN(n2933)
         );
  XOR2_X1 U3433 ( .A(n2935), .B(n2933), .Z(n3403) );
  INV_X1 U3434 ( .A(n2933), .ZN(n2934) );
  NAND2_X1 U3435 ( .A1(n3565), .A2(REG2_REG_10__SCAN_IN), .ZN(n2944) );
  INV_X1 U3436 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2936) );
  OR2_X1 U3437 ( .A1(n3195), .A2(n2936), .ZN(n2943) );
  NOR2_X2 U3438 ( .A1(n2937), .A2(n4602), .ZN(n2951) );
  INV_X1 U3439 ( .A(n2951), .ZN(n2939) );
  NAND2_X1 U3440 ( .A1(n2937), .A2(n4602), .ZN(n2938) );
  NAND2_X1 U3441 ( .A1(n2939), .A2(n2938), .ZN(n5111) );
  OR2_X1 U3442 ( .A1(n2842), .A2(n5111), .ZN(n2942) );
  INV_X1 U3443 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2940) );
  OR2_X1 U3444 ( .A1(n3822), .A2(n2940), .ZN(n2941) );
  OR2_X1 U3445 ( .A1(n2945), .A2(n2761), .ZN(n2946) );
  XNOR2_X1 U3446 ( .A(n2946), .B(IR_REG_10__SCAN_IN), .ZN(n4891) );
  AOI22_X1 U3447 ( .A1(n3665), .A2(n5119), .B1(n3063), .B2(n5102), .ZN(n2947)
         );
  XNOR2_X1 U3448 ( .A(n2947), .B(n2958), .ZN(n2949) );
  AOI22_X1 U3449 ( .A1(n2855), .A2(n5119), .B1(n3665), .B2(n5102), .ZN(n2948)
         );
  XNOR2_X1 U3450 ( .A(n2949), .B(n2948), .ZN(n3449) );
  NOR2_X1 U3451 ( .A1(n2949), .A2(n2948), .ZN(n2950) );
  NAND2_X1 U3452 ( .A1(n3030), .A2(REG0_REG_11__SCAN_IN), .ZN(n2956) );
  OR2_X1 U3453 ( .A1(n3826), .A2(n5139), .ZN(n2955) );
  INV_X1 U3454 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3994) );
  OR2_X1 U3455 ( .A1(n3195), .A2(n3994), .ZN(n2954) );
  NOR2_X1 U3456 ( .A1(n2951), .A2(REG3_REG_11__SCAN_IN), .ZN(n2952) );
  OR2_X1 U3457 ( .A1(n2960), .A2(n2952), .ZN(n3457) );
  OR2_X1 U34580 ( .A1(n2842), .A2(n3457), .ZN(n2953) );
  NAND4_X1 U34590 ( .A1(n2956), .A2(n2955), .A3(n2954), .A4(n2953), .ZN(n3985)
         );
  NAND2_X1 U3460 ( .A1(n2957), .A2(IR_REG_31__SCAN_IN), .ZN(n2967) );
  XNOR2_X1 U3461 ( .A(n2967), .B(IR_REG_11__SCAN_IN), .ZN(n4775) );
  MUX2_X1 U3462 ( .A(DATAI_11_), .B(n4775), .S(n3828), .Z(n5115) );
  AOI22_X1 U3463 ( .A1(n3665), .A2(n3985), .B1(n3063), .B2(n5115), .ZN(n2959)
         );
  INV_X1 U3464 ( .A(n3985), .ZN(n5099) );
  INV_X1 U3465 ( .A(n5115), .ZN(n5122) );
  OAI22_X1 U3466 ( .A1(n3651), .A2(n5099), .B1(n3650), .B2(n5122), .ZN(n3454)
         );
  NAND2_X1 U34670 ( .A1(n3030), .A2(REG0_REG_12__SCAN_IN), .ZN(n2965) );
  INV_X1 U3468 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3427) );
  OR2_X1 U34690 ( .A1(n3826), .A2(n3427), .ZN(n2964) );
  OR2_X1 U3470 ( .A1(n3195), .A2(n5149), .ZN(n2963) );
  NOR2_X1 U34710 ( .A1(n2960), .A2(REG3_REG_12__SCAN_IN), .ZN(n2961) );
  OR2_X1 U3472 ( .A1(n2974), .A2(n2961), .ZN(n3464) );
  OR2_X1 U34730 ( .A1(n2842), .A2(n3464), .ZN(n2962) );
  NAND4_X1 U3474 ( .A1(n2965), .A2(n2964), .A3(n2963), .A4(n2962), .ZN(n5118)
         );
  INV_X1 U34750 ( .A(IR_REG_11__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3476 ( .A1(n2967), .A2(n2966), .ZN(n2968) );
  NAND2_X1 U34770 ( .A1(n2968), .A2(IR_REG_31__SCAN_IN), .ZN(n2969) );
  XNOR2_X1 U3478 ( .A(n2969), .B(IR_REG_12__SCAN_IN), .ZN(n4044) );
  MUX2_X1 U34790 ( .A(DATAI_12_), .B(n4044), .S(n3828), .Z(n3433) );
  AOI22_X1 U3480 ( .A1(n3665), .A2(n5118), .B1(n3063), .B2(n3433), .ZN(n2970)
         );
  XOR2_X1 U34810 ( .A(n2958), .B(n2970), .Z(n2972) );
  INV_X1 U3482 ( .A(n5118), .ZN(n3458) );
  OAI22_X1 U34830 ( .A1(n3651), .A2(n3458), .B1(n3650), .B2(n3467), .ZN(n2971)
         );
  NOR2_X1 U3484 ( .A1(n2972), .A2(n2971), .ZN(n3768) );
  AOI21_X1 U34850 ( .B1(n2972), .B2(n2971), .A(n3768), .ZN(n3463) );
  INV_X1 U3486 ( .A(n3768), .ZN(n2973) );
  NAND2_X1 U34870 ( .A1(n3565), .A2(REG2_REG_13__SCAN_IN), .ZN(n2979) );
  INV_X1 U3488 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4014) );
  OR2_X1 U34890 ( .A1(n3195), .A2(n4014), .ZN(n2978) );
  OAI21_X1 U3490 ( .B1(n2974), .B2(REG3_REG_13__SCAN_IN), .A(n2991), .ZN(n3773) );
  OR2_X1 U34910 ( .A1(n2842), .A2(n3773), .ZN(n2977) );
  INV_X1 U3492 ( .A(REG0_REG_13__SCAN_IN), .ZN(n2975) );
  OR2_X1 U34930 ( .A1(n3822), .A2(n2975), .ZN(n2976) );
  INV_X1 U3494 ( .A(DATAI_13_), .ZN(n4380) );
  INV_X1 U34950 ( .A(n2980), .ZN(n2981) );
  NAND2_X1 U3496 ( .A1(n2981), .A2(IR_REG_31__SCAN_IN), .ZN(n2983) );
  XNOR2_X1 U34970 ( .A(n2983), .B(n2982), .ZN(n4930) );
  MUX2_X1 U3498 ( .A(n4380), .B(n4930), .S(n3828), .Z(n3435) );
  OR2_X1 U34990 ( .A1(n2825), .A2(n3435), .ZN(n2984) );
  OAI21_X1 U3500 ( .B1(n3650), .B2(n3480), .A(n2984), .ZN(n2985) );
  XNOR2_X1 U35010 ( .A(n2985), .B(n2958), .ZN(n2987) );
  OAI22_X1 U3502 ( .A1(n3651), .A2(n3480), .B1(n3650), .B2(n3435), .ZN(n2986)
         );
  OR2_X1 U35030 ( .A1(n2987), .A2(n2986), .ZN(n2989) );
  NAND2_X1 U3504 ( .A1(n2987), .A2(n2986), .ZN(n2988) );
  AND2_X1 U35050 ( .A1(n2989), .A2(n2988), .ZN(n3767) );
  NAND2_X1 U35060 ( .A1(n3030), .A2(REG0_REG_14__SCAN_IN), .ZN(n2995) );
  INV_X1 U35070 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4299) );
  OR2_X1 U35080 ( .A1(n3826), .A2(n4299), .ZN(n2994) );
  INV_X1 U35090 ( .A(REG1_REG_14__SCAN_IN), .ZN(n2990) );
  OR2_X1 U35100 ( .A1(n3195), .A2(n2990), .ZN(n2993) );
  AOI21_X1 U35110 ( .B1(n2991), .B2(n3697), .A(n3007), .ZN(n3696) );
  INV_X1 U35120 ( .A(n3696), .ZN(n4298) );
  OR2_X1 U35130 ( .A1(n2842), .A2(n4298), .ZN(n2992) );
  NAND4_X1 U35140 ( .A1(n2995), .A2(n2994), .A3(n2993), .A4(n2992), .ZN(n5158)
         );
  NAND2_X1 U35150 ( .A1(n2740), .A2(IR_REG_31__SCAN_IN), .ZN(n2997) );
  XNOR2_X1 U35160 ( .A(n2997), .B(IR_REG_14__SCAN_IN), .ZN(n4937) );
  MUX2_X1 U35170 ( .A(DATAI_14_), .B(n4937), .S(n3603), .Z(n3473) );
  AOI22_X1 U35180 ( .A1(n2855), .A2(n5158), .B1(n3665), .B2(n3473), .ZN(n3002)
         );
  OR2_X1 U35190 ( .A1(n2825), .A2(n4290), .ZN(n2998) );
  OAI21_X1 U35200 ( .B1(n3650), .B2(n3775), .A(n2998), .ZN(n2999) );
  XNOR2_X1 U35210 ( .A(n2999), .B(n2958), .ZN(n3000) );
  XNOR2_X1 U35220 ( .A(n3002), .B(n3000), .ZN(n3695) );
  INV_X1 U35230 ( .A(n3000), .ZN(n3001) );
  NAND2_X1 U35240 ( .A1(n3002), .A2(n3001), .ZN(n3003) );
  NAND2_X1 U35250 ( .A1(n3030), .A2(REG0_REG_15__SCAN_IN), .ZN(n3006) );
  NAND2_X1 U35260 ( .A1(n3565), .A2(REG2_REG_15__SCAN_IN), .ZN(n3005) );
  NAND2_X1 U35270 ( .A1(n2843), .A2(REG1_REG_15__SCAN_IN), .ZN(n3004) );
  NAND3_X1 U35280 ( .A1(n3006), .A2(n3005), .A3(n3004), .ZN(n3009) );
  OAI21_X1 U35290 ( .B1(n3007), .B2(REG3_REG_15__SCAN_IN), .A(n3012), .ZN(
        n5176) );
  NOR2_X1 U35300 ( .A1(n5176), .A2(n2842), .ZN(n3008) );
  XNOR2_X1 U35310 ( .A(n3010), .B(IR_REG_15__SCAN_IN), .ZN(n4773) );
  MUX2_X1 U35320 ( .A(DATAI_15_), .B(n4773), .S(n3828), .Z(n5162) );
  AOI22_X1 U35330 ( .A1(n3665), .A2(n4287), .B1(n3063), .B2(n5162), .ZN(n3011)
         );
  OAI22_X1 U35340 ( .A1(n3651), .A2(n4267), .B1(n3650), .B2(n3511), .ZN(n5170)
         );
  AOI21_X1 U35350 ( .B1(n3012), .B2(n4427), .A(n3028), .ZN(n4276) );
  INV_X1 U35360 ( .A(n2842), .ZN(n3013) );
  NAND2_X1 U35370 ( .A1(n4276), .A2(n3013), .ZN(n3017) );
  NAND2_X1 U35380 ( .A1(n3565), .A2(REG2_REG_16__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U35390 ( .A1(n2843), .A2(REG1_REG_16__SCAN_IN), .ZN(n3015) );
  NAND2_X1 U35400 ( .A1(n3030), .A2(REG0_REG_16__SCAN_IN), .ZN(n3014) );
  NAND4_X1 U35410 ( .A1(n3017), .A2(n3016), .A3(n3015), .A4(n3014), .ZN(n5160)
         );
  NAND2_X1 U35420 ( .A1(n3018), .A2(IR_REG_31__SCAN_IN), .ZN(n3019) );
  XNOR2_X1 U35430 ( .A(n3019), .B(IR_REG_16__SCAN_IN), .ZN(n4772) );
  MUX2_X1 U35440 ( .A(DATAI_16_), .B(n4772), .S(n3603), .Z(n4272) );
  AOI22_X1 U35450 ( .A1(n3665), .A2(n5160), .B1(n3063), .B2(n4272), .ZN(n3020)
         );
  XNOR2_X1 U35460 ( .A(n3020), .B(n2958), .ZN(n3022) );
  AOI22_X1 U35470 ( .A1(n2855), .A2(n5160), .B1(n3665), .B2(n4272), .ZN(n3021)
         );
  NAND2_X1 U35480 ( .A1(n3022), .A2(n3021), .ZN(n3026) );
  OAI21_X1 U35490 ( .B1(n3022), .B2(n3021), .A(n3026), .ZN(n3733) );
  INV_X1 U35500 ( .A(n3733), .ZN(n3025) );
  INV_X1 U35510 ( .A(n3023), .ZN(n3024) );
  NAND2_X1 U35520 ( .A1(n3024), .A2(n2516), .ZN(n3729) );
  NAND3_X1 U35530 ( .A1(n3730), .A2(n3025), .A3(n3729), .ZN(n3027) );
  NAND2_X1 U35540 ( .A1(n3027), .A2(n3026), .ZN(n3738) );
  OR2_X1 U35550 ( .A1(n3028), .A2(REG3_REG_17__SCAN_IN), .ZN(n3029) );
  NAND2_X1 U35560 ( .A1(n3028), .A2(REG3_REG_17__SCAN_IN), .ZN(n3041) );
  NAND2_X1 U35570 ( .A1(n3029), .A2(n3041), .ZN(n4257) );
  INV_X1 U35580 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U35590 ( .A1(n3565), .A2(REG2_REG_17__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U35600 ( .A1(n3030), .A2(REG0_REG_17__SCAN_IN), .ZN(n3031) );
  OAI211_X1 U35610 ( .C1(n3195), .C2(n4061), .A(n3032), .B(n3031), .ZN(n3033)
         );
  INV_X1 U35620 ( .A(n3033), .ZN(n3034) );
  XNOR2_X1 U35630 ( .A(n3035), .B(IR_REG_17__SCAN_IN), .ZN(n4771) );
  MUX2_X1 U35640 ( .A(DATAI_17_), .B(n4771), .S(n3828), .Z(n4253) );
  AOI22_X1 U35650 ( .A1(n3665), .A2(n4231), .B1(n3063), .B2(n4253), .ZN(n3036)
         );
  XNOR2_X1 U35660 ( .A(n3036), .B(n2958), .ZN(n3037) );
  INV_X1 U35670 ( .A(n4231), .ZN(n4268) );
  OAI22_X1 U35680 ( .A1(n3651), .A2(n4268), .B1(n3650), .B2(n3742), .ZN(n3038)
         );
  XNOR2_X1 U35690 ( .A(n3037), .B(n3038), .ZN(n3740) );
  INV_X1 U35700 ( .A(n3037), .ZN(n3039) );
  OR2_X1 U35710 ( .A1(n3039), .A2(n3038), .ZN(n3040) );
  NAND2_X1 U35720 ( .A1(n2843), .A2(REG1_REG_18__SCAN_IN), .ZN(n3047) );
  INV_X1 U35730 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4088) );
  OR2_X1 U35740 ( .A1(n3826), .A2(n4088), .ZN(n3046) );
  INV_X1 U35750 ( .A(n3055), .ZN(n3056) );
  OAI21_X1 U35760 ( .B1(REG3_REG_18__SCAN_IN), .B2(n3042), .A(n3056), .ZN(
        n4241) );
  OR2_X1 U35770 ( .A1(n2842), .A2(n4241), .ZN(n3045) );
  INV_X1 U35780 ( .A(REG0_REG_18__SCAN_IN), .ZN(n3043) );
  OR2_X1 U35790 ( .A1(n3822), .A2(n3043), .ZN(n3044) );
  NAND4_X1 U35800 ( .A1(n3047), .A2(n3046), .A3(n3045), .A4(n3044), .ZN(n3983)
         );
  INV_X1 U35810 ( .A(IR_REG_18__SCAN_IN), .ZN(n4665) );
  XNOR2_X1 U3582 ( .A(n3048), .B(n4665), .ZN(n4770) );
  MUX2_X1 U3583 ( .A(DATAI_18_), .B(n4770), .S(n3603), .Z(n4240) );
  AOI22_X1 U3584 ( .A1(n3665), .A2(n3983), .B1(n3063), .B2(n4240), .ZN(n3049)
         );
  XOR2_X1 U3585 ( .A(n2958), .B(n3049), .Z(n3050) );
  INV_X1 U3586 ( .A(n3983), .ZN(n5213) );
  OAI22_X1 U3587 ( .A1(n3651), .A2(n5213), .B1(n4233), .B2(n3650), .ZN(n3051)
         );
  NAND2_X1 U3588 ( .A1(n3050), .A2(n3051), .ZN(n3793) );
  INV_X1 U3589 ( .A(n3050), .ZN(n3053) );
  INV_X1 U3590 ( .A(n3051), .ZN(n3052) );
  NAND2_X1 U3591 ( .A1(n3053), .A2(n3052), .ZN(n3792) );
  NAND2_X1 U3592 ( .A1(n3565), .A2(REG2_REG_19__SCAN_IN), .ZN(n3062) );
  INV_X1 U3593 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3054) );
  OR2_X1 U3594 ( .A1(n3195), .A2(n3054), .ZN(n3061) );
  INV_X1 U3595 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U3596 ( .A1(n3056), .A2(n4608), .ZN(n3057) );
  NAND2_X1 U3597 ( .A1(n3070), .A2(n3057), .ZN(n5223) );
  OR2_X1 U3598 ( .A1(n2842), .A2(n5223), .ZN(n3060) );
  INV_X1 U3599 ( .A(REG0_REG_19__SCAN_IN), .ZN(n3058) );
  OR2_X1 U3600 ( .A1(n3822), .A2(n3058), .ZN(n3059) );
  NAND4_X1 U3601 ( .A1(n3062), .A2(n3061), .A3(n3060), .A4(n3059), .ZN(n4230)
         );
  INV_X1 U3602 ( .A(n5219), .ZN(n3112) );
  MUX2_X1 U3603 ( .A(n3112), .B(DATAI_19_), .S(n2800), .Z(n5215) );
  AOI22_X1 U3604 ( .A1(n3665), .A2(n4230), .B1(n3063), .B2(n5215), .ZN(n3064)
         );
  XNOR2_X1 U3605 ( .A(n3064), .B(n2958), .ZN(n3065) );
  INV_X1 U3606 ( .A(n5215), .ZN(n3499) );
  OAI22_X1 U3607 ( .A1(n3651), .A2(n3762), .B1(n3650), .B2(n3499), .ZN(n3066)
         );
  XNOR2_X1 U3608 ( .A(n3065), .B(n3066), .ZN(n3713) );
  INV_X1 U3609 ( .A(n3065), .ZN(n3067) );
  NAND2_X1 U3610 ( .A1(n2843), .A2(REG1_REG_20__SCAN_IN), .ZN(n3076) );
  INV_X1 U3611 ( .A(REG0_REG_20__SCAN_IN), .ZN(n3068) );
  OR2_X1 U3612 ( .A1(n3822), .A2(n3068), .ZN(n3075) );
  INV_X1 U3613 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U3614 ( .A1(n3070), .A2(n4634), .ZN(n3071) );
  NAND2_X1 U3615 ( .A1(n3082), .A2(n3071), .ZN(n4222) );
  OR2_X1 U3616 ( .A1(n2842), .A2(n4222), .ZN(n3074) );
  INV_X1 U3617 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3072) );
  OR2_X1 U3618 ( .A1(n3826), .A2(n3072), .ZN(n3073) );
  NAND2_X1 U3619 ( .A1(n2800), .A2(DATAI_20_), .ZN(n3519) );
  OAI22_X1 U3620 ( .A1(n5211), .A2(n3650), .B1(n2825), .B2(n3519), .ZN(n3077)
         );
  XNOR2_X1 U3621 ( .A(n3077), .B(n2958), .ZN(n3079) );
  OAI22_X1 U3622 ( .A1(n3651), .A2(n5211), .B1(n3650), .B2(n3519), .ZN(n3078)
         );
  NAND2_X1 U3623 ( .A1(n3079), .A2(n3078), .ZN(n3759) );
  NOR2_X1 U3624 ( .A1(n3079), .A2(n3078), .ZN(n3758) );
  AOI21_X1 U3625 ( .B1(n3757), .B2(n3759), .A(n3758), .ZN(n3117) );
  NAND2_X1 U3626 ( .A1(n3565), .A2(REG2_REG_21__SCAN_IN), .ZN(n3088) );
  INV_X1 U3627 ( .A(REG1_REG_21__SCAN_IN), .ZN(n3080) );
  OR2_X1 U3628 ( .A1(n3195), .A2(n3080), .ZN(n3087) );
  INV_X1 U3629 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U3630 ( .A1(n3082), .A2(n4418), .ZN(n3083) );
  NAND2_X1 U3631 ( .A1(n3129), .A2(n3083), .ZN(n4201) );
  OR2_X1 U3632 ( .A1(n2842), .A2(n4201), .ZN(n3086) );
  INV_X1 U3633 ( .A(REG0_REG_21__SCAN_IN), .ZN(n3084) );
  OR2_X1 U3634 ( .A1(n3822), .A2(n3084), .ZN(n3085) );
  NAND2_X1 U3635 ( .A1(n2800), .A2(DATAI_21_), .ZN(n3538) );
  OR2_X1 U3636 ( .A1(n2825), .A2(n3538), .ZN(n3089) );
  OAI21_X1 U3637 ( .B1(n3650), .B2(n4178), .A(n3089), .ZN(n3090) );
  XNOR2_X1 U3638 ( .A(n3090), .B(n2958), .ZN(n3092) );
  OAI22_X1 U3639 ( .A1(n3651), .A2(n4178), .B1(n3650), .B2(n3538), .ZN(n3091)
         );
  OR2_X1 U3640 ( .A1(n3092), .A2(n3091), .ZN(n3118) );
  NAND2_X1 U3641 ( .A1(n3117), .A2(n3118), .ZN(n3782) );
  INV_X1 U3642 ( .A(n3782), .ZN(n3120) );
  AND2_X1 U3643 ( .A1(n3092), .A2(n3091), .ZN(n3628) );
  INV_X1 U3644 ( .A(n3628), .ZN(n3781) );
  NAND2_X1 U3645 ( .A1(n3140), .A2(B_REG_SCAN_IN), .ZN(n3094) );
  MUX2_X1 U3646 ( .A(n3094), .B(B_REG_SCAN_IN), .S(n3093), .Z(n3095) );
  NOR2_X1 U3647 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_18__SCAN_IN), .ZN(n3099) );
  NOR4_X1 U3648 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n3098) );
  NOR4_X1 U3649 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n3097) );
  NOR4_X1 U3650 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n3096) );
  NAND4_X1 U3651 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3105)
         );
  NOR4_X1 U3652 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n3103) );
  NOR4_X1 U3653 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n3102) );
  NOR4_X1 U3654 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n3101) );
  NOR4_X1 U3655 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n3100) );
  NAND4_X1 U3656 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3104)
         );
  NOR2_X1 U3657 ( .A1(n3105), .A2(n3104), .ZN(n3106) );
  NOR2_X1 U3658 ( .A1(n3150), .A2(n3106), .ZN(n4307) );
  OR2_X1 U3659 ( .A1(n3150), .A2(D_REG_1__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3660 ( .A1(n3108), .A2(n3140), .ZN(n3151) );
  NAND2_X1 U3661 ( .A1(n3107), .A2(n3151), .ZN(n4308) );
  OR2_X1 U3662 ( .A1(n4307), .A2(n4308), .ZN(n3226) );
  INV_X1 U3663 ( .A(n3093), .ZN(n3109) );
  NAND2_X1 U3664 ( .A1(n3109), .A2(n3108), .ZN(n3153) );
  NOR2_X1 U3665 ( .A1(n3226), .A2(n4342), .ZN(n3126) );
  INV_X1 U3666 ( .A(n4311), .ZN(n3115) );
  INV_X1 U3667 ( .A(n3113), .ZN(n3970) );
  NOR2_X1 U3668 ( .A1(n3233), .A2(n3886), .ZN(n3247) );
  INV_X1 U3669 ( .A(n3247), .ZN(n3114) );
  AND3_X1 U3670 ( .A1(n3115), .A2(n5123), .A3(n3114), .ZN(n3116) );
  AOI21_X1 U3671 ( .B1(n3118), .B2(n3781), .A(n3117), .ZN(n3119) );
  AOI211_X1 U3672 ( .C1(n3120), .C2(n3781), .A(n3815), .B(n3119), .ZN(n3139)
         );
  NAND2_X1 U3673 ( .A1(n3167), .A2(n5240), .ZN(n3121) );
  NOR2_X1 U3674 ( .A1(n3743), .A2(n3538), .ZN(n3138) );
  NAND2_X1 U3675 ( .A1(n3113), .A2(n5219), .ZN(n3122) );
  NAND2_X1 U3676 ( .A1(n3122), .A2(n3247), .ZN(n3166) );
  AND2_X1 U3677 ( .A1(n3166), .A2(n2790), .ZN(n3228) );
  OAI211_X1 U3678 ( .C1(n3126), .C2(n4311), .A(n3228), .B(n3158), .ZN(n3123)
         );
  OR2_X1 U3679 ( .A1(n2802), .A2(n3124), .ZN(n3242) );
  INV_X1 U3680 ( .A(n3157), .ZN(n3125) );
  NOR2_X1 U3681 ( .A1(n3242), .A2(n3125), .ZN(n3975) );
  NAND2_X1 U3682 ( .A1(n3126), .A2(n3975), .ZN(n3135) );
  INV_X1 U3683 ( .A(n3127), .ZN(n4807) );
  NAND2_X1 U3684 ( .A1(n3565), .A2(REG2_REG_22__SCAN_IN), .ZN(n3134) );
  INV_X1 U3685 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4332) );
  OR2_X1 U3686 ( .A1(n3195), .A2(n4332), .ZN(n3133) );
  INV_X1 U3687 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U3688 ( .A1(n3129), .A2(n3786), .ZN(n3130) );
  NAND2_X1 U3689 ( .A1(n3177), .A2(n3130), .ZN(n4192) );
  OR2_X1 U3690 ( .A1(n2842), .A2(n4192), .ZN(n3132) );
  INV_X1 U3691 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4353) );
  OR2_X1 U3692 ( .A1(n3822), .A2(n4353), .ZN(n3131) );
  OAI22_X1 U3693 ( .A1(n5177), .A2(n4201), .B1(n3809), .B2(n4205), .ZN(n3137)
         );
  OAI22_X1 U3694 ( .A1(n3810), .A2(n5211), .B1(STATE_REG_SCAN_IN), .B2(n4418), 
        .ZN(n3136) );
  OR4_X1 U3695 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(U3220) );
  INV_X2 U3696 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3697 ( .A(DATAI_25_), .ZN(n3141) );
  MUX2_X1 U3698 ( .A(n3141), .B(n3140), .S(STATE_REG_SCAN_IN), .Z(n3142) );
  INV_X1 U3699 ( .A(n3142), .ZN(U3327) );
  INV_X1 U3700 ( .A(DATAI_27_), .ZN(n3144) );
  MUX2_X1 U3701 ( .A(n3143), .B(n3144), .S(U3149), .Z(n3145) );
  INV_X1 U3702 ( .A(n3145), .ZN(U3325) );
  INV_X1 U3703 ( .A(DATAI_19_), .ZN(n3146) );
  MUX2_X1 U3704 ( .A(n5219), .B(n3146), .S(U3149), .Z(n3147) );
  INV_X1 U3705 ( .A(n3147), .ZN(U3333) );
  INV_X1 U3706 ( .A(DATAI_28_), .ZN(n3148) );
  MUX2_X1 U3707 ( .A(n3148), .B(n3127), .S(STATE_REG_SCAN_IN), .Z(n3149) );
  INV_X1 U3708 ( .A(n3149), .ZN(U3324) );
  NAND2_X1 U3709 ( .A1(n3150), .A2(n3157), .ZN(n4802) );
  INV_X1 U3710 ( .A(D_REG_1__SCAN_IN), .ZN(n4691) );
  INV_X1 U3711 ( .A(n3151), .ZN(n3152) );
  AOI22_X1 U3712 ( .A1(n4802), .A2(n4691), .B1(n4777), .B2(n3152), .ZN(U3459)
         );
  INV_X1 U3713 ( .A(D_REG_0__SCAN_IN), .ZN(n3155) );
  INV_X1 U3714 ( .A(n3153), .ZN(n3154) );
  AOI22_X1 U3715 ( .A1(n4802), .A2(n3155), .B1(n4777), .B2(n3154), .ZN(U3458)
         );
  OR2_X1 U3716 ( .A1(n3158), .A2(U3149), .ZN(n3978) );
  INV_X1 U3717 ( .A(n3978), .ZN(n3156) );
  AND2_X1 U3718 ( .A1(n3247), .A2(n3158), .ZN(n3159) );
  NOR2_X1 U3719 ( .A1(n3159), .A2(n3828), .ZN(n4021) );
  INV_X1 U3720 ( .A(n4021), .ZN(n3160) );
  NOR2_X1 U3721 ( .A1(n4988), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3722 ( .A1(n3984), .A2(DATAO_REG_20__SCAN_IN), .ZN(n3161) );
  OAI21_X1 U3723 ( .B1(n5211), .B2(n3984), .A(n3161), .ZN(U3570) );
  NAND2_X1 U3724 ( .A1(n3984), .A2(DATAO_REG_22__SCAN_IN), .ZN(n3162) );
  OAI21_X1 U3725 ( .B1(n4205), .B2(n3984), .A(n3162), .ZN(U3572) );
  OAI21_X1 U3726 ( .B1(n3165), .B2(n3164), .A(n3163), .ZN(n4974) );
  OAI21_X1 U3727 ( .B1(n3167), .B2(n5135), .A(n3166), .ZN(n3191) );
  AOI22_X1 U3728 ( .A1(n3191), .A2(REG3_REG_0__SCAN_IN), .B1(n5161), .B2(n3237), .ZN(n3169) );
  NAND2_X1 U3729 ( .A1(n5163), .A2(n5004), .ZN(n3168) );
  OAI211_X1 U3730 ( .C1(n4974), .C2(n3815), .A(n3169), .B(n3168), .ZN(U3229)
         );
  OAI211_X1 U3731 ( .C1(n3170), .C2(n3172), .A(n3171), .B(n5172), .ZN(n3175)
         );
  INV_X1 U3732 ( .A(n5010), .ZN(n3248) );
  OAI22_X1 U3733 ( .A1(n3321), .A2(n3810), .B1(n3809), .B2(n3248), .ZN(n3173)
         );
  AOI21_X1 U3734 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3191), .A(n3173), .ZN(n3174)
         );
  OAI211_X1 U3735 ( .C1(n3743), .C2(n3236), .A(n3175), .B(n3174), .ZN(U3219)
         );
  NAND2_X1 U3736 ( .A1(n3565), .A2(REG2_REG_23__SCAN_IN), .ZN(n3183) );
  INV_X1 U3737 ( .A(REG1_REG_23__SCAN_IN), .ZN(n3176) );
  OR2_X1 U3738 ( .A1(n3195), .A2(n3176), .ZN(n3182) );
  INV_X1 U3739 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4603) );
  NAND2_X1 U3740 ( .A1(n3177), .A2(n4603), .ZN(n3178) );
  NAND2_X1 U3741 ( .A1(n3196), .A2(n3178), .ZN(n4170) );
  INV_X1 U3742 ( .A(REG0_REG_23__SCAN_IN), .ZN(n3179) );
  OR2_X1 U3743 ( .A1(n3822), .A2(n3179), .ZN(n3180) );
  NAND2_X1 U3744 ( .A1(n3984), .A2(DATAO_REG_23__SCAN_IN), .ZN(n3184) );
  OAI21_X1 U3745 ( .B1(n4182), .B2(n3984), .A(n3184), .ZN(U3573) );
  AOI21_X1 U3746 ( .B1(n3187), .B2(n3186), .A(n3185), .ZN(n3193) );
  OAI22_X1 U3747 ( .A1(n3266), .A2(n3809), .B1(n3810), .B2(n3188), .ZN(n3190)
         );
  NOR2_X1 U3748 ( .A1(n3743), .A2(n2824), .ZN(n3189) );
  AOI211_X1 U3749 ( .C1(REG3_REG_2__SCAN_IN), .C2(n3191), .A(n3190), .B(n3189), 
        .ZN(n3192) );
  OAI21_X1 U3750 ( .B1(n3193), .B2(n3815), .A(n3192), .ZN(U3234) );
  NAND2_X1 U3751 ( .A1(n3565), .A2(REG2_REG_24__SCAN_IN), .ZN(n3202) );
  INV_X1 U3752 ( .A(REG1_REG_24__SCAN_IN), .ZN(n3194) );
  OR2_X1 U3753 ( .A1(n3195), .A2(n3194), .ZN(n3201) );
  INV_X1 U3754 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3752) );
  NAND2_X1 U3755 ( .A1(n3196), .A2(n3752), .ZN(n3197) );
  NAND2_X1 U3756 ( .A1(n3212), .A2(n3197), .ZN(n4150) );
  INV_X1 U3757 ( .A(REG0_REG_24__SCAN_IN), .ZN(n3198) );
  OR2_X1 U3758 ( .A1(n3822), .A2(n3198), .ZN(n3199) );
  NAND2_X1 U3759 ( .A1(n3984), .A2(DATAO_REG_24__SCAN_IN), .ZN(n3203) );
  OAI21_X1 U3760 ( .B1(n4164), .B2(n3984), .A(n3203), .ZN(U3574) );
  NAND2_X1 U3761 ( .A1(n2843), .A2(REG1_REG_25__SCAN_IN), .ZN(n3208) );
  INV_X1 U3762 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3540) );
  OR2_X1 U3763 ( .A1(n3826), .A2(n3540), .ZN(n3207) );
  INV_X1 U3764 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4617) );
  XNOR2_X1 U3765 ( .A(n3212), .B(n4617), .ZN(n3723) );
  INV_X1 U3766 ( .A(REG0_REG_25__SCAN_IN), .ZN(n3204) );
  OR2_X1 U3767 ( .A1(n3822), .A2(n3204), .ZN(n3205) );
  NAND2_X1 U3768 ( .A1(n3984), .A2(DATAO_REG_25__SCAN_IN), .ZN(n3209) );
  OAI21_X1 U3769 ( .B1(n4141), .B2(n3984), .A(n3209), .ZN(U3575) );
  NAND2_X1 U3770 ( .A1(n3565), .A2(REG2_REG_26__SCAN_IN), .ZN(n3218) );
  INV_X1 U3771 ( .A(REG1_REG_26__SCAN_IN), .ZN(n3210) );
  OR2_X1 U3772 ( .A1(n3195), .A2(n3210), .ZN(n3217) );
  NAND2_X1 U3773 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n3211) );
  INV_X1 U3774 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3808) );
  OAI21_X1 U3775 ( .B1(n3212), .B2(n4617), .A(n3808), .ZN(n3213) );
  NAND2_X1 U3776 ( .A1(n3567), .A2(n3213), .ZN(n4134) );
  INV_X1 U3777 ( .A(REG0_REG_26__SCAN_IN), .ZN(n3214) );
  OR2_X1 U3778 ( .A1(n3822), .A2(n3214), .ZN(n3215) );
  NAND2_X1 U3779 ( .A1(n3984), .A2(DATAO_REG_26__SCAN_IN), .ZN(n3219) );
  OAI21_X1 U3780 ( .B1(n4105), .B2(n3984), .A(n3219), .ZN(U3576) );
  XOR2_X1 U3781 ( .A(n3221), .B(n3220), .Z(n3225) );
  INV_X1 U3782 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U3783 ( .A1(n3796), .A2(n3252), .B1(n5159), .B2(n5010), .ZN(n3224)
         );
  NOR2_X1 U3784 ( .A1(STATE_REG_SCAN_IN), .A2(n3252), .ZN(n4835) );
  INV_X1 U3785 ( .A(n3991), .ZN(n3275) );
  NOR2_X1 U3786 ( .A1(n3809), .A2(n3275), .ZN(n3222) );
  AOI211_X1 U3787 ( .C1(n3285), .C2(n5163), .A(n4835), .B(n3222), .ZN(n3223)
         );
  OAI211_X1 U3788 ( .C1(n3225), .C2(n3815), .A(n3224), .B(n3223), .ZN(U3215)
         );
  INV_X1 U3789 ( .A(n3226), .ZN(n3227) );
  NAND2_X1 U3790 ( .A1(n3227), .A2(n4342), .ZN(n3229) );
  NAND2_X1 U3791 ( .A1(n3228), .A2(n4777), .ZN(n4312) );
  NOR2_X1 U3792 ( .A1(n5029), .A2(n5028), .ZN(n3231) );
  INV_X1 U3793 ( .A(n3231), .ZN(n5031) );
  NAND2_X1 U3794 ( .A1(n3231), .A2(n3239), .ZN(n3296) );
  INV_X1 U3795 ( .A(n3296), .ZN(n3232) );
  AOI211_X1 U3796 ( .C1(n3285), .C2(n5031), .A(n5204), .B(n3232), .ZN(n5052)
         );
  INV_X1 U3797 ( .A(n5052), .ZN(n3255) );
  OR2_X1 U3798 ( .A1(n3113), .A2(n3886), .ZN(n3235) );
  OR2_X1 U3799 ( .A1(n5219), .A2(n3233), .ZN(n3234) );
  NAND2_X1 U3800 ( .A1(n3237), .A2(n3236), .ZN(n3921) );
  INV_X1 U3801 ( .A(n5012), .ZN(n5007) );
  OR2_X1 U3802 ( .A1(n3992), .A2(n3328), .ZN(n3322) );
  INV_X1 U3803 ( .A(n3322), .ZN(n5006) );
  NAND2_X1 U3804 ( .A1(n5007), .A2(n5006), .ZN(n5037) );
  NAND2_X1 U3805 ( .A1(n5037), .A2(n5036), .ZN(n3238) );
  NAND2_X1 U3806 ( .A1(n5010), .A2(n2824), .ZN(n3925) );
  OR2_X1 U3807 ( .A1(n5034), .A2(n3239), .ZN(n3928) );
  NAND2_X1 U3808 ( .A1(n5034), .A2(n3239), .ZN(n3926) );
  NAND2_X1 U3809 ( .A1(n3928), .A2(n3926), .ZN(n3287) );
  INV_X1 U3810 ( .A(n3287), .ZN(n3875) );
  AND2_X1 U3811 ( .A1(n3992), .A2(n5004), .ZN(n5013) );
  NAND2_X1 U3812 ( .A1(n5012), .A2(n5013), .ZN(n5011) );
  NAND2_X1 U3813 ( .A1(n3237), .A2(n5014), .ZN(n3240) );
  OR2_X1 U3814 ( .A1(n5010), .A2(n5028), .ZN(n3241) );
  NAND2_X1 U3815 ( .A1(n5033), .A2(n3241), .ZN(n3288) );
  INV_X1 U3816 ( .A(n3288), .ZN(n3243) );
  NAND2_X1 U3817 ( .A1(n3243), .A2(n5227), .ZN(n3246) );
  AND2_X1 U3818 ( .A1(n5008), .A2(n3923), .ZN(n3244) );
  AOI22_X1 U3819 ( .A1(n3288), .A2(n5227), .B1(n5039), .B2(n3244), .ZN(n3245)
         );
  MUX2_X1 U3820 ( .A(n3246), .B(n3245), .S(n3287), .Z(n3251) );
  NAND2_X1 U3821 ( .A1(n3247), .A2(n3127), .ZN(n5210) );
  OAI22_X1 U3822 ( .A1(n3248), .A2(n5212), .B1(n3275), .B2(n5210), .ZN(n3249)
         );
  AOI21_X1 U3823 ( .B1(n3285), .B2(n5240), .A(n3249), .ZN(n3250) );
  OAI211_X1 U3824 ( .C1(n5217), .C2(n3282), .A(n3251), .B(n3250), .ZN(n5053)
         );
  NAND2_X1 U3825 ( .A1(n5053), .A2(n4242), .ZN(n3254) );
  INV_X2 U3826 ( .A(n4242), .ZN(n5249) );
  AOI22_X1 U3827 ( .A1(n5249), .A2(REG2_REG_3__SCAN_IN), .B1(n5135), .B2(n3252), .ZN(n3253) );
  OAI211_X1 U3828 ( .C1(n4278), .C2(n3255), .A(n3254), .B(n3253), .ZN(U3287)
         );
  NAND2_X1 U3829 ( .A1(n2843), .A2(REG1_REG_29__SCAN_IN), .ZN(n3261) );
  INV_X1 U3830 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3256) );
  OR2_X1 U3831 ( .A1(n3822), .A2(n3256), .ZN(n3260) );
  INV_X1 U3832 ( .A(n3567), .ZN(n3257) );
  NAND2_X1 U3833 ( .A1(n3257), .A2(REG3_REG_27__SCAN_IN), .ZN(n3579) );
  INV_X1 U3834 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4417) );
  OR2_X1 U3835 ( .A1(n2842), .A2(n3620), .ZN(n3259) );
  INV_X1 U3836 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3621) );
  OR2_X1 U3837 ( .A1(n3826), .A2(n3621), .ZN(n3258) );
  NAND2_X1 U3838 ( .A1(n3984), .A2(DATAO_REG_29__SCAN_IN), .ZN(n3262) );
  OAI21_X1 U3839 ( .B1(n3833), .B2(n3984), .A(n3262), .ZN(U3579) );
  AOI211_X1 U3840 ( .C1(n3265), .C2(n3264), .A(n3815), .B(n3263), .ZN(n3271)
         );
  OAI22_X1 U3841 ( .A1(n5177), .A2(n3297), .B1(n3810), .B2(n3266), .ZN(n3270)
         );
  INV_X1 U3842 ( .A(n3309), .ZN(n3281) );
  INV_X1 U3843 ( .A(REG3_REG_4__SCAN_IN), .ZN(n3267) );
  NOR2_X1 U3844 ( .A1(STATE_REG_SCAN_IN), .A2(n3267), .ZN(n4986) );
  AOI21_X1 U3845 ( .B1(n5161), .B2(n3990), .A(n4986), .ZN(n3268) );
  OAI21_X1 U3846 ( .B1(n3743), .B2(n3281), .A(n3268), .ZN(n3269) );
  OR3_X1 U3847 ( .A1(n3271), .A2(n3270), .A3(n3269), .ZN(U3227) );
  OAI21_X1 U3848 ( .B1(n3274), .B2(n3273), .A(n3272), .ZN(n3279) );
  OAI22_X1 U3849 ( .A1(n5177), .A2(n3358), .B1(n3810), .B2(n3275), .ZN(n3278)
         );
  AND2_X1 U3850 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4846) );
  AOI21_X1 U3851 ( .B1(n5161), .B2(n3989), .A(n4846), .ZN(n3276) );
  OAI21_X1 U3852 ( .B1(n3743), .B2(n3903), .A(n3276), .ZN(n3277) );
  AOI211_X1 U3853 ( .C1(n3279), .C2(n5172), .A(n3278), .B(n3277), .ZN(n3280)
         );
  INV_X1 U3854 ( .A(n3280), .ZN(U3224) );
  NAND2_X1 U3855 ( .A1(n3991), .A2(n3281), .ZN(n3932) );
  NAND2_X1 U3856 ( .A1(n3929), .A2(n3932), .ZN(n3289) );
  INV_X1 U3857 ( .A(n3289), .ZN(n3876) );
  INV_X1 U3858 ( .A(n3302), .ZN(n3284) );
  AND3_X1 U3859 ( .A1(n3282), .A2(n3289), .A3(n3928), .ZN(n3283) );
  OAI21_X1 U3860 ( .B1(n3284), .B2(n3283), .A(n5008), .ZN(n3294) );
  AOI22_X1 U3861 ( .A1(n5120), .A2(n5034), .B1(n3990), .B2(n5117), .ZN(n3293)
         );
  NOR2_X1 U3862 ( .A1(n5034), .A2(n3285), .ZN(n3286) );
  OAI211_X1 U3863 ( .C1(n3290), .C2(n3289), .A(n3311), .B(n5227), .ZN(n3292)
         );
  NAND2_X1 U3864 ( .A1(n5240), .A2(n3309), .ZN(n3291) );
  NAND4_X1 U3865 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n5056)
         );
  INV_X1 U3866 ( .A(n5056), .ZN(n3301) );
  INV_X1 U3867 ( .A(n3356), .ZN(n3295) );
  AOI211_X1 U3868 ( .C1(n3309), .C2(n3296), .A(n5204), .B(n3295), .ZN(n5055)
         );
  INV_X1 U3869 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3298) );
  OAI22_X1 U3870 ( .A1(n4242), .A2(n3298), .B1(n3297), .B2(n5224), .ZN(n3299)
         );
  AOI21_X1 U3871 ( .B1(n5055), .B2(n4260), .A(n3299), .ZN(n3300) );
  OAI21_X1 U3872 ( .B1(n3301), .B2(n5249), .A(n3300), .ZN(U3286) );
  INV_X1 U3873 ( .A(n3681), .ZN(n3308) );
  XNOR2_X1 U3874 ( .A(n3990), .B(n3357), .ZN(n3895) );
  NAND2_X1 U3875 ( .A1(n3302), .A2(n2745), .ZN(n3303) );
  NAND2_X1 U3876 ( .A1(n3990), .A2(n3903), .ZN(n3931) );
  NAND2_X1 U3877 ( .A1(n3989), .A2(n3367), .ZN(n3933) );
  INV_X1 U3878 ( .A(n3933), .ZN(n3304) );
  OR2_X1 U3879 ( .A1(n3989), .A2(n3367), .ZN(n3935) );
  OR2_X1 U3880 ( .A1(n3988), .A2(n3308), .ZN(n3936) );
  NAND2_X1 U3881 ( .A1(n3988), .A2(n3308), .ZN(n3904) );
  XNOR2_X1 U3882 ( .A(n3339), .B(n3874), .ZN(n3305) );
  NAND2_X1 U3883 ( .A1(n3305), .A2(n5008), .ZN(n3307) );
  AOI22_X1 U3884 ( .A1(n5120), .A2(n3989), .B1(n3987), .B2(n5117), .ZN(n3306)
         );
  OAI211_X1 U3885 ( .C1(n5123), .C2(n3308), .A(n3307), .B(n3306), .ZN(n5074)
         );
  INV_X1 U3886 ( .A(n5074), .ZN(n3320) );
  NAND2_X1 U3887 ( .A1(n3991), .A2(n3309), .ZN(n3310) );
  OR2_X1 U3888 ( .A1(n3990), .A2(n3357), .ZN(n3312) );
  NAND2_X1 U3889 ( .A1(n3990), .A2(n3357), .ZN(n3313) );
  NAND2_X1 U3890 ( .A1(n3314), .A2(n3313), .ZN(n3363) );
  OR2_X1 U3891 ( .A1(n3989), .A2(n3374), .ZN(n3315) );
  XOR2_X1 U3892 ( .A(n3874), .B(n3338), .Z(n5076) );
  INV_X1 U3893 ( .A(n4282), .ZN(n5201) );
  NAND2_X1 U3894 ( .A1(n5076), .A2(n5201), .ZN(n3319) );
  INV_X1 U3895 ( .A(n3346), .ZN(n3316) );
  AOI211_X1 U3896 ( .C1(n3681), .C2(n3366), .A(n5204), .B(n3316), .ZN(n5075)
         );
  INV_X1 U3897 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4026) );
  OAI22_X1 U3898 ( .A1(n4242), .A2(n4026), .B1(n3677), .B2(n5224), .ZN(n3317)
         );
  AOI21_X1 U3899 ( .B1(n5075), .B2(n4260), .A(n3317), .ZN(n3318) );
  OAI211_X1 U3900 ( .C1(n5249), .C2(n3320), .A(n3319), .B(n3318), .ZN(U3283)
         );
  AOI22_X1 U3901 ( .A1(n4260), .A2(n2504), .B1(n5240), .B2(n4242), .ZN(n3329)
         );
  NOR2_X1 U3902 ( .A1(n5227), .A2(n5008), .ZN(n3323) );
  NAND2_X1 U3903 ( .A1(n3992), .A2(n3328), .ZN(n3922) );
  AND2_X1 U3904 ( .A1(n3322), .A2(n3922), .ZN(n3869) );
  OAI22_X1 U3905 ( .A1(n3323), .A2(n3869), .B1(n3188), .B2(n5210), .ZN(n5001)
         );
  OAI22_X1 U3906 ( .A1(n4242), .A2(n3325), .B1(n3324), .B2(n5224), .ZN(n3326)
         );
  AOI21_X1 U3907 ( .B1(n5140), .B2(n5001), .A(n3326), .ZN(n3327) );
  OAI21_X1 U3908 ( .B1(n3329), .B2(n3328), .A(n3327), .ZN(U3290) );
  XOR2_X1 U3909 ( .A(n3331), .B(n3330), .Z(n3337) );
  INV_X1 U3910 ( .A(n3369), .ZN(n3332) );
  AOI22_X1 U3911 ( .A1(n3796), .A2(n3332), .B1(n5159), .B2(n3990), .ZN(n3336)
         );
  INV_X1 U3912 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3333) );
  NOR2_X1 U3913 ( .A1(STATE_REG_SCAN_IN), .A2(n3333), .ZN(n4848) );
  NOR2_X1 U3914 ( .A1(n3743), .A2(n3367), .ZN(n3334) );
  AOI211_X1 U3915 ( .C1(n5161), .C2(n3988), .A(n4848), .B(n3334), .ZN(n3335)
         );
  OAI211_X1 U3916 ( .C1(n3337), .C2(n3815), .A(n3336), .B(n3335), .ZN(U3236)
         );
  AND2_X1 U3917 ( .A1(n3987), .A2(n3341), .ZN(n3380) );
  INV_X1 U3918 ( .A(n3380), .ZN(n3905) );
  OR2_X1 U3919 ( .A1(n3987), .A2(n3341), .ZN(n3939) );
  AND2_X1 U3920 ( .A1(n3905), .A2(n3939), .ZN(n3867) );
  XOR2_X1 U3921 ( .A(n3867), .B(n3386), .Z(n3345) );
  XOR2_X1 U3922 ( .A(n3867), .B(n3381), .Z(n3343) );
  AOI22_X1 U3923 ( .A1(n5117), .A2(n3986), .B1(n3988), .B2(n5120), .ZN(n3340)
         );
  OAI21_X1 U3924 ( .B1(n5123), .B2(n3341), .A(n3340), .ZN(n3342) );
  AOI21_X1 U3925 ( .B1(n3343), .B2(n5008), .A(n3342), .ZN(n3344) );
  OAI21_X1 U3926 ( .B1(n3345), .B2(n5144), .A(n3344), .ZN(n5081) );
  INV_X1 U3927 ( .A(n5081), .ZN(n3349) );
  AOI211_X1 U3928 ( .C1(n3398), .C2(n3346), .A(n5204), .B(n2524), .ZN(n5080)
         );
  OAI22_X1 U3929 ( .A1(n4242), .A2(n2782), .B1(n3395), .B2(n5224), .ZN(n3347)
         );
  AOI21_X1 U3930 ( .B1(n5080), .B2(n4260), .A(n3347), .ZN(n3348) );
  OAI21_X1 U3931 ( .B1(n3349), .B2(n5249), .A(n3348), .ZN(U3282) );
  INV_X1 U3932 ( .A(n3895), .ZN(n3350) );
  XNOR2_X1 U3933 ( .A(n3351), .B(n3350), .ZN(n5060) );
  NAND2_X1 U3934 ( .A1(n3302), .A2(n3929), .ZN(n3352) );
  XNOR2_X1 U3935 ( .A(n3352), .B(n3895), .ZN(n3353) );
  NAND2_X1 U3936 ( .A1(n3353), .A2(n5008), .ZN(n3355) );
  AOI22_X1 U3937 ( .A1(n5117), .A2(n3989), .B1(n3991), .B2(n5120), .ZN(n3354)
         );
  OAI211_X1 U3938 ( .C1(n5123), .C2(n3903), .A(n3355), .B(n3354), .ZN(n5062)
         );
  NAND2_X1 U3939 ( .A1(n5062), .A2(n4242), .ZN(n3362) );
  NOR2_X2 U3940 ( .A1(n4278), .A2(n5204), .ZN(n5247) );
  AOI21_X1 U3941 ( .B1(n3357), .B2(n3356), .A(n3368), .ZN(n5063) );
  OAI22_X1 U3942 ( .A1(n4242), .A2(n3359), .B1(n3358), .B2(n5224), .ZN(n3360)
         );
  AOI21_X1 U3943 ( .B1(n5247), .B2(n5063), .A(n3360), .ZN(n3361) );
  OAI211_X1 U3944 ( .C1(n4282), .C2(n5060), .A(n3362), .B(n3361), .ZN(U3285)
         );
  INV_X1 U3945 ( .A(n3364), .ZN(n3365) );
  AOI21_X1 U3946 ( .B1(n3873), .B2(n3363), .A(n3365), .ZN(n5068) );
  OAI21_X1 U3947 ( .B1(n3368), .B2(n3367), .A(n3366), .ZN(n5067) );
  INV_X1 U3948 ( .A(n5067), .ZN(n3372) );
  OAI22_X1 U3949 ( .A1(n5140), .A2(n3370), .B1(n3369), .B2(n5224), .ZN(n3371)
         );
  AOI21_X1 U3950 ( .B1(n5247), .B2(n3372), .A(n3371), .ZN(n3379) );
  XNOR2_X1 U3951 ( .A(n3373), .B(n3873), .ZN(n3377) );
  AOI22_X1 U3952 ( .A1(n5120), .A2(n3990), .B1(n3988), .B2(n5117), .ZN(n3376)
         );
  NAND2_X1 U3953 ( .A1(n5240), .A2(n3374), .ZN(n3375) );
  OAI211_X1 U3954 ( .C1(n3377), .C2(n5217), .A(n3376), .B(n3375), .ZN(n5069)
         );
  NAND2_X1 U3955 ( .A1(n5069), .A2(n4242), .ZN(n3378) );
  OAI211_X1 U3956 ( .C1(n5068), .C2(n4282), .A(n3379), .B(n3378), .ZN(U3284)
         );
  OR2_X1 U3957 ( .A1(n3986), .A2(n3406), .ZN(n3938) );
  NAND2_X1 U3958 ( .A1(n3986), .A2(n3406), .ZN(n3945) );
  NAND2_X1 U3959 ( .A1(n3938), .A2(n3945), .ZN(n3411) );
  INV_X1 U3960 ( .A(n3411), .ZN(n3877) );
  XNOR2_X1 U3961 ( .A(n3418), .B(n3877), .ZN(n3384) );
  AOI22_X1 U3962 ( .A1(n5120), .A2(n3987), .B1(n5119), .B2(n5117), .ZN(n3382)
         );
  OAI21_X1 U3963 ( .B1(n5123), .B2(n3406), .A(n3382), .ZN(n3383) );
  AOI21_X1 U3964 ( .B1(n3384), .B2(n5008), .A(n3383), .ZN(n5086) );
  AND2_X1 U3965 ( .A1(n3987), .A2(n3398), .ZN(n3385) );
  XNOR2_X1 U3966 ( .A(n3412), .B(n3411), .ZN(n5089) );
  NAND2_X1 U3967 ( .A1(n5089), .A2(n5201), .ZN(n3392) );
  NOR2_X1 U3968 ( .A1(n2524), .A2(n3406), .ZN(n3387) );
  OR2_X1 U3969 ( .A1(n5093), .A2(n3387), .ZN(n5087) );
  INV_X1 U3970 ( .A(n5087), .ZN(n3390) );
  OAI22_X1 U3971 ( .A1(n4242), .A2(n3388), .B1(n3404), .B2(n5224), .ZN(n3389)
         );
  AOI21_X1 U3972 ( .B1(n3390), .B2(n5247), .A(n3389), .ZN(n3391) );
  OAI211_X1 U3973 ( .C1(n5086), .C2(n5249), .A(n3392), .B(n3391), .ZN(U3281)
         );
  AOI21_X1 U3974 ( .B1(n3394), .B2(n3393), .A(n2518), .ZN(n3401) );
  INV_X1 U3975 ( .A(n3395), .ZN(n3396) );
  AOI22_X1 U3976 ( .A1(n3796), .A2(n3396), .B1(n5159), .B2(n3988), .ZN(n3400)
         );
  NOR2_X1 U3977 ( .A1(STATE_REG_SCAN_IN), .A2(n4416), .ZN(n4870) );
  NOR2_X1 U3978 ( .A1(n3809), .A2(n5100), .ZN(n3397) );
  AOI211_X1 U3979 ( .C1(n3398), .C2(n5163), .A(n4870), .B(n3397), .ZN(n3399)
         );
  OAI211_X1 U3980 ( .C1(n3401), .C2(n3815), .A(n3400), .B(n3399), .ZN(U3218)
         );
  XOR2_X1 U3981 ( .A(n3403), .B(n3402), .Z(n3410) );
  INV_X1 U3982 ( .A(n3404), .ZN(n3405) );
  AOI22_X1 U3983 ( .A1(n3796), .A2(n3405), .B1(n5159), .B2(n3987), .ZN(n3409)
         );
  NOR2_X1 U3984 ( .A1(STATE_REG_SCAN_IN), .A2(n4435), .ZN(n4889) );
  NOR2_X1 U3985 ( .A1(n3743), .A2(n3406), .ZN(n3407) );
  AOI211_X1 U3986 ( .C1(n5161), .C2(n5119), .A(n4889), .B(n3407), .ZN(n3408)
         );
  OAI211_X1 U3987 ( .C1(n3410), .C2(n3815), .A(n3409), .B(n3408), .ZN(U3228)
         );
  OR2_X1 U3988 ( .A1(n3986), .A2(n3413), .ZN(n3414) );
  XNOR2_X1 U3989 ( .A(n5119), .B(n5102), .ZN(n5096) );
  OR2_X1 U3990 ( .A1(n3985), .A2(n5122), .ZN(n3915) );
  NAND2_X1 U3991 ( .A1(n3985), .A2(n5122), .ZN(n3909) );
  NAND2_X1 U3992 ( .A1(n2503), .A2(n3416), .ZN(n5116) );
  OR2_X1 U3993 ( .A1(n3985), .A2(n5115), .ZN(n3417) );
  NAND2_X1 U3994 ( .A1(n5116), .A2(n3417), .ZN(n3432) );
  NAND2_X1 U3995 ( .A1(n5118), .A2(n3467), .ZN(n3477) );
  NAND2_X1 U3996 ( .A1(n3916), .A2(n3477), .ZN(n3431) );
  INV_X1 U3997 ( .A(n3431), .ZN(n3878) );
  XNOR2_X1 U3998 ( .A(n3432), .B(n3878), .ZN(n5145) );
  INV_X1 U3999 ( .A(n3418), .ZN(n3419) );
  NAND2_X1 U4000 ( .A1(n5119), .A2(n5092), .ZN(n3908) );
  NAND2_X1 U4001 ( .A1(n5125), .A2(n5126), .ZN(n3420) );
  INV_X1 U4002 ( .A(n3479), .ZN(n3421) );
  NAND2_X1 U4003 ( .A1(n3421), .A2(n3477), .ZN(n3422) );
  OAI211_X1 U4004 ( .C1(n3878), .C2(n3423), .A(n3422), .B(n5008), .ZN(n3425)
         );
  AOI22_X1 U4005 ( .A1(n4288), .A2(n5117), .B1(n5120), .B2(n3985), .ZN(n3424)
         );
  OAI211_X1 U4006 ( .C1(n5123), .C2(n3467), .A(n3425), .B(n3424), .ZN(n5147)
         );
  NAND2_X1 U4007 ( .A1(n5147), .A2(n4242), .ZN(n3430) );
  AND2_X1 U4008 ( .A1(n5112), .A2(n3433), .ZN(n3426) );
  NOR2_X1 U4009 ( .A1(n3436), .A2(n3426), .ZN(n5148) );
  OAI22_X1 U4010 ( .A1(n4242), .A2(n3427), .B1(n3464), .B2(n5224), .ZN(n3428)
         );
  AOI21_X1 U4011 ( .B1(n5148), .B2(n5247), .A(n3428), .ZN(n3429) );
  OAI211_X1 U4012 ( .C1(n5145), .C2(n4282), .A(n3430), .B(n3429), .ZN(U3278)
         );
  OR2_X1 U4013 ( .A1(n5118), .A2(n3433), .ZN(n3434) );
  XNOR2_X1 U4014 ( .A(n3480), .B(n3777), .ZN(n3890) );
  XNOR2_X1 U4015 ( .A(n3472), .B(n3890), .ZN(n5154) );
  INV_X1 U4016 ( .A(n5154), .ZN(n3446) );
  OAI21_X1 U4017 ( .B1(n3436), .B2(n3435), .A(n5252), .ZN(n3437) );
  NOR2_X1 U4018 ( .A1(n3437), .A2(n4285), .ZN(n5153) );
  INV_X1 U4019 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3438) );
  OAI22_X1 U4020 ( .A1(n5140), .A2(n3438), .B1(n3773), .B2(n5224), .ZN(n3439)
         );
  AOI21_X1 U4021 ( .B1(n5153), .B2(n4260), .A(n3439), .ZN(n3445) );
  NAND2_X1 U4022 ( .A1(n3479), .A2(n3477), .ZN(n3440) );
  XOR2_X1 U4023 ( .A(n3890), .B(n3440), .Z(n3443) );
  OAI22_X1 U4024 ( .A1(n3458), .A2(n5212), .B1(n3775), .B2(n5210), .ZN(n3441)
         );
  AOI21_X1 U4025 ( .B1(n3777), .B2(n5240), .A(n3441), .ZN(n3442) );
  OAI21_X1 U4026 ( .B1(n3443), .B2(n5217), .A(n3442), .ZN(n5152) );
  NAND2_X1 U4027 ( .A1(n5152), .A2(n4242), .ZN(n3444) );
  OAI211_X1 U4028 ( .C1(n3446), .C2(n4282), .A(n3445), .B(n3444), .ZN(U3277)
         );
  AOI211_X1 U4029 ( .C1(n3449), .C2(n3448), .A(n3815), .B(n3447), .ZN(n3453)
         );
  OAI22_X1 U4030 ( .A1(n5177), .A2(n5111), .B1(n3810), .B2(n5100), .ZN(n3452)
         );
  NOR2_X1 U4031 ( .A1(STATE_REG_SCAN_IN), .A2(n4602), .ZN(n4899) );
  AOI21_X1 U4032 ( .B1(n5161), .B2(n3985), .A(n4899), .ZN(n3450) );
  OAI21_X1 U4033 ( .B1(n3743), .B2(n5092), .A(n3450), .ZN(n3451) );
  OR3_X1 U4034 ( .A1(n3453), .A2(n3452), .A3(n3451), .ZN(U3214) );
  XNOR2_X1 U4035 ( .A(n2517), .B(n3454), .ZN(n3455) );
  XNOR2_X1 U4036 ( .A(n3456), .B(n3455), .ZN(n3462) );
  INV_X1 U4037 ( .A(n3457), .ZN(n5136) );
  AOI22_X1 U4038 ( .A1(n3796), .A2(n5136), .B1(n5159), .B2(n5119), .ZN(n3461)
         );
  AND2_X1 U4039 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4911) );
  NOR2_X1 U4040 ( .A1(n3809), .A2(n3458), .ZN(n3459) );
  AOI211_X1 U4041 ( .C1(n5115), .C2(n5163), .A(n4911), .B(n3459), .ZN(n3460)
         );
  OAI211_X1 U4042 ( .C1(n3462), .C2(n3815), .A(n3461), .B(n3460), .ZN(U3233)
         );
  OAI21_X1 U40430 ( .B1(n3463), .B2(n2523), .A(n3771), .ZN(n3470) );
  OAI22_X1 U4044 ( .A1(n5177), .A2(n3464), .B1(n3810), .B2(n5099), .ZN(n3469)
         );
  INV_X1 U4045 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3465) );
  NOR2_X1 U4046 ( .A1(STATE_REG_SCAN_IN), .A2(n3465), .ZN(n4920) );
  AOI21_X1 U4047 ( .B1(n5161), .B2(n4288), .A(n4920), .ZN(n3466) );
  OAI21_X1 U4048 ( .B1(n3743), .B2(n3467), .A(n3466), .ZN(n3468) );
  AOI211_X1 U4049 ( .C1(n3470), .C2(n5172), .A(n3469), .B(n3468), .ZN(n3471)
         );
  INV_X1 U4050 ( .A(n3471), .ZN(U3221) );
  NAND2_X1 U4051 ( .A1(n3775), .A2(n3473), .ZN(n3837) );
  NAND2_X1 U4052 ( .A1(n5158), .A2(n4290), .ZN(n3946) );
  NAND2_X1 U4053 ( .A1(n3475), .A2(n3474), .ZN(n4291) );
  NAND2_X1 U4054 ( .A1(n3775), .A2(n4290), .ZN(n3476) );
  NAND2_X1 U4055 ( .A1(n4291), .A2(n3476), .ZN(n3491) );
  XNOR2_X1 U4056 ( .A(n4287), .B(n3511), .ZN(n3512) );
  XNOR2_X1 U4057 ( .A(n3491), .B(n3512), .ZN(n5181) );
  INV_X1 U4058 ( .A(n5181), .ZN(n3489) );
  OR2_X1 U4059 ( .A1(n3480), .A2(n3777), .ZN(n3478) );
  AND2_X1 U4060 ( .A1(n3478), .A2(n3477), .ZN(n3913) );
  NAND2_X1 U4061 ( .A1(n3480), .A2(n3777), .ZN(n3912) );
  INV_X1 U4062 ( .A(n3512), .ZN(n3896) );
  XNOR2_X1 U4063 ( .A(n3513), .B(n3896), .ZN(n3481) );
  NAND2_X1 U4064 ( .A1(n3481), .A2(n5008), .ZN(n3483) );
  AOI22_X1 U4065 ( .A1(n5160), .A2(n5117), .B1(n5158), .B2(n5120), .ZN(n3482)
         );
  OAI211_X1 U4066 ( .C1(n5123), .C2(n3511), .A(n3483), .B(n3482), .ZN(n5179)
         );
  INV_X1 U4067 ( .A(n4284), .ZN(n3484) );
  OAI21_X1 U4068 ( .B1(n3484), .B2(n3511), .A(n4273), .ZN(n5178) );
  INV_X1 U4069 ( .A(n5247), .ZN(n4303) );
  INV_X1 U4070 ( .A(n5176), .ZN(n3485) );
  AOI22_X1 U4071 ( .A1(n5249), .A2(REG2_REG_15__SCAN_IN), .B1(n5135), .B2(
        n3485), .ZN(n3486) );
  OAI21_X1 U4072 ( .B1(n5178), .B2(n4303), .A(n3486), .ZN(n3487) );
  AOI21_X1 U4073 ( .B1(n5179), .B2(n5140), .A(n3487), .ZN(n3488) );
  OAI21_X1 U4074 ( .B1(n3489), .B2(n4282), .A(n3488), .ZN(U3275) );
  NAND2_X1 U4075 ( .A1(n4287), .A2(n5162), .ZN(n3490) );
  NAND2_X1 U4076 ( .A1(n3491), .A2(n3490), .ZN(n3493) );
  NAND2_X1 U4077 ( .A1(n4267), .A2(n3511), .ZN(n3492) );
  INV_X1 U4078 ( .A(n5160), .ZN(n4247) );
  NAND2_X1 U4079 ( .A1(n3495), .A2(n3742), .ZN(n3497) );
  OR2_X1 U4080 ( .A1(n3983), .A2(n4233), .ZN(n3520) );
  NAND2_X1 U4081 ( .A1(n3983), .A2(n4233), .ZN(n5206) );
  NAND2_X1 U4082 ( .A1(n3520), .A2(n5206), .ZN(n3885) );
  OR2_X1 U4083 ( .A1(n3983), .A2(n4240), .ZN(n3498) );
  NAND2_X1 U4084 ( .A1(n3499), .A2(n4230), .ZN(n3518) );
  NAND2_X1 U4085 ( .A1(n3762), .A2(n5215), .ZN(n3523) );
  NAND2_X1 U4086 ( .A1(n3518), .A2(n3523), .ZN(n5209) );
  NAND2_X1 U4087 ( .A1(n3499), .A2(n3762), .ZN(n3500) );
  AND2_X1 U4088 ( .A1(n5211), .A2(n3519), .ZN(n3502) );
  NOR2_X1 U4089 ( .A1(n4178), .A2(n3538), .ZN(n3503) );
  NAND2_X1 U4090 ( .A1(n4178), .A2(n3538), .ZN(n3504) );
  NAND2_X1 U4091 ( .A1(n2800), .A2(DATAI_22_), .ZN(n4191) );
  INV_X1 U4092 ( .A(n4191), .ZN(n4179) );
  OR2_X1 U4093 ( .A1(n4205), .A2(n4179), .ZN(n3528) );
  INV_X1 U4094 ( .A(n4160), .ZN(n3506) );
  OR2_X1 U4095 ( .A1(n4205), .A2(n4191), .ZN(n3507) );
  NAND2_X1 U4096 ( .A1(n2800), .A2(DATAI_23_), .ZN(n3632) );
  XNOR2_X1 U4097 ( .A(n4182), .B(n4166), .ZN(n4163) );
  OR2_X1 U4098 ( .A1(n4182), .A2(n3632), .ZN(n3558) );
  NAND2_X1 U4099 ( .A1(n2800), .A2(DATAI_24_), .ZN(n4149) );
  NAND2_X1 U4100 ( .A1(n4164), .A2(n4149), .ZN(n3552) );
  NAND2_X1 U4101 ( .A1(n4140), .A2(n3552), .ZN(n3508) );
  OR2_X1 U4102 ( .A1(n4164), .A2(n4149), .ZN(n3548) );
  NAND2_X1 U4103 ( .A1(n2800), .A2(DATAI_25_), .ZN(n3644) );
  NAND2_X1 U4104 ( .A1(n4141), .A2(n3644), .ZN(n3551) );
  NAND2_X1 U4105 ( .A1(n3547), .A2(n3551), .ZN(n3866) );
  INV_X1 U4106 ( .A(n3866), .ZN(n3509) );
  NAND2_X1 U4107 ( .A1(n4287), .A2(n3511), .ZN(n3944) );
  INV_X1 U4108 ( .A(n4272), .ZN(n3514) );
  OR2_X1 U4109 ( .A1(n5160), .A2(n3514), .ZN(n3902) );
  NAND2_X1 U4110 ( .A1(n5160), .A2(n3514), .ZN(n3841) );
  INV_X1 U4111 ( .A(n4246), .ZN(n3515) );
  NAND2_X1 U4112 ( .A1(n3515), .A2(n2526), .ZN(n3516) );
  OR2_X1 U4113 ( .A1(n4231), .A2(n3742), .ZN(n3872) );
  INV_X1 U4114 ( .A(n3520), .ZN(n3517) );
  AND2_X1 U4115 ( .A1(n3518), .A2(n5206), .ZN(n3843) );
  OR2_X1 U4116 ( .A1(n5211), .A2(n4224), .ZN(n3842) );
  NAND2_X1 U4117 ( .A1(n5211), .A2(n4224), .ZN(n3522) );
  NAND2_X1 U4118 ( .A1(n4213), .A2(n4221), .ZN(n3526) );
  NAND2_X1 U4119 ( .A1(n3872), .A2(n3520), .ZN(n3521) );
  NAND2_X1 U4120 ( .A1(n3843), .A2(n3521), .ZN(n3524) );
  NAND3_X1 U4121 ( .A1(n3524), .A2(n3523), .A3(n3522), .ZN(n3525) );
  NAND2_X1 U4122 ( .A1(n3525), .A2(n3842), .ZN(n3846) );
  INV_X1 U4123 ( .A(n3538), .ZN(n4207) );
  AND2_X1 U4124 ( .A1(n4178), .A2(n4207), .ZN(n4157) );
  OR2_X1 U4125 ( .A1(n4160), .A2(n4157), .ZN(n3844) );
  OR2_X1 U4126 ( .A1(n4178), .A2(n4207), .ZN(n4158) );
  OR2_X1 U4127 ( .A1(n4158), .A2(n4160), .ZN(n3530) );
  OR2_X1 U4128 ( .A1(n4182), .A2(n4166), .ZN(n3527) );
  AND2_X1 U4129 ( .A1(n3528), .A2(n3527), .ZN(n3529) );
  NAND2_X1 U4130 ( .A1(n3530), .A2(n3529), .ZN(n3959) );
  NAND2_X1 U4131 ( .A1(n4182), .A2(n4166), .ZN(n3956) );
  NAND2_X1 U4132 ( .A1(n4164), .A2(n4147), .ZN(n3957) );
  INV_X1 U4133 ( .A(n3957), .ZN(n3532) );
  OR2_X1 U4134 ( .A1(n4164), .A2(n4147), .ZN(n3884) );
  INV_X1 U4135 ( .A(n3884), .ZN(n3533) );
  NOR2_X1 U4136 ( .A1(n3576), .A2(n3533), .ZN(n3534) );
  XNOR2_X1 U4137 ( .A(n3534), .B(n3866), .ZN(n3537) );
  NOR2_X1 U4138 ( .A1(n5123), .A2(n3644), .ZN(n3536) );
  OAI22_X1 U4139 ( .A1(n4164), .A2(n5212), .B1(n4105), .B2(n5210), .ZN(n3535)
         );
  AOI211_X1 U4140 ( .C1(n3537), .C2(n5008), .A(n3536), .B(n3535), .ZN(n4321)
         );
  INV_X1 U4141 ( .A(n4321), .ZN(n3543) );
  OAI21_X1 U4142 ( .B1(n4148), .B2(n3644), .A(n5252), .ZN(n3539) );
  OR2_X1 U4143 ( .A1(n3539), .A2(n4133), .ZN(n4320) );
  NOR2_X1 U4144 ( .A1(n4320), .A2(n4278), .ZN(n3542) );
  OAI22_X1 U4145 ( .A1(n5140), .A2(n3540), .B1(n3723), .B2(n5224), .ZN(n3541)
         );
  AOI211_X1 U4146 ( .C1(n3543), .C2(n5140), .A(n3542), .B(n3541), .ZN(n3544)
         );
  OAI21_X1 U4147 ( .B1(n4322), .B2(n4282), .A(n3544), .ZN(U3265) );
  INV_X1 U4148 ( .A(DATAI_20_), .ZN(n3545) );
  MUX2_X1 U4149 ( .A(n3545), .B(n3113), .S(STATE_REG_SCAN_IN), .Z(n3546) );
  INV_X1 U4150 ( .A(n3546), .ZN(U3332) );
  INV_X1 U4151 ( .A(n3551), .ZN(n3550) );
  AND2_X1 U4152 ( .A1(n3548), .A2(n3547), .ZN(n3549) );
  NAND2_X1 U4153 ( .A1(n2800), .A2(DATAI_26_), .ZN(n4132) );
  INV_X1 U4154 ( .A(n4132), .ZN(n3813) );
  NOR2_X1 U4155 ( .A1(n4105), .A2(n3813), .ZN(n3818) );
  NAND2_X1 U4156 ( .A1(n4105), .A2(n3813), .ZN(n3850) );
  INV_X1 U4157 ( .A(n3850), .ZN(n3577) );
  OR2_X1 U4158 ( .A1(n3818), .A2(n3577), .ZN(n4123) );
  AND2_X1 U4159 ( .A1(n4121), .A2(n4123), .ZN(n3557) );
  INV_X1 U4160 ( .A(n3557), .ZN(n3553) );
  AND2_X1 U4161 ( .A1(n4163), .A2(n3556), .ZN(n3554) );
  NAND2_X1 U4162 ( .A1(n4105), .A2(n4132), .ZN(n3555) );
  AND2_X1 U4163 ( .A1(n3554), .A2(n3555), .ZN(n3563) );
  INV_X1 U4164 ( .A(n3555), .ZN(n3562) );
  INV_X1 U4165 ( .A(n3556), .ZN(n3560) );
  AND2_X1 U4166 ( .A1(n3558), .A2(n3557), .ZN(n3559) );
  NAND2_X1 U4167 ( .A1(n3565), .A2(REG2_REG_27__SCAN_IN), .ZN(n3573) );
  INV_X1 U4168 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3566) );
  OR2_X1 U4169 ( .A1(n3195), .A2(n3566), .ZN(n3572) );
  INV_X1 U4170 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U4171 ( .A1(n3567), .A2(n3688), .ZN(n3568) );
  NAND2_X1 U4172 ( .A1(n3579), .A2(n3568), .ZN(n4116) );
  INV_X1 U4173 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3569) );
  OR2_X1 U4174 ( .A1(n3822), .A2(n3569), .ZN(n3570) );
  INV_X1 U4175 ( .A(n4127), .ZN(n3982) );
  NAND2_X1 U4176 ( .A1(n2800), .A2(DATAI_27_), .ZN(n3657) );
  NOR2_X1 U4177 ( .A1(n3982), .A2(n4108), .ZN(n3574) );
  INV_X1 U4178 ( .A(n3644), .ZN(n3726) );
  OR2_X1 U4179 ( .A1(n4141), .A2(n3726), .ZN(n3575) );
  NAND2_X1 U4180 ( .A1(n4141), .A2(n3726), .ZN(n3849) );
  NAND2_X1 U4181 ( .A1(n4127), .A2(n4108), .ZN(n3851) );
  INV_X1 U4182 ( .A(n3851), .ZN(n3588) );
  NOR2_X1 U4183 ( .A1(n4127), .A2(n4108), .ZN(n3819) );
  NOR2_X1 U4184 ( .A1(n4101), .A2(n4115), .ZN(n4104) );
  NAND2_X1 U4185 ( .A1(n5008), .A2(n3851), .ZN(n3578) );
  OAI22_X1 U4186 ( .A1(n3601), .A2(n5144), .B1(n4104), .B2(n3578), .ZN(n3586)
         );
  NAND2_X1 U4187 ( .A1(n2843), .A2(REG1_REG_28__SCAN_IN), .ZN(n3585) );
  INV_X1 U4188 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3597) );
  OR2_X1 U4189 ( .A1(n3826), .A2(n3597), .ZN(n3584) );
  NAND2_X1 U4190 ( .A1(n3579), .A2(n4417), .ZN(n3580) );
  NAND2_X1 U4191 ( .A1(n3620), .A2(n3580), .ZN(n3669) );
  INV_X1 U4192 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3581) );
  OR2_X1 U4193 ( .A1(n3822), .A2(n3581), .ZN(n3582) );
  NAND2_X1 U4194 ( .A1(n2800), .A2(DATAI_28_), .ZN(n3663) );
  NAND2_X1 U4195 ( .A1(n4106), .A2(n3672), .ZN(n3852) );
  OR2_X1 U4196 ( .A1(n4106), .A2(n3672), .ZN(n3817) );
  NAND2_X1 U4197 ( .A1(n3852), .A2(n3817), .ZN(n3889) );
  INV_X1 U4198 ( .A(n3889), .ZN(n3587) );
  NAND3_X1 U4199 ( .A1(n3601), .A2(n5227), .A3(n3587), .ZN(n3594) );
  OAI22_X1 U4200 ( .A1(n3833), .A2(n5210), .B1(n4127), .B2(n5212), .ZN(n3589)
         );
  AOI21_X1 U4201 ( .B1(n3672), .B2(n5240), .A(n3589), .ZN(n3590) );
  INV_X1 U4202 ( .A(n3590), .ZN(n3591) );
  INV_X1 U4203 ( .A(n4099), .ZN(n3596) );
  INV_X1 U4204 ( .A(n3617), .ZN(n3618) );
  OAI211_X1 U4205 ( .C1(n3596), .C2(n3663), .A(n3618), .B(n5252), .ZN(n4313)
         );
  INV_X1 U4206 ( .A(n4313), .ZN(n3599) );
  OAI22_X1 U4207 ( .A1(n5140), .A2(n3597), .B1(n3669), .B2(n5224), .ZN(n3598)
         );
  AOI21_X1 U4208 ( .B1(n3599), .B2(n4260), .A(n3598), .ZN(n3600) );
  OAI21_X1 U4209 ( .B1(n4314), .B2(n5249), .A(n3600), .ZN(U3262) );
  INV_X1 U4210 ( .A(n4106), .ZN(n3981) );
  INV_X1 U4211 ( .A(DATAI_29_), .ZN(n3602) );
  NOR2_X1 U4212 ( .A1(n3603), .A2(n3602), .ZN(n3832) );
  XNOR2_X1 U4213 ( .A(n3833), .B(n3832), .ZN(n3891) );
  NAND2_X1 U4214 ( .A1(n3606), .A2(n3852), .ZN(n3607) );
  INV_X1 U4215 ( .A(n3832), .ZN(n3616) );
  INV_X1 U4216 ( .A(B_REG_SCAN_IN), .ZN(n3608) );
  NOR2_X1 U4217 ( .A1(n3143), .A2(n3608), .ZN(n3609) );
  NOR2_X1 U4218 ( .A1(n5210), .A2(n3609), .ZN(n5230) );
  INV_X1 U4219 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3613) );
  NAND2_X1 U4220 ( .A1(n2843), .A2(REG1_REG_30__SCAN_IN), .ZN(n3612) );
  INV_X1 U4221 ( .A(REG0_REG_30__SCAN_IN), .ZN(n3610) );
  OR2_X1 U4222 ( .A1(n3822), .A2(n3610), .ZN(n3611) );
  OAI211_X1 U4223 ( .C1(n3826), .C2(n3613), .A(n3612), .B(n3611), .ZN(n3980)
         );
  AOI22_X1 U4224 ( .A1(n3981), .A2(n5120), .B1(n5230), .B2(n3980), .ZN(n3614)
         );
  OAI21_X1 U4225 ( .B1(n5123), .B2(n3616), .A(n3614), .ZN(n3615) );
  NAND2_X1 U4226 ( .A1(n3617), .A2(n3616), .ZN(n5244) );
  AOI21_X1 U4227 ( .B1(n3618), .B2(n3832), .A(n5204), .ZN(n3619) );
  NOR2_X1 U4228 ( .A1(n4304), .A2(n4278), .ZN(n3623) );
  OAI22_X1 U4229 ( .A1(n5140), .A2(n3621), .B1(n3620), .B2(n5224), .ZN(n3622)
         );
  AOI211_X1 U4230 ( .C1(n3624), .C2(n5140), .A(n3623), .B(n3622), .ZN(n3625)
         );
  OAI21_X1 U4231 ( .B1(n4306), .B2(n4282), .A(n3625), .ZN(U3354) );
  OR2_X1 U4232 ( .A1(n2825), .A2(n4191), .ZN(n3626) );
  OAI21_X1 U4233 ( .B1(n3650), .B2(n4205), .A(n3626), .ZN(n3627) );
  XNOR2_X1 U4234 ( .A(n3627), .B(n2958), .ZN(n3634) );
  OAI22_X1 U4235 ( .A1(n3651), .A2(n4205), .B1(n3650), .B2(n4191), .ZN(n3633)
         );
  XNOR2_X1 U4236 ( .A(n3634), .B(n3633), .ZN(n3785) );
  NOR2_X1 U4237 ( .A1(n3785), .A2(n3628), .ZN(n3629) );
  NAND2_X1 U4238 ( .A1(n3782), .A2(n3629), .ZN(n3703) );
  OR2_X1 U4239 ( .A1(n2825), .A2(n3632), .ZN(n3630) );
  OAI21_X1 U4240 ( .B1(n3650), .B2(n4182), .A(n3630), .ZN(n3631) );
  XNOR2_X1 U4241 ( .A(n3631), .B(n2958), .ZN(n3637) );
  OAI22_X1 U4242 ( .A1(n3651), .A2(n4182), .B1(n3650), .B2(n3632), .ZN(n3636)
         );
  XNOR2_X1 U4243 ( .A(n3637), .B(n3636), .ZN(n3704) );
  NOR2_X1 U4244 ( .A1(n3634), .A2(n3633), .ZN(n3705) );
  NOR2_X1 U4245 ( .A1(n3704), .A2(n3705), .ZN(n3635) );
  NAND2_X1 U4246 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  OAI22_X1 U4247 ( .A1(n4164), .A2(n3650), .B1(n2825), .B2(n4149), .ZN(n3639)
         );
  XNOR2_X1 U4248 ( .A(n3639), .B(n2958), .ZN(n3640) );
  OR2_X1 U4249 ( .A1(n2825), .A2(n3644), .ZN(n3641) );
  OAI21_X1 U4250 ( .B1(n3650), .B2(n4141), .A(n3641), .ZN(n3643) );
  XNOR2_X1 U4251 ( .A(n3643), .B(n3642), .ZN(n3645) );
  OAI22_X1 U4252 ( .A1(n3651), .A2(n4141), .B1(n3650), .B2(n3644), .ZN(n3646)
         );
  XNOR2_X1 U4253 ( .A(n3645), .B(n3646), .ZN(n3719) );
  NAND2_X1 U4254 ( .A1(n3749), .A2(n3719), .ZN(n3653) );
  INV_X1 U4255 ( .A(n3645), .ZN(n3647) );
  OR2_X1 U4256 ( .A1(n3647), .A2(n3646), .ZN(n3802) );
  OR2_X1 U4257 ( .A1(n2825), .A2(n4132), .ZN(n3648) );
  OAI21_X1 U4258 ( .B1(n3650), .B2(n4105), .A(n3648), .ZN(n3649) );
  XNOR2_X1 U4259 ( .A(n3649), .B(n2958), .ZN(n3655) );
  OAI22_X1 U4260 ( .A1(n3651), .A2(n4105), .B1(n3650), .B2(n4132), .ZN(n3654)
         );
  OR2_X1 U4261 ( .A1(n3655), .A2(n3654), .ZN(n3805) );
  AND2_X1 U4262 ( .A1(n3802), .A2(n3805), .ZN(n3652) );
  NAND2_X1 U4263 ( .A1(n3655), .A2(n3654), .ZN(n3804) );
  NAND2_X1 U4264 ( .A1(n3656), .A2(n3804), .ZN(n3687) );
  OAI22_X1 U4265 ( .A1(n4127), .A2(n3650), .B1(n2825), .B2(n3657), .ZN(n3658)
         );
  XOR2_X1 U4266 ( .A(n2958), .B(n3658), .Z(n3660) );
  AOI22_X1 U4267 ( .A1(n2855), .A2(n3982), .B1(n3665), .B2(n4108), .ZN(n3659)
         );
  NOR2_X1 U4268 ( .A1(n3660), .A2(n3659), .ZN(n3661) );
  AOI21_X1 U4269 ( .B1(n3660), .B2(n3659), .A(n3661), .ZN(n3686) );
  INV_X1 U4270 ( .A(n3661), .ZN(n3662) );
  OAI22_X1 U4271 ( .A1(n4106), .A2(n3650), .B1(n2825), .B2(n3663), .ZN(n3664)
         );
  XNOR2_X1 U4272 ( .A(n3664), .B(n2958), .ZN(n3667) );
  AOI22_X1 U4273 ( .A1(n2855), .A2(n3981), .B1(n3665), .B2(n3672), .ZN(n3666)
         );
  XNOR2_X1 U4274 ( .A(n3667), .B(n3666), .ZN(n3668) );
  OAI22_X1 U4275 ( .A1(n3809), .A2(n3833), .B1(STATE_REG_SCAN_IN), .B2(n4417), 
        .ZN(n3671) );
  OAI22_X1 U4276 ( .A1(n5177), .A2(n3669), .B1(n3810), .B2(n4127), .ZN(n3670)
         );
  AOI211_X1 U4277 ( .C1(n3672), .C2(n5163), .A(n3671), .B(n3670), .ZN(n3673)
         );
  OAI211_X1 U4278 ( .C1(n3676), .C2(n3675), .A(n3674), .B(n5172), .ZN(n3684)
         );
  INV_X1 U4279 ( .A(n3677), .ZN(n3678) );
  AOI22_X1 U4280 ( .A1(n3796), .A2(n3678), .B1(n5159), .B2(n3989), .ZN(n3683)
         );
  AND2_X1 U4281 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4868) );
  NOR2_X1 U4282 ( .A1(n3809), .A2(n3679), .ZN(n3680) );
  AOI211_X1 U4283 ( .C1(n3681), .C2(n5163), .A(n4868), .B(n3680), .ZN(n3682)
         );
  NAND3_X1 U4284 ( .A1(n3684), .A2(n3683), .A3(n3682), .ZN(U3210) );
  OAI211_X1 U4285 ( .C1(n3687), .C2(n3686), .A(n3685), .B(n5172), .ZN(n3692)
         );
  OAI22_X1 U4286 ( .A1(n3809), .A2(n4106), .B1(STATE_REG_SCAN_IN), .B2(n3688), 
        .ZN(n3690) );
  OAI22_X1 U4287 ( .A1(n5177), .A2(n4116), .B1(n3810), .B2(n4105), .ZN(n3689)
         );
  AOI211_X1 U4288 ( .C1(n4108), .C2(n5163), .A(n3690), .B(n3689), .ZN(n3691)
         );
  NAND2_X1 U4289 ( .A1(n3692), .A2(n3691), .ZN(U3211) );
  OAI21_X1 U4290 ( .B1(n3695), .B2(n3694), .A(n3693), .ZN(n3701) );
  AOI22_X1 U4291 ( .A1(n3796), .A2(n3696), .B1(n5159), .B2(n4288), .ZN(n3699)
         );
  NOR2_X1 U4292 ( .A1(STATE_REG_SCAN_IN), .A2(n3697), .ZN(n4934) );
  AOI21_X1 U4293 ( .B1(n5161), .B2(n4287), .A(n4934), .ZN(n3698) );
  OAI211_X1 U4294 ( .C1(n3743), .C2(n4290), .A(n3699), .B(n3698), .ZN(n3700)
         );
  AOI21_X1 U4295 ( .B1(n3701), .B2(n5172), .A(n3700), .ZN(n3702) );
  INV_X1 U4296 ( .A(n3702), .ZN(U3212) );
  INV_X1 U4297 ( .A(n3703), .ZN(n3783) );
  OAI21_X1 U4298 ( .B1(n3783), .B2(n3705), .A(n3704), .ZN(n3707) );
  NAND3_X1 U4299 ( .A1(n3707), .A2(n5172), .A3(n3706), .ZN(n3711) );
  OAI22_X1 U4300 ( .A1(n3810), .A2(n4205), .B1(STATE_REG_SCAN_IN), .B2(n4603), 
        .ZN(n3709) );
  OAI22_X1 U4301 ( .A1(n5177), .A2(n4170), .B1(n3809), .B2(n4164), .ZN(n3708)
         );
  AOI211_X1 U4302 ( .C1(n4166), .C2(n5163), .A(n3709), .B(n3708), .ZN(n3710)
         );
  NAND2_X1 U4303 ( .A1(n3711), .A2(n3710), .ZN(U3213) );
  XOR2_X1 U4304 ( .A(n3713), .B(n3712), .Z(n3717) );
  NAND2_X1 U4305 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4094) );
  OAI21_X1 U4306 ( .B1(n3810), .B2(n5213), .A(n4094), .ZN(n3715) );
  OAI22_X1 U4307 ( .A1(n5177), .A2(n5223), .B1(n3809), .B2(n5211), .ZN(n3714)
         );
  AOI211_X1 U4308 ( .C1(n5215), .C2(n5163), .A(n3715), .B(n3714), .ZN(n3716)
         );
  OAI21_X1 U4309 ( .B1(n3717), .B2(n3815), .A(n3716), .ZN(U3216) );
  INV_X1 U4310 ( .A(n3803), .ZN(n3722) );
  AOI21_X1 U4311 ( .B1(n3720), .B2(n3749), .A(n3719), .ZN(n3721) );
  OAI21_X1 U4312 ( .B1(n3722), .B2(n3721), .A(n5172), .ZN(n3728) );
  OAI22_X1 U4313 ( .A1(n3810), .A2(n4164), .B1(STATE_REG_SCAN_IN), .B2(n4617), 
        .ZN(n3725) );
  OAI22_X1 U4314 ( .A1(n5177), .A2(n3723), .B1(n3809), .B2(n4105), .ZN(n3724)
         );
  AOI211_X1 U4315 ( .C1(n3726), .C2(n5163), .A(n3725), .B(n3724), .ZN(n3727)
         );
  NAND2_X1 U4316 ( .A1(n3728), .A2(n3727), .ZN(U3222) );
  NAND2_X1 U4317 ( .A1(n3730), .A2(n3729), .ZN(n3732) );
  NOR2_X1 U4318 ( .A1(n3732), .A2(n3733), .ZN(n3731) );
  AOI21_X1 U4319 ( .B1(n3733), .B2(n3732), .A(n3731), .ZN(n3737) );
  AOI22_X1 U4320 ( .A1(n3796), .A2(n4276), .B1(n5161), .B2(n4231), .ZN(n3736)
         );
  NOR2_X1 U4321 ( .A1(STATE_REG_SCAN_IN), .A2(n4427), .ZN(n4054) );
  NOR2_X1 U4322 ( .A1(n3810), .A2(n4267), .ZN(n3734) );
  AOI211_X1 U4323 ( .C1(n4272), .C2(n5163), .A(n4054), .B(n3734), .ZN(n3735)
         );
  OAI211_X1 U4324 ( .C1(n3737), .C2(n3815), .A(n3736), .B(n3735), .ZN(U3223)
         );
  OAI21_X1 U4325 ( .B1(n3740), .B2(n3738), .A(n3739), .ZN(n3746) );
  OAI22_X1 U4326 ( .A1(n5177), .A2(n4257), .B1(n3809), .B2(n5213), .ZN(n3745)
         );
  AND2_X1 U4327 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4071) );
  AOI21_X1 U4328 ( .B1(n5159), .B2(n5160), .A(n4071), .ZN(n3741) );
  OAI21_X1 U4329 ( .B1(n3743), .B2(n3742), .A(n3741), .ZN(n3744) );
  AOI211_X1 U4330 ( .C1(n3746), .C2(n5172), .A(n3745), .B(n3744), .ZN(n3747)
         );
  INV_X1 U4331 ( .A(n3747), .ZN(U3225) );
  NAND2_X1 U4332 ( .A1(n3748), .A2(n3749), .ZN(n3750) );
  XOR2_X1 U4333 ( .A(n3751), .B(n3750), .Z(n3756) );
  OAI22_X1 U4334 ( .A1(n3810), .A2(n4182), .B1(STATE_REG_SCAN_IN), .B2(n3752), 
        .ZN(n3754) );
  OAI22_X1 U4335 ( .A1(n5177), .A2(n4150), .B1(n3809), .B2(n4141), .ZN(n3753)
         );
  AOI211_X1 U4336 ( .C1(n4147), .C2(n5163), .A(n3754), .B(n3753), .ZN(n3755)
         );
  OAI21_X1 U4337 ( .B1(n3756), .B2(n3815), .A(n3755), .ZN(U3226) );
  INV_X1 U4338 ( .A(n3758), .ZN(n3760) );
  NAND2_X1 U4339 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  XNOR2_X1 U4340 ( .A(n3757), .B(n3761), .ZN(n3766) );
  OAI22_X1 U4341 ( .A1(n3810), .A2(n3762), .B1(STATE_REG_SCAN_IN), .B2(n4634), 
        .ZN(n3764) );
  OAI22_X1 U4342 ( .A1(n5177), .A2(n4222), .B1(n3809), .B2(n4178), .ZN(n3763)
         );
  AOI211_X1 U4343 ( .C1(n4224), .C2(n5163), .A(n3764), .B(n3763), .ZN(n3765)
         );
  OAI21_X1 U4344 ( .B1(n3766), .B2(n3815), .A(n3765), .ZN(U3230) );
  NOR2_X1 U4345 ( .A1(n3768), .A2(n3767), .ZN(n3772) );
  INV_X1 U4346 ( .A(n3769), .ZN(n3770) );
  AOI21_X1 U4347 ( .B1(n3772), .B2(n3771), .A(n3770), .ZN(n3780) );
  INV_X1 U4348 ( .A(n3773), .ZN(n3774) );
  AOI22_X1 U4349 ( .A1(n3796), .A2(n3774), .B1(n5159), .B2(n5118), .ZN(n3779)
         );
  INV_X1 U4350 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4633) );
  NOR2_X1 U4351 ( .A1(STATE_REG_SCAN_IN), .A2(n4633), .ZN(n4932) );
  NOR2_X1 U4352 ( .A1(n3809), .A2(n3775), .ZN(n3776) );
  AOI211_X1 U4353 ( .C1(n3777), .C2(n5163), .A(n4932), .B(n3776), .ZN(n3778)
         );
  OAI211_X1 U4354 ( .C1(n3780), .C2(n3815), .A(n3779), .B(n3778), .ZN(U3231)
         );
  NAND2_X1 U4355 ( .A1(n3782), .A2(n3781), .ZN(n3784) );
  AOI21_X1 U4356 ( .B1(n3785), .B2(n3784), .A(n3783), .ZN(n3790) );
  OAI22_X1 U4357 ( .A1(n3810), .A2(n4178), .B1(STATE_REG_SCAN_IN), .B2(n3786), 
        .ZN(n3788) );
  OAI22_X1 U4358 ( .A1(n5177), .A2(n4192), .B1(n3809), .B2(n4182), .ZN(n3787)
         );
  AOI211_X1 U4359 ( .C1(n4179), .C2(n5163), .A(n3788), .B(n3787), .ZN(n3789)
         );
  OAI21_X1 U4360 ( .B1(n3790), .B2(n3815), .A(n3789), .ZN(U3232) );
  NAND2_X1 U4361 ( .A1(n3793), .A2(n3792), .ZN(n3794) );
  XNOR2_X1 U4362 ( .A(n3791), .B(n3794), .ZN(n3801) );
  INV_X1 U4363 ( .A(n4241), .ZN(n3795) );
  AOI22_X1 U4364 ( .A1(n3796), .A2(n3795), .B1(n5161), .B2(n4230), .ZN(n3800)
         );
  INV_X1 U4365 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3797) );
  NOR2_X1 U4366 ( .A1(STATE_REG_SCAN_IN), .A2(n3797), .ZN(n4961) );
  NOR2_X1 U4367 ( .A1(n3810), .A2(n4268), .ZN(n3798) );
  AOI211_X1 U4368 ( .C1(n4240), .C2(n5163), .A(n4961), .B(n3798), .ZN(n3799)
         );
  OAI211_X1 U4369 ( .C1(n3801), .C2(n3815), .A(n3800), .B(n3799), .ZN(U3235)
         );
  NAND2_X1 U4370 ( .A1(n3803), .A2(n3802), .ZN(n3807) );
  NAND2_X1 U4371 ( .A1(n3805), .A2(n3804), .ZN(n3806) );
  XNOR2_X1 U4372 ( .A(n3807), .B(n3806), .ZN(n3816) );
  OAI22_X1 U4373 ( .A1(n3809), .A2(n4127), .B1(STATE_REG_SCAN_IN), .B2(n3808), 
        .ZN(n3812) );
  OAI22_X1 U4374 ( .A1(n5177), .A2(n4134), .B1(n3810), .B2(n4141), .ZN(n3811)
         );
  AOI211_X1 U4375 ( .C1(n3813), .C2(n5163), .A(n3812), .B(n3811), .ZN(n3814)
         );
  OAI21_X1 U4376 ( .B1(n3816), .B2(n3815), .A(n3814), .ZN(U3237) );
  OAI21_X1 U4377 ( .B1(n3833), .B2(n3832), .A(n3817), .ZN(n3834) );
  NOR3_X1 U4378 ( .A1(n3819), .A2(n3818), .A3(n3834), .ZN(n3962) );
  INV_X1 U4379 ( .A(n3962), .ZN(n3858) );
  INV_X1 U4380 ( .A(DATAI_30_), .ZN(n3820) );
  OR2_X1 U4381 ( .A1(n3828), .A2(n3820), .ZN(n5233) );
  OR2_X1 U4382 ( .A1(n3980), .A2(n5233), .ZN(n3830) );
  INV_X1 U4383 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U4384 ( .A1(n2843), .A2(REG1_REG_31__SCAN_IN), .ZN(n3824) );
  INV_X1 U4385 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3821) );
  OR2_X1 U4386 ( .A1(n3822), .A2(n3821), .ZN(n3823) );
  OAI211_X1 U4387 ( .C1(n3826), .C2(n3825), .A(n3824), .B(n3823), .ZN(n5231)
         );
  INV_X1 U4388 ( .A(DATAI_31_), .ZN(n3827) );
  OR2_X1 U4389 ( .A1(n3828), .A2(n3827), .ZN(n3861) );
  NAND2_X1 U4390 ( .A1(n5231), .A2(n3861), .ZN(n3829) );
  AND2_X1 U4391 ( .A1(n3830), .A2(n3829), .ZN(n3887) );
  INV_X1 U4392 ( .A(n3887), .ZN(n3831) );
  AOI21_X1 U4393 ( .B1(n3833), .B2(n3832), .A(n3831), .ZN(n3853) );
  OAI221_X1 U4394 ( .B1(n3852), .B2(n3834), .C1(n3851), .C2(n3834), .A(n3853), 
        .ZN(n3835) );
  INV_X1 U4395 ( .A(n3835), .ZN(n3967) );
  NAND2_X1 U4396 ( .A1(n4267), .A2(n5162), .ZN(n3838) );
  NAND2_X1 U4397 ( .A1(n3838), .A2(n3837), .ZN(n3917) );
  NOR2_X1 U4398 ( .A1(n3836), .A2(n3917), .ZN(n3840) );
  INV_X1 U4399 ( .A(n3838), .ZN(n3839) );
  OAI21_X1 U4400 ( .B1(n3839), .B2(n3946), .A(n3944), .ZN(n3950) );
  OAI21_X1 U4401 ( .B1(n3840), .B2(n3950), .A(n3902), .ZN(n3847) );
  AND4_X1 U4402 ( .A1(n3843), .A2(n2526), .A3(n3842), .A4(n3841), .ZN(n3954)
         );
  INV_X1 U4403 ( .A(n3844), .ZN(n3845) );
  NAND2_X1 U4404 ( .A1(n3846), .A2(n3845), .ZN(n3952) );
  AOI21_X1 U4405 ( .B1(n3847), .B2(n3954), .A(n3952), .ZN(n3848) );
  OAI211_X1 U4406 ( .C1(n3848), .C2(n3959), .A(n3957), .B(n3956), .ZN(n3855)
         );
  NAND2_X1 U4407 ( .A1(n3850), .A2(n3849), .ZN(n3963) );
  NAND3_X1 U4408 ( .A1(n3853), .A2(n3852), .A3(n3851), .ZN(n3854) );
  AOI211_X1 U4409 ( .C1(n3856), .C2(n3855), .A(n3963), .B(n3854), .ZN(n3857)
         );
  AOI21_X1 U4410 ( .B1(n3858), .B2(n3967), .A(n3857), .ZN(n3860) );
  NOR2_X1 U4411 ( .A1(n5231), .A2(n5233), .ZN(n3859) );
  OAI21_X1 U4412 ( .B1(n3860), .B2(n3859), .A(n4769), .ZN(n3864) );
  INV_X1 U4413 ( .A(n3861), .ZN(n5245) );
  OR2_X1 U4414 ( .A1(n5231), .A2(n3861), .ZN(n3863) );
  NAND2_X1 U4415 ( .A1(n3980), .A2(n5233), .ZN(n3862) );
  NAND2_X1 U4416 ( .A1(n3863), .A2(n3862), .ZN(n3966) );
  AOI22_X1 U4417 ( .A1(n3864), .A2(n3970), .B1(n5245), .B2(n3966), .ZN(n3972)
         );
  INV_X1 U4418 ( .A(n4157), .ZN(n3865) );
  AND2_X1 U4419 ( .A1(n3865), .A2(n4158), .ZN(n4204) );
  INV_X1 U4420 ( .A(n3966), .ZN(n3868) );
  NAND4_X1 U4421 ( .A1(n4204), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3871)
         );
  NAND4_X1 U4422 ( .A1(n4221), .A2(n4293), .A3(n5126), .A4(n3869), .ZN(n3870)
         );
  NOR2_X1 U4423 ( .A1(n3871), .A2(n3870), .ZN(n3883) );
  INV_X1 U4424 ( .A(n4123), .ZN(n4125) );
  AND2_X1 U4425 ( .A1(n2526), .A2(n3872), .ZN(n4251) );
  AND4_X1 U4426 ( .A1(n4125), .A2(n4251), .A3(n3873), .A4(n4266), .ZN(n3882)
         );
  NAND4_X1 U4427 ( .A1(n4186), .A2(n3874), .A3(n5032), .A4(n5007), .ZN(n3880)
         );
  NAND4_X1 U4428 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3879)
         );
  NOR2_X1 U4429 ( .A1(n3880), .A2(n3879), .ZN(n3881) );
  NAND4_X1 U4430 ( .A1(n3883), .A2(n3882), .A3(n5096), .A4(n3881), .ZN(n3901)
         );
  NAND2_X1 U4431 ( .A1(n3884), .A2(n3957), .ZN(n4142) );
  NOR2_X1 U4432 ( .A1(n4115), .A2(n4142), .ZN(n3894) );
  INV_X1 U4433 ( .A(n3885), .ZN(n4228) );
  NAND2_X1 U4434 ( .A1(n3887), .A2(n3886), .ZN(n3888) );
  NOR2_X1 U4435 ( .A1(n3889), .A2(n3888), .ZN(n3893) );
  NOR2_X1 U4436 ( .A1(n3891), .A2(n3890), .ZN(n3892) );
  NAND4_X1 U4437 ( .A1(n3894), .A2(n4228), .A3(n3893), .A4(n3892), .ZN(n3899)
         );
  INV_X1 U4438 ( .A(n4163), .ZN(n3897) );
  NAND3_X1 U4439 ( .A1(n3897), .A2(n3896), .A3(n3895), .ZN(n3898) );
  OR2_X1 U4440 ( .A1(n3899), .A2(n3898), .ZN(n3900) );
  NOR3_X1 U4441 ( .A1(n3901), .A2(n3900), .A3(n5209), .ZN(n3971) );
  INV_X1 U4442 ( .A(n3902), .ZN(n3955) );
  NOR4_X1 U4443 ( .A1(n2588), .A2(n3304), .A3(n3990), .A4(n3903), .ZN(n3907)
         );
  AND2_X1 U4444 ( .A1(n3905), .A2(n3904), .ZN(n3941) );
  INV_X1 U4445 ( .A(n5119), .ZN(n3906) );
  AOI22_X1 U4446 ( .A1(n3907), .A2(n3941), .B1(n3906), .B2(n5102), .ZN(n3911)
         );
  AND2_X1 U4447 ( .A1(n3909), .A2(n3908), .ZN(n3910) );
  NAND2_X1 U4448 ( .A1(n3913), .A2(n3910), .ZN(n3943) );
  NOR2_X1 U4449 ( .A1(n3911), .A2(n3943), .ZN(n3920) );
  INV_X1 U4450 ( .A(n3912), .ZN(n3919) );
  INV_X1 U4451 ( .A(n3913), .ZN(n3914) );
  AOI21_X1 U4452 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3918) );
  NOR4_X1 U4453 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3951)
         );
  OAI211_X1 U4454 ( .C1(n5006), .C2(n4769), .A(n3922), .B(n3921), .ZN(n3924)
         );
  NAND3_X1 U4455 ( .A1(n3924), .A2(n3923), .A3(n5036), .ZN(n3927) );
  NAND3_X1 U4456 ( .A1(n3927), .A2(n3926), .A3(n3925), .ZN(n3930) );
  NAND3_X1 U4457 ( .A1(n3930), .A2(n3929), .A3(n3928), .ZN(n3934) );
  NAND4_X1 U4458 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3937)
         );
  NAND3_X1 U4459 ( .A1(n3937), .A2(n3936), .A3(n3935), .ZN(n3942) );
  INV_X1 U4460 ( .A(n3938), .ZN(n3940) );
  AOI211_X1 U4461 ( .C1(n3942), .C2(n3941), .A(n3940), .B(n2646), .ZN(n3949)
         );
  INV_X1 U4462 ( .A(n3943), .ZN(n3947) );
  NAND4_X1 U4463 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3948)
         );
  OAI22_X1 U4464 ( .A1(n3951), .A2(n3950), .B1(n3949), .B2(n3948), .ZN(n3953)
         );
  AOI221_X1 U4465 ( .B1(n3955), .B2(n3954), .C1(n3953), .C2(n3954), .A(n3952), 
        .ZN(n3961) );
  AND2_X1 U4466 ( .A1(n3957), .A2(n3956), .ZN(n3960) );
  AOI221_X1 U4467 ( .B1(n3961), .B2(n3960), .C1(n3959), .C2(n3960), .A(n3958), 
        .ZN(n3964) );
  OAI21_X1 U4468 ( .B1(n3964), .B2(n3963), .A(n3962), .ZN(n3968) );
  INV_X1 U4469 ( .A(n5231), .ZN(n3965) );
  AOI22_X1 U4470 ( .A1(n3968), .A2(n3967), .B1(n3966), .B2(n3965), .ZN(n3969)
         );
  OAI22_X1 U4471 ( .A1(n3972), .A2(n3971), .B1(n3970), .B2(n3969), .ZN(n3973)
         );
  XNOR2_X1 U4472 ( .A(n3973), .B(n5219), .ZN(n3979) );
  OR2_X1 U4473 ( .A1(n3143), .A2(n3127), .ZN(n4970) );
  INV_X1 U4474 ( .A(n4970), .ZN(n3974) );
  NAND2_X1 U4475 ( .A1(n3975), .A2(n3974), .ZN(n3976) );
  OAI211_X1 U4476 ( .C1(n4768), .C2(n3978), .A(n3976), .B(B_REG_SCAN_IN), .ZN(
        n3977) );
  OAI21_X1 U4477 ( .B1(n3979), .B2(n3978), .A(n3977), .ZN(U3239) );
  MUX2_X1 U4478 ( .A(n5231), .B(DATAO_REG_31__SCAN_IN), .S(n3984), .Z(U3581)
         );
  MUX2_X1 U4479 ( .A(n3980), .B(DATAO_REG_30__SCAN_IN), .S(n3984), .Z(U3580)
         );
  MUX2_X1 U4480 ( .A(DATAO_REG_28__SCAN_IN), .B(n3981), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4481 ( .A(DATAO_REG_27__SCAN_IN), .B(n3982), .S(U4043), .Z(U3577)
         );
  INV_X1 U4482 ( .A(n4178), .ZN(n4215) );
  MUX2_X1 U4483 ( .A(DATAO_REG_21__SCAN_IN), .B(n4215), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4484 ( .A(DATAO_REG_19__SCAN_IN), .B(n4230), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4485 ( .A(DATAO_REG_18__SCAN_IN), .B(n3983), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4486 ( .A(n4231), .B(DATAO_REG_17__SCAN_IN), .S(n3984), .Z(U3567)
         );
  MUX2_X1 U4487 ( .A(DATAO_REG_16__SCAN_IN), .B(n5160), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4488 ( .A(n4287), .B(DATAO_REG_15__SCAN_IN), .S(n3984), .Z(U3565)
         );
  MUX2_X1 U4489 ( .A(n5158), .B(DATAO_REG_14__SCAN_IN), .S(n3984), .Z(U3564)
         );
  MUX2_X1 U4490 ( .A(DATAO_REG_13__SCAN_IN), .B(n4288), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4491 ( .A(DATAO_REG_12__SCAN_IN), .B(n5118), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4492 ( .A(DATAO_REG_11__SCAN_IN), .B(n3985), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4493 ( .A(DATAO_REG_10__SCAN_IN), .B(n5119), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4494 ( .A(DATAO_REG_9__SCAN_IN), .B(n3986), .S(U4043), .Z(U3559) );
  MUX2_X1 U4495 ( .A(DATAO_REG_8__SCAN_IN), .B(n3987), .S(U4043), .Z(U3558) );
  MUX2_X1 U4496 ( .A(DATAO_REG_7__SCAN_IN), .B(n3988), .S(U4043), .Z(U3557) );
  MUX2_X1 U4497 ( .A(DATAO_REG_6__SCAN_IN), .B(n3989), .S(U4043), .Z(U3556) );
  MUX2_X1 U4498 ( .A(DATAO_REG_5__SCAN_IN), .B(n3990), .S(U4043), .Z(U3555) );
  MUX2_X1 U4499 ( .A(DATAO_REG_4__SCAN_IN), .B(n3991), .S(U4043), .Z(U3554) );
  MUX2_X1 U4500 ( .A(DATAO_REG_3__SCAN_IN), .B(n5034), .S(U4043), .Z(U3553) );
  MUX2_X1 U4501 ( .A(DATAO_REG_2__SCAN_IN), .B(n5010), .S(U4043), .Z(U3552) );
  MUX2_X1 U4502 ( .A(DATAO_REG_1__SCAN_IN), .B(n3237), .S(U4043), .Z(U3551) );
  MUX2_X1 U4503 ( .A(DATAO_REG_0__SCAN_IN), .B(n3992), .S(U4043), .Z(U3550) );
  INV_X1 U4504 ( .A(n4772), .ZN(n4056) );
  NAND2_X1 U4505 ( .A1(n4773), .A2(REG1_REG_15__SCAN_IN), .ZN(n4019) );
  NOR2_X1 U4506 ( .A1(n4773), .A2(REG1_REG_15__SCAN_IN), .ZN(n3993) );
  AOI21_X1 U4507 ( .B1(REG1_REG_15__SCAN_IN), .B2(n4773), .A(n3993), .ZN(n4945) );
  INV_X1 U4508 ( .A(n4044), .ZN(n5143) );
  INV_X1 U4509 ( .A(n4775), .ZN(n4909) );
  NOR2_X1 U4510 ( .A1(n4909), .A2(n3994), .ZN(n3995) );
  AOI21_X1 U4511 ( .B1(n3994), .B2(n4909), .A(n3995), .ZN(n4902) );
  INV_X1 U4512 ( .A(n4025), .ZN(n5085) );
  MUX2_X1 U4513 ( .A(REG1_REG_9__SCAN_IN), .B(n3996), .S(n4025), .Z(n4881) );
  NAND2_X1 U4514 ( .A1(n4776), .A2(REG1_REG_7__SCAN_IN), .ZN(n4007) );
  MUX2_X1 U4515 ( .A(REG1_REG_7__SCAN_IN), .B(n5077), .S(n4776), .Z(n4859) );
  INV_X1 U4516 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5064) );
  MUX2_X1 U4517 ( .A(REG1_REG_5__SCAN_IN), .B(n5064), .S(n4027), .Z(n4838) );
  INV_X1 U4518 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3997) );
  MUX2_X1 U4519 ( .A(n3997), .B(REG1_REG_1__SCAN_IN), .S(n5003), .Z(n4818) );
  NAND3_X1 U4520 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .A3(n4818), .ZN(n4817) );
  OR2_X1 U4521 ( .A1(n5003), .A2(n3997), .ZN(n3998) );
  NAND2_X1 U4522 ( .A1(n4817), .A2(n3998), .ZN(n4978) );
  MUX2_X1 U4523 ( .A(REG1_REG_2__SCAN_IN), .B(n3999), .S(n4975), .Z(n4977) );
  NAND2_X1 U4524 ( .A1(n4028), .A2(n4000), .ZN(n4001) );
  NAND2_X1 U4525 ( .A1(n4989), .A2(n4002), .ZN(n4003) );
  INV_X1 U4526 ( .A(n4989), .ZN(n4033) );
  XNOR2_X1 U4527 ( .A(n4002), .B(n4033), .ZN(n4993) );
  NAND2_X1 U4528 ( .A1(REG1_REG_4__SCAN_IN), .A2(n4993), .ZN(n4991) );
  NAND2_X1 U4529 ( .A1(n4003), .A2(n4991), .ZN(n4839) );
  NAND2_X1 U4530 ( .A1(n4838), .A2(n4839), .ZN(n4837) );
  NAND2_X1 U4531 ( .A1(n4851), .A2(n4005), .ZN(n4006) );
  NAND2_X1 U4532 ( .A1(n4006), .A2(n4852), .ZN(n4860) );
  NAND2_X1 U4533 ( .A1(n4859), .A2(n4860), .ZN(n4858) );
  NAND2_X1 U4534 ( .A1(n4873), .A2(n4008), .ZN(n4009) );
  INV_X1 U4535 ( .A(n4873), .ZN(n4039) );
  XNOR2_X1 U4536 ( .A(n4008), .B(n4039), .ZN(n4872) );
  NAND2_X1 U4537 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U4538 ( .A1(n4009), .A2(n4871), .ZN(n4882) );
  NAND2_X1 U4539 ( .A1(n4881), .A2(n4882), .ZN(n4880) );
  NAND2_X1 U4540 ( .A1(n4891), .A2(n4010), .ZN(n4011) );
  NAND2_X1 U4541 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U4542 ( .A1(n4044), .A2(n4012), .ZN(n4013) );
  NAND2_X1 U4543 ( .A1(n4937), .A2(n4017), .ZN(n4018) );
  INV_X1 U4544 ( .A(n4937), .ZN(n4016) );
  NOR2_X1 U4545 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4020), .ZN(n4065) );
  AOI21_X1 U4546 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4020), .A(n4065), .ZN(n4060) );
  NAND2_X1 U4547 ( .A1(n4022), .A2(n4021), .ZN(n4815) );
  INV_X1 U4548 ( .A(n4815), .ZN(n4053) );
  NAND2_X1 U4549 ( .A1(n4053), .A2(n3143), .ZN(n4816) );
  NAND2_X1 U4550 ( .A1(n4773), .A2(REG2_REG_15__SCAN_IN), .ZN(n4050) );
  INV_X1 U4551 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4024) );
  INV_X1 U4552 ( .A(n4773), .ZN(n4948) );
  INV_X1 U4553 ( .A(n4050), .ZN(n4023) );
  AOI21_X1 U4554 ( .B1(n4024), .B2(n4948), .A(n4023), .ZN(n4952) );
  INV_X1 U4555 ( .A(REG2_REG_11__SCAN_IN), .ZN(n5139) );
  AOI22_X1 U4556 ( .A1(n4775), .A2(REG2_REG_11__SCAN_IN), .B1(n5139), .B2(
        n4909), .ZN(n4905) );
  AOI22_X1 U4557 ( .A1(n4025), .A2(REG2_REG_9__SCAN_IN), .B1(n3388), .B2(n5085), .ZN(n4884) );
  NAND2_X1 U4558 ( .A1(n4776), .A2(REG2_REG_7__SCAN_IN), .ZN(n4037) );
  INV_X1 U4559 ( .A(n4776), .ZN(n4866) );
  AOI22_X1 U4560 ( .A1(n4776), .A2(REG2_REG_7__SCAN_IN), .B1(n4026), .B2(n4866), .ZN(n4862) );
  AOI22_X1 U4561 ( .A1(n4027), .A2(REG2_REG_5__SCAN_IN), .B1(n3359), .B2(n5059), .ZN(n4841) );
  INV_X1 U4562 ( .A(REG2_REG_2__SCAN_IN), .ZN(n5049) );
  AOI22_X1 U4563 ( .A1(n4975), .A2(REG2_REG_2__SCAN_IN), .B1(n5049), .B2(n5027), .ZN(n4981) );
  INV_X1 U4564 ( .A(REG2_REG_1__SCAN_IN), .ZN(n5024) );
  NAND3_X1 U4565 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .A3(n4822), .ZN(n4821) );
  OAI21_X1 U4566 ( .B1(n5024), .B2(n5003), .A(n4821), .ZN(n4980) );
  NAND2_X1 U4567 ( .A1(n4981), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U4568 ( .A1(n4028), .A2(n4030), .ZN(n4031) );
  NAND2_X1 U4569 ( .A1(n4989), .A2(n4032), .ZN(n4034) );
  NAND2_X1 U4570 ( .A1(REG2_REG_4__SCAN_IN), .A2(n4996), .ZN(n4994) );
  NAND2_X1 U4571 ( .A1(n4851), .A2(n4035), .ZN(n4036) );
  NAND2_X1 U4572 ( .A1(n4873), .A2(n4038), .ZN(n4040) );
  NAND2_X1 U4573 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4875), .ZN(n4874) );
  NAND2_X1 U4574 ( .A1(n4040), .A2(n4874), .ZN(n4885) );
  NAND2_X1 U4575 ( .A1(n4884), .A2(n4885), .ZN(n4883) );
  NAND2_X1 U4576 ( .A1(n4891), .A2(n4042), .ZN(n4043) );
  NAND2_X1 U4577 ( .A1(n4044), .A2(n4045), .ZN(n4046) );
  NAND2_X1 U4578 ( .A1(n4930), .A2(REG2_REG_13__SCAN_IN), .ZN(n4047) );
  OAI21_X1 U4579 ( .B1(n4930), .B2(REG2_REG_13__SCAN_IN), .A(n4047), .ZN(n4926) );
  NAND2_X1 U4580 ( .A1(n4937), .A2(n4048), .ZN(n4049) );
  NAND2_X1 U4581 ( .A1(REG2_REG_14__SCAN_IN), .A2(n4939), .ZN(n4938) );
  NOR2_X1 U4582 ( .A1(REG2_REG_16__SCAN_IN), .A2(n4051), .ZN(n4073) );
  AOI21_X1 U4583 ( .B1(REG2_REG_16__SCAN_IN), .B2(n4051), .A(n4073), .ZN(n4052) );
  INV_X1 U4584 ( .A(n4052), .ZN(n4058) );
  NOR2_X2 U4585 ( .A1(n4815), .A2(n4970), .ZN(n4995) );
  NAND2_X1 U4586 ( .A1(n4053), .A2(n3127), .ZN(n4958) );
  AOI21_X1 U4587 ( .B1(n4988), .B2(ADDR_REG_16__SCAN_IN), .A(n4054), .ZN(n4055) );
  OAI21_X1 U4588 ( .B1(n4958), .B2(n4056), .A(n4055), .ZN(n4057) );
  AOI21_X1 U4589 ( .B1(n4058), .B2(n4995), .A(n4057), .ZN(n4059) );
  OAI21_X1 U4590 ( .B1(n4060), .B2(n4816), .A(n4059), .ZN(U3256) );
  OR2_X1 U4591 ( .A1(n4771), .A2(n4061), .ZN(n4063) );
  NAND2_X1 U4592 ( .A1(n4771), .A2(n4061), .ZN(n4062) );
  AND2_X1 U4593 ( .A1(n4063), .A2(n4062), .ZN(n4069) );
  NOR2_X1 U4594 ( .A1(n4772), .A2(n4064), .ZN(n4066) );
  INV_X1 U4595 ( .A(n4082), .ZN(n4067) );
  AOI21_X1 U4596 ( .B1(n4069), .B2(n4068), .A(n4067), .ZN(n4081) );
  INV_X1 U4597 ( .A(n4771), .ZN(n4087) );
  NOR2_X1 U4598 ( .A1(n4958), .A2(n4087), .ZN(n4070) );
  AOI211_X1 U4599 ( .C1(n4988), .C2(ADDR_REG_17__SCAN_IN), .A(n4071), .B(n4070), .ZN(n4080) );
  NOR2_X1 U4600 ( .A1(n4772), .A2(n4072), .ZN(n4074) );
  INV_X1 U4601 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4258) );
  OR2_X1 U4602 ( .A1(n4771), .A2(n4258), .ZN(n4075) );
  OAI21_X1 U4603 ( .B1(n4087), .B2(REG2_REG_17__SCAN_IN), .A(n4075), .ZN(n4077) );
  NAND2_X1 U4604 ( .A1(n4771), .A2(REG2_REG_17__SCAN_IN), .ZN(n4076) );
  OAI211_X1 U4605 ( .C1(n4771), .C2(REG2_REG_17__SCAN_IN), .A(n4078), .B(n4076), .ZN(n4086) );
  OAI211_X1 U4606 ( .C1(n4078), .C2(n4077), .A(n4086), .B(n4995), .ZN(n4079)
         );
  OAI211_X1 U4607 ( .C1(n4081), .C2(n4816), .A(n4080), .B(n4079), .ZN(U3257)
         );
  NOR2_X1 U4608 ( .A1(n4770), .A2(REG1_REG_18__SCAN_IN), .ZN(n4083) );
  OAI21_X1 U4609 ( .B1(n4771), .B2(REG1_REG_17__SCAN_IN), .A(n4082), .ZN(n4956) );
  AOI21_X1 U4610 ( .B1(n4770), .B2(REG1_REG_18__SCAN_IN), .A(n4960), .ZN(n4085) );
  MUX2_X1 U4611 ( .A(REG1_REG_19__SCAN_IN), .B(n3054), .S(n5219), .Z(n4084) );
  XNOR2_X1 U4612 ( .A(n4085), .B(n4084), .ZN(n4098) );
  INV_X1 U4613 ( .A(n4770), .ZN(n4959) );
  OAI21_X1 U4614 ( .B1(n4258), .B2(n4087), .A(n4086), .ZN(n4963) );
  NOR2_X1 U4615 ( .A1(n4959), .A2(n4088), .ZN(n4089) );
  AOI21_X1 U4616 ( .B1(n4959), .B2(n4088), .A(n4089), .ZN(n4964) );
  NAND2_X1 U4617 ( .A1(n4963), .A2(n4964), .ZN(n4962) );
  OAI21_X1 U4618 ( .B1(n4959), .B2(n4088), .A(n4962), .ZN(n4092) );
  INV_X1 U4619 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4090) );
  MUX2_X1 U4620 ( .A(REG2_REG_19__SCAN_IN), .B(n4090), .S(n5219), .Z(n4091) );
  XNOR2_X1 U4621 ( .A(n4092), .B(n4091), .ZN(n4096) );
  NAND2_X1 U4622 ( .A1(n4988), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4093) );
  OAI211_X1 U4623 ( .C1(n4958), .C2(n5219), .A(n4094), .B(n4093), .ZN(n4095)
         );
  AOI21_X1 U4624 ( .B1(n4096), .B2(n4995), .A(n4095), .ZN(n4097) );
  OAI21_X1 U4625 ( .B1(n4098), .B2(n4816), .A(n4097), .ZN(U3259) );
  AOI21_X1 U4626 ( .B1(n4131), .B2(n4108), .A(n5204), .ZN(n4100) );
  NAND2_X1 U4627 ( .A1(n4100), .A2(n4099), .ZN(n4315) );
  INV_X1 U4628 ( .A(n4111), .ZN(n4103) );
  INV_X1 U4629 ( .A(n4101), .ZN(n4102) );
  OAI22_X1 U4630 ( .A1(n4103), .A2(n5144), .B1(n5217), .B2(n4102), .ZN(n4114)
         );
  INV_X1 U4631 ( .A(n4104), .ZN(n4110) );
  OAI22_X1 U4632 ( .A1(n4106), .A2(n5210), .B1(n4105), .B2(n5212), .ZN(n4107)
         );
  AOI21_X1 U4633 ( .B1(n4108), .B2(n5240), .A(n4107), .ZN(n4109) );
  OAI21_X1 U4634 ( .B1(n4110), .B2(n5217), .A(n4109), .ZN(n4113) );
  NOR3_X1 U4635 ( .A1(n4111), .A2(n5144), .A3(n4115), .ZN(n4112) );
  AOI211_X1 U4636 ( .C1(n4115), .C2(n4114), .A(n4113), .B(n4112), .ZN(n4316)
         );
  OR2_X1 U4637 ( .A1(n4316), .A2(n5249), .ZN(n4119) );
  INV_X1 U4638 ( .A(n4116), .ZN(n4117) );
  AOI22_X1 U4639 ( .A1(n5249), .A2(REG2_REG_27__SCAN_IN), .B1(n4117), .B2(
        n5135), .ZN(n4118) );
  OAI211_X1 U4640 ( .C1(n4315), .C2(n4278), .A(n4119), .B(n4118), .ZN(U3263)
         );
  NAND2_X1 U4641 ( .A1(n4140), .A2(n4120), .ZN(n4122) );
  NAND2_X1 U4642 ( .A1(n4122), .A2(n4121), .ZN(n4124) );
  XNOR2_X1 U4643 ( .A(n4124), .B(n4123), .ZN(n4319) );
  XNOR2_X1 U4644 ( .A(n4126), .B(n4125), .ZN(n4130) );
  NOR2_X1 U4645 ( .A1(n5123), .A2(n4132), .ZN(n4129) );
  OAI22_X1 U4646 ( .A1(n4141), .A2(n5212), .B1(n4127), .B2(n5210), .ZN(n4128)
         );
  AOI211_X1 U4647 ( .C1(n4130), .C2(n5008), .A(n4129), .B(n4128), .ZN(n4318)
         );
  INV_X1 U4648 ( .A(n4318), .ZN(n4138) );
  OAI211_X1 U4649 ( .C1(n4133), .C2(n4132), .A(n5252), .B(n4131), .ZN(n4317)
         );
  INV_X1 U4650 ( .A(n4134), .ZN(n4135) );
  AOI22_X1 U4651 ( .A1(n5249), .A2(REG2_REG_26__SCAN_IN), .B1(n4135), .B2(
        n5135), .ZN(n4136) );
  OAI21_X1 U4652 ( .B1(n4317), .B2(n4278), .A(n4136), .ZN(n4137) );
  AOI21_X1 U4653 ( .B1(n4138), .B2(n4242), .A(n4137), .ZN(n4139) );
  OAI21_X1 U4654 ( .B1(n4319), .B2(n4282), .A(n4139), .ZN(U3264) );
  XNOR2_X1 U4655 ( .A(n4140), .B(n4142), .ZN(n4325) );
  OAI22_X1 U4656 ( .A1(n4141), .A2(n5210), .B1(n4182), .B2(n5212), .ZN(n4146)
         );
  XNOR2_X1 U4657 ( .A(n4143), .B(n4142), .ZN(n4144) );
  NOR2_X1 U4658 ( .A1(n4144), .A2(n5217), .ZN(n4145) );
  AOI211_X1 U4659 ( .C1(n5240), .C2(n4147), .A(n4146), .B(n4145), .ZN(n4324)
         );
  INV_X1 U4660 ( .A(n4324), .ZN(n4154) );
  OAI211_X1 U4661 ( .C1(n2501), .C2(n4149), .A(n2620), .B(n5252), .ZN(n4323)
         );
  INV_X1 U4662 ( .A(n4150), .ZN(n4151) );
  AOI22_X1 U4663 ( .A1(n5249), .A2(REG2_REG_24__SCAN_IN), .B1(n4151), .B2(
        n5135), .ZN(n4152) );
  OAI21_X1 U4664 ( .B1(n4323), .B2(n4278), .A(n4152), .ZN(n4153) );
  AOI21_X1 U4665 ( .B1(n4154), .B2(n5140), .A(n4153), .ZN(n4155) );
  OAI21_X1 U4666 ( .B1(n4325), .B2(n4282), .A(n4155), .ZN(U3266) );
  AOI211_X1 U4667 ( .C1(n4166), .C2(n4190), .A(n5204), .B(n2501), .ZN(n4326)
         );
  INV_X1 U4668 ( .A(n4326), .ZN(n4174) );
  NAND2_X1 U4669 ( .A1(n4159), .A2(n4158), .ZN(n4175) );
  NOR2_X1 U4670 ( .A1(n4177), .A2(n4160), .ZN(n4161) );
  XOR2_X1 U4671 ( .A(n4163), .B(n4161), .Z(n4169) );
  OAI211_X1 U4672 ( .C1(n3564), .C2(n4163), .A(n4162), .B(n5227), .ZN(n4168)
         );
  OAI22_X1 U4673 ( .A1(n4205), .A2(n5212), .B1(n4164), .B2(n5210), .ZN(n4165)
         );
  AOI21_X1 U4674 ( .B1(n4166), .B2(n5240), .A(n4165), .ZN(n4167) );
  OAI211_X1 U4675 ( .C1(n5217), .C2(n4169), .A(n4168), .B(n4167), .ZN(n4327)
         );
  NAND2_X1 U4676 ( .A1(n4327), .A2(n4242), .ZN(n4173) );
  INV_X1 U4677 ( .A(n4170), .ZN(n4171) );
  AOI22_X1 U4678 ( .A1(n5249), .A2(REG2_REG_23__SCAN_IN), .B1(n4171), .B2(
        n5135), .ZN(n4172) );
  OAI211_X1 U4679 ( .C1(n4174), .C2(n4278), .A(n4173), .B(n4172), .ZN(U3267)
         );
  AND2_X1 U4680 ( .A1(n4175), .A2(n2682), .ZN(n4176) );
  OAI21_X1 U4681 ( .B1(n4177), .B2(n4176), .A(n5008), .ZN(n4185) );
  OR2_X1 U4682 ( .A1(n4178), .A2(n5212), .ZN(n4181) );
  NAND2_X1 U4683 ( .A1(n5240), .A2(n4179), .ZN(n4180) );
  OAI211_X1 U4684 ( .C1(n4182), .C2(n5210), .A(n4181), .B(n4180), .ZN(n4183)
         );
  INV_X1 U4685 ( .A(n4183), .ZN(n4184) );
  NAND2_X1 U4686 ( .A1(n4187), .A2(n4186), .ZN(n4188) );
  AND2_X1 U4687 ( .A1(n4189), .A2(n4188), .ZN(n4331) );
  NAND2_X1 U4688 ( .A1(n4331), .A2(n5201), .ZN(n4197) );
  OAI211_X1 U4689 ( .C1(n4200), .C2(n4191), .A(n5252), .B(n4190), .ZN(n4328)
         );
  INV_X1 U4690 ( .A(n4328), .ZN(n4195) );
  INV_X1 U4691 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4193) );
  OAI22_X1 U4692 ( .A1(n5140), .A2(n4193), .B1(n4192), .B2(n5224), .ZN(n4194)
         );
  AOI21_X1 U4693 ( .B1(n4195), .B2(n4260), .A(n4194), .ZN(n4196) );
  OAI211_X1 U4694 ( .C1(n5249), .C2(n4329), .A(n4197), .B(n4196), .ZN(U3268)
         );
  XOR2_X1 U4695 ( .A(n4204), .B(n4198), .Z(n4337) );
  INV_X1 U4696 ( .A(n4199), .ZN(n4339) );
  AOI21_X1 U4697 ( .B1(n4207), .B2(n4339), .A(n4200), .ZN(n4335) );
  INV_X1 U4698 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4202) );
  OAI22_X1 U4699 ( .A1(n5140), .A2(n4202), .B1(n4201), .B2(n5224), .ZN(n4203)
         );
  AOI21_X1 U4700 ( .B1(n4335), .B2(n5247), .A(n4203), .ZN(n4211) );
  XOR2_X1 U4701 ( .A(n4204), .B(n4156), .Z(n4209) );
  OAI22_X1 U4702 ( .A1(n4205), .A2(n5210), .B1(n5211), .B2(n5212), .ZN(n4206)
         );
  AOI21_X1 U4703 ( .B1(n4207), .B2(n5240), .A(n4206), .ZN(n4208) );
  OAI21_X1 U4704 ( .B1(n4209), .B2(n5217), .A(n4208), .ZN(n4334) );
  NAND2_X1 U4705 ( .A1(n4334), .A2(n4242), .ZN(n4210) );
  OAI211_X1 U4706 ( .C1(n4337), .C2(n4282), .A(n4211), .B(n4210), .ZN(U3269)
         );
  INV_X1 U4707 ( .A(n4213), .ZN(n4214) );
  OAI22_X1 U4708 ( .A1(n4212), .A2(n5144), .B1(n5217), .B2(n4214), .ZN(n4220)
         );
  AOI22_X1 U4709 ( .A1(n4212), .A2(n5227), .B1(n4214), .B2(n5008), .ZN(n4218)
         );
  AOI22_X1 U4710 ( .A1(n4215), .A2(n5117), .B1(n5120), .B2(n4230), .ZN(n4217)
         );
  NAND2_X1 U4711 ( .A1(n5240), .A2(n4224), .ZN(n4216) );
  OAI211_X1 U4712 ( .C1(n4218), .C2(n4221), .A(n4217), .B(n4216), .ZN(n4219)
         );
  AOI21_X1 U4713 ( .B1(n4221), .B2(n4220), .A(n4219), .ZN(n4341) );
  INV_X1 U4714 ( .A(n4222), .ZN(n4223) );
  AOI22_X1 U4715 ( .A1(n5249), .A2(REG2_REG_20__SCAN_IN), .B1(n4223), .B2(
        n5135), .ZN(n4226) );
  NAND2_X1 U4716 ( .A1(n5202), .A2(n4224), .ZN(n4338) );
  NAND3_X1 U4717 ( .A1(n4339), .A2(n5247), .A3(n4338), .ZN(n4225) );
  OAI211_X1 U4718 ( .C1(n4341), .C2(n5249), .A(n4226), .B(n4225), .ZN(U3270)
         );
  XNOR2_X1 U4719 ( .A(n4227), .B(n4228), .ZN(n4237) );
  XNOR2_X1 U4720 ( .A(n4229), .B(n4228), .ZN(n4235) );
  AOI22_X1 U4721 ( .A1(n4231), .A2(n5120), .B1(n5117), .B2(n4230), .ZN(n4232)
         );
  OAI21_X1 U4722 ( .B1(n4233), .B2(n5123), .A(n4232), .ZN(n4234) );
  AOI21_X1 U4723 ( .B1(n4235), .B2(n5008), .A(n4234), .ZN(n4236) );
  OAI21_X1 U4724 ( .B1(n4237), .B2(n5144), .A(n4236), .ZN(n5196) );
  INV_X1 U4725 ( .A(n5196), .ZN(n4245) );
  INV_X1 U4726 ( .A(n4256), .ZN(n4239) );
  INV_X1 U4727 ( .A(n5205), .ZN(n4238) );
  AOI211_X1 U4728 ( .C1(n4240), .C2(n4239), .A(n5204), .B(n4238), .ZN(n5197)
         );
  OAI22_X1 U4729 ( .A1(n4242), .A2(n4088), .B1(n4241), .B2(n5224), .ZN(n4243)
         );
  AOI21_X1 U4730 ( .B1(n5197), .B2(n4260), .A(n4243), .ZN(n4244) );
  OAI21_X1 U4731 ( .B1(n4245), .B2(n5249), .A(n4244), .ZN(U3272) );
  XNOR2_X1 U4732 ( .A(n4246), .B(n4251), .ZN(n4250) );
  OAI22_X1 U4733 ( .A1(n4247), .A2(n5212), .B1(n5213), .B2(n5210), .ZN(n4248)
         );
  AOI21_X1 U4734 ( .B1(n4253), .B2(n5240), .A(n4248), .ZN(n4249) );
  OAI21_X1 U4735 ( .B1(n4250), .B2(n5217), .A(n4249), .ZN(n5191) );
  INV_X1 U4736 ( .A(n5191), .ZN(n4263) );
  XNOR2_X1 U4737 ( .A(n4252), .B(n4251), .ZN(n5193) );
  NAND2_X1 U4738 ( .A1(n5193), .A2(n5201), .ZN(n4262) );
  NAND2_X1 U4739 ( .A1(n4275), .A2(n4253), .ZN(n4254) );
  NAND2_X1 U4740 ( .A1(n4254), .A2(n5252), .ZN(n4255) );
  NOR2_X1 U4741 ( .A1(n4256), .A2(n4255), .ZN(n5192) );
  OAI22_X1 U4742 ( .A1(n5140), .A2(n4258), .B1(n4257), .B2(n5224), .ZN(n4259)
         );
  AOI21_X1 U4743 ( .B1(n5192), .B2(n4260), .A(n4259), .ZN(n4261) );
  OAI211_X1 U4744 ( .C1(n5249), .C2(n4263), .A(n4262), .B(n4261), .ZN(U3273)
         );
  XNOR2_X1 U4745 ( .A(n4264), .B(n4266), .ZN(n5187) );
  INV_X1 U4746 ( .A(n5187), .ZN(n4283) );
  XNOR2_X1 U4747 ( .A(n4265), .B(n4266), .ZN(n4271) );
  OAI22_X1 U4748 ( .A1(n4268), .A2(n5210), .B1(n4267), .B2(n5212), .ZN(n4269)
         );
  AOI21_X1 U4749 ( .B1(n4272), .B2(n5240), .A(n4269), .ZN(n4270) );
  OAI21_X1 U4750 ( .B1(n4271), .B2(n5217), .A(n4270), .ZN(n5185) );
  AOI21_X1 U4751 ( .B1(n4273), .B2(n4272), .A(n5204), .ZN(n4274) );
  AND2_X1 U4752 ( .A1(n4275), .A2(n4274), .ZN(n5186) );
  INV_X1 U4753 ( .A(n5186), .ZN(n4279) );
  AOI22_X1 U4754 ( .A1(n5249), .A2(REG2_REG_16__SCAN_IN), .B1(n4276), .B2(
        n5135), .ZN(n4277) );
  OAI21_X1 U4755 ( .B1(n4279), .B2(n4278), .A(n4277), .ZN(n4280) );
  AOI21_X1 U4756 ( .B1(n5185), .B2(n5140), .A(n4280), .ZN(n4281) );
  OAI21_X1 U4757 ( .B1(n4283), .B2(n4282), .A(n4281), .ZN(U3274) );
  OAI21_X1 U4758 ( .B1(n4285), .B2(n4290), .A(n4284), .ZN(n4760) );
  OAI21_X1 U4759 ( .B1(n4293), .B2(n3836), .A(n4286), .ZN(n4297) );
  AOI22_X1 U4760 ( .A1(n4288), .A2(n5120), .B1(n5117), .B2(n4287), .ZN(n4289)
         );
  OAI21_X1 U4761 ( .B1(n4290), .B2(n5123), .A(n4289), .ZN(n4296) );
  NAND2_X1 U4762 ( .A1(n4292), .A2(n4293), .ZN(n4294) );
  AOI21_X1 U4763 ( .B1(n4291), .B2(n4294), .A(n5144), .ZN(n4295) );
  AOI211_X1 U4764 ( .C1(n5008), .C2(n4297), .A(n4296), .B(n4295), .ZN(n4759)
         );
  OAI21_X1 U4765 ( .B1(n4298), .B2(n5224), .A(n4759), .ZN(n4301) );
  NOR2_X1 U4766 ( .A1(n5140), .A2(n4299), .ZN(n4300) );
  AOI21_X1 U4767 ( .B1(n4301), .B2(n5140), .A(n4300), .ZN(n4302) );
  OAI21_X1 U4768 ( .B1(n4760), .B2(n4303), .A(n4302), .ZN(U3276) );
  INV_X1 U4769 ( .A(n4307), .ZN(n4309) );
  NAND2_X1 U4770 ( .A1(n4309), .A2(n4308), .ZN(n4310) );
  INV_X2 U4771 ( .A(n5254), .ZN(n5256) );
  MUX2_X1 U4772 ( .A(REG1_REG_29__SCAN_IN), .B(n4345), .S(n5256), .Z(U3547) );
  NAND2_X1 U4773 ( .A1(n4314), .A2(n4313), .ZN(n4346) );
  MUX2_X1 U4774 ( .A(REG1_REG_28__SCAN_IN), .B(n4346), .S(n5256), .Z(U3546) );
  NAND2_X1 U4775 ( .A1(n4316), .A2(n4315), .ZN(n4347) );
  MUX2_X1 U4776 ( .A(REG1_REG_27__SCAN_IN), .B(n4347), .S(n5256), .Z(U3545) );
  OAI211_X1 U4777 ( .C1(n4319), .C2(n5144), .A(n4318), .B(n4317), .ZN(n4348)
         );
  MUX2_X1 U4778 ( .A(REG1_REG_26__SCAN_IN), .B(n4348), .S(n5256), .Z(U3544) );
  OAI211_X1 U4779 ( .C1(n4322), .C2(n5144), .A(n4321), .B(n4320), .ZN(n4349)
         );
  MUX2_X1 U4780 ( .A(REG1_REG_25__SCAN_IN), .B(n4349), .S(n5256), .Z(U3543) );
  OAI211_X1 U4781 ( .C1(n4325), .C2(n5144), .A(n4324), .B(n4323), .ZN(n4350)
         );
  MUX2_X1 U4782 ( .A(REG1_REG_24__SCAN_IN), .B(n4350), .S(n5256), .Z(U3542) );
  OR2_X1 U4783 ( .A1(n4327), .A2(n4326), .ZN(n4351) );
  MUX2_X1 U4784 ( .A(n4351), .B(REG1_REG_23__SCAN_IN), .S(n5254), .Z(U3541) );
  NAND2_X1 U4785 ( .A1(n4329), .A2(n4328), .ZN(n4330) );
  AOI21_X1 U4786 ( .B1(n4331), .B2(n5227), .A(n4330), .ZN(n4352) );
  MUX2_X1 U4787 ( .A(n4332), .B(n4352), .S(n5256), .Z(n4333) );
  INV_X1 U4788 ( .A(n4333), .ZN(U3540) );
  AOI21_X1 U4789 ( .B1(n5252), .B2(n4335), .A(n4334), .ZN(n4336) );
  OAI21_X1 U4790 ( .B1(n4337), .B2(n5144), .A(n4336), .ZN(n4355) );
  MUX2_X1 U4791 ( .A(REG1_REG_21__SCAN_IN), .B(n4355), .S(n5256), .Z(U3539) );
  NAND3_X1 U4792 ( .A1(n4339), .A2(n4338), .A3(n5252), .ZN(n4340) );
  NAND2_X1 U4793 ( .A1(n4341), .A2(n4340), .ZN(n4356) );
  MUX2_X1 U4794 ( .A(REG1_REG_20__SCAN_IN), .B(n4356), .S(n5256), .Z(U3538) );
  INV_X1 U4795 ( .A(n4342), .ZN(n4343) );
  MUX2_X1 U4796 ( .A(REG0_REG_29__SCAN_IN), .B(n4345), .S(n5259), .Z(U3515) );
  MUX2_X1 U4797 ( .A(REG0_REG_28__SCAN_IN), .B(n4346), .S(n5259), .Z(U3514) );
  MUX2_X1 U4798 ( .A(REG0_REG_27__SCAN_IN), .B(n4347), .S(n5259), .Z(U3513) );
  MUX2_X1 U4799 ( .A(REG0_REG_26__SCAN_IN), .B(n4348), .S(n5259), .Z(U3512) );
  MUX2_X1 U4800 ( .A(REG0_REG_25__SCAN_IN), .B(n4349), .S(n5259), .Z(U3511) );
  MUX2_X1 U4801 ( .A(REG0_REG_24__SCAN_IN), .B(n4350), .S(n5259), .Z(U3510) );
  MUX2_X1 U4802 ( .A(n4351), .B(REG0_REG_23__SCAN_IN), .S(n5257), .Z(U3509) );
  MUX2_X1 U4803 ( .A(n4353), .B(n4352), .S(n5259), .Z(n4354) );
  INV_X1 U4804 ( .A(n4354), .ZN(U3508) );
  MUX2_X1 U4805 ( .A(REG0_REG_21__SCAN_IN), .B(n4355), .S(n5259), .Z(U3507) );
  MUX2_X1 U4806 ( .A(REG0_REG_20__SCAN_IN), .B(n4356), .S(n5259), .Z(U3506) );
  XOR2_X1 U4807 ( .A(DATAI_28_), .B(keyinput_3), .Z(n4360) );
  XOR2_X1 U4808 ( .A(DATAI_27_), .B(keyinput_4), .Z(n4359) );
  XOR2_X1 U4809 ( .A(DATAI_26_), .B(keyinput_5), .Z(n4358) );
  XOR2_X1 U4810 ( .A(DATAI_30_), .B(keyinput_1), .Z(n4357) );
  NAND4_X1 U4811 ( .A1(n4360), .A2(n4359), .A3(n4358), .A4(n4357), .ZN(n4364)
         );
  XNOR2_X1 U4812 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n4363) );
  XNOR2_X1 U4813 ( .A(DATAI_31_), .B(keyinput_0), .ZN(n4362) );
  XNOR2_X1 U4814 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n4361) );
  NOR4_X1 U4815 ( .A1(n4364), .A2(n4363), .A3(n4362), .A4(n4361), .ZN(n4367)
         );
  XOR2_X1 U4816 ( .A(DATAI_24_), .B(keyinput_7), .Z(n4366) );
  XNOR2_X1 U4817 ( .A(DATAI_23_), .B(keyinput_8), .ZN(n4365) );
  NOR3_X1 U4818 ( .A1(n4367), .A2(n4366), .A3(n4365), .ZN(n4370) );
  XNOR2_X1 U4819 ( .A(DATAI_22_), .B(keyinput_9), .ZN(n4369) );
  XNOR2_X1 U4820 ( .A(DATAI_21_), .B(keyinput_10), .ZN(n4368) );
  NOR3_X1 U4821 ( .A1(n4370), .A2(n4369), .A3(n4368), .ZN(n4373) );
  XNOR2_X1 U4822 ( .A(DATAI_20_), .B(keyinput_11), .ZN(n4372) );
  XOR2_X1 U4823 ( .A(DATAI_19_), .B(keyinput_12), .Z(n4371) );
  OAI21_X1 U4824 ( .B1(n4373), .B2(n4372), .A(n4371), .ZN(n4376) );
  XOR2_X1 U4825 ( .A(DATAI_18_), .B(keyinput_13), .Z(n4375) );
  XOR2_X1 U4826 ( .A(DATAI_17_), .B(keyinput_14), .Z(n4374) );
  AOI21_X1 U4827 ( .B1(n4376), .B2(n4375), .A(n4374), .ZN(n4379) );
  XOR2_X1 U4828 ( .A(DATAI_15_), .B(keyinput_16), .Z(n4378) );
  XNOR2_X1 U4829 ( .A(DATAI_16_), .B(keyinput_15), .ZN(n4377) );
  NOR3_X1 U4830 ( .A1(n4379), .A2(n4378), .A3(n4377), .ZN(n4390) );
  XOR2_X1 U4831 ( .A(DATAI_14_), .B(keyinput_17), .Z(n4389) );
  XNOR2_X1 U4832 ( .A(n4380), .B(keyinput_18), .ZN(n4384) );
  XNOR2_X1 U4833 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n4383) );
  XNOR2_X1 U4834 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n4382) );
  XNOR2_X1 U4835 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n4381) );
  NAND4_X1 U4836 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), .ZN(n4387)
         );
  XNOR2_X1 U4837 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n4386) );
  XNOR2_X1 U4838 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n4385) );
  NOR3_X1 U4839 ( .A1(n4387), .A2(n4386), .A3(n4385), .ZN(n4388) );
  OAI21_X1 U4840 ( .B1(n4390), .B2(n4389), .A(n4388), .ZN(n4397) );
  XNOR2_X1 U4841 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n4394) );
  XNOR2_X1 U4842 ( .A(DATAI_5_), .B(keyinput_26), .ZN(n4393) );
  XNOR2_X1 U4843 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n4392) );
  XNOR2_X1 U4844 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n4391) );
  NOR4_X1 U4845 ( .A1(n4394), .A2(n4393), .A3(n4392), .A4(n4391), .ZN(n4396)
         );
  INV_X1 U4846 ( .A(DATAI_3_), .ZN(n5051) );
  XNOR2_X1 U4847 ( .A(n5051), .B(keyinput_28), .ZN(n4395) );
  AOI21_X1 U4848 ( .B1(n4397), .B2(n4396), .A(n4395), .ZN(n4400) );
  INV_X1 U4849 ( .A(DATAI_2_), .ZN(n5026) );
  XNOR2_X1 U4850 ( .A(n5026), .B(keyinput_29), .ZN(n4399) );
  XNOR2_X1 U4851 ( .A(n2849), .B(keyinput_30), .ZN(n4398) );
  OAI21_X1 U4852 ( .B1(n4400), .B2(n4399), .A(n4398), .ZN(n4403) );
  INV_X1 U4853 ( .A(DATAI_0_), .ZN(n4966) );
  XNOR2_X1 U4854 ( .A(n4966), .B(keyinput_31), .ZN(n4402) );
  XNOR2_X1 U4855 ( .A(U3149), .B(keyinput_32), .ZN(n4401) );
  NAND3_X1 U4856 ( .A1(n4403), .A2(n4402), .A3(n4401), .ZN(n4406) );
  XOR2_X1 U4857 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .Z(n4405) );
  XNOR2_X1 U4858 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_34), .ZN(n4404) );
  AOI21_X1 U4859 ( .B1(n4406), .B2(n4405), .A(n4404), .ZN(n4413) );
  XNOR2_X1 U4860 ( .A(n4603), .B(keyinput_36), .ZN(n4410) );
  XNOR2_X1 U4861 ( .A(n4602), .B(keyinput_37), .ZN(n4409) );
  XNOR2_X1 U4862 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_38), .ZN(n4408) );
  XNOR2_X1 U4863 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_35), .ZN(n4407) );
  NAND4_X1 U4864 ( .A1(n4410), .A2(n4409), .A3(n4408), .A4(n4407), .ZN(n4412)
         );
  XNOR2_X1 U4865 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .ZN(n4411) );
  OAI21_X1 U4866 ( .B1(n4413), .B2(n4412), .A(n4411), .ZN(n4431) );
  AOI22_X1 U4867 ( .A1(keyinput_41), .A2(n4416), .B1(n4418), .B2(keyinput_43), 
        .ZN(n4430) );
  AOI22_X1 U4868 ( .A1(n4617), .A2(keyinput_45), .B1(keyinput_42), .B2(
        REG3_REG_1__SCAN_IN), .ZN(n4429) );
  NAND2_X1 U4869 ( .A1(n4417), .A2(keyinput_40), .ZN(n4423) );
  OAI22_X1 U4870 ( .A1(n4427), .A2(keyinput_46), .B1(keyinput_44), .B2(
        REG3_REG_12__SCAN_IN), .ZN(n4415) );
  OAI22_X1 U4871 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_47), .B1(
        REG3_REG_1__SCAN_IN), .B2(keyinput_42), .ZN(n4414) );
  NOR2_X1 U4872 ( .A1(n4415), .A2(n4414), .ZN(n4422) );
  OAI22_X1 U4873 ( .A1(n4416), .A2(keyinput_41), .B1(n4617), .B2(keyinput_45), 
        .ZN(n4420) );
  OAI22_X1 U4874 ( .A1(n4418), .A2(keyinput_43), .B1(n4417), .B2(keyinput_40), 
        .ZN(n4419) );
  NOR2_X1 U4875 ( .A1(n4420), .A2(n4419), .ZN(n4421) );
  NAND3_X1 U4876 ( .A1(n4423), .A2(n4422), .A3(n4421), .ZN(n4426) );
  AOI22_X1 U4877 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_44), .B1(
        REG3_REG_5__SCAN_IN), .B2(keyinput_47), .ZN(n4424) );
  INV_X1 U4878 ( .A(n4424), .ZN(n4425) );
  AOI211_X1 U4879 ( .C1(keyinput_46), .C2(n4427), .A(n4426), .B(n4425), .ZN(
        n4428) );
  NAND4_X1 U4880 ( .A1(n4431), .A2(n4430), .A3(n4429), .A4(n4428), .ZN(n4434)
         );
  XOR2_X1 U4881 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_48), .Z(n4433) );
  XNOR2_X1 U4882 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_49), .ZN(n4432) );
  AOI21_X1 U4883 ( .B1(n4434), .B2(n4433), .A(n4432), .ZN(n4438) );
  XOR2_X1 U4884 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .Z(n4437) );
  XNOR2_X1 U4885 ( .A(n4435), .B(keyinput_51), .ZN(n4436) );
  OAI21_X1 U4886 ( .B1(n4438), .B2(n4437), .A(n4436), .ZN(n4440) );
  XNOR2_X1 U4887 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .ZN(n4439) );
  NAND2_X1 U4888 ( .A1(n4440), .A2(n4439), .ZN(n4444) );
  XOR2_X1 U4889 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .Z(n4443) );
  XNOR2_X1 U4890 ( .A(n4633), .B(keyinput_54), .ZN(n4442) );
  XNOR2_X1 U4891 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .ZN(n4441) );
  NAND4_X1 U4892 ( .A1(n4444), .A2(n4443), .A3(n4442), .A4(n4441), .ZN(n4449)
         );
  XOR2_X1 U4893 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .Z(n4448) );
  XNOR2_X1 U4894 ( .A(n4445), .B(keyinput_57), .ZN(n4447) );
  XNOR2_X1 U4895 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_58), .ZN(n4446) );
  AOI211_X1 U4896 ( .C1(n4449), .C2(n4448), .A(n4447), .B(n4446), .ZN(n4452)
         );
  XNOR2_X1 U4897 ( .A(n2748), .B(keyinput_59), .ZN(n4451) );
  XNOR2_X1 U4898 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4450) );
  NOR3_X1 U4899 ( .A1(n4452), .A2(n4451), .A3(n4450), .ZN(n4460) );
  INV_X1 U4900 ( .A(keyinput_63), .ZN(n4453) );
  XNOR2_X1 U4901 ( .A(n4453), .B(IR_REG_8__SCAN_IN), .ZN(n4457) );
  XNOR2_X1 U4902 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .ZN(n4456) );
  XNOR2_X1 U4903 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n4455) );
  XNOR2_X1 U4904 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n4454) );
  NAND4_X1 U4905 ( .A1(n4457), .A2(n4456), .A3(n4455), .A4(n4454), .ZN(n4459)
         );
  XNOR2_X1 U4906 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_65), .ZN(n4458) );
  OAI21_X1 U4907 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(n4463) );
  XOR2_X1 U4908 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_67), .Z(n4462) );
  XNOR2_X1 U4909 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_66), .ZN(n4461) );
  NAND3_X1 U4910 ( .A1(n4463), .A2(n4462), .A3(n4461), .ZN(n4468) );
  XNOR2_X1 U4911 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_68), .ZN(n4467) );
  XNOR2_X1 U4912 ( .A(n4464), .B(keyinput_69), .ZN(n4466) );
  XNOR2_X1 U4913 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_70), .ZN(n4465) );
  AOI211_X1 U4914 ( .C1(n4468), .C2(n4467), .A(n4466), .B(n4465), .ZN(n4471)
         );
  XOR2_X1 U4915 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_71), .Z(n4470) );
  XOR2_X1 U4916 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_72), .Z(n4469) );
  OAI21_X1 U4917 ( .B1(n4471), .B2(n4470), .A(n4469), .ZN(n4474) );
  XNOR2_X1 U4918 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_73), .ZN(n4473) );
  XNOR2_X1 U4919 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_74), .ZN(n4472) );
  NAND3_X1 U4920 ( .A1(n4474), .A2(n4473), .A3(n4472), .ZN(n4479) );
  XNOR2_X1 U4921 ( .A(n4475), .B(keyinput_76), .ZN(n4478) );
  XNOR2_X1 U4922 ( .A(n4669), .B(keyinput_75), .ZN(n4477) );
  XNOR2_X1 U4923 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_77), .ZN(n4476) );
  NAND4_X1 U4924 ( .A1(n4479), .A2(n4478), .A3(n4477), .A4(n4476), .ZN(n4483)
         );
  XNOR2_X1 U4925 ( .A(n4480), .B(keyinput_78), .ZN(n4482) );
  XNOR2_X1 U4926 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_79), .ZN(n4481) );
  NAND3_X1 U4927 ( .A1(n4483), .A2(n4482), .A3(n4481), .ZN(n4486) );
  XNOR2_X1 U4928 ( .A(n2759), .B(keyinput_80), .ZN(n4485) );
  XNOR2_X1 U4929 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_81), .ZN(n4484) );
  AOI21_X1 U4930 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(n4494) );
  XNOR2_X1 U4931 ( .A(n4680), .B(keyinput_85), .ZN(n4491) );
  XNOR2_X1 U4932 ( .A(n4681), .B(keyinput_83), .ZN(n4490) );
  XNOR2_X1 U4933 ( .A(n4487), .B(keyinput_82), .ZN(n4489) );
  XNOR2_X1 U4934 ( .A(n4682), .B(keyinput_84), .ZN(n4488) );
  NAND4_X1 U4935 ( .A1(n4491), .A2(n4490), .A3(n4489), .A4(n4488), .ZN(n4493)
         );
  XNOR2_X1 U4936 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .ZN(n4492) );
  OAI21_X1 U4937 ( .B1(n4494), .B2(n4493), .A(n4492), .ZN(n4498) );
  XNOR2_X1 U4938 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .ZN(n4497) );
  XNOR2_X1 U4939 ( .A(D_REG_0__SCAN_IN), .B(keyinput_87), .ZN(n4496) );
  XNOR2_X1 U4940 ( .A(D_REG_2__SCAN_IN), .B(keyinput_89), .ZN(n4495) );
  NAND4_X1 U4941 ( .A1(n4498), .A2(n4497), .A3(n4496), .A4(n4495), .ZN(n4501)
         );
  INV_X1 U4942 ( .A(D_REG_3__SCAN_IN), .ZN(n4780) );
  XNOR2_X1 U4943 ( .A(n4780), .B(keyinput_90), .ZN(n4500) );
  XNOR2_X1 U4944 ( .A(D_REG_4__SCAN_IN), .B(keyinput_91), .ZN(n4499) );
  AOI21_X1 U4945 ( .B1(n4501), .B2(n4500), .A(n4499), .ZN(n4504) );
  XNOR2_X1 U4946 ( .A(D_REG_6__SCAN_IN), .B(keyinput_93), .ZN(n4503) );
  XNOR2_X1 U4947 ( .A(D_REG_5__SCAN_IN), .B(keyinput_92), .ZN(n4502) );
  NOR3_X1 U4948 ( .A1(n4504), .A2(n4503), .A3(n4502), .ZN(n4508) );
  INV_X1 U4949 ( .A(D_REG_7__SCAN_IN), .ZN(n4784) );
  XNOR2_X1 U4950 ( .A(n4784), .B(keyinput_94), .ZN(n4507) );
  INV_X1 U4951 ( .A(D_REG_9__SCAN_IN), .ZN(n4785) );
  XNOR2_X1 U4952 ( .A(n4785), .B(keyinput_96), .ZN(n4506) );
  XNOR2_X1 U4953 ( .A(D_REG_8__SCAN_IN), .B(keyinput_95), .ZN(n4505) );
  NOR4_X1 U4954 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), .ZN(n4511)
         );
  INV_X1 U4955 ( .A(D_REG_10__SCAN_IN), .ZN(n4786) );
  XNOR2_X1 U4956 ( .A(n4786), .B(keyinput_97), .ZN(n4510) );
  INV_X1 U4957 ( .A(D_REG_11__SCAN_IN), .ZN(n4787) );
  XNOR2_X1 U4958 ( .A(n4787), .B(keyinput_98), .ZN(n4509) );
  NOR3_X1 U4959 ( .A1(n4511), .A2(n4510), .A3(n4509), .ZN(n4518) );
  INV_X1 U4960 ( .A(D_REG_12__SCAN_IN), .ZN(n4788) );
  XNOR2_X1 U4961 ( .A(n4788), .B(keyinput_99), .ZN(n4517) );
  INV_X1 U4962 ( .A(D_REG_13__SCAN_IN), .ZN(n4789) );
  XNOR2_X1 U4963 ( .A(n4789), .B(keyinput_100), .ZN(n4515) );
  INV_X1 U4964 ( .A(D_REG_14__SCAN_IN), .ZN(n4790) );
  XNOR2_X1 U4965 ( .A(n4790), .B(keyinput_101), .ZN(n4514) );
  XNOR2_X1 U4966 ( .A(D_REG_16__SCAN_IN), .B(keyinput_103), .ZN(n4513) );
  XNOR2_X1 U4967 ( .A(D_REG_15__SCAN_IN), .B(keyinput_102), .ZN(n4512) );
  NOR4_X1 U4968 ( .A1(n4515), .A2(n4514), .A3(n4513), .A4(n4512), .ZN(n4516)
         );
  OAI21_X1 U4969 ( .B1(n4518), .B2(n4517), .A(n4516), .ZN(n4521) );
  INV_X1 U4970 ( .A(D_REG_17__SCAN_IN), .ZN(n4791) );
  XNOR2_X1 U4971 ( .A(n4791), .B(keyinput_104), .ZN(n4520) );
  INV_X1 U4972 ( .A(D_REG_18__SCAN_IN), .ZN(n4792) );
  XNOR2_X1 U4973 ( .A(n4792), .B(keyinput_105), .ZN(n4519) );
  NAND3_X1 U4974 ( .A1(n4521), .A2(n4520), .A3(n4519), .ZN(n4524) );
  XNOR2_X1 U4975 ( .A(D_REG_19__SCAN_IN), .B(keyinput_106), .ZN(n4523) );
  XNOR2_X1 U4976 ( .A(D_REG_20__SCAN_IN), .B(keyinput_107), .ZN(n4522) );
  AOI21_X1 U4977 ( .B1(n4524), .B2(n4523), .A(n4522), .ZN(n4530) );
  INV_X1 U4978 ( .A(D_REG_21__SCAN_IN), .ZN(n4795) );
  XNOR2_X1 U4979 ( .A(n4795), .B(keyinput_108), .ZN(n4529) );
  INV_X1 U4980 ( .A(D_REG_24__SCAN_IN), .ZN(n4797) );
  XNOR2_X1 U4981 ( .A(n4797), .B(keyinput_111), .ZN(n4527) );
  XNOR2_X1 U4982 ( .A(D_REG_22__SCAN_IN), .B(keyinput_109), .ZN(n4526) );
  XNOR2_X1 U4983 ( .A(D_REG_23__SCAN_IN), .B(keyinput_110), .ZN(n4525) );
  NOR3_X1 U4984 ( .A1(n4527), .A2(n4526), .A3(n4525), .ZN(n4528) );
  OAI21_X1 U4985 ( .B1(n4530), .B2(n4529), .A(n4528), .ZN(n4533) );
  INV_X1 U4986 ( .A(D_REG_25__SCAN_IN), .ZN(n4798) );
  XNOR2_X1 U4987 ( .A(n4798), .B(keyinput_112), .ZN(n4532) );
  XNOR2_X1 U4988 ( .A(D_REG_26__SCAN_IN), .B(keyinput_113), .ZN(n4531) );
  AOI21_X1 U4989 ( .B1(n4533), .B2(n4532), .A(n4531), .ZN(n4536) );
  INV_X1 U4990 ( .A(D_REG_27__SCAN_IN), .ZN(n4800) );
  XNOR2_X1 U4991 ( .A(n4800), .B(keyinput_114), .ZN(n4535) );
  INV_X1 U4992 ( .A(D_REG_28__SCAN_IN), .ZN(n4801) );
  XNOR2_X1 U4993 ( .A(n4801), .B(keyinput_115), .ZN(n4534) );
  OAI21_X1 U4994 ( .B1(n4536), .B2(n4535), .A(n4534), .ZN(n4539) );
  XOR2_X1 U4995 ( .A(D_REG_29__SCAN_IN), .B(keyinput_116), .Z(n4538) );
  XNOR2_X1 U4996 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n4537) );
  NAND3_X1 U4997 ( .A1(n4539), .A2(n4538), .A3(n4537), .ZN(n4542) );
  XNOR2_X1 U4998 ( .A(n4737), .B(keyinput_119), .ZN(n4541) );
  XNOR2_X1 U4999 ( .A(D_REG_31__SCAN_IN), .B(keyinput_118), .ZN(n4540) );
  NAND3_X1 U5000 ( .A1(n4542), .A2(n4541), .A3(n4540), .ZN(n4548) );
  XOR2_X1 U5001 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .Z(n4547) );
  XNOR2_X1 U5002 ( .A(n4742), .B(keyinput_123), .ZN(n4545) );
  XNOR2_X1 U5003 ( .A(n4741), .B(keyinput_122), .ZN(n4544) );
  XNOR2_X1 U5004 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n4543) );
  NAND3_X1 U5005 ( .A1(n4545), .A2(n4544), .A3(n4543), .ZN(n4546) );
  AOI21_X1 U5006 ( .B1(n4548), .B2(n4547), .A(n4546), .ZN(n4551) );
  XNOR2_X1 U5007 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .ZN(n4550) );
  XNOR2_X1 U5008 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .ZN(n4549) );
  NOR3_X1 U5009 ( .A1(n4551), .A2(n4550), .A3(n4549), .ZN(n4758) );
  XOR2_X1 U5010 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .Z(n4757) );
  XOR2_X1 U5011 ( .A(DATAI_28_), .B(keyinput_131), .Z(n4555) );
  XOR2_X1 U5012 ( .A(DATAI_26_), .B(keyinput_133), .Z(n4554) );
  XNOR2_X1 U5013 ( .A(DATAI_25_), .B(keyinput_134), .ZN(n4553) );
  XNOR2_X1 U5014 ( .A(DATAI_31_), .B(keyinput_128), .ZN(n4552) );
  NOR4_X1 U5015 ( .A1(n4555), .A2(n4554), .A3(n4553), .A4(n4552), .ZN(n4559)
         );
  XOR2_X1 U5016 ( .A(DATAI_30_), .B(keyinput_129), .Z(n4558) );
  XNOR2_X1 U5017 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n4557) );
  XNOR2_X1 U5018 ( .A(DATAI_29_), .B(keyinput_130), .ZN(n4556) );
  NAND4_X1 U5019 ( .A1(n4559), .A2(n4558), .A3(n4557), .A4(n4556), .ZN(n4562)
         );
  XOR2_X1 U5020 ( .A(DATAI_23_), .B(keyinput_136), .Z(n4561) );
  XOR2_X1 U5021 ( .A(DATAI_24_), .B(keyinput_135), .Z(n4560) );
  NAND3_X1 U5022 ( .A1(n4562), .A2(n4561), .A3(n4560), .ZN(n4565) );
  XOR2_X1 U5023 ( .A(DATAI_21_), .B(keyinput_138), .Z(n4564) );
  XNOR2_X1 U5024 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n4563) );
  NAND3_X1 U5025 ( .A1(n4565), .A2(n4564), .A3(n4563), .ZN(n4568) );
  XNOR2_X1 U5026 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4567) );
  XNOR2_X1 U5027 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n4566) );
  AOI21_X1 U5028 ( .B1(n4568), .B2(n4567), .A(n4566), .ZN(n4571) );
  XOR2_X1 U5029 ( .A(DATAI_18_), .B(keyinput_141), .Z(n4570) );
  XOR2_X1 U5030 ( .A(DATAI_17_), .B(keyinput_142), .Z(n4569) );
  OAI21_X1 U5031 ( .B1(n4571), .B2(n4570), .A(n4569), .ZN(n4574) );
  XNOR2_X1 U5032 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n4573) );
  XNOR2_X1 U5033 ( .A(DATAI_15_), .B(keyinput_144), .ZN(n4572) );
  NAND3_X1 U5034 ( .A1(n4574), .A2(n4573), .A3(n4572), .ZN(n4584) );
  XNOR2_X1 U5035 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n4583) );
  XOR2_X1 U5036 ( .A(DATAI_10_), .B(keyinput_149), .Z(n4578) );
  XOR2_X1 U5037 ( .A(DATAI_11_), .B(keyinput_148), .Z(n4577) );
  XNOR2_X1 U5038 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n4576) );
  XNOR2_X1 U5039 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n4575) );
  NOR4_X1 U5040 ( .A1(n4578), .A2(n4577), .A3(n4576), .A4(n4575), .ZN(n4581)
         );
  XOR2_X1 U5041 ( .A(DATAI_8_), .B(keyinput_151), .Z(n4580) );
  INV_X1 U5042 ( .A(DATAI_9_), .ZN(n5084) );
  XNOR2_X1 U5043 ( .A(n5084), .B(keyinput_150), .ZN(n4579) );
  NAND3_X1 U5044 ( .A1(n4581), .A2(n4580), .A3(n4579), .ZN(n4582) );
  AOI21_X1 U5045 ( .B1(n4584), .B2(n4583), .A(n4582), .ZN(n4592) );
  INV_X1 U5046 ( .A(keyinput_154), .ZN(n4585) );
  XNOR2_X1 U5047 ( .A(n4585), .B(DATAI_5_), .ZN(n4589) );
  XNOR2_X1 U5048 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n4588) );
  XNOR2_X1 U5049 ( .A(DATAI_7_), .B(keyinput_152), .ZN(n4587) );
  XNOR2_X1 U5050 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n4586) );
  NAND4_X1 U5051 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4591)
         );
  XNOR2_X1 U5052 ( .A(n5051), .B(keyinput_156), .ZN(n4590) );
  OAI21_X1 U5053 ( .B1(n4592), .B2(n4591), .A(n4590), .ZN(n4595) );
  XNOR2_X1 U5054 ( .A(n5026), .B(keyinput_157), .ZN(n4594) );
  XNOR2_X1 U5055 ( .A(n2849), .B(keyinput_158), .ZN(n4593) );
  AOI21_X1 U5056 ( .B1(n4595), .B2(n4594), .A(n4593), .ZN(n4598) );
  XNOR2_X1 U5057 ( .A(n4966), .B(keyinput_159), .ZN(n4597) );
  XNOR2_X1 U5058 ( .A(STATE_REG_SCAN_IN), .B(keyinput_160), .ZN(n4596) );
  NOR3_X1 U5059 ( .A1(n4598), .A2(n4597), .A3(n4596), .ZN(n4601) );
  XNOR2_X1 U5060 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .ZN(n4600) );
  XNOR2_X1 U5061 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_162), .ZN(n4599) );
  OAI21_X1 U5062 ( .B1(n4601), .B2(n4600), .A(n4599), .ZN(n4611) );
  XOR2_X1 U5063 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_163), .Z(n4607) );
  XOR2_X1 U5064 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_166), .Z(n4606) );
  XNOR2_X1 U5065 ( .A(n4602), .B(keyinput_165), .ZN(n4605) );
  XNOR2_X1 U5066 ( .A(n4603), .B(keyinput_164), .ZN(n4604) );
  NOR4_X1 U5067 ( .A1(n4607), .A2(n4606), .A3(n4605), .A4(n4604), .ZN(n4610)
         );
  XNOR2_X1 U5068 ( .A(n4608), .B(keyinput_167), .ZN(n4609) );
  AOI21_X1 U5069 ( .B1(n4611), .B2(n4610), .A(n4609), .ZN(n4624) );
  XNOR2_X1 U5070 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_169), .ZN(n4615) );
  XNOR2_X1 U5071 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_171), .ZN(n4614) );
  XNOR2_X1 U5072 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .ZN(n4613) );
  XNOR2_X1 U5073 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_168), .ZN(n4612) );
  NAND4_X1 U5074 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4623)
         );
  XOR2_X1 U5075 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_174), .Z(n4621) );
  XOR2_X1 U5076 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_172), .Z(n4620) );
  XNOR2_X1 U5077 ( .A(n4616), .B(keyinput_175), .ZN(n4619) );
  XNOR2_X1 U5078 ( .A(n4617), .B(keyinput_173), .ZN(n4618) );
  NAND4_X1 U5079 ( .A1(n4621), .A2(n4620), .A3(n4619), .A4(n4618), .ZN(n4622)
         );
  NOR3_X1 U5080 ( .A1(n4624), .A2(n4623), .A3(n4622), .ZN(n4627) );
  XNOR2_X1 U5081 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_176), .ZN(n4626) );
  XNOR2_X1 U5082 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_177), .ZN(n4625) );
  OAI21_X1 U5083 ( .B1(n4627), .B2(n4626), .A(n4625), .ZN(n4630) );
  XNOR2_X1 U5084 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n4629) );
  XNOR2_X1 U5085 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_179), .ZN(n4628) );
  AOI21_X1 U5086 ( .B1(n4630), .B2(n4629), .A(n4628), .ZN(n4632) );
  XNOR2_X1 U5087 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .ZN(n4631) );
  NOR2_X1 U5088 ( .A1(n4632), .A2(n4631), .ZN(n4638) );
  XNOR2_X1 U5089 ( .A(n4633), .B(keyinput_182), .ZN(n4637) );
  XNOR2_X1 U5090 ( .A(n4634), .B(keyinput_181), .ZN(n4636) );
  XNOR2_X1 U5091 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .ZN(n4635) );
  NOR4_X1 U5092 ( .A1(n4638), .A2(n4637), .A3(n4636), .A4(n4635), .ZN(n4642)
         );
  XNOR2_X1 U5093 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .ZN(n4641) );
  XNOR2_X1 U5094 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_185), .ZN(n4640) );
  XNOR2_X1 U5095 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_186), .ZN(n4639) );
  OAI211_X1 U5096 ( .C1(n4642), .C2(n4641), .A(n4640), .B(n4639), .ZN(n4646)
         );
  XNOR2_X1 U5097 ( .A(n4643), .B(keyinput_188), .ZN(n4645) );
  XNOR2_X1 U5098 ( .A(n2748), .B(keyinput_187), .ZN(n4644) );
  NAND3_X1 U5099 ( .A1(n4646), .A2(n4645), .A3(n4644), .ZN(n4654) );
  XOR2_X1 U5100 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_192), .Z(n4651) );
  XOR2_X1 U5101 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_189), .Z(n4650) );
  XNOR2_X1 U5102 ( .A(n4647), .B(keyinput_190), .ZN(n4649) );
  XNOR2_X1 U5103 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_191), .ZN(n4648) );
  NOR4_X1 U5104 ( .A1(n4651), .A2(n4650), .A3(n4649), .A4(n4648), .ZN(n4653)
         );
  XNOR2_X1 U5105 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_193), .ZN(n4652) );
  AOI21_X1 U5106 ( .B1(n4654), .B2(n4653), .A(n4652), .ZN(n4657) );
  XOR2_X1 U5107 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_195), .Z(n4656) );
  XNOR2_X1 U5108 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_194), .ZN(n4655) );
  NOR3_X1 U5109 ( .A1(n4657), .A2(n4656), .A3(n4655), .ZN(n4661) );
  XNOR2_X1 U5110 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_196), .ZN(n4660) );
  XNOR2_X1 U5111 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n4659) );
  XNOR2_X1 U5112 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n4658) );
  OAI211_X1 U5113 ( .C1(n4661), .C2(n4660), .A(n4659), .B(n4658), .ZN(n4664)
         );
  XOR2_X1 U5114 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_199), .Z(n4663) );
  XOR2_X1 U5115 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_200), .Z(n4662) );
  AOI21_X1 U5116 ( .B1(n4664), .B2(n4663), .A(n4662), .ZN(n4668) );
  XNOR2_X1 U5117 ( .A(n4665), .B(keyinput_201), .ZN(n4667) );
  XNOR2_X1 U5118 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_202), .ZN(n4666) );
  NOR3_X1 U5119 ( .A1(n4668), .A2(n4667), .A3(n4666), .ZN(n4673) );
  XNOR2_X1 U5120 ( .A(n4669), .B(keyinput_203), .ZN(n4672) );
  XNOR2_X1 U5121 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_205), .ZN(n4671) );
  XNOR2_X1 U5122 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n4670) );
  NOR4_X1 U5123 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4676)
         );
  XNOR2_X1 U5124 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_207), .ZN(n4675) );
  XNOR2_X1 U5125 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_206), .ZN(n4674) );
  NOR3_X1 U5126 ( .A1(n4676), .A2(n4675), .A3(n4674), .ZN(n4679) );
  XNOR2_X1 U5127 ( .A(n2759), .B(keyinput_208), .ZN(n4678) );
  XNOR2_X1 U5128 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_209), .ZN(n4677) );
  OAI21_X1 U5129 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(n4689) );
  XNOR2_X1 U5130 ( .A(n4680), .B(keyinput_213), .ZN(n4686) );
  XNOR2_X1 U5131 ( .A(n4681), .B(keyinput_211), .ZN(n4685) );
  XNOR2_X1 U5132 ( .A(n4682), .B(keyinput_212), .ZN(n4684) );
  XNOR2_X1 U5133 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_210), .ZN(n4683) );
  NOR4_X1 U5134 ( .A1(n4686), .A2(n4685), .A3(n4684), .A4(n4683), .ZN(n4688)
         );
  XOR2_X1 U5135 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .Z(n4687) );
  AOI21_X1 U5136 ( .B1(n4689), .B2(n4688), .A(n4687), .ZN(n4697) );
  INV_X1 U5137 ( .A(keyinput_217), .ZN(n4694) );
  INV_X1 U5138 ( .A(D_REG_2__SCAN_IN), .ZN(n4779) );
  OAI22_X1 U5139 ( .A1(n4691), .A2(keyinput_216), .B1(n4779), .B2(keyinput_217), .ZN(n4690) );
  AOI21_X1 U5140 ( .B1(n4691), .B2(keyinput_216), .A(n4690), .ZN(n4693) );
  XNOR2_X1 U5141 ( .A(D_REG_0__SCAN_IN), .B(keyinput_215), .ZN(n4692) );
  OAI211_X1 U5142 ( .C1(D_REG_2__SCAN_IN), .C2(n4694), .A(n4693), .B(n4692), 
        .ZN(n4696) );
  XNOR2_X1 U5143 ( .A(D_REG_3__SCAN_IN), .B(keyinput_218), .ZN(n4695) );
  OAI21_X1 U5144 ( .B1(n4697), .B2(n4696), .A(n4695), .ZN(n4701) );
  XNOR2_X1 U5145 ( .A(D_REG_4__SCAN_IN), .B(keyinput_219), .ZN(n4700) );
  INV_X1 U5146 ( .A(D_REG_6__SCAN_IN), .ZN(n4783) );
  XNOR2_X1 U5147 ( .A(n4783), .B(keyinput_221), .ZN(n4699) );
  INV_X1 U5148 ( .A(D_REG_5__SCAN_IN), .ZN(n4782) );
  XNOR2_X1 U5149 ( .A(n4782), .B(keyinput_220), .ZN(n4698) );
  AOI211_X1 U5150 ( .C1(n4701), .C2(n4700), .A(n4699), .B(n4698), .ZN(n4705)
         );
  XNOR2_X1 U5151 ( .A(n4785), .B(keyinput_224), .ZN(n4704) );
  XNOR2_X1 U5152 ( .A(n4784), .B(keyinput_222), .ZN(n4703) );
  XOR2_X1 U5153 ( .A(D_REG_8__SCAN_IN), .B(keyinput_223), .Z(n4702) );
  NOR4_X1 U5154 ( .A1(n4705), .A2(n4704), .A3(n4703), .A4(n4702), .ZN(n4708)
         );
  XNOR2_X1 U5155 ( .A(D_REG_11__SCAN_IN), .B(keyinput_226), .ZN(n4707) );
  XNOR2_X1 U5156 ( .A(D_REG_10__SCAN_IN), .B(keyinput_225), .ZN(n4706) );
  NOR3_X1 U5157 ( .A1(n4708), .A2(n4707), .A3(n4706), .ZN(n4715) );
  XNOR2_X1 U5158 ( .A(D_REG_12__SCAN_IN), .B(keyinput_227), .ZN(n4714) );
  XNOR2_X1 U5159 ( .A(D_REG_16__SCAN_IN), .B(keyinput_231), .ZN(n4712) );
  XNOR2_X1 U5160 ( .A(D_REG_15__SCAN_IN), .B(keyinput_230), .ZN(n4711) );
  XNOR2_X1 U5161 ( .A(D_REG_13__SCAN_IN), .B(keyinput_228), .ZN(n4710) );
  XNOR2_X1 U5162 ( .A(D_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n4709) );
  NOR4_X1 U5163 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4713)
         );
  OAI21_X1 U5164 ( .B1(n4715), .B2(n4714), .A(n4713), .ZN(n4718) );
  XNOR2_X1 U5165 ( .A(D_REG_18__SCAN_IN), .B(keyinput_233), .ZN(n4717) );
  XNOR2_X1 U5166 ( .A(D_REG_17__SCAN_IN), .B(keyinput_232), .ZN(n4716) );
  NAND3_X1 U5167 ( .A1(n4718), .A2(n4717), .A3(n4716), .ZN(n4721) );
  INV_X1 U5168 ( .A(D_REG_19__SCAN_IN), .ZN(n4793) );
  XNOR2_X1 U5169 ( .A(n4793), .B(keyinput_234), .ZN(n4720) );
  INV_X1 U5170 ( .A(D_REG_20__SCAN_IN), .ZN(n4794) );
  XNOR2_X1 U5171 ( .A(n4794), .B(keyinput_235), .ZN(n4719) );
  AOI21_X1 U5172 ( .B1(n4721), .B2(n4720), .A(n4719), .ZN(n4727) );
  XNOR2_X1 U5173 ( .A(n4795), .B(keyinput_236), .ZN(n4726) );
  INV_X1 U5174 ( .A(D_REG_23__SCAN_IN), .ZN(n4796) );
  XNOR2_X1 U5175 ( .A(n4796), .B(keyinput_238), .ZN(n4724) );
  XNOR2_X1 U5176 ( .A(D_REG_22__SCAN_IN), .B(keyinput_237), .ZN(n4723) );
  XNOR2_X1 U5177 ( .A(D_REG_24__SCAN_IN), .B(keyinput_239), .ZN(n4722) );
  NOR3_X1 U5178 ( .A1(n4724), .A2(n4723), .A3(n4722), .ZN(n4725) );
  OAI21_X1 U5179 ( .B1(n4727), .B2(n4726), .A(n4725), .ZN(n4730) );
  XNOR2_X1 U5180 ( .A(D_REG_25__SCAN_IN), .B(keyinput_240), .ZN(n4729) );
  XNOR2_X1 U5181 ( .A(D_REG_26__SCAN_IN), .B(keyinput_241), .ZN(n4728) );
  AOI21_X1 U5182 ( .B1(n4730), .B2(n4729), .A(n4728), .ZN(n4733) );
  XNOR2_X1 U5183 ( .A(D_REG_27__SCAN_IN), .B(keyinput_242), .ZN(n4732) );
  XNOR2_X1 U5184 ( .A(n4801), .B(keyinput_243), .ZN(n4731) );
  OAI21_X1 U5185 ( .B1(n4733), .B2(n4732), .A(n4731), .ZN(n4736) );
  XOR2_X1 U5186 ( .A(D_REG_29__SCAN_IN), .B(keyinput_244), .Z(n4735) );
  XNOR2_X1 U5187 ( .A(D_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n4734) );
  NAND3_X1 U5188 ( .A1(n4736), .A2(n4735), .A3(n4734), .ZN(n4740) );
  INV_X1 U5189 ( .A(D_REG_31__SCAN_IN), .ZN(n4804) );
  XNOR2_X1 U5190 ( .A(n4804), .B(keyinput_246), .ZN(n4739) );
  XNOR2_X1 U5191 ( .A(n4737), .B(keyinput_247), .ZN(n4738) );
  NAND3_X1 U5192 ( .A1(n4740), .A2(n4739), .A3(n4738), .ZN(n4748) );
  XNOR2_X1 U5193 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .ZN(n4747) );
  XNOR2_X1 U5194 ( .A(n4741), .B(keyinput_250), .ZN(n4745) );
  XNOR2_X1 U5195 ( .A(n4742), .B(keyinput_251), .ZN(n4744) );
  XNOR2_X1 U5196 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .ZN(n4743) );
  NAND3_X1 U5197 ( .A1(n4745), .A2(n4744), .A3(n4743), .ZN(n4746) );
  AOI21_X1 U5198 ( .B1(n4748), .B2(n4747), .A(n4746), .ZN(n4751) );
  XOR2_X1 U5199 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .Z(n4750) );
  XOR2_X1 U5200 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .Z(n4749) );
  NOR3_X1 U5201 ( .A1(n4751), .A2(n4750), .A3(n4749), .ZN(n4754) );
  XNOR2_X1 U5202 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .ZN(n4753) );
  XOR2_X1 U5203 ( .A(keyinput_127), .B(keyinput_255), .Z(n4752) );
  OAI21_X1 U5204 ( .B1(n4754), .B2(n4753), .A(n4752), .ZN(n4756) );
  XOR2_X1 U5205 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .Z(n4755) );
  OAI211_X1 U5206 ( .C1(n4758), .C2(n4757), .A(n4756), .B(n4755), .ZN(n4762)
         );
  OAI21_X1 U5207 ( .B1(n5204), .B2(n4760), .A(n4759), .ZN(n5156) );
  MUX2_X1 U5208 ( .A(REG0_REG_14__SCAN_IN), .B(n5156), .S(n5259), .Z(n4761) );
  XNOR2_X1 U5209 ( .A(n4762), .B(n4761), .ZN(U3495) );
  NOR3_X1 U5210 ( .A1(n4763), .A2(IR_REG_30__SCAN_IN), .A3(n2761), .ZN(n4764)
         );
  MUX2_X1 U5211 ( .A(DATAI_31_), .B(n4764), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5212 ( .A(DATAI_30_), .B(n4765), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5213 ( .A(n4766), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5214 ( .A(n4767), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5215 ( .A(DATAI_24_), .B(n3093), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5216 ( .A(n4768), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5217 ( .A(n4769), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5218 ( .A(DATAI_18_), .B(n4770), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5219 ( .A(DATAI_17_), .B(n4771), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U5220 ( .A(n4772), .B(DATAI_16_), .S(U3149), .Z(U3336) );
  MUX2_X1 U5221 ( .A(n4773), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5222 ( .A(DATAI_14_), .B(n4937), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  INV_X1 U5223 ( .A(n4930), .ZN(n4774) );
  MUX2_X1 U5224 ( .A(DATAI_13_), .B(n4774), .S(STATE_REG_SCAN_IN), .Z(U3339)
         );
  MUX2_X1 U5225 ( .A(DATAI_11_), .B(n4775), .S(STATE_REG_SCAN_IN), .Z(U3341)
         );
  MUX2_X1 U5226 ( .A(n4891), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5227 ( .A(DATAI_8_), .B(n4873), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5228 ( .A(DATAI_7_), .B(n4776), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5229 ( .A(DATAI_6_), .B(n4851), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5230 ( .A(DATAI_4_), .B(n4989), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  INV_X1 U5231 ( .A(DATAI_23_), .ZN(n4778) );
  AOI21_X1 U5232 ( .B1(U3149), .B2(n4778), .A(n4777), .ZN(U3329) );
  INV_X2 U5233 ( .A(n4802), .ZN(n4805) );
  NOR2_X1 U5234 ( .A1(n4805), .A2(n4779), .ZN(U3320) );
  NOR2_X1 U5235 ( .A1(n4805), .A2(n4780), .ZN(U3319) );
  INV_X1 U5236 ( .A(D_REG_4__SCAN_IN), .ZN(n4781) );
  NOR2_X1 U5237 ( .A1(n4805), .A2(n4781), .ZN(U3318) );
  NOR2_X1 U5238 ( .A1(n4805), .A2(n4782), .ZN(U3317) );
  NOR2_X1 U5239 ( .A1(n4805), .A2(n4783), .ZN(U3316) );
  NOR2_X1 U5240 ( .A1(n4805), .A2(n4784), .ZN(U3315) );
  AND2_X1 U5241 ( .A1(n4802), .A2(D_REG_8__SCAN_IN), .ZN(U3314) );
  NOR2_X1 U5242 ( .A1(n4805), .A2(n4785), .ZN(U3313) );
  NOR2_X1 U5243 ( .A1(n4805), .A2(n4786), .ZN(U3312) );
  NOR2_X1 U5244 ( .A1(n4805), .A2(n4787), .ZN(U3311) );
  NOR2_X1 U5245 ( .A1(n4805), .A2(n4788), .ZN(U3310) );
  NOR2_X1 U5246 ( .A1(n4805), .A2(n4789), .ZN(U3309) );
  NOR2_X1 U5247 ( .A1(n4805), .A2(n4790), .ZN(U3308) );
  AND2_X1 U5248 ( .A1(n4802), .A2(D_REG_15__SCAN_IN), .ZN(U3307) );
  AND2_X1 U5249 ( .A1(n4802), .A2(D_REG_16__SCAN_IN), .ZN(U3306) );
  NOR2_X1 U5250 ( .A1(n4805), .A2(n4791), .ZN(U3305) );
  NOR2_X1 U5251 ( .A1(n4805), .A2(n4792), .ZN(U3304) );
  NOR2_X1 U5252 ( .A1(n4805), .A2(n4793), .ZN(U3303) );
  NOR2_X1 U5253 ( .A1(n4805), .A2(n4794), .ZN(U3302) );
  NOR2_X1 U5254 ( .A1(n4805), .A2(n4795), .ZN(U3301) );
  AND2_X1 U5255 ( .A1(n4802), .A2(D_REG_22__SCAN_IN), .ZN(U3300) );
  NOR2_X1 U5256 ( .A1(n4805), .A2(n4796), .ZN(U3299) );
  NOR2_X1 U5257 ( .A1(n4805), .A2(n4797), .ZN(U3298) );
  NOR2_X1 U5258 ( .A1(n4805), .A2(n4798), .ZN(U3297) );
  INV_X1 U5259 ( .A(D_REG_26__SCAN_IN), .ZN(n4799) );
  NOR2_X1 U5260 ( .A1(n4805), .A2(n4799), .ZN(U3296) );
  NOR2_X1 U5261 ( .A1(n4805), .A2(n4800), .ZN(U3295) );
  NOR2_X1 U5262 ( .A1(n4805), .A2(n4801), .ZN(U3294) );
  AND2_X1 U5263 ( .A1(n4802), .A2(D_REG_29__SCAN_IN), .ZN(U3293) );
  INV_X1 U5264 ( .A(D_REG_30__SCAN_IN), .ZN(n4803) );
  NOR2_X1 U5265 ( .A1(n4805), .A2(n4803), .ZN(U3292) );
  NOR2_X1 U5266 ( .A1(n4805), .A2(n4804), .ZN(U3291) );
  OR2_X1 U5267 ( .A1(n3143), .A2(REG2_REG_0__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U5268 ( .A1(n4807), .A2(n4806), .ZN(n4811) );
  INV_X1 U5269 ( .A(n4811), .ZN(n4808) );
  NAND2_X1 U5270 ( .A1(n3143), .A2(n2837), .ZN(n4809) );
  NAND2_X1 U5271 ( .A1(n4808), .A2(n4809), .ZN(n4810) );
  MUX2_X1 U5272 ( .A(n4810), .B(n4809), .S(n4967), .Z(n4812) );
  NAND2_X1 U5273 ( .A1(n4811), .A2(n4967), .ZN(n4969) );
  NAND2_X1 U5274 ( .A1(n4812), .A2(n4969), .ZN(n4814) );
  AOI22_X1 U5275 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4988), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4813) );
  OAI21_X1 U5276 ( .B1(n4815), .B2(n4814), .A(n4813), .ZN(U3240) );
  AOI22_X1 U5277 ( .A1(ADDR_REG_1__SCAN_IN), .A2(n4988), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4827) );
  NOR2_X1 U5278 ( .A1(n4967), .A2(n2837), .ZN(n4819) );
  OAI211_X1 U5279 ( .C1(n4819), .C2(n4818), .A(n4992), .B(n4817), .ZN(n4826)
         );
  NAND2_X1 U5280 ( .A1(n4990), .A2(n4820), .ZN(n4825) );
  NAND2_X1 U5281 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4971) );
  INV_X1 U5282 ( .A(n4971), .ZN(n4823) );
  OAI211_X1 U5283 ( .C1(n4823), .C2(n4822), .A(n4995), .B(n4821), .ZN(n4824)
         );
  NAND4_X1 U5284 ( .A1(n4827), .A2(n4826), .A3(n4825), .A4(n4824), .ZN(U3241)
         );
  OAI211_X1 U5285 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4829), .A(n4992), .B(n4828), 
        .ZN(n4833) );
  OAI211_X1 U5286 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4831), .A(n4995), .B(n4830), 
        .ZN(n4832) );
  OAI211_X1 U5287 ( .C1(n4958), .C2(n4029), .A(n4833), .B(n4832), .ZN(n4834)
         );
  AOI211_X1 U5288 ( .C1(n4988), .C2(ADDR_REG_3__SCAN_IN), .A(n4835), .B(n4834), 
        .ZN(n4836) );
  INV_X1 U5289 ( .A(n4836), .ZN(U3243) );
  OAI211_X1 U5290 ( .C1(n4839), .C2(n4838), .A(n4992), .B(n4837), .ZN(n4844)
         );
  OAI211_X1 U5291 ( .C1(n4842), .C2(n4841), .A(n4995), .B(n4840), .ZN(n4843)
         );
  OAI211_X1 U5292 ( .C1(n4958), .C2(n5059), .A(n4844), .B(n4843), .ZN(n4845)
         );
  AOI211_X1 U5293 ( .C1(n4988), .C2(ADDR_REG_5__SCAN_IN), .A(n4846), .B(n4845), 
        .ZN(n4847) );
  INV_X1 U5294 ( .A(n4847), .ZN(U3245) );
  AOI21_X1 U5295 ( .B1(n4988), .B2(ADDR_REG_6__SCAN_IN), .A(n4848), .ZN(n4857)
         );
  OAI211_X1 U5296 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4850), .A(n4995), .B(n4849), 
        .ZN(n4856) );
  NAND2_X1 U5297 ( .A1(n4990), .A2(n4851), .ZN(n4855) );
  OAI211_X1 U5298 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4853), .A(n4992), .B(n4852), 
        .ZN(n4854) );
  NAND4_X1 U5299 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(U3246)
         );
  OAI211_X1 U5300 ( .C1(n4860), .C2(n4859), .A(n4992), .B(n4858), .ZN(n4865)
         );
  OAI211_X1 U5301 ( .C1(n4863), .C2(n4862), .A(n4995), .B(n4861), .ZN(n4864)
         );
  OAI211_X1 U5302 ( .C1(n4958), .C2(n4866), .A(n4865), .B(n4864), .ZN(n4867)
         );
  AOI211_X1 U5303 ( .C1(n4988), .C2(ADDR_REG_7__SCAN_IN), .A(n4868), .B(n4867), 
        .ZN(n4869) );
  INV_X1 U5304 ( .A(n4869), .ZN(U3247) );
  AOI21_X1 U5305 ( .B1(n4988), .B2(ADDR_REG_8__SCAN_IN), .A(n4870), .ZN(n4879)
         );
  OAI211_X1 U5306 ( .C1(n4872), .C2(REG1_REG_8__SCAN_IN), .A(n4992), .B(n4871), 
        .ZN(n4878) );
  NAND2_X1 U5307 ( .A1(n4990), .A2(n4873), .ZN(n4877) );
  OAI211_X1 U5308 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4875), .A(n4995), .B(n4874), 
        .ZN(n4876) );
  NAND4_X1 U5309 ( .A1(n4879), .A2(n4878), .A3(n4877), .A4(n4876), .ZN(U3248)
         );
  OAI211_X1 U5310 ( .C1(n4882), .C2(n4881), .A(n4992), .B(n4880), .ZN(n4887)
         );
  OAI211_X1 U5311 ( .C1(n4885), .C2(n4884), .A(n4995), .B(n4883), .ZN(n4886)
         );
  OAI211_X1 U5312 ( .C1(n4958), .C2(n5085), .A(n4887), .B(n4886), .ZN(n4888)
         );
  AOI211_X1 U5313 ( .C1(n4988), .C2(ADDR_REG_9__SCAN_IN), .A(n4889), .B(n4888), 
        .ZN(n4890) );
  INV_X1 U5314 ( .A(n4890), .ZN(U3249) );
  OAI211_X1 U5315 ( .C1(n4893), .C2(REG2_REG_10__SCAN_IN), .A(n4995), .B(n4892), .ZN(n4897) );
  OAI211_X1 U5316 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4895), .A(n4992), .B(n4894), .ZN(n4896) );
  OAI211_X1 U5317 ( .C1(n4958), .C2(n4041), .A(n4897), .B(n4896), .ZN(n4898)
         );
  AOI211_X1 U5318 ( .C1(n4988), .C2(ADDR_REG_10__SCAN_IN), .A(n4899), .B(n4898), .ZN(n4900) );
  INV_X1 U5319 ( .A(n4900), .ZN(U3250) );
  OAI211_X1 U5320 ( .C1(n4903), .C2(n4902), .A(n4992), .B(n4901), .ZN(n4908)
         );
  OAI211_X1 U5321 ( .C1(n4906), .C2(n4905), .A(n4995), .B(n4904), .ZN(n4907)
         );
  OAI211_X1 U5322 ( .C1(n4958), .C2(n4909), .A(n4908), .B(n4907), .ZN(n4910)
         );
  AOI211_X1 U5323 ( .C1(n4988), .C2(ADDR_REG_11__SCAN_IN), .A(n4911), .B(n4910), .ZN(n4912) );
  INV_X1 U5324 ( .A(n4912), .ZN(U3251) );
  OAI211_X1 U5325 ( .C1(n4914), .C2(REG2_REG_12__SCAN_IN), .A(n4995), .B(n4913), .ZN(n4918) );
  OAI211_X1 U5326 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4916), .A(n4992), .B(n4915), .ZN(n4917) );
  OAI211_X1 U5327 ( .C1(n4958), .C2(n5143), .A(n4918), .B(n4917), .ZN(n4919)
         );
  AOI211_X1 U5328 ( .C1(n4988), .C2(ADDR_REG_12__SCAN_IN), .A(n4920), .B(n4919), .ZN(n4921) );
  INV_X1 U5329 ( .A(n4921), .ZN(U3252) );
  OAI211_X1 U5330 ( .C1(n4924), .C2(n4923), .A(n4922), .B(n4992), .ZN(n4929)
         );
  OAI211_X1 U5331 ( .C1(n4927), .C2(n4926), .A(n4925), .B(n4995), .ZN(n4928)
         );
  OAI211_X1 U5332 ( .C1(n4958), .C2(n4930), .A(n4929), .B(n4928), .ZN(n4931)
         );
  AOI211_X1 U5333 ( .C1(n4988), .C2(ADDR_REG_13__SCAN_IN), .A(n4932), .B(n4931), .ZN(n4933) );
  INV_X1 U5334 ( .A(n4933), .ZN(U3253) );
  AOI21_X1 U5335 ( .B1(n4988), .B2(ADDR_REG_14__SCAN_IN), .A(n4934), .ZN(n4943) );
  OAI211_X1 U5336 ( .C1(n4936), .C2(REG1_REG_14__SCAN_IN), .A(n4992), .B(n4935), .ZN(n4942) );
  NAND2_X1 U5337 ( .A1(n4990), .A2(n4937), .ZN(n4941) );
  OAI211_X1 U5338 ( .C1(REG2_REG_14__SCAN_IN), .C2(n4939), .A(n4995), .B(n4938), .ZN(n4940) );
  NAND4_X1 U5339 ( .A1(n4943), .A2(n4942), .A3(n4941), .A4(n4940), .ZN(U3254)
         );
  AND2_X1 U5340 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n5164) );
  OAI211_X1 U5341 ( .C1(n4946), .C2(n4945), .A(n4992), .B(n4944), .ZN(n4947)
         );
  OAI21_X1 U5342 ( .B1(n4958), .B2(n4948), .A(n4947), .ZN(n4949) );
  AOI211_X1 U5343 ( .C1(n4988), .C2(ADDR_REG_15__SCAN_IN), .A(n5164), .B(n4949), .ZN(n4954) );
  OAI211_X1 U5344 ( .C1(n4952), .C2(n4951), .A(n4995), .B(n4950), .ZN(n4953)
         );
  NAND2_X1 U5345 ( .A1(n4954), .A2(n4953), .ZN(U3255) );
  NAND2_X1 U5346 ( .A1(n4959), .A2(REG1_REG_18__SCAN_IN), .ZN(n4955) );
  OAI211_X1 U5347 ( .C1(n4959), .C2(REG1_REG_18__SCAN_IN), .A(n4956), .B(n4955), .ZN(n4957) );
  OAI211_X1 U5348 ( .C1(n4964), .C2(n4963), .A(n4995), .B(n4962), .ZN(n4965)
         );
  AOI22_X1 U5349 ( .A1(STATE_REG_SCAN_IN), .A2(n4967), .B1(n4966), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5350 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4988), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4985) );
  INV_X1 U5351 ( .A(n3143), .ZN(n4968) );
  NOR2_X1 U5352 ( .A1(n4968), .A2(n3127), .ZN(n4973) );
  OAI211_X1 U5353 ( .C1(n4971), .C2(n4970), .A(U4043), .B(n4969), .ZN(n4972)
         );
  AOI21_X1 U5354 ( .B1(n4974), .B2(n4973), .A(n4972), .ZN(n4987) );
  AOI21_X1 U5355 ( .B1(n4990), .B2(n4975), .A(n4987), .ZN(n4984) );
  OAI211_X1 U5356 ( .C1(n4978), .C2(n4977), .A(n4992), .B(n4976), .ZN(n4983)
         );
  OAI211_X1 U5357 ( .C1(n4981), .C2(n4980), .A(n4995), .B(n4979), .ZN(n4982)
         );
  NAND4_X1 U5358 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(U3242)
         );
  AOI211_X1 U5359 ( .C1(n4988), .C2(ADDR_REG_4__SCAN_IN), .A(n4987), .B(n4986), 
        .ZN(n5000) );
  NAND2_X1 U5360 ( .A1(n4990), .A2(n4989), .ZN(n4999) );
  OAI211_X1 U5361 ( .C1(REG1_REG_4__SCAN_IN), .C2(n4993), .A(n4992), .B(n4991), 
        .ZN(n4998) );
  OAI211_X1 U5362 ( .C1(REG2_REG_4__SCAN_IN), .C2(n4996), .A(n4995), .B(n4994), 
        .ZN(n4997) );
  NAND4_X1 U5363 ( .A1(n5000), .A2(n4999), .A3(n4998), .A4(n4997), .ZN(U3244)
         );
  AOI21_X1 U5364 ( .B1(n2504), .B2(n5004), .A(n5001), .ZN(n5002) );
  AOI22_X1 U5365 ( .A1(n5256), .A2(n5002), .B1(n2837), .B2(n5254), .ZN(U3518)
         );
  AOI22_X1 U5366 ( .A1(n5259), .A2(n5002), .B1(n4737), .B2(n5257), .ZN(U3467)
         );
  AOI22_X1 U5367 ( .A1(STATE_REG_SCAN_IN), .A2(n5003), .B1(n2849), .B2(U3149), 
        .ZN(U3351) );
  NAND2_X1 U5368 ( .A1(n5014), .A2(n5004), .ZN(n5005) );
  AND2_X1 U5369 ( .A1(n5029), .A2(n5005), .ZN(n5022) );
  OAI21_X1 U5370 ( .B1(n5007), .B2(n5006), .A(n5037), .ZN(n5009) );
  NAND2_X1 U5371 ( .A1(n5009), .A2(n5008), .ZN(n5018) );
  AOI22_X1 U5372 ( .A1(n5120), .A2(n3992), .B1(n5010), .B2(n5117), .ZN(n5017)
         );
  OAI211_X1 U5373 ( .C1(n5013), .C2(n5012), .A(n5227), .B(n5011), .ZN(n5016)
         );
  NAND2_X1 U5374 ( .A1(n5240), .A2(n5014), .ZN(n5015) );
  AND4_X1 U5375 ( .A1(n5018), .A2(n5017), .A3(n5016), .A4(n5015), .ZN(n5025)
         );
  INV_X1 U5376 ( .A(n5025), .ZN(n5019) );
  AOI21_X1 U5377 ( .B1(n5252), .B2(n5022), .A(n5019), .ZN(n5021) );
  AOI22_X1 U5378 ( .A1(n5256), .A2(n5021), .B1(n3997), .B2(n5254), .ZN(U3519)
         );
  AOI22_X1 U5379 ( .A1(n5259), .A2(n5021), .B1(n5020), .B2(n5257), .ZN(U3469)
         );
  AOI22_X1 U5380 ( .A1(n5247), .A2(n5022), .B1(REG3_REG_1__SCAN_IN), .B2(n5135), .ZN(n5023) );
  OAI221_X1 U5381 ( .B1(n5249), .B2(n5025), .C1(n5140), .C2(n5024), .A(n5023), 
        .ZN(U3289) );
  AOI22_X1 U5382 ( .A1(STATE_REG_SCAN_IN), .A2(n5027), .B1(n5026), .B2(U3149), 
        .ZN(U3350) );
  NAND2_X1 U5383 ( .A1(n5029), .A2(n5028), .ZN(n5030) );
  NAND2_X1 U5384 ( .A1(n5031), .A2(n5030), .ZN(n5046) );
  OAI21_X1 U5385 ( .B1(n2747), .B2(n2565), .A(n5033), .ZN(n5042) );
  AOI22_X1 U5386 ( .A1(n5117), .A2(n5034), .B1(n3237), .B2(n5120), .ZN(n5035)
         );
  OAI21_X1 U5387 ( .B1(n5123), .B2(n2824), .A(n5035), .ZN(n5041) );
  NAND3_X1 U5388 ( .A1(n5037), .A2(n2565), .A3(n5036), .ZN(n5038) );
  AOI21_X1 U5389 ( .B1(n5039), .B2(n5038), .A(n5217), .ZN(n5040) );
  AOI211_X1 U5390 ( .C1(n5227), .C2(n5042), .A(n5041), .B(n5040), .ZN(n5050)
         );
  OAI21_X1 U5391 ( .B1(n5204), .B2(n5046), .A(n5050), .ZN(n5043) );
  INV_X1 U5392 ( .A(n5043), .ZN(n5045) );
  AOI22_X1 U5393 ( .A1(n5256), .A2(n5045), .B1(n3999), .B2(n5254), .ZN(U3520)
         );
  AOI22_X1 U5394 ( .A1(n5259), .A2(n5045), .B1(n5044), .B2(n5257), .ZN(U3471)
         );
  INV_X1 U5395 ( .A(n5046), .ZN(n5047) );
  AOI22_X1 U5396 ( .A1(n5247), .A2(n5047), .B1(REG3_REG_2__SCAN_IN), .B2(n5135), .ZN(n5048) );
  OAI221_X1 U5397 ( .B1(n5249), .B2(n5050), .C1(n5140), .C2(n5049), .A(n5048), 
        .ZN(U3288) );
  AOI22_X1 U5398 ( .A1(STATE_REG_SCAN_IN), .A2(n4029), .B1(n5051), .B2(U3149), 
        .ZN(U3349) );
  NOR2_X1 U5399 ( .A1(n5053), .A2(n5052), .ZN(n5054) );
  AOI22_X1 U5400 ( .A1(n5256), .A2(n5054), .B1(n2863), .B2(n5254), .ZN(U3521)
         );
  AOI22_X1 U5401 ( .A1(n5259), .A2(n5054), .B1(n4741), .B2(n5257), .ZN(U3473)
         );
  NOR2_X1 U5402 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  AOI22_X1 U5403 ( .A1(n5256), .A2(n5057), .B1(n2875), .B2(n5254), .ZN(U3522)
         );
  AOI22_X1 U5404 ( .A1(n5259), .A2(n5057), .B1(n4742), .B2(n5257), .ZN(U3475)
         );
  INV_X1 U5405 ( .A(DATAI_5_), .ZN(n5058) );
  AOI22_X1 U5406 ( .A1(STATE_REG_SCAN_IN), .A2(n5059), .B1(n5058), .B2(U3149), 
        .ZN(U3347) );
  NOR2_X1 U5407 ( .A1(n5060), .A2(n5144), .ZN(n5061) );
  AOI211_X1 U5408 ( .C1(n5252), .C2(n5063), .A(n5062), .B(n5061), .ZN(n5066)
         );
  AOI22_X1 U5409 ( .A1(n5256), .A2(n5066), .B1(n5064), .B2(n5254), .ZN(U3523)
         );
  AOI22_X1 U5410 ( .A1(n5259), .A2(n5066), .B1(n5065), .B2(n5257), .ZN(U3477)
         );
  OAI22_X1 U5411 ( .A1(n5068), .A2(n5144), .B1(n5204), .B2(n5067), .ZN(n5070)
         );
  NOR2_X1 U5412 ( .A1(n5070), .A2(n5069), .ZN(n5073) );
  INV_X1 U5413 ( .A(REG1_REG_6__SCAN_IN), .ZN(n5071) );
  AOI22_X1 U5414 ( .A1(n5256), .A2(n5073), .B1(n5071), .B2(n5254), .ZN(U3524)
         );
  AOI22_X1 U5415 ( .A1(n5259), .A2(n5073), .B1(n5072), .B2(n5257), .ZN(U3479)
         );
  AOI211_X1 U5416 ( .C1(n5076), .C2(n5227), .A(n5075), .B(n5074), .ZN(n5079)
         );
  INV_X1 U5417 ( .A(REG1_REG_7__SCAN_IN), .ZN(n5077) );
  AOI22_X1 U5418 ( .A1(n5256), .A2(n5079), .B1(n5077), .B2(n5254), .ZN(U3525)
         );
  AOI22_X1 U5419 ( .A1(n5259), .A2(n5079), .B1(n5078), .B2(n5257), .ZN(U3481)
         );
  NOR2_X1 U5420 ( .A1(n5081), .A2(n5080), .ZN(n5083) );
  AOI22_X1 U5421 ( .A1(n5256), .A2(n5083), .B1(n2783), .B2(n5254), .ZN(U3526)
         );
  INV_X1 U5422 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U5423 ( .A1(n5259), .A2(n5083), .B1(n5082), .B2(n5257), .ZN(U3483)
         );
  AOI22_X1 U5424 ( .A1(STATE_REG_SCAN_IN), .A2(n5085), .B1(n5084), .B2(U3149), 
        .ZN(U3343) );
  OAI21_X1 U5425 ( .B1(n5204), .B2(n5087), .A(n5086), .ZN(n5088) );
  AOI21_X1 U5426 ( .B1(n5227), .B2(n5089), .A(n5088), .ZN(n5091) );
  AOI22_X1 U5427 ( .A1(n5256), .A2(n5091), .B1(n3996), .B2(n5254), .ZN(U3527)
         );
  INV_X1 U5428 ( .A(REG0_REG_9__SCAN_IN), .ZN(n5090) );
  AOI22_X1 U5429 ( .A1(n5259), .A2(n5091), .B1(n5090), .B2(n5257), .ZN(U3485)
         );
  OR2_X1 U5430 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  AND2_X1 U5431 ( .A1(n5114), .A2(n5094), .ZN(n5107) );
  XNOR2_X1 U5432 ( .A(n5095), .B(n5096), .ZN(n5105) );
  INV_X1 U5433 ( .A(n5096), .ZN(n5098) );
  OAI211_X1 U5434 ( .C1(n2529), .C2(n5098), .A(n5227), .B(n5097), .ZN(n5104)
         );
  OAI22_X1 U5435 ( .A1(n5100), .A2(n5212), .B1(n5099), .B2(n5210), .ZN(n5101)
         );
  AOI21_X1 U5436 ( .B1(n5102), .B2(n5240), .A(n5101), .ZN(n5103) );
  OAI211_X1 U5437 ( .C1(n5217), .C2(n5105), .A(n5104), .B(n5103), .ZN(n5108)
         );
  AOI21_X1 U5438 ( .B1(n5252), .B2(n5107), .A(n5108), .ZN(n5106) );
  AOI22_X1 U5439 ( .A1(n5256), .A2(n5106), .B1(n2936), .B2(n5254), .ZN(U3528)
         );
  AOI22_X1 U5440 ( .A1(n5259), .A2(n5106), .B1(n2940), .B2(n5257), .ZN(U3487)
         );
  AOI22_X1 U5441 ( .A1(n5107), .A2(n5247), .B1(REG2_REG_10__SCAN_IN), .B2(
        n5249), .ZN(n5110) );
  NAND2_X1 U5442 ( .A1(n5140), .A2(n5108), .ZN(n5109) );
  OAI211_X1 U5443 ( .C1(n5224), .C2(n5111), .A(n5110), .B(n5109), .ZN(U3280)
         );
  INV_X1 U5444 ( .A(n5112), .ZN(n5113) );
  AOI21_X1 U5445 ( .B1(n5115), .B2(n5114), .A(n5113), .ZN(n5137) );
  INV_X1 U5446 ( .A(n5116), .ZN(n5131) );
  AOI22_X1 U5447 ( .A1(n5120), .A2(n5119), .B1(n5118), .B2(n5117), .ZN(n5121)
         );
  OAI21_X1 U5448 ( .B1(n5123), .B2(n5122), .A(n5121), .ZN(n5130) );
  INV_X1 U5449 ( .A(n5125), .ZN(n5124) );
  NOR2_X1 U5450 ( .A1(n5124), .A2(n5217), .ZN(n5128) );
  OAI22_X1 U5451 ( .A1(n2503), .A2(n5144), .B1(n5217), .B2(n5125), .ZN(n5127)
         );
  MUX2_X1 U5452 ( .A(n5128), .B(n5127), .S(n5126), .Z(n5129) );
  AOI211_X1 U5453 ( .C1(n5131), .C2(n5227), .A(n5130), .B(n5129), .ZN(n5141)
         );
  INV_X1 U5454 ( .A(n5141), .ZN(n5132) );
  AOI21_X1 U5455 ( .B1(n5252), .B2(n5137), .A(n5132), .ZN(n5134) );
  AOI22_X1 U5456 ( .A1(n5256), .A2(n5134), .B1(n3994), .B2(n5254), .ZN(U3529)
         );
  INV_X1 U5457 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5133) );
  AOI22_X1 U5458 ( .A1(n5259), .A2(n5134), .B1(n5133), .B2(n5257), .ZN(U3489)
         );
  AOI22_X1 U5459 ( .A1(n5137), .A2(n5247), .B1(n5136), .B2(n5135), .ZN(n5138)
         );
  OAI221_X1 U5460 ( .B1(n5249), .B2(n5141), .C1(n5140), .C2(n5139), .A(n5138), 
        .ZN(U3279) );
  INV_X1 U5461 ( .A(DATAI_12_), .ZN(n5142) );
  AOI22_X1 U5462 ( .A1(STATE_REG_SCAN_IN), .A2(n5143), .B1(n5142), .B2(U3149), 
        .ZN(U3340) );
  NOR2_X1 U5463 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  AOI211_X1 U5464 ( .C1(n5252), .C2(n5148), .A(n5147), .B(n5146), .ZN(n5151)
         );
  INV_X1 U5465 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5149) );
  AOI22_X1 U5466 ( .A1(n5256), .A2(n5151), .B1(n5149), .B2(n5254), .ZN(U3530)
         );
  INV_X1 U5467 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5150) );
  AOI22_X1 U5468 ( .A1(n5259), .A2(n5151), .B1(n5150), .B2(n5257), .ZN(U3491)
         );
  AOI211_X1 U5469 ( .C1(n5227), .C2(n5154), .A(n5153), .B(n5152), .ZN(n5155)
         );
  AOI22_X1 U5470 ( .A1(n5256), .A2(n5155), .B1(n4014), .B2(n5254), .ZN(U3531)
         );
  AOI22_X1 U5471 ( .A1(n5259), .A2(n5155), .B1(n2975), .B2(n5257), .ZN(U3493)
         );
  OAI22_X1 U5472 ( .A1(n5254), .A2(n5156), .B1(REG1_REG_14__SCAN_IN), .B2(
        n5256), .ZN(n5157) );
  INV_X1 U5473 ( .A(n5157), .ZN(U3532) );
  NAND2_X1 U5474 ( .A1(n5159), .A2(n5158), .ZN(n5168) );
  NAND2_X1 U5475 ( .A1(n5161), .A2(n5160), .ZN(n5167) );
  NAND2_X1 U5476 ( .A1(n5163), .A2(n5162), .ZN(n5166) );
  INV_X1 U5477 ( .A(n5164), .ZN(n5165) );
  AND4_X1 U5478 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n5175)
         );
  NAND2_X1 U5479 ( .A1(n3729), .A2(n5169), .ZN(n5171) );
  XNOR2_X1 U5480 ( .A(n5171), .B(n5170), .ZN(n5173) );
  NAND2_X1 U5481 ( .A1(n5173), .A2(n5172), .ZN(n5174) );
  OAI211_X1 U5482 ( .C1(n5177), .C2(n5176), .A(n5175), .B(n5174), .ZN(U3238)
         );
  NOR2_X1 U5483 ( .A1(n5178), .A2(n5204), .ZN(n5180) );
  AOI211_X1 U5484 ( .C1(n5181), .C2(n5227), .A(n5180), .B(n5179), .ZN(n5184)
         );
  INV_X1 U5485 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5182) );
  AOI22_X1 U5486 ( .A1(n5256), .A2(n5184), .B1(n5182), .B2(n5254), .ZN(U3533)
         );
  INV_X1 U5487 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5183) );
  AOI22_X1 U5488 ( .A1(n5259), .A2(n5184), .B1(n5183), .B2(n5257), .ZN(U3497)
         );
  AOI211_X1 U5489 ( .C1(n5187), .C2(n5227), .A(n5186), .B(n5185), .ZN(n5190)
         );
  INV_X1 U5490 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5188) );
  AOI22_X1 U5491 ( .A1(n5256), .A2(n5190), .B1(n5188), .B2(n5254), .ZN(U3534)
         );
  INV_X1 U5492 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5189) );
  AOI22_X1 U5493 ( .A1(n5259), .A2(n5190), .B1(n5189), .B2(n5257), .ZN(U3499)
         );
  AOI211_X1 U5494 ( .C1(n5193), .C2(n5227), .A(n5192), .B(n5191), .ZN(n5195)
         );
  AOI22_X1 U5495 ( .A1(n5256), .A2(n5195), .B1(n4061), .B2(n5254), .ZN(U3535)
         );
  INV_X1 U5496 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5194) );
  AOI22_X1 U5497 ( .A1(n5259), .A2(n5195), .B1(n5194), .B2(n5257), .ZN(U3501)
         );
  NOR2_X1 U5498 ( .A1(n5197), .A2(n5196), .ZN(n5199) );
  INV_X1 U5499 ( .A(REG1_REG_18__SCAN_IN), .ZN(n5198) );
  AOI22_X1 U5500 ( .A1(n5256), .A2(n5199), .B1(n5198), .B2(n5254), .ZN(U3536)
         );
  AOI22_X1 U5501 ( .A1(n5259), .A2(n5199), .B1(n3043), .B2(n5257), .ZN(U3503)
         );
  XNOR2_X1 U5502 ( .A(n5200), .B(n5209), .ZN(n5228) );
  AOI22_X1 U5503 ( .A1(n5228), .A2(n5201), .B1(REG2_REG_19__SCAN_IN), .B2(
        n5249), .ZN(n5222) );
  INV_X1 U5504 ( .A(n5202), .ZN(n5203) );
  AOI211_X1 U5505 ( .C1(n5215), .C2(n5205), .A(n5204), .B(n5203), .ZN(n5226)
         );
  NAND2_X1 U5506 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  XOR2_X1 U5507 ( .A(n5209), .B(n5208), .Z(n5218) );
  OAI22_X1 U5508 ( .A1(n5213), .A2(n5212), .B1(n5211), .B2(n5210), .ZN(n5214)
         );
  AOI21_X1 U5509 ( .B1(n5215), .B2(n5240), .A(n5214), .ZN(n5216) );
  OAI21_X1 U5510 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n5225) );
  AOI21_X1 U5511 ( .B1(n5226), .B2(n5219), .A(n5225), .ZN(n5220) );
  OR2_X1 U5512 ( .A1(n5220), .A2(n5249), .ZN(n5221) );
  OAI211_X1 U5513 ( .C1(n5224), .C2(n5223), .A(n5222), .B(n5221), .ZN(U3271)
         );
  AOI211_X1 U5514 ( .C1(n5228), .C2(n5227), .A(n5226), .B(n5225), .ZN(n5229)
         );
  AOI22_X1 U5515 ( .A1(n5256), .A2(n5229), .B1(n3054), .B2(n5254), .ZN(U3537)
         );
  AOI22_X1 U5516 ( .A1(n5259), .A2(n5229), .B1(n3058), .B2(n5257), .ZN(U3505)
         );
  INV_X1 U5517 ( .A(n5233), .ZN(n5243) );
  NAND2_X1 U5518 ( .A1(n5240), .A2(n5243), .ZN(n5232) );
  NAND2_X1 U5519 ( .A1(n5231), .A2(n5230), .ZN(n5241) );
  AND2_X1 U5520 ( .A1(n5232), .A2(n5241), .ZN(n5235) );
  XNOR2_X1 U5521 ( .A(n5244), .B(n5233), .ZN(n5237) );
  AOI22_X1 U5522 ( .A1(n5237), .A2(n5247), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5249), .ZN(n5234) );
  OAI21_X1 U5523 ( .B1(n5249), .B2(n5235), .A(n5234), .ZN(U3261) );
  INV_X1 U5524 ( .A(n5235), .ZN(n5236) );
  AOI21_X1 U5525 ( .B1(n5237), .B2(n5252), .A(n5236), .ZN(n5239) );
  INV_X1 U5526 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5238) );
  AOI22_X1 U5527 ( .A1(n5256), .A2(n5239), .B1(n5238), .B2(n5254), .ZN(U3548)
         );
  AOI22_X1 U5528 ( .A1(n5259), .A2(n5239), .B1(n3610), .B2(n5257), .ZN(U3516)
         );
  NAND2_X1 U5529 ( .A1(n5240), .A2(n5245), .ZN(n5242) );
  AND2_X1 U5530 ( .A1(n5242), .A2(n5241), .ZN(n5250) );
  NOR2_X1 U5531 ( .A1(n5244), .A2(n5243), .ZN(n5246) );
  XNOR2_X1 U5532 ( .A(n5246), .B(n5245), .ZN(n5253) );
  AOI22_X1 U5533 ( .A1(n5253), .A2(n5247), .B1(n5249), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5248) );
  OAI21_X1 U5534 ( .B1(n5249), .B2(n5250), .A(n5248), .ZN(U3260) );
  INV_X1 U5535 ( .A(n5250), .ZN(n5251) );
  AOI21_X1 U5536 ( .B1(n5253), .B2(n5252), .A(n5251), .ZN(n5258) );
  INV_X1 U5537 ( .A(REG1_REG_31__SCAN_IN), .ZN(n5255) );
  AOI22_X1 U5538 ( .A1(n5256), .A2(n5258), .B1(n5255), .B2(n5254), .ZN(U3549)
         );
  AOI22_X1 U5539 ( .A1(n5259), .A2(n5258), .B1(n3821), .B2(n5257), .ZN(U3517)
         );
  CLKBUF_X1 U2593 ( .A(n2840), .Z(n3822) );
  CLKBUF_X1 U2935 ( .A(n3111), .Z(n5252) );
endmodule

