

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11151, n11152, n11154, n11155, n11156, n11157, n11159, n11161,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22598, n22599, n22600, n22601;

  AND2_X1 U11258 ( .A1(n13667), .A2(n13666), .ZN(n13715) );
  INV_X1 U11260 ( .A(n20864), .ZN(n21065) );
  NOR2_X1 U11261 ( .A1(n13015), .A2(n11699), .ZN(n13017) );
  XNOR2_X1 U11262 ( .A(n12477), .B(n21909), .ZN(n14331) );
  AND2_X1 U11263 ( .A1(n12903), .A2(n12890), .ZN(n12983) );
  AND2_X1 U11264 ( .A1(n12907), .A2(n12890), .ZN(n15644) );
  NAND2_X1 U11265 ( .A1(n11991), .A2(n11990), .ZN(n15118) );
  BUF_X1 U11266 ( .A(n14387), .Z(n18071) );
  AND2_X1 U11267 ( .A1(n15926), .A2(n12761), .ZN(n16061) );
  AND2_X1 U11268 ( .A1(n12727), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12952) );
  AND2_X1 U11269 ( .A1(n15926), .A2(n14282), .ZN(n16060) );
  AND2_X1 U11270 ( .A1(n16135), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12772) );
  AND2_X1 U11271 ( .A1(n15953), .A2(n14603), .ZN(n16059) );
  CLKBUF_X2 U11272 ( .A(n12078), .Z(n11182) );
  INV_X1 U11273 ( .A(n15925), .ZN(n12754) );
  CLKBUF_X2 U11274 ( .A(n12108), .Z(n13698) );
  CLKBUF_X2 U11275 ( .A(n11883), .Z(n11183) );
  CLKBUF_X2 U11276 ( .A(n11869), .Z(n11184) );
  INV_X1 U11277 ( .A(n12390), .ZN(n11902) );
  CLKBUF_X2 U11278 ( .A(n11803), .Z(n12394) );
  INV_X2 U11279 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n15635) );
  CLKBUF_X2 U11280 ( .A(n13189), .Z(n19060) );
  NOR2_X1 U11281 ( .A1(n12809), .A2(n12743), .ZN(n12806) );
  CLKBUF_X1 U11282 ( .A(n14440), .Z(n18095) );
  INV_X1 U11283 ( .A(n14351), .ZN(n18149) );
  CLKBUF_X1 U11284 ( .A(n14396), .Z(n11168) );
  INV_X1 U11285 ( .A(n12740), .ZN(n13188) );
  INV_X1 U11286 ( .A(n11214), .ZN(n18127) );
  CLKBUF_X2 U11287 ( .A(n14440), .Z(n18128) );
  OR2_X1 U11288 ( .A1(n15905), .A2(n20676), .ZN(n17909) );
  NOR2_X2 U11289 ( .A1(n20676), .A2(n14337), .ZN(n14455) );
  INV_X1 U11290 ( .A(n11860), .ZN(n11836) );
  INV_X2 U11291 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21310) );
  AND4_X1 U11292 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11746) );
  AND4_X1 U11293 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n11747) );
  CLKBUF_X2 U11294 ( .A(n12237), .Z(n12333) );
  AND2_X1 U11295 ( .A1(n11720), .A2(n11719), .ZN(n11803) );
  AND2_X1 U11296 ( .A1(n11720), .A2(n16830), .ZN(n11883) );
  AND2_X1 U11297 ( .A1(n11712), .A2(n13935), .ZN(n12053) );
  AND2_X1 U11298 ( .A1(n11711), .A2(n11712), .ZN(n11954) );
  AND2_X1 U11299 ( .A1(n11712), .A2(n14191), .ZN(n11949) );
  AND2_X2 U11300 ( .A1(n11711), .A2(n11718), .ZN(n12108) );
  AND2_X1 U11301 ( .A1(n11702), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11720) );
  CLKBUF_X1 U11302 ( .A(n20180), .Z(n11151) );
  NOR3_X1 U11303 ( .A1(n15753), .A2(n22169), .A3(n19799), .ZN(n20180) );
  CLKBUF_X1 U11304 ( .A(n22475), .Z(n11152) );
  NOR2_X1 U11305 ( .A1(n16270), .A2(n20496), .ZN(n22475) );
  INV_X1 U11307 ( .A(n22599), .ZN(n11154) );
  INV_X1 U11309 ( .A(n17493), .ZN(n11155) );
  INV_X1 U11310 ( .A(n11155), .ZN(n11156) );
  INV_X1 U11311 ( .A(n11155), .ZN(n11157) );
  INV_X1 U11313 ( .A(n22598), .ZN(n11159) );
  INV_X1 U11315 ( .A(n22601), .ZN(n11161) );
  INV_X1 U11317 ( .A(n22600), .ZN(n11163) );
  AND2_X1 U11318 ( .A1(n11712), .A2(n11720), .ZN(n11869) );
  INV_X1 U11319 ( .A(n12520), .ZN(n16779) );
  AND4_X1 U11320 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11727) );
  NAND2_X2 U11321 ( .A1(n21296), .A2(n21310), .ZN(n20676) );
  NOR2_X1 U11322 ( .A1(n15325), .A2(n15444), .ZN(n15442) );
  AND4_X2 U11324 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11838) );
  BUF_X1 U11325 ( .A(n12872), .Z(n13112) );
  NAND2_X1 U11326 ( .A1(n16922), .A2(n11612), .ZN(n16090) );
  OR2_X1 U11327 ( .A1(n13619), .A2(n13618), .ZN(n17106) );
  NOR2_X1 U11328 ( .A1(n18356), .A2(n21658), .ZN(n18361) );
  INV_X1 U11329 ( .A(n18106), .ZN(n20700) );
  OR2_X1 U11330 ( .A1(n16975), .A2(n13645), .ZN(n13719) );
  AND2_X1 U11331 ( .A1(n13719), .A2(n13646), .ZN(n19015) );
  AND2_X1 U11332 ( .A1(n16992), .A2(n16981), .ZN(n16983) );
  NAND4_X1 U11333 ( .A1(n21262), .A2(P3_EAX_REG_10__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n21158), .ZN(n21258) );
  INV_X1 U11334 ( .A(n18607), .ZN(n18619) );
  NAND2_X1 U11335 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21294) );
  INV_X1 U11336 ( .A(n22110), .ZN(n22128) );
  INV_X2 U11337 ( .A(n17750), .ZN(n22203) );
  INV_X1 U11338 ( .A(n18446), .ZN(n18397) );
  NAND2_X1 U11339 ( .A1(n21835), .A2(n21341), .ZN(n18623) );
  NOR4_X1 U11340 ( .A1(n21649), .A2(n21730), .A3(n21648), .A4(n21647), .ZN(
        n21654) );
  AND4_X1 U11341 ( .A1(n11807), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(
        n11164) );
  NAND3_X2 U11342 ( .A1(n12975), .A2(n12974), .A3(n13222), .ZN(n11347) );
  INV_X1 U11343 ( .A(n11661), .ZN(n12872) );
  AND2_X1 U11345 ( .A1(n11838), .A2(n11832), .ZN(n13823) );
  OR2_X4 U11346 ( .A1(n12830), .A2(n11402), .ZN(n13180) );
  NAND2_X2 U11347 ( .A1(n11434), .A2(n12862), .ZN(n12880) );
  NAND2_X2 U11348 ( .A1(n11327), .A2(n12843), .ZN(n11434) );
  NAND2_X1 U11349 ( .A1(n12745), .A2(n20069), .ZN(n12832) );
  NAND2_X2 U11350 ( .A1(n12888), .A2(n12889), .ZN(n11327) );
  NAND2_X4 U11351 ( .A1(n12687), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16124) );
  AOI22_X2 U11352 ( .A1(n13180), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12877), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12821) );
  NOR2_X2 U11353 ( .A1(n13655), .A2(n13653), .ZN(n13744) );
  AOI21_X2 U11354 ( .B1(n11673), .B2(n13593), .A(n17049), .ZN(n13655) );
  INV_X2 U11355 ( .A(n13112), .ZN(n11165) );
  NAND2_X1 U11356 ( .A1(n11428), .A2(n12859), .ZN(n11661) );
  XNOR2_X2 U11357 ( .A(n21275), .B(n21390), .ZN(n18611) );
  NOR2_X4 U11358 ( .A1(n13423), .A2(n13419), .ZN(n13451) );
  AND2_X2 U11359 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12687) );
  NOR2_X2 U11360 ( .A1(n12738), .A2(n12826), .ZN(n12820) );
  NAND2_X2 U11361 ( .A1(n12676), .A2(n12675), .ZN(n13381) );
  INV_X2 U11364 ( .A(n21351), .ZN(n17448) );
  AOI211_X1 U11365 ( .C1(n14569), .C2(n22256), .A(n15378), .B(n15348), .ZN(
        n15121) );
  MUX2_X2 U11366 ( .A(n12625), .B(n12624), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13189) );
  AND2_X4 U11367 ( .A1(n12761), .A2(n17422), .ZN(n16134) );
  NAND2_X2 U11368 ( .A1(n15215), .A2(n13192), .ZN(n13722) );
  BUF_X2 U11369 ( .A(n16007), .Z(n11166) );
  BUF_X4 U11370 ( .A(n16007), .Z(n11167) );
  NOR2_X1 U11371 ( .A1(n14341), .A2(n14340), .ZN(n14396) );
  NAND2_X1 U11372 ( .A1(n17636), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19107) );
  AND2_X1 U11373 ( .A1(n13080), .A2(n11308), .ZN(n17099) );
  NOR2_X1 U11374 ( .A1(n13719), .A2(n13718), .ZN(n13724) );
  NAND2_X1 U11375 ( .A1(n18340), .A2(n18224), .ZN(n18282) );
  AND2_X1 U11376 ( .A1(n17000), .A2(n16990), .ZN(n16992) );
  NOR2_X1 U11377 ( .A1(n18267), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18235) );
  NAND2_X1 U11378 ( .A1(n18494), .A2(n11296), .ZN(n18267) );
  AND2_X1 U11379 ( .A1(n13532), .A2(n17585), .ZN(n11674) );
  NOR3_X2 U11380 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18607), .A3(n20664), 
        .ZN(n18446) );
  CLKBUF_X1 U11381 ( .A(n12990), .Z(n19777) );
  CLKBUF_X1 U11382 ( .A(n12981), .Z(n19798) );
  NOR2_X2 U11383 ( .A1(n12905), .A2(n12904), .ZN(n12993) );
  NAND2_X1 U11384 ( .A1(n13214), .A2(n13213), .ZN(n11635) );
  CLKBUF_X2 U11385 ( .A(n20652), .Z(n20661) );
  NAND3_X1 U11386 ( .A1(n14296), .A2(n12828), .A3(n11690), .ZN(n14606) );
  AND2_X1 U11387 ( .A1(n13380), .A2(n12814), .ZN(n15204) );
  INV_X4 U11388 ( .A(n13479), .ZN(n13448) );
  INV_X2 U11389 ( .A(n21338), .ZN(n21342) );
  NAND4_X1 U11390 ( .A1(n15212), .A2(n13188), .A3(n15649), .A4(n19967), .ZN(
        n12831) );
  INV_X2 U11391 ( .A(n15294), .ZN(n11828) );
  CLKBUF_X2 U11393 ( .A(n12053), .Z(n12282) );
  CLKBUF_X2 U11394 ( .A(n11949), .Z(n13691) );
  BUF_X2 U11395 ( .A(n11954), .Z(n12307) );
  CLKBUF_X2 U11396 ( .A(n14388), .Z(n18116) );
  CLKBUF_X2 U11397 ( .A(n11864), .Z(n13692) );
  CLKBUF_X2 U11398 ( .A(n20376), .Z(n21841) );
  BUF_X2 U11399 ( .A(n12656), .Z(n12726) );
  INV_X2 U11400 ( .A(n11214), .ZN(n11169) );
  AND2_X2 U11401 ( .A1(n13935), .A2(n16830), .ZN(n12030) );
  INV_X4 U11402 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21772) );
  INV_X1 U11403 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14603) );
  NOR2_X1 U11404 ( .A1(n17264), .A2(n17107), .ZN(n17111) );
  OR3_X1 U11405 ( .A1(n17264), .A2(n17263), .A3(n17608), .ZN(n11682) );
  AND2_X1 U11406 ( .A1(n13621), .A2(n17274), .ZN(n17263) );
  NOR2_X1 U11407 ( .A1(n13621), .A2(n17274), .ZN(n17264) );
  NAND2_X1 U11408 ( .A1(n17106), .A2(n13620), .ZN(n13621) );
  OR2_X1 U11409 ( .A1(n16278), .A2(n20496), .ZN(n13714) );
  NOR2_X1 U11410 ( .A1(n17075), .A2(n17191), .ZN(n17072) );
  NAND2_X1 U11411 ( .A1(n13081), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17086) );
  OAI21_X1 U11412 ( .B1(n16912), .B2(n11617), .A(n11615), .ZN(n11614) );
  NAND2_X1 U11413 ( .A1(n11343), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17621) );
  INV_X1 U11414 ( .A(n17216), .ZN(n13081) );
  AOI221_X1 U11415 ( .B1(n19108), .B2(n19107), .C1(n19106), .C2(n19107), .A(
        n19105), .ZN(n19127) );
  INV_X1 U11416 ( .A(n11616), .ZN(n11615) );
  AND2_X1 U11417 ( .A1(n16091), .A2(n11617), .ZN(n11613) );
  OAI21_X2 U11418 ( .B1(n16634), .B2(n11424), .A(n16779), .ZN(n16604) );
  NAND2_X1 U11419 ( .A1(n11678), .A2(n13078), .ZN(n17579) );
  OR2_X1 U11420 ( .A1(n17132), .A2(n17131), .ZN(n17333) );
  NAND3_X1 U11421 ( .A1(n11565), .A2(n20516), .A3(n11324), .ZN(n16603) );
  NAND2_X1 U11422 ( .A1(n11566), .A2(n12537), .ZN(n16634) );
  AND2_X1 U11423 ( .A1(n13650), .A2(n13649), .ZN(n13651) );
  NAND2_X1 U11424 ( .A1(n17584), .A2(n11674), .ZN(n13559) );
  OAI21_X1 U11425 ( .B1(n11194), .B2(n11681), .A(n17265), .ZN(n11680) );
  NAND2_X1 U11426 ( .A1(n17166), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17152) );
  CLKBUF_X1 U11427 ( .A(n16939), .Z(n16946) );
  NAND2_X1 U11428 ( .A1(n11398), .A2(n13057), .ZN(n17166) );
  AND2_X1 U11429 ( .A1(n11221), .A2(n17568), .ZN(n11194) );
  AND2_X1 U11430 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  INV_X1 U11431 ( .A(n13056), .ZN(n13057) );
  OAI21_X1 U11432 ( .B1(n13055), .B2(n13058), .A(n13054), .ZN(n13056) );
  NAND2_X1 U11433 ( .A1(n18352), .A2(n18356), .ZN(n18351) );
  INV_X1 U11434 ( .A(n19015), .ZN(n16247) );
  XNOR2_X1 U11435 ( .A(n13719), .B(n13718), .ZN(n19034) );
  AND2_X1 U11436 ( .A1(n13053), .A2(n13051), .ZN(n11396) );
  XNOR2_X1 U11437 ( .A(n13076), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17568) );
  OR2_X1 U11438 ( .A1(n12533), .A2(n11568), .ZN(n11567) );
  NAND2_X1 U11439 ( .A1(n20475), .A2(n12495), .ZN(n20483) );
  NAND2_X1 U11440 ( .A1(n18416), .A2(n18456), .ZN(n18340) );
  NAND2_X1 U11441 ( .A1(n15508), .A2(n12979), .ZN(n13053) );
  INV_X1 U11442 ( .A(n21215), .ZN(n21211) );
  OR2_X1 U11443 ( .A1(n16983), .A2(n16982), .ZN(n18995) );
  OAI21_X1 U11444 ( .B1(n11423), .B2(n12514), .A(n12526), .ZN(n11421) );
  NOR2_X1 U11445 ( .A1(n15106), .A2(n15107), .ZN(n14671) );
  NAND2_X1 U11446 ( .A1(n18475), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n21520) );
  OAI211_X1 U11447 ( .C1(n12536), .C2(n20516), .A(n16650), .B(n16639), .ZN(
        n11568) );
  OR2_X1 U11448 ( .A1(n16778), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16781) );
  AND2_X1 U11449 ( .A1(n16665), .A2(n16662), .ZN(n16650) );
  AND2_X1 U11450 ( .A1(n12535), .A2(n16653), .ZN(n16639) );
  AND2_X1 U11451 ( .A1(n17016), .A2(n11642), .ZN(n17000) );
  OR2_X1 U11452 ( .A1(n12506), .A2(n12516), .ZN(n12512) );
  OR2_X1 U11453 ( .A1(n12487), .A2(n12516), .ZN(n12493) );
  NAND2_X1 U11454 ( .A1(n18211), .A2(n18523), .ZN(n21472) );
  NAND2_X1 U11455 ( .A1(n12519), .A2(n12518), .ZN(n12520) );
  NAND2_X1 U11456 ( .A1(n21255), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21244) );
  XNOR2_X1 U11457 ( .A(n12519), .B(n12069), .ZN(n12505) );
  NAND2_X1 U11458 ( .A1(n13046), .A2(n13045), .ZN(n13048) );
  NAND2_X1 U11459 ( .A1(n12038), .A2(n11410), .ZN(n12519) );
  AND4_X1 U11460 ( .A1(n13553), .A2(n13552), .A3(n17108), .A4(n17122), .ZN(
        n13558) );
  OR2_X1 U11461 ( .A1(n13033), .A2(n13032), .ZN(n13046) );
  AND2_X1 U11462 ( .A1(n17278), .A2(n17277), .ZN(n17280) );
  INV_X1 U11463 ( .A(n18549), .ZN(n18624) );
  NOR2_X1 U11464 ( .A1(n17315), .A2(n11637), .ZN(n17278) );
  OAI211_X1 U11465 ( .C1(n19824), .C2(n12919), .A(n12918), .B(n19060), .ZN(
        n12920) );
  NAND2_X1 U11466 ( .A1(n18829), .A2(n17313), .ZN(n17315) );
  NOR2_X1 U11467 ( .A1(n18544), .A2(n21456), .ZN(n18206) );
  NAND2_X1 U11468 ( .A1(n11932), .A2(n11918), .ZN(n16820) );
  AND2_X1 U11469 ( .A1(n18791), .A2(n11269), .ZN(n18829) );
  NAND2_X1 U11470 ( .A1(n18538), .A2(n18176), .ZN(n18526) );
  INV_X1 U11471 ( .A(n12002), .ZN(n11412) );
  NAND2_X1 U11472 ( .A1(n14036), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14169) );
  NAND2_X1 U11473 ( .A1(n21809), .A2(n20667), .ZN(n20811) );
  NAND2_X1 U11474 ( .A1(n18539), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18538) );
  NOR2_X2 U11475 ( .A1(n18792), .A2(n18793), .ZN(n18791) );
  OR2_X1 U11476 ( .A1(n13576), .A2(n13574), .ZN(n13579) );
  AND2_X1 U11477 ( .A1(n15118), .A2(n12025), .ZN(n11411) );
  AND2_X1 U11478 ( .A1(n13510), .A2(n13509), .ZN(n17629) );
  AOI22_X1 U11479 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12993), .B1(
        n12994), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12908) );
  AND2_X1 U11480 ( .A1(n14205), .A2(n14157), .ZN(n14162) );
  XNOR2_X1 U11481 ( .A(n18232), .B(n11607), .ZN(n18539) );
  NAND2_X1 U11482 ( .A1(n14161), .A2(n14160), .ZN(n14212) );
  AND2_X1 U11483 ( .A1(n14254), .A2(n14131), .ZN(n12903) );
  NAND2_X1 U11484 ( .A1(n17391), .A2(n11653), .ZN(n18792) );
  NOR2_X2 U11485 ( .A1(n12905), .A2(n12900), .ZN(n12992) );
  INV_X1 U11486 ( .A(n12900), .ZN(n12890) );
  NOR2_X2 U11487 ( .A1(n21777), .A2(n20609), .ZN(n20670) );
  NOR2_X1 U11488 ( .A1(n21269), .A2(n21270), .ZN(n21153) );
  NOR2_X1 U11489 ( .A1(n21105), .A2(n21269), .ZN(n21278) );
  NAND2_X1 U11490 ( .A1(n15419), .A2(n22153), .ZN(n11991) );
  NOR2_X2 U11491 ( .A1(n21732), .A2(n21754), .ZN(n21613) );
  CLKBUF_X1 U11492 ( .A(n16273), .Z(n16543) );
  NAND2_X1 U11493 ( .A1(n11367), .A2(n11370), .ZN(n11931) );
  OAI21_X1 U11494 ( .B1(n21104), .B2(n21103), .A(n21832), .ZN(n21269) );
  AND2_X1 U11495 ( .A1(n11946), .A2(n11973), .ZN(n11947) );
  OR2_X1 U11496 ( .A1(n14605), .A2(n19069), .ZN(n12900) );
  OR2_X1 U11497 ( .A1(n11945), .A2(n11944), .ZN(n11946) );
  NAND2_X1 U11498 ( .A1(n12885), .A2(n12887), .ZN(n14605) );
  NAND2_X2 U11499 ( .A1(n16523), .A2(n14100), .ZN(n16553) );
  XNOR2_X1 U11500 ( .A(n14154), .B(n14155), .ZN(n14207) );
  XNOR2_X1 U11501 ( .A(n11925), .B(n11426), .ZN(n14520) );
  NAND2_X1 U11502 ( .A1(n11323), .A2(n11911), .ZN(n11925) );
  OAI21_X1 U11503 ( .B1(n14615), .B2(n14661), .A(n14104), .ZN(n14154) );
  NOR2_X2 U11504 ( .A1(n19661), .A2(n20174), .ZN(n15675) );
  NOR2_X2 U11505 ( .A1(n20016), .A2(n20174), .ZN(n20017) );
  NOR2_X2 U11506 ( .A1(n19861), .A2(n20174), .ZN(n15648) );
  NOR2_X2 U11507 ( .A1(n19911), .A2(n20174), .ZN(n19912) );
  NAND2_X1 U11508 ( .A1(n21291), .A2(n21311), .ZN(n17474) );
  NAND2_X2 U11509 ( .A1(n16451), .A2(n15092), .ZN(n16425) );
  AND2_X1 U11510 ( .A1(n13504), .A2(n11268), .ZN(n13516) );
  AND2_X1 U11511 ( .A1(n11658), .A2(n12871), .ZN(n12881) );
  NAND2_X1 U11512 ( .A1(n18578), .A2(n18168), .ZN(n18170) );
  NAND2_X1 U11513 ( .A1(n11322), .A2(n11321), .ZN(n11895) );
  NOR2_X1 U11514 ( .A1(n20661), .A2(n20617), .ZN(n20660) );
  NOR2_X2 U11515 ( .A1(n13857), .A2(n16097), .ZN(n13858) );
  AOI21_X1 U11516 ( .B1(n13783), .B2(n13208), .A(n13207), .ZN(n13212) );
  OR2_X1 U11517 ( .A1(n13472), .A2(n13471), .ZN(n13513) );
  NAND2_X2 U11518 ( .A1(n11385), .A2(n12594), .ZN(n15095) );
  NAND2_X1 U11519 ( .A1(n11446), .A2(n12863), .ZN(n12869) );
  INV_X2 U11520 ( .A(n13109), .ZN(n13730) );
  NAND2_X1 U11521 ( .A1(n12813), .A2(n12848), .ZN(n12876) );
  AND2_X1 U11522 ( .A1(n13082), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12836) );
  CLKBUF_X1 U11523 ( .A(n13082), .Z(n13109) );
  AND2_X1 U11524 ( .A1(n12846), .A2(n12845), .ZN(n12854) );
  NAND2_X1 U11525 ( .A1(n18598), .A2(n18165), .ZN(n18166) );
  CLKBUF_X1 U11526 ( .A(n12864), .Z(n13097) );
  AND2_X1 U11527 ( .A1(n15193), .A2(n15192), .ZN(n13204) );
  NOR2_X1 U11528 ( .A1(n13459), .A2(n11471), .ZN(n11470) );
  AND2_X1 U11529 ( .A1(n13815), .A2(n11830), .ZN(n14050) );
  NAND2_X1 U11530 ( .A1(n11344), .A2(n12805), .ZN(n12844) );
  NOR2_X2 U11531 ( .A1(n17639), .A2(n18864), .ZN(n17652) );
  NOR2_X1 U11532 ( .A1(n12829), .A2(n18721), .ZN(n11429) );
  OR2_X1 U11533 ( .A1(n12810), .A2(n12806), .ZN(n13385) );
  AND2_X1 U11534 ( .A1(n15094), .A2(n13823), .ZN(n11312) );
  INV_X2 U11535 ( .A(n21197), .ZN(n21263) );
  NAND2_X1 U11536 ( .A1(n12831), .A2(n12745), .ZN(n12805) );
  NAND2_X1 U11537 ( .A1(n19325), .A2(n17448), .ZN(n17463) );
  OR2_X1 U11538 ( .A1(n11840), .A2(n14098), .ZN(n13820) );
  INV_X1 U11539 ( .A(n12546), .ZN(n12579) );
  OAI21_X1 U11540 ( .B1(n13823), .B2(n14565), .A(n11311), .ZN(n11316) );
  INV_X1 U11541 ( .A(n21160), .ZN(n19325) );
  NAND2_X1 U11542 ( .A1(n11223), .A2(n11522), .ZN(n21160) );
  INV_X2 U11543 ( .A(n15657), .ZN(n16261) );
  NAND3_X1 U11544 ( .A1(n14413), .A2(n14412), .A3(n14411), .ZN(n21338) );
  OR2_X1 U11545 ( .A1(n12785), .A2(n12784), .ZN(n13218) );
  NAND2_X1 U11546 ( .A1(n16097), .A2(n20177), .ZN(n12823) );
  NAND2_X1 U11547 ( .A1(n12549), .A2(n11948), .ZN(n12582) );
  OR2_X1 U11548 ( .A1(n12938), .A2(n12937), .ZN(n13410) );
  NOR2_X1 U11549 ( .A1(n12449), .A2(n13838), .ZN(n14077) );
  AND2_X2 U11550 ( .A1(n14245), .A2(n15294), .ZN(n16206) );
  INV_X1 U11551 ( .A(n11832), .ZN(n14532) );
  INV_X1 U11552 ( .A(n20069), .ZN(n12793) );
  OR2_X1 U11553 ( .A1(n14401), .A2(n11525), .ZN(n11524) );
  OR2_X2 U11554 ( .A1(n11787), .A2(n11786), .ZN(n15092) );
  INV_X2 U11555 ( .A(U212), .ZN(n11170) );
  AND2_X2 U11556 ( .A1(n11701), .A2(n11700), .ZN(n14565) );
  OR2_X2 U11557 ( .A1(n11797), .A2(n11796), .ZN(n12449) );
  AND4_X1 U11558 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11768) );
  NAND2_X2 U11559 ( .A1(U214), .A2(n20531), .ZN(n20597) );
  AND2_X1 U11560 ( .A1(n12626), .A2(n14603), .ZN(n12628) );
  AND2_X1 U11561 ( .A1(n11441), .A2(n11440), .ZN(n12668) );
  AND4_X1 U11562 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11767) );
  AND4_X1 U11563 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11766) );
  AND4_X1 U11564 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11765) );
  AND4_X1 U11565 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11193) );
  AND4_X1 U11566 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11827) );
  AND4_X1 U11567 ( .A1(n11744), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(
        n11745) );
  AND4_X1 U11569 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11825) );
  AND4_X1 U11570 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11824) );
  AND4_X1 U11571 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11728) );
  AND4_X1 U11572 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11726) );
  AND4_X1 U11573 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11748) );
  AND4_X1 U11574 ( .A1(n11724), .A2(n11723), .A3(n11722), .A4(n11721), .ZN(
        n11725) );
  AND3_X1 U11575 ( .A1(n12632), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n12631), .ZN(n12635) );
  INV_X1 U11576 ( .A(n11180), .ZN(n11171) );
  INV_X2 U11577 ( .A(n20416), .ZN(n11172) );
  NAND2_X2 U11578 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22203), .ZN(n17744) );
  BUF_X2 U11579 ( .A(n14387), .Z(n18155) );
  NAND2_X2 U11580 ( .A1(n22203), .A2(n22205), .ZN(n17745) );
  CLKBUF_X1 U11581 ( .A(n13918), .Z(n15750) );
  BUF_X2 U11582 ( .A(n14396), .Z(n18157) );
  BUF_X2 U11583 ( .A(n18108), .Z(n18158) );
  INV_X1 U11584 ( .A(n14351), .ZN(n18082) );
  INV_X2 U11585 ( .A(n11192), .ZN(n18067) );
  INV_X1 U11586 ( .A(n11218), .ZN(n18156) );
  INV_X1 U11587 ( .A(n22172), .ZN(n17493) );
  AND2_X2 U11588 ( .A1(n12755), .A2(n14603), .ZN(n12773) );
  BUF_X4 U11589 ( .A(n12030), .Z(n12326) );
  INV_X2 U11590 ( .A(n18279), .ZN(n11173) );
  AND2_X2 U11591 ( .A1(n11711), .A2(n16830), .ZN(n11180) );
  OR2_X1 U11592 ( .A1(n14339), .A2(n15905), .ZN(n11192) );
  BUF_X4 U11593 ( .A(n14455), .Z(n11174) );
  AND2_X2 U11594 ( .A1(n14608), .A2(n14598), .ZN(n16007) );
  NAND2_X2 U11595 ( .A1(n22225), .A2(n18692), .ZN(n17479) );
  INV_X2 U11596 ( .A(n19154), .ZN(n19003) );
  BUF_X4 U11597 ( .A(n14472), .Z(n11175) );
  OR2_X1 U11599 ( .A1(n15905), .A2(n14340), .ZN(n11218) );
  AND2_X1 U11600 ( .A1(n14593), .A2(n11328), .ZN(n12656) );
  AND2_X1 U11601 ( .A1(n11328), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14608) );
  AND2_X1 U11602 ( .A1(n16832), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11712) );
  NAND2_X1 U11603 ( .A1(n21333), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14341) );
  BUF_X2 U11604 ( .A(n12030), .Z(n11177) );
  AND2_X1 U11605 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14191) );
  AND2_X2 U11606 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16830) );
  AND2_X1 U11607 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13933) );
  NOR2_X1 U11608 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14593) );
  INV_X1 U11609 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16832) );
  INV_X1 U11610 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14598) );
  AND2_X1 U11611 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11439) );
  AND2_X1 U11612 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14282) );
  BUF_X2 U11613 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n17422) );
  NOR2_X1 U11614 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12761) );
  AND2_X1 U11615 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15229) );
  OAI21_X1 U11616 ( .B1(n17077), .B2(n11671), .A(n13588), .ZN(n11673) );
  AND2_X1 U11617 ( .A1(n11711), .A2(n11719), .ZN(n11181) );
  NOR2_X2 U11618 ( .A1(n16323), .A2(n20431), .ZN(n16302) );
  NOR2_X2 U11619 ( .A1(n14258), .A2(n11626), .ZN(n15108) );
  NOR2_X2 U11620 ( .A1(n16313), .A2(n16314), .ZN(n12446) );
  NAND3_X2 U11621 ( .A1(n14350), .A2(n14349), .A3(n14348), .ZN(n21197) );
  NAND2_X2 U11622 ( .A1(n11560), .A2(n11562), .ZN(n16576) );
  NOR2_X2 U11623 ( .A1(n16584), .A2(n11258), .ZN(n11561) );
  NAND2_X1 U11624 ( .A1(n11846), .A2(n11829), .ZN(n13828) );
  NOR2_X1 U11625 ( .A1(n15292), .A2(n11829), .ZN(n15302) );
  AOI21_X1 U11626 ( .B1(n11844), .B2(n14245), .A(n11843), .ZN(n11855) );
  AND3_X1 U11627 ( .A1(n14245), .A2(n11890), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12546) );
  INV_X2 U11628 ( .A(n14245), .ZN(n11829) );
  NAND4_X1 U11629 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11178) );
  OR2_X2 U11630 ( .A1(n14254), .A2(n14131), .ZN(n12901) );
  NAND2_X4 U11631 ( .A1(n16676), .A2(n12527), .ZN(n16638) );
  NOR2_X2 U11632 ( .A1(n15625), .A2(n11621), .ZN(n15815) );
  NAND2_X2 U11633 ( .A1(n11850), .A2(n11371), .ZN(n11938) );
  NAND2_X2 U11634 ( .A1(n16603), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16584) );
  INV_X1 U11635 ( .A(n11183), .ZN(n11179) );
  NAND2_X2 U11636 ( .A1(n11829), .A2(n11828), .ZN(n15284) );
  NOR2_X4 U11638 ( .A1(n15080), .A2(n11569), .ZN(n17546) );
  OAI21_X2 U11639 ( .B1(n17224), .B2(n11358), .A(n11356), .ZN(n17077) );
  NOR2_X2 U11640 ( .A1(n21534), .A2(n21525), .ZN(n21517) );
  AND2_X1 U11641 ( .A1(n11711), .A2(n11719), .ZN(n12078) );
  NOR2_X4 U11642 ( .A1(n15497), .A2(n15496), .ZN(n15619) );
  NAND2_X4 U11643 ( .A1(n11937), .A2(n15377), .ZN(n15410) );
  NAND2_X2 U11644 ( .A1(n11559), .A2(n11895), .ZN(n15377) );
  INV_X1 U11645 ( .A(n16124), .ZN(n11185) );
  INV_X1 U11646 ( .A(n16124), .ZN(n11186) );
  AOI21_X1 U11647 ( .B1(n16236), .B2(n15635), .A(n11508), .ZN(n11187) );
  AOI21_X1 U11648 ( .B1(n16236), .B2(n15635), .A(n11508), .ZN(n11188) );
  AOI21_X4 U11649 ( .B1(n16236), .B2(n15635), .A(n11508), .ZN(n17412) );
  NAND2_X1 U11650 ( .A1(n21280), .A2(n21197), .ZN(n11189) );
  AND2_X2 U11651 ( .A1(n16099), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12951) );
  NOR2_X1 U11652 ( .A1(n21336), .A2(n17448), .ZN(n21293) );
  NAND2_X1 U11653 ( .A1(n12805), .A2(n12745), .ZN(n11350) );
  NAND2_X1 U11654 ( .A1(n22476), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12442) );
  INV_X1 U11655 ( .A(n13688), .ZN(n13710) );
  NAND2_X1 U11656 ( .A1(n11372), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11371) );
  NOR2_X1 U11657 ( .A1(n17422), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15926) );
  NOR2_X1 U11658 ( .A1(n13189), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13192) );
  AND2_X1 U11659 ( .A1(n11252), .A2(n11457), .ZN(n11456) );
  INV_X1 U11660 ( .A(n15898), .ZN(n11457) );
  INV_X1 U11661 ( .A(n16941), .ZN(n11449) );
  OR2_X1 U11662 ( .A1(n11242), .A2(n11640), .ZN(n11639) );
  INV_X1 U11663 ( .A(n15818), .ZN(n11640) );
  INV_X1 U11664 ( .A(n11680), .ZN(n11679) );
  NAND2_X1 U11665 ( .A1(n17164), .A2(n17165), .ZN(n11670) );
  OAI21_X1 U11666 ( .B1(n12827), .B2(n12826), .A(n12825), .ZN(n12828) );
  NOR2_X1 U11667 ( .A1(n14337), .A2(n21294), .ZN(n18109) );
  NOR2_X1 U11668 ( .A1(n20665), .A2(n21338), .ZN(n21352) );
  AOI22_X1 U11669 ( .A1(n17446), .A2(n17445), .B1(n17444), .B2(n17463), .ZN(
        n17457) );
  AND2_X1 U11670 ( .A1(n13808), .A2(n13807), .ZN(n15085) );
  NOR2_X1 U11671 ( .A1(n20437), .A2(n20433), .ZN(n11374) );
  NAND2_X1 U11672 ( .A1(n15842), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15292) );
  INV_X1 U11673 ( .A(n12442), .ZN(n16281) );
  NAND2_X1 U11674 ( .A1(n11307), .A2(n11425), .ZN(n11424) );
  NOR2_X1 U11675 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11425) );
  NOR3_X1 U11676 ( .A1(n16337), .A2(n11490), .A3(n11486), .ZN(n16295) );
  OR2_X1 U11677 ( .A1(n11487), .A2(n16316), .ZN(n11486) );
  INV_X1 U11678 ( .A(n16293), .ZN(n11490) );
  NAND2_X1 U11679 ( .A1(n11488), .A2(n16303), .ZN(n11487) );
  OR2_X1 U11680 ( .A1(n16349), .A2(n16339), .ZN(n16337) );
  OR2_X1 U11681 ( .A1(n20516), .A2(n21960), .ZN(n12527) );
  NAND2_X1 U11682 ( .A1(n16261), .A2(n14072), .ZN(n16210) );
  INV_X1 U11683 ( .A(n22162), .ZN(n14093) );
  AND2_X1 U11684 ( .A1(n16820), .A2(n14520), .ZN(n15353) );
  INV_X1 U11685 ( .A(n12592), .ZN(n11386) );
  NOR2_X1 U11686 ( .A1(n16901), .A2(n13642), .ZN(n13726) );
  INV_X1 U11687 ( .A(n11434), .ZN(n11433) );
  AND2_X1 U11688 ( .A1(n13479), .A2(n12815), .ZN(n15215) );
  NAND2_X1 U11689 ( .A1(n14252), .A2(n14229), .ZN(n14235) );
  AND2_X1 U11690 ( .A1(n14228), .A2(n14227), .ZN(n14229) );
  AND2_X1 U11691 ( .A1(n12801), .A2(n19160), .ZN(n13605) );
  NAND3_X1 U11692 ( .A1(n19325), .A2(n18052), .A3(n17457), .ZN(n17451) );
  CLKBUF_X3 U11693 ( .A(n14414), .Z(n18129) );
  INV_X1 U11694 ( .A(n16670), .ZN(n20514) );
  AND2_X1 U11695 ( .A1(n16670), .A2(n12601), .ZN(n20505) );
  XNOR2_X1 U11696 ( .A(n13644), .B(n13725), .ZN(n19029) );
  NAND2_X1 U11697 ( .A1(n12753), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U11698 ( .A1(n12856), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n12835) );
  NAND2_X1 U11699 ( .A1(n12638), .A2(n12609), .ZN(n12615) );
  XNOR2_X1 U11700 ( .A(n14603), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12614) );
  OAI21_X1 U11701 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21772), .A(
        n14372), .ZN(n14373) );
  OR2_X1 U11702 ( .A1(n14376), .A2(n14377), .ZN(n14372) );
  NAND2_X1 U11703 ( .A1(n12038), .A2(n12037), .ZN(n12065) );
  OR2_X1 U11704 ( .A1(n11889), .A2(n11888), .ZN(n12521) );
  INV_X1 U11705 ( .A(n11838), .ZN(n11890) );
  NAND2_X1 U11706 ( .A1(n11838), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12549) );
  AND2_X1 U11707 ( .A1(n11890), .A2(n15092), .ZN(n11798) );
  INV_X1 U11708 ( .A(n11798), .ZN(n11314) );
  INV_X1 U11709 ( .A(n12642), .ZN(n12643) );
  INV_X1 U11710 ( .A(n12864), .ZN(n13082) );
  NAND2_X1 U11711 ( .A1(n11427), .A2(n11662), .ZN(n12859) );
  NOR2_X1 U11712 ( .A1(n12832), .A2(n15635), .ZN(n11662) );
  INV_X1 U11713 ( .A(n14606), .ZN(n11427) );
  OR2_X1 U11714 ( .A1(n17078), .A2(n17088), .ZN(n13577) );
  NAND2_X1 U11715 ( .A1(n11402), .A2(n11246), .ZN(n12864) );
  NAND2_X1 U11716 ( .A1(n11348), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12813) );
  INV_X1 U11717 ( .A(n16092), .ZN(n16085) );
  NAND2_X1 U11718 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11441) );
  NAND2_X1 U11719 ( .A1(n12753), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11440) );
  AOI22_X1 U11720 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12673) );
  NAND2_X1 U11721 ( .A1(n18145), .A2(n21143), .ZN(n18169) );
  INV_X1 U11722 ( .A(n11408), .ZN(n18190) );
  AOI21_X1 U11723 ( .B1(n21784), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14371), .ZN(n14377) );
  AND2_X1 U11724 ( .A1(n17459), .A2(n17460), .ZN(n14371) );
  AND2_X1 U11725 ( .A1(n11860), .A2(n11832), .ZN(n14098) );
  NOR2_X1 U11726 ( .A1(n11576), .A2(n16336), .ZN(n11575) );
  NAND2_X1 U11727 ( .A1(n16347), .A2(n11577), .ZN(n11576) );
  INV_X1 U11728 ( .A(n16430), .ZN(n11577) );
  NAND2_X1 U11729 ( .A1(n11580), .A2(n11581), .ZN(n11579) );
  INV_X1 U11730 ( .A(n16437), .ZN(n11580) );
  NOR2_X1 U11731 ( .A1(n11582), .A2(n11583), .ZN(n11581) );
  INV_X1 U11732 ( .A(n16372), .ZN(n11582) );
  NAND2_X1 U11733 ( .A1(n16442), .A2(n11584), .ZN(n11583) );
  AND2_X1 U11734 ( .A1(n12018), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12042) );
  NAND2_X1 U11735 ( .A1(n11412), .A2(n15118), .ZN(n12024) );
  NOR2_X1 U11736 ( .A1(n11482), .A2(n11485), .ZN(n11481) );
  INV_X1 U11737 ( .A(n16383), .ZN(n11485) );
  INV_X1 U11738 ( .A(n11483), .ZN(n11482) );
  INV_X1 U11739 ( .A(n15662), .ZN(n11502) );
  AND2_X1 U11740 ( .A1(n15608), .A2(n20488), .ZN(n11318) );
  OR2_X1 U11741 ( .A1(n11960), .A2(n11959), .ZN(n12464) );
  NAND2_X1 U11742 ( .A1(n11798), .A2(n14098), .ZN(n11839) );
  INV_X1 U11743 ( .A(n12463), .ZN(n15127) );
  OR2_X1 U11744 ( .A1(n13521), .A2(n13519), .ZN(n13529) );
  NAND2_X1 U11745 ( .A1(n13516), .A2(n13515), .ZN(n13521) );
  INV_X1 U11746 ( .A(n13490), .ZN(n11476) );
  NOR2_X1 U11747 ( .A1(n13494), .A2(n11478), .ZN(n11477) );
  INV_X1 U11748 ( .A(n13503), .ZN(n11478) );
  INV_X1 U11749 ( .A(n15744), .ZN(n11622) );
  OR2_X1 U11750 ( .A1(n13043), .A2(n13042), .ZN(n13449) );
  NOR2_X1 U11751 ( .A1(n11298), .A2(n11645), .ZN(n11644) );
  INV_X1 U11752 ( .A(n17018), .ZN(n11645) );
  INV_X1 U11753 ( .A(n15853), .ZN(n11458) );
  OR2_X1 U11754 ( .A1(n17570), .A2(n17156), .ZN(n13467) );
  NOR2_X1 U11755 ( .A1(n18773), .A2(n11655), .ZN(n11654) );
  INV_X1 U11756 ( .A(n17390), .ZN(n11655) );
  INV_X1 U11757 ( .A(n13112), .ZN(n13727) );
  NAND2_X1 U11758 ( .A1(n13099), .A2(n11445), .ZN(n11444) );
  INV_X1 U11759 ( .A(n14230), .ZN(n11445) );
  NAND2_X1 U11760 ( .A1(n13058), .A2(n15685), .ZN(n11339) );
  AND2_X1 U11761 ( .A1(n12751), .A2(n12750), .ZN(n13379) );
  NAND2_X1 U11762 ( .A1(n12736), .A2(n12735), .ZN(n13604) );
  NAND2_X1 U11763 ( .A1(n13386), .A2(n13389), .ZN(n11344) );
  AOI221_X1 U11764 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12613), 
        .C1(n19065), .C2(n12613), .A(n12612), .ZN(n12790) );
  NAND2_X1 U11765 ( .A1(n12892), .A2(n12891), .ZN(n12898) );
  INV_X1 U11766 ( .A(n12659), .ZN(n11355) );
  AND2_X1 U11767 ( .A1(n14254), .A2(n15322), .ZN(n12907) );
  INV_X1 U11768 ( .A(n12898), .ZN(n12899) );
  NAND2_X1 U11769 ( .A1(n14403), .A2(n14402), .ZN(n11523) );
  AND2_X1 U11770 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11525) );
  AND2_X1 U11771 ( .A1(n11606), .A2(n11605), .ZN(n11604) );
  NAND2_X1 U11772 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11605) );
  INV_X1 U11773 ( .A(n18113), .ZN(n11597) );
  NAND2_X1 U11774 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11595) );
  NAND2_X1 U11775 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11596) );
  NAND2_X1 U11776 ( .A1(n18112), .A2(n11601), .ZN(n11600) );
  AOI21_X1 U11777 ( .B1(n18106), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n11602), .ZN(n11601) );
  NAND2_X1 U11778 ( .A1(n11603), .A2(n11230), .ZN(n11602) );
  INV_X1 U11779 ( .A(n21336), .ZN(n17449) );
  INV_X1 U11780 ( .A(n18243), .ZN(n11538) );
  NAND2_X1 U11781 ( .A1(n18235), .A2(n18178), .ZN(n11611) );
  NAND2_X1 U11782 ( .A1(n18174), .A2(n18552), .ZN(n18232) );
  NOR2_X1 U11783 ( .A1(n17463), .A2(n18051), .ZN(n17452) );
  AND3_X1 U11784 ( .A1(n18052), .A2(n21344), .A3(n21293), .ZN(n18050) );
  NOR2_X1 U11785 ( .A1(n22123), .A2(n22107), .ZN(n16362) );
  AND2_X1 U11786 ( .A1(n12293), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16280) );
  NOR2_X1 U11787 ( .A1(n16291), .A2(n11591), .ZN(n11590) );
  INV_X1 U11788 ( .A(n12447), .ZN(n11591) );
  AND2_X1 U11789 ( .A1(n16257), .A2(n13710), .ZN(n13711) );
  AND2_X1 U11790 ( .A1(n12263), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12264) );
  NAND2_X1 U11791 ( .A1(n14311), .A2(n14310), .ZN(n14309) );
  INV_X1 U11792 ( .A(n14314), .ZN(n11971) );
  OAI21_X1 U11793 ( .B1(n13661), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11197), .ZN(n11415) );
  AOI21_X1 U11794 ( .B1(n20516), .B2(n11418), .A(n11417), .ZN(n11416) );
  NOR2_X1 U11795 ( .A1(n16706), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11417) );
  NOR3_X1 U11796 ( .A1(n16337), .A2(n11489), .A3(n11491), .ZN(n16305) );
  NOR2_X1 U11797 ( .A1(n20516), .A2(n11564), .ZN(n11563) );
  AND2_X1 U11798 ( .A1(n16444), .A2(n16377), .ZN(n16434) );
  OR2_X1 U11799 ( .A1(n16638), .A2(n16652), .ZN(n11366) );
  OR2_X1 U11800 ( .A1(n12520), .A2(n21873), .ZN(n16653) );
  NAND2_X1 U11801 ( .A1(n11365), .A2(n11364), .ZN(n16677) );
  NAND2_X1 U11802 ( .A1(n16638), .A2(n16779), .ZN(n11365) );
  NAND2_X1 U11803 ( .A1(n11359), .A2(n12478), .ZN(n20469) );
  AND2_X1 U11804 ( .A1(n13837), .A2(n16831), .ZN(n15088) );
  AOI21_X1 U11805 ( .B1(n14048), .B2(n14047), .A(n22162), .ZN(n14066) );
  AND2_X1 U11806 ( .A1(n14046), .A2(n14045), .ZN(n14047) );
  INV_X1 U11807 ( .A(n11924), .ZN(n11426) );
  NAND2_X1 U11808 ( .A1(n11978), .A2(n11977), .ZN(n15165) );
  AND2_X1 U11809 ( .A1(n14569), .A2(n12463), .ZN(n14688) );
  INV_X1 U11810 ( .A(n22290), .ZN(n15381) );
  NOR2_X1 U11811 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14531), .ZN(n15699) );
  AOI21_X1 U11812 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n15376), .A(n22479), 
        .ZN(n15379) );
  INV_X1 U11813 ( .A(n15699), .ZN(n22479) );
  NAND2_X1 U11814 ( .A1(n16948), .A2(n11259), .ZN(n16926) );
  INV_X1 U11815 ( .A(n16924), .ZN(n11447) );
  NAND2_X1 U11816 ( .A1(n16931), .A2(n16930), .ZN(n16929) );
  NAND2_X1 U11817 ( .A1(n11636), .A2(n11630), .ZN(n11633) );
  AND2_X1 U11818 ( .A1(n11634), .A2(n15197), .ZN(n11630) );
  INV_X1 U11819 ( .A(n15201), .ZN(n11634) );
  OAI21_X1 U11820 ( .B1(n13722), .B2(n12850), .A(n13194), .ZN(n15192) );
  AND2_X2 U11821 ( .A1(n12722), .A2(n12723), .ZN(n14153) );
  OR2_X1 U11822 ( .A1(n13060), .A2(n13507), .ZN(n13076) );
  NAND2_X1 U11823 ( .A1(n13075), .A2(n17152), .ZN(n11677) );
  NAND2_X1 U11824 ( .A1(n11665), .A2(n11228), .ZN(n11666) );
  AND2_X1 U11825 ( .A1(n13466), .A2(n13465), .ZN(n17571) );
  NOR2_X1 U11826 ( .A1(n14275), .A2(n14276), .ZN(n14319) );
  INV_X1 U11827 ( .A(n13738), .ZN(n13741) );
  AND2_X1 U11828 ( .A1(n13081), .A2(n11212), .ZN(n13716) );
  OR3_X1 U11829 ( .A1(n18942), .A2(n13507), .A3(n17232), .ZN(n17096) );
  NAND2_X1 U11830 ( .A1(n16948), .A2(n16949), .ZN(n16950) );
  NAND2_X1 U11831 ( .A1(n13080), .A2(n13079), .ZN(n17113) );
  INV_X1 U11832 ( .A(n15797), .ZN(n11641) );
  NAND2_X1 U11833 ( .A1(n13615), .A2(n17642), .ZN(n17304) );
  INV_X1 U11834 ( .A(n18827), .ZN(n11646) );
  NAND2_X1 U11835 ( .A1(n17579), .A2(n17334), .ZN(n17356) );
  INV_X1 U11836 ( .A(n13020), .ZN(n13051) );
  XNOR2_X1 U11837 ( .A(n14212), .B(n14210), .ZN(n14163) );
  NAND2_X1 U11838 ( .A1(n14162), .A2(n14163), .ZN(n14214) );
  AOI21_X1 U11839 ( .B1(n14605), .B2(n14215), .A(n14152), .ZN(n14206) );
  NAND2_X1 U11840 ( .A1(n14206), .A2(n14207), .ZN(n14205) );
  AND2_X1 U11841 ( .A1(n19690), .A2(n20170), .ZN(n17424) );
  OR2_X1 U11842 ( .A1(n19690), .A2(n20170), .ZN(n19718) );
  NAND2_X1 U11843 ( .A1(n15637), .A2(n15638), .ZN(n19846) );
  NAND2_X1 U11844 ( .A1(n19162), .A2(n15635), .ZN(n15637) );
  NAND2_X1 U11845 ( .A1(n19846), .A2(n19788), .ZN(n19799) );
  NAND2_X1 U11846 ( .A1(n21352), .A2(n17447), .ZN(n20611) );
  AOI21_X1 U11847 ( .B1(n18442), .B2(n11542), .A(n11541), .ZN(n11540) );
  OR2_X1 U11848 ( .A1(n18442), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11544) );
  NOR2_X1 U11849 ( .A1(n11545), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11541) );
  INV_X1 U11850 ( .A(n21353), .ZN(n21359) );
  NOR2_X1 U11851 ( .A1(n18557), .A2(n20742), .ZN(n18540) );
  XNOR2_X1 U11852 ( .A(n18204), .B(n11403), .ZN(n18559) );
  INV_X1 U11853 ( .A(n18203), .ZN(n11403) );
  NAND2_X1 U11854 ( .A1(n18559), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18558) );
  NAND2_X1 U11855 ( .A1(n18553), .A2(n18554), .ZN(n18552) );
  NAND2_X1 U11856 ( .A1(n14370), .A2(n11391), .ZN(n11390) );
  NOR2_X1 U11857 ( .A1(n18545), .A2(n18546), .ZN(n18544) );
  AND2_X1 U11858 ( .A1(n17456), .A2(n11199), .ZN(n21328) );
  NAND2_X1 U11859 ( .A1(n17458), .A2(n19407), .ZN(n11373) );
  NOR2_X1 U11860 ( .A1(n14434), .A2(n14433), .ZN(n21351) );
  NAND2_X1 U11861 ( .A1(n15095), .A2(n13810), .ZN(n13976) );
  NOR2_X1 U11862 ( .A1(n22125), .A2(n20435), .ZN(n11378) );
  NAND2_X1 U11863 ( .A1(n22118), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U11864 ( .A1(n22124), .A2(n11306), .ZN(n16333) );
  NAND2_X1 U11865 ( .A1(n22124), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16354) );
  INV_X1 U11866 ( .A(n22134), .ZN(n22113) );
  AND2_X1 U11867 ( .A1(n15302), .A2(n15295), .ZN(n22118) );
  XNOR2_X1 U11868 ( .A(n16212), .B(n16211), .ZN(n16418) );
  NAND2_X1 U11869 ( .A1(n22141), .A2(n12598), .ZN(n16670) );
  NAND2_X1 U11870 ( .A1(n15095), .A2(n12597), .ZN(n22141) );
  INV_X1 U11871 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15376) );
  NAND2_X1 U11872 ( .A1(n11368), .A2(n11931), .ZN(n11932) );
  INV_X1 U11873 ( .A(n11947), .ZN(n16826) );
  NAND2_X1 U11874 ( .A1(n14650), .A2(n19160), .ZN(n19174) );
  AND2_X1 U11875 ( .A1(n16975), .A2(n16974), .ZN(n19000) );
  INV_X1 U11876 ( .A(n19009), .ZN(n19037) );
  AND2_X1 U11877 ( .A1(n13644), .A2(n13643), .ZN(n16252) );
  NAND2_X1 U11878 ( .A1(n14324), .A2(n11627), .ZN(n11626) );
  INV_X1 U11879 ( .A(n11628), .ZN(n11627) );
  INV_X1 U11880 ( .A(n18976), .ZN(n17198) );
  AOI21_X1 U11881 ( .B1(n19029), .B2(n19103), .A(n11651), .ZN(n11650) );
  NAND2_X1 U11882 ( .A1(n11695), .A2(n11652), .ZN(n11651) );
  AND2_X1 U11883 ( .A1(n13402), .A2(n17034), .ZN(n11652) );
  OAI21_X1 U11884 ( .B1(n17204), .B2(n19134), .A(n11461), .ZN(n11460) );
  AOI21_X1 U11885 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17208), .A(
        n11462), .ZN(n11461) );
  NOR2_X1 U11886 ( .A1(n17210), .A2(n17202), .ZN(n11462) );
  OAI21_X1 U11887 ( .B1(n11400), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17113), .ZN(n17286) );
  NOR2_X1 U11888 ( .A1(n17300), .A2(n17293), .ZN(n11400) );
  INV_X1 U11889 ( .A(n19138), .ZN(n19091) );
  AND2_X1 U11890 ( .A1(n13605), .A2(n14633), .ZN(n19138) );
  INV_X1 U11891 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19819) );
  INV_X1 U11892 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19786) );
  INV_X1 U11893 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19733) );
  INV_X1 U11894 ( .A(n21077), .ZN(n11558) );
  OR2_X1 U11895 ( .A1(n21080), .A2(n21068), .ZN(n11556) );
  OAI21_X1 U11896 ( .B1(n21004), .B2(n20864), .A(n11528), .ZN(n21027) );
  AOI21_X1 U11897 ( .B1(n21065), .B2(n11530), .A(n11529), .ZN(n11528) );
  INV_X1 U11898 ( .A(n21005), .ZN(n11530) );
  INV_X1 U11899 ( .A(n21021), .ZN(n11529) );
  NAND2_X1 U11900 ( .A1(n21003), .A2(n21065), .ZN(n21004) );
  NAND2_X1 U11901 ( .A1(n21004), .A2(n21005), .ZN(n21019) );
  INV_X1 U11902 ( .A(n21075), .ZN(n21092) );
  NAND2_X1 U11903 ( .A1(n21226), .A2(n11213), .ZN(n21215) );
  NOR3_X1 U11904 ( .A1(n21237), .A2(n21197), .A3(n11384), .ZN(n21198) );
  NAND2_X1 U11905 ( .A1(n21153), .A2(P3_EAX_REG_2__SCAN_IN), .ZN(n21152) );
  NAND2_X1 U11906 ( .A1(n21283), .A2(n21280), .ZN(n21274) );
  INV_X1 U11907 ( .A(n21274), .ZN(n21277) );
  INV_X1 U11908 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20671) );
  OAI21_X1 U11909 ( .B1(n11407), .B2(n21644), .A(n11406), .ZN(n21614) );
  OR2_X1 U11910 ( .A1(n21605), .A2(n21700), .ZN(n11406) );
  INV_X1 U11911 ( .A(n21604), .ZN(n11407) );
  OR2_X1 U11912 ( .A1(n21648), .A2(n11265), .ZN(n11405) );
  NOR2_X2 U11913 ( .A1(n21747), .A2(n21463), .ZN(n21765) );
  XNOR2_X1 U11914 ( .A(n13188), .B(n15649), .ZN(n12747) );
  NAND2_X1 U11915 ( .A1(n16134), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11334) );
  AOI22_X1 U11916 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U11917 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12731) );
  OR2_X1 U11918 ( .A1(n11876), .A2(n11875), .ZN(n12454) );
  NOR2_X1 U11919 ( .A1(n12066), .A2(n12039), .ZN(n11410) );
  INV_X1 U11920 ( .A(n12454), .ZN(n11892) );
  AND2_X2 U11921 ( .A1(n11419), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11718) );
  INV_X1 U11922 ( .A(n11850), .ZN(n11934) );
  OR2_X1 U11923 ( .A1(n11989), .A2(n11988), .ZN(n12480) );
  AND2_X1 U11924 ( .A1(n13603), .A2(n12641), .ZN(n13411) );
  AND2_X1 U11925 ( .A1(n11468), .A2(n11467), .ZN(n16106) );
  NAND2_X1 U11926 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11467) );
  NAND2_X1 U11927 ( .A1(n15953), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11468) );
  AND2_X1 U11928 ( .A1(n11466), .A2(n11465), .ZN(n15958) );
  NAND2_X1 U11929 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11465) );
  NAND2_X1 U11930 ( .A1(n15953), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U11931 ( .A1(n12835), .A2(n12834), .ZN(n12837) );
  AND2_X1 U11932 ( .A1(n13385), .A2(n12811), .ZN(n12846) );
  INV_X1 U11933 ( .A(n12913), .ZN(n12917) );
  AOI22_X1 U11934 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12984), .B1(
        n12993), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12913) );
  AND4_X1 U11935 ( .A1(n12924), .A2(n12923), .A3(n12922), .A4(n12921), .ZN(
        n12925) );
  NAND2_X1 U11936 ( .A1(n12804), .A2(n12803), .ZN(n13386) );
  AOI21_X1 U11937 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19786), .A(
        n12611), .ZN(n12613) );
  NOR2_X1 U11938 ( .A1(n12610), .A2(n12614), .ZN(n12611) );
  INV_X1 U11939 ( .A(n16124), .ZN(n15953) );
  NAND2_X1 U11940 ( .A1(n12608), .A2(n12607), .ZN(n12640) );
  NAND2_X1 U11941 ( .A1(n18109), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11603) );
  AND2_X1 U11942 ( .A1(n21147), .A2(n18191), .ZN(n18145) );
  OR2_X1 U11943 ( .A1(n18195), .A2(n21151), .ZN(n11408) );
  NAND2_X1 U11944 ( .A1(n11575), .A2(n16327), .ZN(n11574) );
  INV_X1 U11945 ( .A(n13685), .ZN(n13707) );
  INV_X1 U11946 ( .A(n11589), .ZN(n11588) );
  OAI21_X1 U11947 ( .B1(n15762), .B2(n15824), .A(n15656), .ZN(n11589) );
  AND2_X1 U11948 ( .A1(n15656), .A2(n15762), .ZN(n11587) );
  NAND2_X1 U11949 ( .A1(n12119), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12124) );
  AND2_X1 U11950 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11992), .ZN(
        n12018) );
  INV_X1 U11951 ( .A(n16328), .ZN(n11488) );
  INV_X1 U11952 ( .A(n16705), .ZN(n11418) );
  OR2_X1 U11953 ( .A1(n16316), .A2(n16328), .ZN(n11489) );
  INV_X1 U11954 ( .A(n13659), .ZN(n11564) );
  INV_X1 U11955 ( .A(n16427), .ZN(n11503) );
  NOR2_X1 U11956 ( .A1(n11505), .A2(n16365), .ZN(n11504) );
  INV_X1 U11957 ( .A(n16433), .ZN(n11505) );
  NOR2_X1 U11958 ( .A1(n16393), .A2(n11484), .ZN(n11483) );
  INV_X1 U11959 ( .A(n16407), .ZN(n11484) );
  NAND2_X1 U11960 ( .A1(n16206), .A2(n15657), .ZN(n16205) );
  NOR2_X1 U11961 ( .A1(n11495), .A2(n14682), .ZN(n11494) );
  INV_X1 U11962 ( .A(n16205), .ZN(n11479) );
  OR2_X1 U11963 ( .A1(n14677), .A2(n11496), .ZN(n11495) );
  INV_X1 U11964 ( .A(n15103), .ZN(n11496) );
  NAND2_X1 U11965 ( .A1(n16261), .A2(n16206), .ZN(n16199) );
  AND2_X1 U11966 ( .A1(n11832), .A2(n11178), .ZN(n12557) );
  NOR2_X1 U11967 ( .A1(n12549), .A2(n11896), .ZN(n12515) );
  NAND2_X1 U11968 ( .A1(n11894), .A2(n11915), .ZN(n11369) );
  NAND2_X1 U11969 ( .A1(n11314), .A2(n16272), .ZN(n11313) );
  NAND2_X1 U11970 ( .A1(n11839), .A2(n12449), .ZN(n11317) );
  INV_X1 U11971 ( .A(n11316), .ZN(n11315) );
  INV_X1 U11972 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17523) );
  INV_X1 U11973 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17517) );
  AOI21_X1 U11974 ( .B1(n15279), .B2(n22152), .A(n22156), .ZN(n14531) );
  AND2_X1 U11975 ( .A1(n12596), .A2(n13825), .ZN(n13834) );
  NAND2_X1 U11976 ( .A1(n12546), .A2(n12557), .ZN(n12593) );
  NOR2_X1 U11977 ( .A1(n13586), .A2(n13585), .ZN(n11469) );
  NOR2_X1 U11978 ( .A1(n13579), .A2(n13578), .ZN(n13581) );
  NAND2_X1 U11979 ( .A1(n13581), .A2(n13580), .ZN(n13586) );
  NOR2_X1 U11980 ( .A1(n13562), .A2(n11473), .ZN(n11472) );
  INV_X1 U11981 ( .A(n13524), .ZN(n11473) );
  NOR2_X1 U11982 ( .A1(n13448), .A2(n13475), .ZN(n13511) );
  INV_X1 U11983 ( .A(n13450), .ZN(n11471) );
  NAND2_X1 U11984 ( .A1(n13451), .A2(n13450), .ZN(n13460) );
  OAI21_X1 U11985 ( .B1(n13417), .B2(n13479), .A(n11474), .ZN(n13426) );
  NAND2_X1 U11986 ( .A1(n13479), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11474) );
  NOR2_X1 U11987 ( .A1(n11620), .A2(n16963), .ZN(n11619) );
  INV_X1 U11988 ( .A(n11697), .ZN(n11620) );
  NAND2_X1 U11989 ( .A1(n11638), .A2(n11288), .ZN(n11637) );
  INV_X1 U11990 ( .A(n11639), .ZN(n11638) );
  NAND2_X1 U11991 ( .A1(n11246), .A2(n14153), .ZN(n16092) );
  NOR2_X1 U11992 ( .A1(n17092), .A2(n11516), .ZN(n11515) );
  INV_X1 U11993 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11516) );
  AND2_X1 U11994 ( .A1(n13079), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11675) );
  NOR2_X1 U11995 ( .A1(n17120), .A2(n11512), .ZN(n11511) );
  INV_X1 U11996 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11512) );
  NOR2_X1 U11997 ( .A1(n17615), .A2(n17130), .ZN(n17632) );
  AND2_X1 U11998 ( .A1(n14319), .A2(n11451), .ZN(n15272) );
  AND2_X1 U11999 ( .A1(n11251), .A2(n11452), .ZN(n11451) );
  INV_X1 U12000 ( .A(n15273), .ZN(n11452) );
  NAND2_X1 U12001 ( .A1(n11520), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11519) );
  INV_X1 U12002 ( .A(n11521), .ZN(n11520) );
  NOR2_X1 U12003 ( .A1(n15110), .A2(n11454), .ZN(n11453) );
  INV_X1 U12004 ( .A(n14320), .ZN(n11454) );
  NAND2_X1 U12005 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11521) );
  OAI211_X1 U12006 ( .C1(n13097), .C2(n12868), .A(n12867), .B(n12866), .ZN(
        n12870) );
  NAND2_X1 U12007 ( .A1(n12876), .A2(n17422), .ZN(n11446) );
  NAND2_X1 U12008 ( .A1(n11346), .A2(n11345), .ZN(n11658) );
  INV_X1 U12009 ( .A(n12869), .ZN(n11346) );
  INV_X1 U12010 ( .A(n12870), .ZN(n11345) );
  AND2_X1 U12011 ( .A1(n13451), .A2(n11196), .ZN(n13746) );
  NAND2_X1 U12012 ( .A1(n11469), .A2(n11295), .ZN(n13745) );
  NAND2_X1 U12013 ( .A1(n11672), .A2(n13583), .ZN(n11671) );
  INV_X1 U12014 ( .A(n13577), .ZN(n11672) );
  AND2_X1 U12015 ( .A1(n11207), .A2(n16934), .ZN(n11448) );
  NOR2_X1 U12016 ( .A1(n11648), .A2(n17350), .ZN(n11647) );
  INV_X1 U12017 ( .A(n17363), .ZN(n11648) );
  AND2_X1 U12018 ( .A1(n11254), .A2(n17585), .ZN(n11438) );
  OR2_X1 U12019 ( .A1(n18789), .A2(n13507), .ZN(n13540) );
  XNOR2_X1 U12020 ( .A(n13060), .B(n13507), .ZN(n13073) );
  NAND2_X1 U12021 ( .A1(n12879), .A2(n12878), .ZN(n13090) );
  NAND2_X1 U12022 ( .A1(n12856), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n12874) );
  NOR2_X1 U12023 ( .A1(n13437), .A2(n13426), .ZN(n13424) );
  NAND2_X1 U12024 ( .A1(n13425), .A2(n13424), .ZN(n13423) );
  AND4_X1 U12025 ( .A1(n12797), .A2(n14297), .A3(n13622), .A4(n12796), .ZN(
        n12798) );
  NAND2_X1 U12026 ( .A1(n12819), .A2(n12818), .ZN(n12830) );
  NAND2_X1 U12027 ( .A1(n19069), .A2(n11220), .ZN(n12902) );
  INV_X1 U12028 ( .A(n12902), .ZN(n12906) );
  NAND2_X1 U12029 ( .A1(n12701), .A2(n14603), .ZN(n11660) );
  NAND2_X1 U12030 ( .A1(n12674), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12675) );
  NAND2_X1 U12031 ( .A1(n19819), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12642) );
  AND2_X1 U12032 ( .A1(n15635), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14215) );
  NOR2_X1 U12033 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21310), .ZN(
        n17459) );
  NAND3_X1 U12034 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20684) );
  NOR2_X1 U12035 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21316), .ZN(
        n14414) );
  NAND2_X1 U12036 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21772), .ZN(
        n14337) );
  NAND2_X1 U12037 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21310), .ZN(
        n14339) );
  NOR2_X1 U12038 ( .A1(n14339), .A2(n14338), .ZN(n14387) );
  NAND2_X1 U12039 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21296), .ZN(
        n14340) );
  NOR2_X1 U12040 ( .A1(n11546), .A2(n11550), .ZN(n11545) );
  INV_X1 U12041 ( .A(n11547), .ZN(n11546) );
  NOR2_X1 U12042 ( .A1(n11543), .A2(n11549), .ZN(n11542) );
  INV_X1 U12043 ( .A(n11545), .ZN(n11543) );
  NOR2_X1 U12044 ( .A1(n20671), .A2(n11548), .ZN(n11547) );
  INV_X1 U12045 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11548) );
  NOR2_X1 U12046 ( .A1(n20941), .A2(n11555), .ZN(n11554) );
  INV_X1 U12047 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11555) );
  AOI21_X1 U12048 ( .B1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18129), .A(
        n11392), .ZN(n11391) );
  INV_X1 U12049 ( .A(n14369), .ZN(n11392) );
  AOI22_X1 U12050 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18128), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14369) );
  AOI22_X1 U12051 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14370) );
  AND2_X1 U12052 ( .A1(n21472), .A2(n18234), .ZN(n18475) );
  NAND2_X1 U12053 ( .A1(n18587), .A2(n18198), .ZN(n18199) );
  NAND2_X1 U12054 ( .A1(n11409), .A2(n11408), .ZN(n18192) );
  NAND2_X1 U12055 ( .A1(n18191), .A2(n21276), .ZN(n11409) );
  AOI21_X1 U12056 ( .B1(n14377), .B2(n14376), .A(n14375), .ZN(n18047) );
  AND2_X1 U12057 ( .A1(n14378), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14380) );
  NAND2_X1 U12058 ( .A1(n17484), .A2(n20611), .ZN(n17485) );
  INV_X1 U12059 ( .A(n21314), .ZN(n21291) );
  NAND2_X1 U12060 ( .A1(n18048), .A2(n21328), .ZN(n21314) );
  NAND2_X1 U12061 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15905) );
  INV_X1 U12062 ( .A(n15284), .ZN(n15094) );
  NOR2_X1 U12063 ( .A1(n20425), .A2(n11382), .ZN(n11381) );
  INV_X1 U12064 ( .A(n16613), .ZN(n22109) );
  NAND2_X1 U12065 ( .A1(n22106), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n22107) );
  NAND2_X1 U12066 ( .A1(n11829), .A2(n15294), .ZN(n15283) );
  AND2_X1 U12067 ( .A1(n14268), .A2(n14267), .ZN(n14328) );
  NAND2_X1 U12068 ( .A1(n14312), .A2(n11972), .ZN(n14266) );
  AND2_X1 U12069 ( .A1(n14244), .A2(n14243), .ZN(n20356) );
  NOR2_X1 U12070 ( .A1(n13664), .A2(n13663), .ZN(n13668) );
  NOR2_X1 U12071 ( .A1(n12369), .A2(n16597), .ZN(n12370) );
  INV_X1 U12072 ( .A(n11575), .ZN(n11573) );
  NAND2_X1 U12073 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12320) );
  NAND2_X1 U12074 ( .A1(n11219), .A2(n11568), .ZN(n11565) );
  NAND2_X1 U12075 ( .A1(n11219), .A2(n16638), .ZN(n11324) );
  NOR2_X1 U12076 ( .A1(n12298), .A2(n16624), .ZN(n12299) );
  AND2_X1 U12077 ( .A1(n12281), .A2(n12280), .ZN(n16372) );
  AND2_X1 U12078 ( .A1(n12266), .A2(n12265), .ZN(n16442) );
  INV_X1 U12079 ( .A(n11568), .ZN(n12537) );
  NAND2_X1 U12080 ( .A1(n16638), .A2(n12533), .ZN(n11566) );
  NOR2_X1 U12081 ( .A1(n12232), .A2(n12231), .ZN(n12263) );
  NAND2_X1 U12082 ( .A1(n12199), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12232) );
  OR2_X1 U12083 ( .A1(n16455), .A2(n16405), .ZN(n16403) );
  AND2_X1 U12084 ( .A1(n12184), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12214) );
  AND2_X1 U12085 ( .A1(n12179), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12184) );
  NOR2_X1 U12086 ( .A1(n12164), .A2(n12140), .ZN(n12179) );
  INV_X1 U12087 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U12088 ( .A1(n12125), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12164) );
  NOR2_X1 U12089 ( .A1(n12094), .A2(n12093), .ZN(n12119) );
  INV_X1 U12090 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12093) );
  AND3_X1 U12091 ( .A1(n12092), .A2(n12091), .A3(n12090), .ZN(n15444) );
  CLKBUF_X1 U12092 ( .A(n15442), .Z(n15443) );
  INV_X1 U12093 ( .A(n12070), .ZN(n12071) );
  NAND2_X1 U12094 ( .A1(n12071), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12094) );
  AOI21_X1 U12095 ( .B1(n12496), .B2(n12226), .A(n12062), .ZN(n15220) );
  AND2_X1 U12096 ( .A1(n12042), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12060) );
  AOI21_X1 U12097 ( .B1(n12479), .B2(n12226), .A(n12023), .ZN(n15107) );
  OAI21_X1 U12098 ( .B1(n12463), .B2(n12182), .A(n11968), .ZN(n11969) );
  NAND2_X1 U12099 ( .A1(n11923), .A2(n11922), .ZN(n14145) );
  NAND2_X1 U12100 ( .A1(n16570), .A2(n16706), .ZN(n16153) );
  NOR2_X1 U12101 ( .A1(n16337), .A2(n11489), .ZN(n16315) );
  NAND2_X1 U12102 ( .A1(n16434), .A2(n16433), .ZN(n16436) );
  NAND2_X1 U12103 ( .A1(n16434), .A2(n11504), .ZN(n16428) );
  AND2_X1 U12104 ( .A1(n16459), .A2(n11264), .ZN(n16444) );
  INV_X1 U12105 ( .A(n16446), .ZN(n11480) );
  NAND2_X1 U12106 ( .A1(n16459), .A2(n11481), .ZN(n16445) );
  NAND2_X1 U12107 ( .A1(n16459), .A2(n16407), .ZN(n16408) );
  NOR2_X1 U12108 ( .A1(n16461), .A2(n16460), .ZN(n16459) );
  INV_X1 U12109 ( .A(n16638), .ZN(n16641) );
  NAND2_X1 U12110 ( .A1(n15868), .A2(n15867), .ZN(n16460) );
  NAND2_X1 U12111 ( .A1(n11499), .A2(n11497), .ZN(n15876) );
  NOR2_X1 U12112 ( .A1(n11200), .A2(n11498), .ZN(n11497) );
  INV_X1 U12113 ( .A(n15875), .ZN(n11498) );
  NOR2_X1 U12114 ( .A1(n15838), .A2(n15876), .ZN(n15868) );
  AOI21_X1 U12115 ( .B1(n16638), .B2(n16664), .A(n16663), .ZN(n16801) );
  NOR2_X1 U12116 ( .A1(n15598), .A2(n11200), .ZN(n15874) );
  NAND2_X1 U12117 ( .A1(n11499), .A2(n11500), .ZN(n15768) );
  NOR2_X1 U12118 ( .A1(n15598), .A2(n15599), .ZN(n15663) );
  INV_X1 U12119 ( .A(n11421), .ZN(n11420) );
  NAND2_X1 U12120 ( .A1(n20489), .A2(n11318), .ZN(n11422) );
  NOR2_X1 U12121 ( .A1(n15452), .A2(n15451), .ZN(n15454) );
  NAND2_X1 U12122 ( .A1(n20483), .A2(n20482), .ZN(n20481) );
  NOR2_X1 U12123 ( .A1(n14676), .A2(n11492), .ZN(n15331) );
  INV_X1 U12124 ( .A(n11494), .ZN(n11492) );
  OR2_X1 U12125 ( .A1(n14676), .A2(n11495), .ZN(n15104) );
  OR2_X1 U12126 ( .A1(n20525), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12602) );
  NAND2_X1 U12127 ( .A1(n14309), .A2(n12470), .ZN(n14330) );
  NAND2_X1 U12128 ( .A1(n14330), .A2(n14331), .ZN(n11359) );
  NOR2_X1 U12129 ( .A1(n16215), .A2(n21932), .ZN(n21877) );
  AND2_X1 U12130 ( .A1(n21850), .A2(n21855), .ZN(n21932) );
  AND2_X1 U12131 ( .A1(n14065), .A2(n14064), .ZN(n21880) );
  XNOR2_X1 U12132 ( .A(n13957), .B(n12460), .ZN(n14036) );
  MUX2_X1 U12133 ( .A(n16261), .B(n14072), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n14074) );
  NAND2_X1 U12134 ( .A1(n13958), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13957) );
  AND2_X1 U12135 ( .A1(n14062), .A2(n11853), .ZN(n11320) );
  AOI21_X1 U12136 ( .B1(n11925), .B2(n11924), .A(n12515), .ZN(n11915) );
  INV_X1 U12137 ( .A(n11369), .ZN(n11368) );
  NAND2_X1 U12138 ( .A1(n11931), .A2(n11894), .ZN(n11917) );
  NAND2_X1 U12139 ( .A1(n11369), .A2(n11931), .ZN(n11963) );
  AOI21_X1 U12140 ( .B1(n11947), .B2(n22153), .A(n11413), .ZN(n11962) );
  INV_X1 U12141 ( .A(n11961), .ZN(n11413) );
  AND2_X1 U12142 ( .A1(n15337), .A2(n16824), .ZN(n15338) );
  NOR2_X1 U12143 ( .A1(n14569), .A2(n15127), .ZN(n15342) );
  AND2_X1 U12144 ( .A1(n16270), .A2(n20519), .ZN(n22474) );
  AND2_X1 U12145 ( .A1(n15293), .A2(n15297), .ZN(n17544) );
  AND2_X1 U12146 ( .A1(n15288), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17549) );
  NAND2_X1 U12147 ( .A1(n12823), .A2(n13603), .ZN(n14296) );
  INV_X1 U12148 ( .A(n11469), .ZN(n13598) );
  NAND2_X1 U12149 ( .A1(n13525), .A2(n11201), .ZN(n13567) );
  INV_X1 U12150 ( .A(n13484), .ZN(n11475) );
  NAND2_X1 U12151 ( .A1(n13504), .A2(n11248), .ZN(n13492) );
  NAND2_X1 U12152 ( .A1(n13504), .A2(n11477), .ZN(n13496) );
  NAND2_X1 U12153 ( .A1(n13504), .A2(n13503), .ZN(n13506) );
  AND2_X1 U12154 ( .A1(n15225), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11508) );
  NAND2_X1 U12155 ( .A1(n15791), .A2(n11456), .ZN(n15901) );
  NAND2_X1 U12156 ( .A1(n16912), .A2(n16091), .ZN(n11618) );
  NAND2_X1 U12157 ( .A1(n17016), .A2(n11644), .ZN(n17008) );
  OAI21_X2 U12158 ( .B1(n16939), .B2(n16940), .A(n11273), .ZN(n16931) );
  NAND2_X1 U12159 ( .A1(n17016), .A2(n17018), .ZN(n17017) );
  NAND2_X1 U12160 ( .A1(n11206), .A2(n15790), .ZN(n11621) );
  INV_X1 U12161 ( .A(n11633), .ZN(n11632) );
  INV_X1 U12162 ( .A(n12824), .ZN(n15211) );
  INV_X1 U12163 ( .A(n12654), .ZN(n13865) );
  AND2_X1 U12164 ( .A1(n13864), .A2(n18722), .ZN(n17709) );
  INV_X1 U12165 ( .A(n13918), .ZN(n15753) );
  AND2_X1 U12166 ( .A1(n17056), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17042) );
  NOR2_X1 U12167 ( .A1(n17067), .A2(n18997), .ZN(n17056) );
  NAND2_X1 U12168 ( .A1(n17669), .A2(n11514), .ZN(n17067) );
  AND2_X1 U12169 ( .A1(n11204), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11514) );
  NOR2_X1 U12170 ( .A1(n16926), .A2(n13172), .ZN(n16908) );
  NAND2_X1 U12171 ( .A1(n17669), .A2(n11204), .ZN(n17081) );
  NAND2_X1 U12172 ( .A1(n17669), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17668) );
  NOR2_X1 U12173 ( .A1(n17661), .A2(n18940), .ZN(n17669) );
  NAND2_X1 U12174 ( .A1(n17662), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17661) );
  AND2_X1 U12175 ( .A1(n17652), .A2(n11510), .ZN(n17662) );
  AND2_X1 U12176 ( .A1(n11203), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11510) );
  NAND2_X1 U12177 ( .A1(n17652), .A2(n11203), .ZN(n17114) );
  AND2_X1 U12178 ( .A1(n15791), .A2(n11267), .ZN(n16959) );
  INV_X1 U12179 ( .A(n13632), .ZN(n11455) );
  NAND2_X1 U12180 ( .A1(n17652), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17651) );
  NAND2_X1 U12181 ( .A1(n17632), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17639) );
  NAND2_X1 U12182 ( .A1(n17616), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17615) );
  NOR2_X1 U12183 ( .A1(n15550), .A2(n17614), .ZN(n17616) );
  NAND2_X1 U12184 ( .A1(n15558), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15550) );
  NAND2_X1 U12185 ( .A1(n15272), .A2(n13128), .ZN(n15545) );
  INV_X1 U12186 ( .A(n15490), .ZN(n13128) );
  NOR2_X1 U12187 ( .A1(n15553), .A2(n11518), .ZN(n15558) );
  OR2_X1 U12188 ( .A1(n11519), .A2(n18801), .ZN(n11518) );
  NAND2_X1 U12189 ( .A1(n14319), .A2(n11251), .ZN(n15274) );
  NOR2_X1 U12190 ( .A1(n15553), .A2(n11521), .ZN(n15555) );
  NOR2_X1 U12191 ( .A1(n15553), .A2(n17578), .ZN(n15557) );
  NAND2_X1 U12192 ( .A1(n14319), .A2(n14320), .ZN(n15109) );
  NAND2_X1 U12193 ( .A1(n15554), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15553) );
  NOR2_X1 U12194 ( .A1(n15551), .A2(n17167), .ZN(n15554) );
  NAND2_X1 U12195 ( .A1(n15226), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15551) );
  INV_X1 U12196 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15510) );
  INV_X1 U12197 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U12198 ( .A1(n11625), .A2(n11624), .ZN(n12891) );
  INV_X1 U12199 ( .A(n12889), .ZN(n11624) );
  AND2_X1 U12200 ( .A1(n13597), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13739) );
  AND2_X1 U12201 ( .A1(n11644), .A2(n11643), .ZN(n11642) );
  INV_X1 U12202 ( .A(n16999), .ZN(n11643) );
  AND2_X1 U12203 ( .A1(n13591), .A2(n13590), .ZN(n17088) );
  NAND2_X1 U12204 ( .A1(n17225), .A2(n11357), .ZN(n11356) );
  NOR2_X1 U12205 ( .A1(n17225), .A2(n11357), .ZN(n11358) );
  NAND2_X1 U12206 ( .A1(n16948), .A2(n11448), .ZN(n16936) );
  NAND2_X1 U12207 ( .A1(n15791), .A2(n11252), .ZN(n15899) );
  NOR2_X1 U12208 ( .A1(n19107), .A2(n13625), .ZN(n17645) );
  AOI21_X1 U12209 ( .B1(n13612), .B2(n13610), .A(n11431), .ZN(n11430) );
  INV_X1 U12210 ( .A(n13612), .ZN(n11432) );
  INV_X1 U12211 ( .A(n13613), .ZN(n11431) );
  NAND2_X1 U12212 ( .A1(n15791), .A2(n15792), .ZN(n15854) );
  AND2_X1 U12213 ( .A1(n15628), .A2(n15730), .ZN(n15791) );
  NAND2_X1 U12214 ( .A1(n18791), .A2(n11249), .ZN(n18828) );
  INV_X1 U12215 ( .A(n17356), .ZN(n11343) );
  OR3_X1 U12216 ( .A1(n13544), .A2(n13507), .A3(n17348), .ZN(n17342) );
  NAND2_X1 U12217 ( .A1(n18791), .A2(n17363), .ZN(n17362) );
  AND2_X1 U12218 ( .A1(n11654), .A2(n17377), .ZN(n11653) );
  AOI21_X1 U12219 ( .B1(n13467), .B2(n17156), .A(n17571), .ZN(n11667) );
  NOR2_X1 U12220 ( .A1(n11664), .A2(n17155), .ZN(n11663) );
  INV_X1 U12221 ( .A(n13467), .ZN(n11664) );
  NAND2_X1 U12222 ( .A1(n11677), .A2(n11194), .ZN(n11678) );
  AND2_X1 U12223 ( .A1(n17391), .A2(n11654), .ZN(n18771) );
  NAND2_X1 U12224 ( .A1(n17391), .A2(n17390), .ZN(n18772) );
  AOI21_X1 U12225 ( .B1(n13022), .B2(n15685), .A(n11396), .ZN(n13059) );
  NAND2_X1 U12226 ( .A1(n11442), .A2(n11231), .ZN(n14275) );
  INV_X1 U12227 ( .A(n11444), .ZN(n11443) );
  NOR2_X1 U12228 ( .A1(n14237), .A2(n11444), .ZN(n14261) );
  OAI21_X1 U12229 ( .B1(n13022), .B2(n11396), .A(n11395), .ZN(n11398) );
  NAND2_X1 U12230 ( .A1(n12856), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13096) );
  OR2_X1 U12231 ( .A1(n14237), .A2(n14236), .ZN(n14239) );
  AND2_X1 U12232 ( .A1(n14127), .A2(n19106), .ZN(n15469) );
  INV_X1 U12233 ( .A(n12974), .ZN(n11394) );
  XNOR2_X1 U12234 ( .A(n13204), .B(n13198), .ZN(n13779) );
  NAND2_X1 U12235 ( .A1(n14214), .A2(n14213), .ZN(n14251) );
  NOR2_X1 U12236 ( .A1(n17691), .A2(n20060), .ZN(n19825) );
  INV_X1 U12237 ( .A(n19718), .ZN(n19821) );
  AND2_X1 U12238 ( .A1(n17691), .A2(n17686), .ZN(n19719) );
  INV_X1 U12239 ( .A(n17424), .ZN(n19729) );
  OR2_X1 U12240 ( .A1(n19690), .A2(n19674), .ZN(n19755) );
  OAI21_X1 U12241 ( .B1(n11353), .B2(n11352), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11342) );
  OAI21_X1 U12242 ( .B1(n11355), .B2(n11354), .A(n14603), .ZN(n11341) );
  INV_X1 U12243 ( .A(n12663), .ZN(n11353) );
  NAND2_X1 U12244 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19846), .ZN(n20176) );
  INV_X1 U12245 ( .A(n11151), .ZN(n20065) );
  NAND2_X1 U12247 ( .A1(n19690), .A2(n19674), .ZN(n19750) );
  NAND2_X1 U12248 ( .A1(n17691), .A2(n20060), .ZN(n19691) );
  CLKBUF_X1 U12249 ( .A(n12820), .Z(n14665) );
  NOR2_X1 U12250 ( .A1(n20666), .A2(n20665), .ZN(n17487) );
  NOR2_X1 U12251 ( .A1(n18049), .A2(n17485), .ZN(n21777) );
  INV_X1 U12252 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20798) );
  INV_X1 U12253 ( .A(n20674), .ZN(n20667) );
  NOR2_X1 U12254 ( .A1(n21220), .A2(n20629), .ZN(n11380) );
  NOR2_X1 U12255 ( .A1(n11524), .A2(n11523), .ZN(n11522) );
  CLKBUF_X3 U12256 ( .A(n14484), .Z(n18134) );
  NAND3_X1 U12257 ( .A1(n11233), .A2(n11599), .A3(n11598), .ZN(n18193) );
  NOR2_X1 U12258 ( .A1(n11229), .A2(n11600), .ZN(n11599) );
  NOR3_X1 U12259 ( .A1(n17484), .A2(n21339), .A3(n20609), .ZN(n18672) );
  NAND2_X1 U12260 ( .A1(n18442), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18408) );
  NOR2_X1 U12261 ( .A1(n18394), .A2(n21016), .ZN(n18364) );
  AND2_X1 U12262 ( .A1(n18219), .A2(n11553), .ZN(n18331) );
  AND2_X1 U12263 ( .A1(n11205), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11553) );
  NAND2_X1 U12264 ( .A1(n18219), .A2(n11205), .ZN(n18313) );
  NOR2_X1 U12265 ( .A1(n18451), .A2(n20913), .ZN(n18219) );
  NOR2_X1 U12266 ( .A1(n11536), .A2(n18497), .ZN(n18453) );
  NAND2_X1 U12267 ( .A1(n11534), .A2(n11537), .ZN(n18451) );
  NOR2_X1 U12268 ( .A1(n18497), .A2(n11535), .ZN(n11534) );
  INV_X1 U12269 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11535) );
  NOR2_X1 U12270 ( .A1(n18497), .A2(n20826), .ZN(n18255) );
  OAI21_X1 U12271 ( .B1(n20671), .B2(n18407), .A(n19324), .ZN(n18363) );
  NOR2_X1 U12272 ( .A1(n21733), .A2(n21487), .ZN(n18474) );
  NAND2_X1 U12273 ( .A1(n11539), .A2(n11195), .ZN(n18229) );
  INV_X1 U12274 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18470) );
  INV_X1 U12275 ( .A(n18363), .ZN(n18406) );
  NAND2_X1 U12276 ( .A1(n21832), .A2(n21801), .ZN(n18212) );
  NAND2_X1 U12277 ( .A1(n11552), .A2(n11260), .ZN(n18557) );
  INV_X1 U12278 ( .A(n18581), .ZN(n11552) );
  NAND2_X1 U12279 ( .A1(n18563), .A2(n18172), .ZN(n18553) );
  XNOR2_X1 U12280 ( .A(n18199), .B(n21419), .ZN(n18576) );
  NAND2_X1 U12281 ( .A1(n18576), .A2(n18575), .ZN(n18574) );
  NAND2_X1 U12282 ( .A1(n18591), .A2(n18167), .ZN(n18579) );
  NAND2_X1 U12283 ( .A1(n18611), .A2(n18618), .ZN(n18609) );
  OAI211_X1 U12284 ( .C1(n18373), .C2(n21573), .A(n18372), .B(n18390), .ZN(
        n18374) );
  INV_X1 U12285 ( .A(n18373), .ZN(n18391) );
  NOR2_X1 U12286 ( .A1(n21292), .A2(n21290), .ZN(n21357) );
  INV_X1 U12287 ( .A(n11610), .ZN(n11609) );
  AOI22_X1 U12288 ( .A1(n18179), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n18492), .B2(n21722), .ZN(n11610) );
  NAND2_X1 U12289 ( .A1(n18526), .A2(n18527), .ZN(n18525) );
  NAND2_X1 U12290 ( .A1(n18558), .A2(n18205), .ZN(n18545) );
  INV_X1 U12291 ( .A(n18175), .ZN(n11607) );
  XNOR2_X1 U12292 ( .A(n18170), .B(n11608), .ZN(n18564) );
  INV_X1 U12293 ( .A(n18171), .ZN(n11608) );
  NAND2_X1 U12294 ( .A1(n18564), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18563) );
  XNOR2_X1 U12295 ( .A(n18166), .B(n21420), .ZN(n18593) );
  NAND2_X1 U12296 ( .A1(n18593), .A2(n18592), .ZN(n18591) );
  NAND2_X1 U12297 ( .A1(n18588), .A2(n18589), .ZN(n18587) );
  INV_X1 U12298 ( .A(n21759), .ZN(n21742) );
  XNOR2_X1 U12299 ( .A(n18192), .B(n21399), .ZN(n18604) );
  AOI211_X1 U12300 ( .C1(n11176), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n14410), .B(n14409), .ZN(n14411) );
  INV_X1 U12301 ( .A(n21644), .ZN(n21780) );
  INV_X1 U12302 ( .A(n17474), .ZN(n18049) );
  NOR2_X1 U12303 ( .A1(n14394), .A2(n14393), .ZN(n19407) );
  NOR2_X1 U12304 ( .A1(n14424), .A2(n14423), .ZN(n21336) );
  INV_X1 U12305 ( .A(n19366), .ZN(n19532) );
  OAI22_X1 U12306 ( .A1(n21349), .A2(n21721), .B1(n21781), .B2(n21644), .ZN(
        n21801) );
  NOR2_X1 U12307 ( .A1(n21341), .A2(n17451), .ZN(n21808) );
  AND2_X1 U12308 ( .A1(n15284), .A2(n16261), .ZN(n13818) );
  AND3_X1 U12309 ( .A1(n14242), .A2(n13976), .A3(n13816), .ZN(n21838) );
  NAND2_X1 U12310 ( .A1(n16302), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16298) );
  OR2_X1 U12311 ( .A1(n16333), .A2(n20430), .ZN(n16323) );
  AND2_X1 U12312 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n16256), .ZN(n22124) );
  NOR2_X1 U12313 ( .A1(n22094), .A2(n22000), .ZN(n22106) );
  NOR2_X1 U12314 ( .A1(n16412), .A2(n20413), .ZN(n16397) );
  NAND2_X1 U12315 ( .A1(n16397), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n22094) );
  NOR2_X1 U12316 ( .A1(n20408), .A2(n22087), .ZN(n16413) );
  NOR2_X1 U12317 ( .A1(n15859), .A2(n21853), .ZN(n15861) );
  AND2_X1 U12318 ( .A1(n15302), .A2(n17544), .ZN(n22024) );
  NAND2_X1 U12319 ( .A1(n22024), .A2(n11389), .ZN(n15859) );
  AND2_X1 U12320 ( .A1(n22071), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n11389) );
  AND2_X1 U12321 ( .A1(n15842), .A2(n15446), .ZN(n22100) );
  INV_X1 U12322 ( .A(n22118), .ZN(n22131) );
  OR2_X1 U12323 ( .A1(n15290), .A2(n22137), .ZN(n22030) );
  INV_X1 U12324 ( .A(n22024), .ZN(n22073) );
  XNOR2_X1 U12325 ( .A(n16264), .B(n16263), .ZN(n16684) );
  NAND2_X2 U12326 ( .A1(n14080), .A2(n14079), .ZN(n16451) );
  INV_X1 U12327 ( .A(n16523), .ZN(n16549) );
  NOR2_X1 U12328 ( .A1(n16549), .A2(n14100), .ZN(n16551) );
  NAND2_X1 U12329 ( .A1(n14097), .A2(n14096), .ZN(n16523) );
  INV_X1 U12330 ( .A(n16279), .ZN(n11592) );
  OR2_X1 U12331 ( .A1(n20522), .A2(n22069), .ZN(n11363) );
  NAND2_X1 U12332 ( .A1(n15609), .A2(n15608), .ZN(n15607) );
  NAND2_X1 U12333 ( .A1(n20487), .A2(n12514), .ZN(n15609) );
  INV_X1 U12334 ( .A(n11415), .ZN(n11414) );
  OR2_X1 U12335 ( .A1(n16295), .A2(n16294), .ZN(n16700) );
  NAND2_X1 U12336 ( .A1(n11366), .A2(n16651), .ZN(n16654) );
  XNOR2_X1 U12337 ( .A(n16814), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20493) );
  INV_X1 U12338 ( .A(n22004), .ZN(n22018) );
  NAND2_X1 U12339 ( .A1(n11895), .A2(n11319), .ZN(n14523) );
  INV_X1 U12340 ( .A(n14520), .ZN(n14687) );
  INV_X1 U12341 ( .A(n22253), .ZN(n22290) );
  INV_X1 U12342 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U12343 ( .A1(n15527), .A2(n15526), .ZN(n22495) );
  OAI21_X1 U12344 ( .B1(n22260), .B2(n22508), .A(n22297), .ZN(n22510) );
  OR3_X1 U12345 ( .A1(n15171), .A2(n15170), .A3(n15169), .ZN(n22517) );
  INV_X1 U12346 ( .A(n22527), .ZN(n22530) );
  OAI211_X1 U12347 ( .C1(n22535), .C2(n22280), .A(n22279), .B(n22278), .ZN(
        n22538) );
  OAI22_X1 U12348 ( .A1(n15721), .A2(n15722), .B1(n22274), .B2(n22288), .ZN(
        n22549) );
  AND2_X1 U12349 ( .A1(n14688), .A2(n15382), .ZN(n22548) );
  NAND2_X1 U12350 ( .A1(n14688), .A2(n15352), .ZN(n22553) );
  INV_X1 U12351 ( .A(n22553), .ZN(n22556) );
  INV_X1 U12352 ( .A(n22573), .ZN(n16887) );
  INV_X1 U12353 ( .A(n22563), .ZN(n16893) );
  NAND2_X1 U12354 ( .A1(n14688), .A2(n15353), .ZN(n22567) );
  OAI211_X1 U12355 ( .C1(n16860), .C2(n12293), .A(n22297), .B(n16859), .ZN(
        n22564) );
  NOR2_X1 U12356 ( .A1(n14536), .A2(n22479), .ZN(n22325) );
  NOR2_X1 U12357 ( .A1(n14562), .A2(n22479), .ZN(n22354) );
  OAI211_X1 U12358 ( .C1(n22298), .C2(n22575), .A(n22297), .B(n22296), .ZN(
        n22578) );
  INV_X1 U12359 ( .A(n22355), .ZN(n22341) );
  INV_X1 U12360 ( .A(n22378), .ZN(n22370) );
  OR2_X1 U12361 ( .A1(n15388), .A2(n14521), .ZN(n22235) );
  NOR2_X1 U12362 ( .A1(n13829), .A2(n22280), .ZN(n22156) );
  INV_X1 U12363 ( .A(n15095), .ZN(n13829) );
  INV_X1 U12364 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22280) );
  NOR2_X1 U12365 ( .A1(n14638), .A2(n13798), .ZN(n13859) );
  OAI21_X1 U12366 ( .B1(n19002), .B2(n19001), .A(n17412), .ZN(n19005) );
  NAND2_X1 U12367 ( .A1(n18979), .A2(n18980), .ZN(n19001) );
  NAND2_X1 U12368 ( .A1(n18948), .A2(n18949), .ZN(n11506) );
  AND2_X1 U12369 ( .A1(n16942), .A2(n11450), .ZN(n18945) );
  INV_X1 U12370 ( .A(n19040), .ZN(n19013) );
  NAND2_X1 U12371 ( .A1(n11187), .A2(n18887), .ZN(n11507) );
  NAND2_X1 U12372 ( .A1(n11507), .A2(n18888), .ZN(n18899) );
  INV_X1 U12373 ( .A(n19041), .ZN(n19011) );
  INV_X1 U12374 ( .A(n19045), .ZN(n19008) );
  AND2_X1 U12375 ( .A1(n15246), .A2(n15245), .ZN(n19009) );
  INV_X1 U12376 ( .A(n14615), .ZN(n19069) );
  AND2_X1 U12377 ( .A1(n15246), .A2(n15244), .ZN(n19045) );
  XNOR2_X1 U12378 ( .A(n13732), .B(n13731), .ZN(n16894) );
  OR2_X1 U12379 ( .A1(n13317), .A2(n13316), .ZN(n15621) );
  NAND2_X1 U12380 ( .A1(n11693), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11628) );
  OR2_X1 U12381 ( .A1(n13248), .A2(n13247), .ZN(n14324) );
  OR2_X1 U12382 ( .A1(n14258), .A2(n11629), .ZN(n14321) );
  INV_X1 U12383 ( .A(n17691), .ZN(n19795) );
  INV_X2 U12384 ( .A(n16952), .ZN(n16966) );
  INV_X1 U12385 ( .A(n11327), .ZN(n12886) );
  INV_X1 U12386 ( .A(n16968), .ZN(n15746) );
  XNOR2_X1 U12387 ( .A(n13724), .B(n13723), .ZN(n19052) );
  AND2_X1 U12388 ( .A1(n20162), .A2(n15215), .ZN(n19955) );
  NOR2_X1 U12389 ( .A1(n11633), .A2(n11631), .ZN(n15232) );
  INV_X1 U12390 ( .A(n11635), .ZN(n11631) );
  NOR2_X1 U12391 ( .A1(n14154), .A2(n14106), .ZN(n20170) );
  BUF_X1 U12393 ( .A(n17725), .Z(n17733) );
  NOR2_X1 U12394 ( .A1(n17709), .A2(n17733), .ZN(n17722) );
  XNOR2_X1 U12395 ( .A(n11509), .B(n15224), .ZN(n16236) );
  NAND2_X1 U12396 ( .A1(n17042), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11509) );
  NOR2_X1 U12397 ( .A1(n17286), .A2(n17676), .ZN(n13637) );
  AND2_X1 U12398 ( .A1(n11677), .A2(n11221), .ZN(n17569) );
  NAND2_X1 U12399 ( .A1(n11666), .A2(n13463), .ZN(n17574) );
  INV_X1 U12400 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17167) );
  INV_X1 U12401 ( .A(n17640), .ZN(n17681) );
  NAND2_X1 U12402 ( .A1(n19174), .A2(n13627), .ZN(n17633) );
  CLKBUF_X1 U12403 ( .A(n14254), .Z(n14255) );
  AND2_X1 U12404 ( .A1(n17633), .A2(n17494), .ZN(n17673) );
  OR2_X1 U12405 ( .A1(n19174), .A2(n19060), .ZN(n17676) );
  INV_X1 U12406 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13967) );
  AND2_X1 U12407 ( .A1(n17633), .A2(n13954), .ZN(n17640) );
  OR2_X1 U12408 ( .A1(n19174), .A2(n16097), .ZN(n17608) );
  INV_X1 U12409 ( .A(n17676), .ZN(n17664) );
  INV_X1 U12410 ( .A(n17673), .ZN(n17657) );
  AOI21_X1 U12411 ( .B1(n16252), .B2(n19103), .A(n17043), .ZN(n13650) );
  AOI211_X1 U12412 ( .C1(n19129), .C2(n19000), .A(n17175), .B(n17174), .ZN(
        n17178) );
  OR2_X1 U12413 ( .A1(n17210), .A2(n13407), .ZN(n17184) );
  NAND2_X1 U12414 ( .A1(n13561), .A2(n13560), .ZN(n11657) );
  NAND2_X1 U12415 ( .A1(n17304), .A2(n17301), .ZN(n17121) );
  NOR2_X1 U12416 ( .A1(n17315), .A2(n11242), .ZN(n15817) );
  NAND2_X1 U12417 ( .A1(n17132), .A2(n13611), .ZN(n17630) );
  OR2_X1 U12418 ( .A1(n13053), .A2(n13051), .ZN(n11397) );
  INV_X1 U12419 ( .A(n19103), .ZN(n19133) );
  INV_X1 U12420 ( .A(n19119), .ZN(n19129) );
  AND2_X1 U12421 ( .A1(n14214), .A2(n14164), .ZN(n20060) );
  OR2_X1 U12422 ( .A1(n14163), .A2(n14162), .ZN(n14164) );
  AND2_X1 U12423 ( .A1(n11635), .A2(n11636), .ZN(n15199) );
  INV_X1 U12424 ( .A(n20170), .ZN(n19674) );
  OAI21_X1 U12425 ( .B1(n14207), .B2(n14206), .A(n14205), .ZN(n19690) );
  INV_X1 U12426 ( .A(n20060), .ZN(n17686) );
  AND2_X1 U12427 ( .A1(n14646), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19162) );
  CLKBUF_X1 U12428 ( .A(n12818), .Z(n19062) );
  OAI21_X1 U12429 ( .B1(n19850), .B2(n19849), .A(n19848), .ZN(n20285) );
  NOR2_X1 U12430 ( .A1(n19691), .A2(n19729), .ZN(n20155) );
  INV_X1 U12431 ( .A(n20276), .ZN(n20053) );
  AND2_X1 U12432 ( .A1(n19825), .A2(n19821), .ZN(n20282) );
  OAI21_X1 U12433 ( .B1(n17434), .B2(n17433), .A(n17432), .ZN(n20252) );
  NOR2_X1 U12434 ( .A1(n19766), .A2(n19750), .ZN(n20138) );
  AND2_X1 U12435 ( .A1(n19719), .A2(n19821), .ZN(n20225) );
  INV_X1 U12436 ( .A(n20223), .ZN(n20212) );
  OR3_X1 U12437 ( .A1(n19712), .A2(n20174), .A3(n19711), .ZN(n20214) );
  OAI21_X1 U12438 ( .B1(n19715), .B2(n19714), .A(n19713), .ZN(n20213) );
  INV_X1 U12439 ( .A(n20217), .ZN(n20130) );
  OR2_X1 U12440 ( .A1(n15642), .A2(n15641), .ZN(n20201) );
  INV_X1 U12441 ( .A(n20272), .ZN(n20283) );
  INV_X1 U12442 ( .A(n20160), .ZN(n20150) );
  OAI22_X1 U12443 ( .A1(n20569), .A2(n22599), .B1(n20066), .B2(n20065), .ZN(
        n20100) );
  INV_X1 U12444 ( .A(n20058), .ZN(n20045) );
  OAI22_X1 U12445 ( .A1(n20573), .A2(n22599), .B1(n19964), .B2(n20065), .ZN(
        n19999) );
  AOI21_X1 U12446 ( .B1(n20185), .B2(n19846), .A(n19686), .ZN(n20187) );
  INV_X1 U12447 ( .A(n20290), .ZN(n20267) );
  AND2_X1 U12448 ( .A1(n19060), .A2(n17431), .ZN(n20154) );
  INV_X1 U12449 ( .A(n20103), .ZN(n20105) );
  INV_X1 U12450 ( .A(n20036), .ZN(n20055) );
  INV_X1 U12451 ( .A(n20002), .ZN(n20004) );
  INV_X1 U12452 ( .A(n19902), .ZN(n19892) );
  INV_X1 U12453 ( .A(n19864), .ZN(n19898) );
  NOR2_X2 U12454 ( .A1(n19691), .A2(n19750), .ZN(n20186) );
  INV_X1 U12455 ( .A(n20155), .ZN(n20289) );
  INV_X1 U12456 ( .A(n19171), .ZN(n19160) );
  OR2_X1 U12457 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n17492), .ZN(n17750) );
  NAND2_X1 U12458 ( .A1(n21832), .A2(n21795), .ZN(n20609) );
  INV_X1 U12459 ( .A(n18212), .ZN(n21835) );
  OAI21_X1 U12460 ( .B1(n20930), .B2(n20864), .A(n11531), .ZN(n20953) );
  AOI21_X1 U12461 ( .B1(n21065), .B2(n11533), .A(n11532), .ZN(n11531) );
  INV_X1 U12462 ( .A(n20946), .ZN(n11532) );
  INV_X1 U12463 ( .A(n20931), .ZN(n11533) );
  NAND2_X1 U12464 ( .A1(n20944), .A2(n21065), .ZN(n20945) );
  NAND2_X1 U12465 ( .A1(n20929), .A2(n21065), .ZN(n20930) );
  NAND2_X1 U12466 ( .A1(n20930), .A2(n20931), .ZN(n20944) );
  INV_X1 U12467 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20705) );
  INV_X1 U12468 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18060) );
  INV_X1 U12469 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18107) );
  INV_X2 U12470 ( .A(n18037), .ZN(n18034) );
  NAND2_X1 U12471 ( .A1(n21226), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21225) );
  NAND2_X1 U12472 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(P3_EAX_REG_25__SCAN_IN), 
        .ZN(n11383) );
  NOR3_X1 U12473 ( .A1(n21197), .A2(n21244), .A3(n21159), .ZN(n21189) );
  INV_X1 U12474 ( .A(n18193), .ZN(n21275) );
  NOR2_X1 U12475 ( .A1(n21102), .A2(n21101), .ZN(n21103) );
  CLKBUF_X1 U12476 ( .A(n18681), .Z(n21770) );
  CLKBUF_X1 U12477 ( .A(n18685), .Z(n18689) );
  NOR3_X1 U12478 ( .A1(n21807), .A2(n21343), .A3(n20611), .ZN(n20652) );
  NOR2_X1 U12480 ( .A1(n21590), .A2(n21603), .ZN(n21646) );
  NOR2_X1 U12481 ( .A1(n18368), .A2(n21039), .ZN(n18442) );
  OR2_X1 U12482 ( .A1(n18623), .A2(n21353), .ZN(n18484) );
  NAND2_X1 U12483 ( .A1(n18219), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18302) );
  NOR2_X1 U12484 ( .A1(n18465), .A2(n21355), .ZN(n18359) );
  NAND2_X1 U12485 ( .A1(n21696), .A2(n18521), .ZN(n18465) );
  NAND2_X1 U12486 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18474), .ZN(
        n21525) );
  OAI21_X1 U12487 ( .B1(n18624), .B2(n18213), .A(n11527), .ZN(n18521) );
  INV_X1 U12488 ( .A(n21472), .ZN(n18213) );
  OR2_X1 U12489 ( .A1(n18484), .A2(n21469), .ZN(n11527) );
  NOR2_X2 U12490 ( .A1(n21359), .A2(n18623), .ZN(n18535) );
  INV_X1 U12491 ( .A(n18484), .ZN(n18536) );
  AND3_X1 U12492 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20717) );
  INV_X1 U12493 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18583) );
  NAND2_X1 U12494 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18581) );
  XNOR2_X1 U12495 ( .A(n18422), .B(n18421), .ZN(n21629) );
  OAI21_X2 U12496 ( .B1(n21357), .B2(n21315), .A(n21328), .ZN(n21754) );
  NAND2_X1 U12497 ( .A1(n21759), .A2(n21601), .ZN(n21732) );
  INV_X1 U12498 ( .A(n21636), .ZN(n21463) );
  INV_X1 U12499 ( .A(n21613), .ZN(n21721) );
  INV_X1 U12500 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21791) );
  CLKBUF_X1 U12501 ( .A(n19529), .Z(n19487) );
  NOR2_X1 U12502 ( .A1(n16286), .A2(n11375), .ZN(n16287) );
  NAND2_X1 U12503 ( .A1(n11377), .A2(n11376), .ZN(n11375) );
  AOI21_X1 U12504 ( .B1(n16559), .B2(n20519), .A(n16558), .ZN(n16560) );
  OR2_X1 U12505 ( .A1(n16478), .A2(n20496), .ZN(n11688) );
  OAI21_X1 U12506 ( .B1(n16713), .B2(n22141), .A(n12604), .ZN(n12605) );
  OAI21_X1 U12507 ( .B1(n20493), .B2(n22141), .A(n11360), .ZN(P1_U2988) );
  AOI21_X1 U12508 ( .B1(n22066), .B2(n20519), .A(n11361), .ZN(n11360) );
  NAND2_X1 U12509 ( .A1(n11363), .A2(n11362), .ZN(n11361) );
  AOI21_X1 U12510 ( .B1(n20514), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20494), .ZN(n11362) );
  AOI211_X1 U12511 ( .C1(n16225), .C2(n22017), .A(n16555), .B(n16224), .ZN(
        n16232) );
  INV_X1 U12512 ( .A(n11649), .ZN(n11685) );
  OAI21_X1 U12513 ( .B1(n19034), .B2(n19119), .A(n11650), .ZN(n11649) );
  NAND2_X1 U12514 ( .A1(n11463), .A2(n11459), .ZN(P2_U3020) );
  NAND2_X1 U12515 ( .A1(n17203), .A2(n19138), .ZN(n11463) );
  NOR2_X1 U12516 ( .A1(n17201), .A2(n11460), .ZN(n11459) );
  OAI21_X1 U12517 ( .B1(n11436), .B2(n17263), .A(n11435), .ZN(P2_U3026) );
  INV_X1 U12518 ( .A(n11399), .ZN(n11435) );
  OAI21_X1 U12519 ( .B1(n17286), .B2(n19134), .A(n11232), .ZN(n11399) );
  AOI21_X1 U12520 ( .B1(n11557), .B2(n21069), .A(n11556), .ZN(n21072) );
  XNOR2_X1 U12521 ( .A(n21076), .B(n11558), .ZN(n11557) );
  NAND2_X1 U12522 ( .A1(n21019), .A2(n21065), .ZN(n21020) );
  NOR2_X1 U12523 ( .A1(n21237), .A2(n21197), .ZN(n21232) );
  NAND2_X1 U12524 ( .A1(n11404), .A2(n21712), .ZN(n21607) );
  OAI21_X1 U12525 ( .B1(n21614), .B2(n11405), .A(n21757), .ZN(n11404) );
  OR2_X1 U12526 ( .A1(n20531), .A2(n20584), .ZN(U212) );
  BUF_X2 U12527 ( .A(n13188), .Z(n13479) );
  NOR2_X1 U12528 ( .A1(n16358), .A2(n16430), .ZN(n16346) );
  OR2_X1 U12529 ( .A1(n16382), .A2(n16381), .ZN(n11190) );
  NAND2_X1 U12530 ( .A1(n11578), .A2(n11581), .ZN(n16371) );
  INV_X1 U12531 ( .A(n11585), .ZN(n15831) );
  OR3_X1 U12532 ( .A1(n18465), .A2(n21594), .A3(n11305), .ZN(n11191) );
  INV_X1 U12533 ( .A(n15625), .ZN(n11623) );
  NOR2_X1 U12534 ( .A1(n14340), .A2(n14337), .ZN(n14472) );
  NAND2_X1 U12535 ( .A1(n11544), .A2(n11540), .ZN(n20864) );
  AND2_X1 U12536 ( .A1(n17546), .A2(n14245), .ZN(n13809) );
  AND2_X1 U12537 ( .A1(n15890), .A2(n11276), .ZN(n16945) );
  NAND2_X1 U12538 ( .A1(n15890), .A2(n11697), .ZN(n16044) );
  AND2_X1 U12539 ( .A1(n20863), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11195) );
  AND2_X1 U12540 ( .A1(n11470), .A2(n13461), .ZN(n11196) );
  AND2_X1 U12541 ( .A1(n16562), .A2(n11416), .ZN(n11197) );
  INV_X1 U12542 ( .A(n22066), .ZN(n20495) );
  NAND2_X1 U12543 ( .A1(n12820), .A2(n15241), .ZN(n13797) );
  INV_X1 U12544 ( .A(n13797), .ZN(n11402) );
  OR2_X1 U12545 ( .A1(n16358), .A2(n11576), .ZN(n11198) );
  AND3_X1 U12546 ( .A1(n17468), .A2(n17457), .A3(n11373), .ZN(n11199) );
  OR2_X1 U12547 ( .A1(n11501), .A2(n15769), .ZN(n11200) );
  AND2_X1 U12548 ( .A1(n11472), .A2(n13564), .ZN(n11201) );
  NAND2_X1 U12549 ( .A1(n11623), .A2(n15627), .ZN(n15743) );
  OR2_X1 U12550 ( .A1(n19535), .A2(n20665), .ZN(n11202) );
  AND2_X1 U12551 ( .A1(n11511), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11203) );
  AND2_X1 U12552 ( .A1(n11515), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11204) );
  AND2_X1 U12553 ( .A1(n11554), .A2(n11261), .ZN(n11205) );
  NAND2_X1 U12554 ( .A1(n11635), .A2(n11279), .ZN(n15200) );
  AND2_X1 U12555 ( .A1(n15627), .A2(n11622), .ZN(n11206) );
  AND2_X1 U12556 ( .A1(n11449), .A2(n16949), .ZN(n11207) );
  INV_X1 U12557 ( .A(n12039), .ZN(n12037) );
  AND2_X1 U12558 ( .A1(n11201), .A2(n11287), .ZN(n11208) );
  OR2_X1 U12559 ( .A1(n16966), .A2(n15212), .ZN(n16968) );
  AND2_X1 U12560 ( .A1(n11281), .A2(n11588), .ZN(n11209) );
  AND2_X1 U12561 ( .A1(n11504), .A2(n11503), .ZN(n11210) );
  AND2_X1 U12562 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11211) );
  AND2_X1 U12563 ( .A1(n11211), .A2(n13401), .ZN(n11212) );
  AND2_X1 U12564 ( .A1(n11380), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n11213) );
  OR2_X1 U12565 ( .A1(n20676), .A2(n14338), .ZN(n11214) );
  OR3_X1 U12566 ( .A1(n21237), .A2(n11383), .A3(n21197), .ZN(n11215) );
  INV_X1 U12567 ( .A(n11192), .ZN(n18133) );
  NAND2_X1 U12568 ( .A1(n11433), .A2(n12862), .ZN(n12885) );
  NAND2_X1 U12569 ( .A1(n13080), .A2(n11675), .ZN(n17098) );
  NAND2_X1 U12570 ( .A1(n13801), .A2(n11312), .ZN(n13815) );
  AND2_X1 U12571 ( .A1(n13933), .A2(n11713), .ZN(n11864) );
  NAND2_X1 U12572 ( .A1(n15593), .A2(n11587), .ZN(n15761) );
  AND2_X1 U12573 ( .A1(n12903), .A2(n12899), .ZN(n13027) );
  OR2_X1 U12574 ( .A1(n13639), .A2(n13716), .ZN(n11216) );
  AND2_X1 U12575 ( .A1(n21226), .A2(n11380), .ZN(n11217) );
  AND4_X1 U12576 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11860) );
  INV_X1 U12577 ( .A(n11836), .ZN(n11571) );
  NOR2_X1 U12578 ( .A1(n21333), .A2(n20684), .ZN(n18058) );
  INV_X1 U12579 ( .A(n18058), .ZN(n14351) );
  AND2_X1 U12580 ( .A1(n11567), .A2(n12538), .ZN(n11219) );
  NAND2_X1 U12581 ( .A1(n16584), .A2(n16604), .ZN(n13658) );
  NAND2_X1 U12582 ( .A1(n11665), .A2(n13454), .ZN(n17157) );
  AND2_X2 U12583 ( .A1(n12903), .A2(n12906), .ZN(n12985) );
  NAND2_X1 U12584 ( .A1(n12862), .A2(n12843), .ZN(n11220) );
  NAND2_X1 U12585 ( .A1(n11340), .A2(n11397), .ZN(n15681) );
  NAND2_X1 U12586 ( .A1(n11656), .A2(n17096), .ZN(n17224) );
  OR2_X1 U12587 ( .A1(n13074), .A2(n17153), .ZN(n11221) );
  AND2_X1 U12588 ( .A1(n13559), .A2(n13558), .ZN(n17240) );
  NAND2_X1 U12589 ( .A1(n12975), .A2(n12974), .ZN(n11222) );
  NAND2_X1 U12590 ( .A1(n18407), .A2(n18397), .ZN(n18613) );
  AND4_X1 U12591 ( .A1(n14400), .A2(n14399), .A3(n14398), .A4(n14397), .ZN(
        n11223) );
  XNOR2_X1 U12592 ( .A(n11593), .B(n11592), .ZN(n16278) );
  AND2_X1 U12593 ( .A1(n11668), .A2(n11438), .ZN(n11224) );
  AND2_X1 U12594 ( .A1(n17630), .A2(n13612), .ZN(n11225) );
  NAND2_X1 U12595 ( .A1(n16948), .A2(n11207), .ZN(n11450) );
  AND4_X1 U12596 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11226) );
  AND2_X1 U12597 ( .A1(n13454), .A2(n11663), .ZN(n11227) );
  AND2_X1 U12598 ( .A1(n13454), .A2(n11669), .ZN(n11228) );
  NAND2_X2 U12599 ( .A1(n11660), .A2(n11659), .ZN(n13389) );
  AND2_X1 U12600 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11229) );
  OR2_X1 U12601 ( .A1(n14351), .A2(n18107), .ZN(n11230) );
  AND2_X1 U12602 ( .A1(n11443), .A2(n14260), .ZN(n11231) );
  AND2_X1 U12603 ( .A1(n11464), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12762) );
  NOR2_X1 U12604 ( .A1(n17285), .A2(n17284), .ZN(n11232) );
  NAND2_X1 U12605 ( .A1(n18315), .A2(n18619), .ZN(n18407) );
  INV_X1 U12606 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11702) );
  INV_X1 U12607 ( .A(n11347), .ZN(n13018) );
  INV_X1 U12608 ( .A(n16382), .ZN(n11578) );
  NOR2_X1 U12609 ( .A1(n16358), .A2(n11573), .ZN(n16325) );
  NOR2_X1 U12610 ( .A1(n16382), .A2(n11583), .ZN(n16370) );
  AND2_X1 U12611 ( .A1(n11604), .A2(n18110), .ZN(n11233) );
  INV_X1 U12612 ( .A(n15608), .ZN(n11423) );
  INV_X1 U12613 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17578) );
  OR2_X1 U12614 ( .A1(n16240), .A2(n17676), .ZN(n11234) );
  INV_X1 U12615 ( .A(n18048), .ZN(n21315) );
  AOI21_X1 U12616 ( .B1(n17453), .B2(n17452), .A(n17485), .ZN(n18048) );
  AND2_X1 U12617 ( .A1(n14224), .A2(n14228), .ZN(n14250) );
  AND2_X1 U12618 ( .A1(n11862), .A2(n11320), .ZN(n11235) );
  AND2_X1 U12619 ( .A1(n13525), .A2(n11472), .ZN(n11236) );
  AND2_X1 U12620 ( .A1(n15092), .A2(n11838), .ZN(n11237) );
  NAND2_X1 U12621 ( .A1(n12579), .A2(n13802), .ZN(n11238) );
  INV_X1 U12622 ( .A(n13603), .ZN(n15234) );
  INV_X1 U12623 ( .A(n13078), .ZN(n11681) );
  OR2_X1 U12624 ( .A1(n13060), .A2(n13077), .ZN(n13078) );
  INV_X1 U12625 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11328) );
  NOR2_X1 U12626 ( .A1(n16638), .A2(n20516), .ZN(n11239) );
  AND2_X2 U12627 ( .A1(n11719), .A2(n14191), .ZN(n11870) );
  AND2_X2 U12628 ( .A1(n16134), .A2(n14603), .ZN(n12944) );
  INV_X1 U12629 ( .A(n13455), .ZN(n13507) );
  NAND2_X1 U12630 ( .A1(n13236), .A2(n13235), .ZN(n17391) );
  AND2_X2 U12631 ( .A1(n12449), .A2(n11178), .ZN(n15657) );
  AND2_X1 U12632 ( .A1(n11623), .A2(n11206), .ZN(n11240) );
  INV_X1 U12633 ( .A(n12832), .ZN(n13380) );
  NOR2_X1 U12634 ( .A1(n17026), .A2(n17239), .ZN(n17016) );
  AND2_X1 U12635 ( .A1(n16434), .A2(n11210), .ZN(n11241) );
  OR2_X1 U12636 ( .A1(n15749), .A2(n11641), .ZN(n11242) );
  NAND2_X1 U12637 ( .A1(n22124), .A2(n11381), .ZN(n11243) );
  OR2_X1 U12638 ( .A1(n18985), .A2(n13507), .ZN(n11244) );
  AND2_X1 U12639 ( .A1(n17652), .A2(n11511), .ZN(n11245) );
  AND2_X1 U12640 ( .A1(n19060), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11246) );
  OR2_X1 U12641 ( .A1(n17315), .A2(n15749), .ZN(n11247) );
  NOR2_X2 U12642 ( .A1(n21359), .A2(n21637), .ZN(n18492) );
  INV_X1 U12643 ( .A(n18492), .ZN(n18416) );
  AND2_X1 U12644 ( .A1(n11477), .A2(n11476), .ZN(n11248) );
  AND2_X1 U12645 ( .A1(n11647), .A2(n15561), .ZN(n11249) );
  AND2_X1 U12646 ( .A1(n15615), .A2(n15629), .ZN(n15628) );
  AND2_X1 U12647 ( .A1(n15546), .A2(n15616), .ZN(n15615) );
  NOR2_X1 U12648 ( .A1(n15545), .A2(n15544), .ZN(n15546) );
  AND2_X1 U12649 ( .A1(n15890), .A2(n11619), .ZN(n16955) );
  AND2_X1 U12650 ( .A1(n16459), .A2(n11483), .ZN(n11250) );
  AND2_X1 U12651 ( .A1(n11453), .A2(n15265), .ZN(n11251) );
  AND2_X1 U12652 ( .A1(n11458), .A2(n15792), .ZN(n11252) );
  AND2_X1 U12653 ( .A1(n11668), .A2(n11667), .ZN(n17143) );
  INV_X1 U12654 ( .A(n16779), .ZN(n16778) );
  AND2_X1 U12655 ( .A1(n13451), .A2(n11470), .ZN(n11253) );
  AND2_X1 U12656 ( .A1(n11667), .A2(n17144), .ZN(n11254) );
  XNOR2_X1 U12657 ( .A(n16929), .B(n16081), .ZN(n16921) );
  OR2_X1 U12658 ( .A1(n15553), .A2(n11519), .ZN(n11255) );
  OR2_X1 U12659 ( .A1(n16337), .A2(n16328), .ZN(n11256) );
  OR2_X1 U12660 ( .A1(n21101), .A2(n21807), .ZN(n11257) );
  NAND2_X1 U12661 ( .A1(n12449), .A2(n14565), .ZN(n13821) );
  INV_X1 U12662 ( .A(n13821), .ZN(n11570) );
  NAND2_X1 U12663 ( .A1(n14060), .A2(n14059), .ZN(n14267) );
  NAND2_X1 U12664 ( .A1(n15593), .A2(n11209), .ZN(n11585) );
  OR2_X1 U12665 ( .A1(n16779), .A2(n16726), .ZN(n11258) );
  INV_X1 U12666 ( .A(n11586), .ZN(n15763) );
  NAND2_X1 U12667 ( .A1(n15593), .A2(n15656), .ZN(n11586) );
  AND2_X1 U12668 ( .A1(n11448), .A2(n11447), .ZN(n11259) );
  AND2_X1 U12669 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11260) );
  AND2_X1 U12670 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11261) );
  INV_X1 U12671 ( .A(n11537), .ZN(n11536) );
  AND2_X1 U12672 ( .A1(n11195), .A2(n11538), .ZN(n11537) );
  INV_X1 U12673 ( .A(n11501), .ZN(n11500) );
  OR2_X1 U12674 ( .A1(n15599), .A2(n11502), .ZN(n11501) );
  INV_X1 U12675 ( .A(n17155), .ZN(n11669) );
  NAND2_X1 U12676 ( .A1(n13566), .A2(n17232), .ZN(n11262) );
  AND2_X1 U12677 ( .A1(n14319), .A2(n11453), .ZN(n11263) );
  AND2_X1 U12678 ( .A1(n16959), .A2(n16958), .ZN(n16948) );
  INV_X1 U12679 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11419) );
  AND2_X1 U12680 ( .A1(n11481), .A2(n11480), .ZN(n11264) );
  AND2_X1 U12681 ( .A1(n21721), .A2(n21606), .ZN(n11265) );
  AND2_X1 U12682 ( .A1(n17122), .A2(n17301), .ZN(n11266) );
  AND2_X1 U12683 ( .A1(n11456), .A2(n11455), .ZN(n11267) );
  AND2_X1 U12684 ( .A1(n11248), .A2(n11475), .ZN(n11268) );
  AND2_X1 U12685 ( .A1(n11249), .A2(n11646), .ZN(n11269) );
  AND2_X1 U12686 ( .A1(n11438), .A2(n13607), .ZN(n11270) );
  OR2_X1 U12687 ( .A1(n17315), .A2(n11639), .ZN(n11271) );
  INV_X1 U12688 ( .A(n14035), .ZN(n14091) );
  NOR2_X2 U12689 ( .A1(n14028), .A2(n11828), .ZN(n11272) );
  OR2_X1 U12690 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13688) );
  INV_X1 U12691 ( .A(n13507), .ZN(n13749) );
  NAND2_X1 U12692 ( .A1(n16071), .A2(n16097), .ZN(n11273) );
  AND2_X1 U12693 ( .A1(n18219), .A2(n11554), .ZN(n11274) );
  AND2_X1 U12694 ( .A1(n18791), .A2(n11647), .ZN(n15560) );
  AND2_X1 U12695 ( .A1(n12756), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13303) );
  INV_X1 U12696 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19787) );
  NOR2_X1 U12697 ( .A1(n14606), .A2(n12832), .ZN(n13181) );
  AND2_X1 U12698 ( .A1(n17669), .A2(n11515), .ZN(n11275) );
  NAND2_X1 U12699 ( .A1(n13232), .A2(n13231), .ZN(n17403) );
  OR2_X1 U12700 ( .A1(n13212), .A2(n13209), .ZN(n14136) );
  AND2_X1 U12701 ( .A1(n11619), .A2(n16957), .ZN(n11276) );
  AND2_X1 U12702 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11277) );
  AND2_X1 U12703 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11278) );
  OR3_X1 U12704 ( .A1(n11390), .A2(n14368), .A3(n14367), .ZN(n21341) );
  NOR2_X1 U12705 ( .A1(n14258), .A2(n11628), .ZN(n14322) );
  NAND2_X1 U12706 ( .A1(n15454), .A2(n15453), .ZN(n15598) );
  INV_X1 U12707 ( .A(n15598), .ZN(n11499) );
  AND2_X1 U12708 ( .A1(n11636), .A2(n15197), .ZN(n11279) );
  OR2_X1 U12709 ( .A1(n16210), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11280) );
  AND2_X1 U12710 ( .A1(n15832), .A2(n15827), .ZN(n11281) );
  OR2_X1 U12711 ( .A1(n12768), .A2(n12767), .ZN(n13222) );
  INV_X1 U12712 ( .A(n14236), .ZN(n13099) );
  AND2_X1 U12713 ( .A1(n11209), .A2(n15851), .ZN(n11282) );
  AND2_X1 U12714 ( .A1(n11276), .A2(n16947), .ZN(n11283) );
  AND2_X1 U12715 ( .A1(n11210), .A2(n16350), .ZN(n11284) );
  NOR2_X1 U12716 ( .A1(n14676), .A2(n14677), .ZN(n11285) );
  AND2_X1 U12717 ( .A1(n11837), .A2(n15092), .ZN(n11286) );
  BUF_X1 U12718 ( .A(n11167), .Z(n16099) );
  OR2_X1 U12719 ( .A1(n13448), .A2(n16932), .ZN(n11287) );
  NAND2_X1 U12720 ( .A1(n13355), .A2(n13354), .ZN(n11288) );
  AND2_X1 U12721 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11289) );
  AND2_X1 U12722 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11290) );
  AND2_X1 U12723 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11291) );
  AND2_X1 U12724 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11292) );
  AND2_X1 U12725 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11293) );
  AND2_X1 U12726 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11294) );
  OR2_X1 U12727 ( .A1(n13448), .A2(n13594), .ZN(n11295) );
  AND3_X1 U12728 ( .A1(n18504), .A2(n18268), .A3(n21484), .ZN(n11296) );
  INV_X1 U12729 ( .A(n16381), .ZN(n11584) );
  AND2_X1 U12730 ( .A1(n21538), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11297) );
  AND2_X1 U12731 ( .A1(n13365), .A2(n13364), .ZN(n11298) );
  NAND2_X1 U12732 ( .A1(n18442), .A2(n11547), .ZN(n11551) );
  AND2_X1 U12733 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11299) );
  AND2_X1 U12734 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11300) );
  AND2_X1 U12735 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11301) );
  INV_X1 U12736 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19807) );
  INV_X1 U12737 ( .A(n20519), .ZN(n20496) );
  AND2_X1 U12738 ( .A1(n12448), .A2(n15381), .ZN(n20519) );
  AND2_X1 U12739 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11302) );
  AND2_X1 U12740 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11303) );
  AND2_X1 U12741 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U12742 ( .A1(n20806), .A2(n18540), .ZN(n18497) );
  INV_X1 U12743 ( .A(n18497), .ZN(n11539) );
  OR3_X1 U12744 ( .A1(n21355), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n21602), .ZN(n11305) );
  AND2_X1 U12745 ( .A1(n11381), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n11306) );
  AND2_X1 U12746 ( .A1(n16615), .A2(n21995), .ZN(n11307) );
  INV_X1 U12747 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11357) );
  AND2_X1 U12748 ( .A1(n11675), .A2(n17231), .ZN(n11308) );
  AND2_X1 U12749 ( .A1(n11212), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11309) );
  INV_X1 U12750 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11464) );
  AND2_X1 U12751 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11310) );
  INV_X1 U12752 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11549) );
  INV_X1 U12753 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n11382) );
  INV_X1 U12754 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n11384) );
  INV_X1 U12755 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11550) );
  INV_X1 U12756 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11513) );
  INV_X1 U12757 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11517) );
  NOR2_X1 U12758 ( .A1(n11202), .A2(n11257), .ZN(n18039) );
  NOR2_X1 U12759 ( .A1(n14361), .A2(n14360), .ZN(n19535) );
  INV_X1 U12760 ( .A(n21341), .ZN(n20665) );
  AOI22_X1 U12761 ( .A1(n21348), .A2(n18050), .B1(n17452), .B2(n14435), .ZN(
        n21101) );
  AOI21_X1 U12762 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11302), .ZN(n16127) );
  AOI21_X1 U12763 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n11303), .ZN(n16137) );
  AOI21_X1 U12764 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n11304), .ZN(n16114) );
  AOI21_X1 U12765 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n11289), .ZN(n16022) );
  AOI21_X1 U12766 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n11290), .ZN(n16029) );
  AOI21_X1 U12767 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n11291), .ZN(n16005) );
  AOI21_X1 U12768 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n11292), .ZN(n16013) );
  AOI21_X1 U12769 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n11293), .ZN(n15996) );
  AOI21_X1 U12770 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n11294), .ZN(n15988) );
  AOI21_X1 U12771 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n11277), .ZN(n15968) );
  AOI21_X1 U12772 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n11278), .ZN(n15976) );
  AOI21_X1 U12773 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n11299), .ZN(n15951) );
  AOI21_X1 U12774 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n11300), .ZN(n15934) );
  AOI21_X1 U12775 ( .B1(n15970), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n11301), .ZN(n15941) );
  INV_X1 U12776 ( .A(n21269), .ZN(n21280) );
  AOI22_X2 U12777 ( .A1(DATAI_28_), .A2(n11152), .B1(BUF1_REG_28__SCAN_IN), 
        .B2(n22474), .ZN(n22432) );
  AOI22_X2 U12778 ( .A1(DATAI_22_), .A2(n11152), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n22474), .ZN(n22473) );
  AOI22_X2 U12779 ( .A1(DATAI_23_), .A2(n11152), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n22474), .ZN(n22581) );
  AOI22_X2 U12780 ( .A1(DATAI_16_), .A2(n11152), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n22474), .ZN(n22302) );
  AOI22_X2 U12781 ( .A1(DATAI_19_), .A2(n11152), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n22474), .ZN(n22382) );
  AOI22_X2 U12782 ( .A1(DATAI_18_), .A2(n11152), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n22474), .ZN(n22359) );
  NOR4_X2 U12783 ( .A1(n17472), .A2(n21104), .A3(n17471), .A4(n21345), .ZN(
        n21789) );
  AOI21_X1 U12784 ( .B1(n17474), .B2(n20611), .A(n21343), .ZN(n21104) );
  NAND2_X1 U12785 ( .A1(n19532), .A2(n19241), .ZN(n19324) );
  AOI22_X2 U12786 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n11151), .ZN(n19853) );
  NAND2_X1 U12787 ( .A1(n11337), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U12788 ( .A1(n11337), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U12789 ( .A1(n11337), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n13170) );
  NAND2_X1 U12790 ( .A1(n11337), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n13164) );
  NAND2_X1 U12791 ( .A1(n11337), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13084) );
  NAND2_X1 U12792 ( .A1(n11337), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n13160) );
  NAND2_X1 U12793 ( .A1(n11337), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13153) );
  NAND2_X1 U12794 ( .A1(n11337), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U12795 ( .A1(n11337), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13141) );
  NAND2_X1 U12796 ( .A1(n11337), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U12797 ( .A1(n11337), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13147) );
  NAND2_X1 U12798 ( .A1(n11337), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13126) );
  NAND2_X1 U12799 ( .A1(n11337), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13122) );
  NAND2_X1 U12800 ( .A1(n11337), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13117) );
  NAND2_X1 U12801 ( .A1(n11337), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U12802 ( .A1(n11337), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13114) );
  NAND2_X1 U12803 ( .A1(n11337), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13101) );
  AOI22_X2 U12804 ( .A1(DATAI_21_), .A2(n11152), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n22474), .ZN(n22459) );
  NAND3_X1 U12805 ( .A1(n11836), .A2(n11832), .A3(n14565), .ZN(n11311) );
  AND3_X2 U12806 ( .A1(n11317), .A2(n11315), .A3(n11313), .ZN(n13801) );
  NAND2_X1 U12807 ( .A1(n11836), .A2(n15092), .ZN(n16272) );
  NAND2_X2 U12808 ( .A1(n20481), .A2(n12504), .ZN(n20489) );
  NAND2_X1 U12809 ( .A1(n14169), .A2(n12462), .ZN(n12469) );
  NAND3_X1 U12810 ( .A1(n11319), .A2(n11895), .A3(n22153), .ZN(n11323) );
  NAND2_X1 U12811 ( .A1(n11854), .A2(n11235), .ZN(n11319) );
  NAND2_X1 U12812 ( .A1(n11862), .A2(n14062), .ZN(n11321) );
  NAND2_X1 U12813 ( .A1(n11854), .A2(n11853), .ZN(n11322) );
  NAND2_X2 U12814 ( .A1(n15772), .A2(n15771), .ZN(n16676) );
  AND2_X2 U12815 ( .A1(n11326), .A2(n13661), .ZN(n16570) );
  OAI21_X1 U12816 ( .B1(n16576), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11326), .ZN(n16733) );
  OAI21_X1 U12817 ( .B1(n11326), .B2(n11418), .A(n20516), .ZN(n16152) );
  OAI211_X1 U12818 ( .C1(n11326), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11414), .B(n11325), .ZN(n13662) );
  NAND2_X1 U12819 ( .A1(n11326), .A2(n20516), .ZN(n11325) );
  NAND2_X2 U12820 ( .A1(n16576), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U12821 ( .A1(n12891), .A2(n11327), .ZN(n14615) );
  NAND3_X2 U12822 ( .A1(n11328), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16131) );
  MUX2_X1 U12823 ( .A(n14617), .B(n14618), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14619) );
  NAND2_X1 U12824 ( .A1(n11329), .A2(n12912), .ZN(n12974) );
  OAI21_X1 U12825 ( .B1(n11331), .B2(n11330), .A(n19060), .ZN(n11329) );
  NAND4_X1 U12826 ( .A1(n12910), .A2(n12894), .A3(n12908), .A4(n12909), .ZN(
        n11330) );
  NAND4_X1 U12827 ( .A1(n12896), .A2(n12911), .A3(n12897), .A4(n12895), .ZN(
        n11331) );
  NAND2_X1 U12828 ( .A1(n11332), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12734) );
  NAND3_X1 U12829 ( .A1(n12724), .A2(n11226), .A3(n12725), .ZN(n11332) );
  NAND2_X1 U12830 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U12831 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11336) );
  CLKBUF_X1 U12832 ( .A(n12856), .Z(n11337) );
  NAND2_X1 U12833 ( .A1(n11338), .A2(n11339), .ZN(n11395) );
  NAND3_X1 U12834 ( .A1(n13053), .A2(n13051), .A3(n13058), .ZN(n11338) );
  INV_X1 U12835 ( .A(n11396), .ZN(n11340) );
  AND2_X2 U12836 ( .A1(n11342), .A2(n11341), .ZN(n20069) );
  NAND2_X2 U12837 ( .A1(n12880), .A2(n12881), .ZN(n11401) );
  NAND3_X1 U12838 ( .A1(n13385), .A2(n11349), .A3(n12811), .ZN(n11348) );
  NAND3_X1 U12839 ( .A1(n11351), .A2(n15234), .A3(n11350), .ZN(n11349) );
  NAND3_X1 U12840 ( .A1(n12804), .A2(n12805), .A3(n12803), .ZN(n11351) );
  AND2_X2 U12841 ( .A1(n11668), .A2(n11254), .ZN(n17584) );
  NAND2_X2 U12842 ( .A1(n11670), .A2(n11227), .ZN(n11668) );
  NAND3_X1 U12843 ( .A1(n12661), .A2(n12662), .A3(n12664), .ZN(n11352) );
  NAND3_X1 U12844 ( .A1(n12660), .A2(n12657), .A3(n12658), .ZN(n11354) );
  NOR2_X1 U12845 ( .A1(n17077), .A2(n13577), .ZN(n17050) );
  NAND3_X1 U12846 ( .A1(n13019), .A2(n13507), .A3(n13049), .ZN(n13422) );
  AND2_X1 U12847 ( .A1(n13019), .A2(n13049), .ZN(n13020) );
  OAI21_X1 U12848 ( .B1(n14330), .B2(n14331), .A(n11359), .ZN(n21903) );
  NAND2_X1 U12849 ( .A1(n16676), .A2(n16778), .ZN(n11364) );
  NAND2_X1 U12850 ( .A1(n12453), .A2(n11893), .ZN(n11894) );
  INV_X1 U12851 ( .A(n12453), .ZN(n11367) );
  INV_X1 U12852 ( .A(n11893), .ZN(n11370) );
  NAND2_X1 U12853 ( .A1(n11842), .A2(n15283), .ZN(n11843) );
  NAND2_X4 U12854 ( .A1(n11193), .A2(n11164), .ZN(n14245) );
  NAND3_X1 U12855 ( .A1(n11855), .A2(n13828), .A3(n11845), .ZN(n11372) );
  NAND2_X1 U12856 ( .A1(n16302), .A2(n11374), .ZN(n11379) );
  NAND2_X1 U12857 ( .A1(n11379), .A2(n11378), .ZN(n11377) );
  INV_X1 U12858 ( .A(n21198), .ZN(n21231) );
  NAND2_X1 U12859 ( .A1(n11387), .A2(n11386), .ZN(n11385) );
  NAND2_X1 U12860 ( .A1(n11388), .A2(n11238), .ZN(n11387) );
  NAND2_X1 U12861 ( .A1(n12581), .A2(n12580), .ZN(n11388) );
  NAND3_X1 U12862 ( .A1(n11193), .A2(n11164), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11948) );
  XNOR2_X2 U12863 ( .A(n11394), .B(n12975), .ZN(n15466) );
  AND2_X2 U12864 ( .A1(n11393), .A2(n12964), .ZN(n12975) );
  NAND3_X1 U12865 ( .A1(n12927), .A2(n12925), .A3(n12926), .ZN(n11393) );
  NAND2_X2 U12866 ( .A1(n11401), .A2(n11658), .ZN(n13089) );
  NAND2_X2 U12867 ( .A1(n12884), .A2(n11401), .ZN(n15322) );
  AND2_X4 U12868 ( .A1(n12762), .A2(n14598), .ZN(n12753) );
  AOI22_X1 U12869 ( .A1(n12753), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n12756), .ZN(n12664) );
  NOR2_X2 U12870 ( .A1(n19113), .A2(n17316), .ZN(n17636) );
  NOR2_X2 U12871 ( .A1(n21520), .A2(n21534), .ZN(n21698) );
  NAND2_X1 U12872 ( .A1(n11412), .A2(n11411), .ZN(n12040) );
  AND2_X4 U12873 ( .A1(n14191), .A2(n11718), .ZN(n11769) );
  NAND2_X1 U12874 ( .A1(n11837), .A2(n11237), .ZN(n11840) );
  AND2_X1 U12875 ( .A1(n11286), .A2(n12595), .ZN(n13825) );
  NAND2_X2 U12876 ( .A1(n11422), .A2(n11420), .ZN(n15772) );
  NAND2_X1 U12877 ( .A1(n20489), .A2(n20488), .ZN(n20487) );
  OAI21_X2 U12878 ( .B1(n12830), .B2(n11429), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11428) );
  OAI21_X1 U12879 ( .B1(n17132), .B2(n11432), .A(n11430), .ZN(n17644) );
  INV_X1 U12880 ( .A(n17644), .ZN(n13614) );
  OR2_X1 U12881 ( .A1(n19091), .A2(n17264), .ZN(n11436) );
  NAND2_X1 U12882 ( .A1(n17304), .A2(n11266), .ZN(n13617) );
  NAND2_X1 U12883 ( .A1(n11668), .A2(n11270), .ZN(n11437) );
  NAND2_X1 U12884 ( .A1(n11437), .A2(n13608), .ZN(n17345) );
  NAND2_X1 U12885 ( .A1(n13089), .A2(n13088), .ZN(n13094) );
  AND2_X4 U12886 ( .A1(n11439), .A2(n11464), .ZN(n12756) );
  INV_X1 U12887 ( .A(n14237), .ZN(n11442) );
  INV_X1 U12888 ( .A(n11450), .ZN(n16933) );
  NAND3_X1 U12889 ( .A1(n13451), .A2(n11196), .A3(n13470), .ZN(n13472) );
  NAND2_X1 U12890 ( .A1(n13525), .A2(n11208), .ZN(n13576) );
  NAND2_X1 U12891 ( .A1(n13525), .A2(n13524), .ZN(n13563) );
  MUX2_X1 U12892 ( .A(n13218), .B(n12786), .S(n13603), .Z(n13417) );
  NAND3_X1 U12893 ( .A1(n16206), .A2(n15657), .A3(n14147), .ZN(n14060) );
  NAND2_X1 U12894 ( .A1(n11479), .A2(n16432), .ZN(n16188) );
  NAND2_X1 U12895 ( .A1(n11479), .A2(n16422), .ZN(n16198) );
  NAND2_X1 U12896 ( .A1(n11479), .A2(n14329), .ZN(n14272) );
  NAND2_X1 U12897 ( .A1(n11479), .A2(n15588), .ZN(n14681) );
  NAND2_X1 U12898 ( .A1(n11479), .A2(n15462), .ZN(n15450) );
  NAND2_X1 U12899 ( .A1(n11479), .A2(n15695), .ZN(n15660) );
  NAND2_X1 U12900 ( .A1(n11479), .A2(n22078), .ZN(n15836) );
  NAND2_X1 U12901 ( .A1(n11479), .A2(n15878), .ZN(n15866) );
  NAND2_X1 U12902 ( .A1(n11479), .A2(n16452), .ZN(n16174) );
  NAND2_X1 U12903 ( .A1(n11479), .A2(n16448), .ZN(n16168) );
  INV_X1 U12904 ( .A(n16303), .ZN(n11491) );
  INV_X1 U12905 ( .A(n14676), .ZN(n11493) );
  NAND3_X1 U12906 ( .A1(n11493), .A2(n15330), .A3(n11494), .ZN(n15452) );
  NAND2_X1 U12907 ( .A1(n16434), .A2(n11284), .ZN(n16349) );
  NAND2_X1 U12908 ( .A1(n11506), .A2(n17412), .ZN(n18956) );
  OAI211_X1 U12909 ( .C1(n18948), .C2(n18949), .A(n11506), .B(n19003), .ZN(
        n18950) );
  OAI211_X1 U12910 ( .C1(n11507), .C2(n18888), .A(n18899), .B(n19003), .ZN(
        n18889) );
  NOR2_X2 U12911 ( .A1(n17448), .A2(n19325), .ZN(n21283) );
  AND2_X2 U12912 ( .A1(n17474), .A2(n18048), .ZN(n21759) );
  NAND2_X1 U12913 ( .A1(n18431), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11526) );
  OR3_X1 U12914 ( .A1(n18465), .A2(n21355), .A3(n21594), .ZN(n18429) );
  NAND2_X1 U12915 ( .A1(n11191), .A2(n11526), .ZN(n18432) );
  NAND2_X2 U12916 ( .A1(n21613), .A2(n20665), .ZN(n21644) );
  INV_X1 U12917 ( .A(n11551), .ZN(n18443) );
  AND2_X1 U12918 ( .A1(n21065), .A2(n21064), .ZN(n21076) );
  NAND2_X1 U12919 ( .A1(n21059), .A2(n21060), .ZN(n21064) );
  OR2_X2 U12920 ( .A1(n11559), .A2(n11895), .ZN(n11937) );
  NOR2_X1 U12921 ( .A1(n14523), .A2(n11559), .ZN(n15349) );
  XNOR2_X2 U12922 ( .A(n11851), .B(n11934), .ZN(n11559) );
  NOR2_X4 U12923 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11719) );
  AND2_X2 U12924 ( .A1(n11719), .A2(n13935), .ZN(n12237) );
  NOR2_X4 U12925 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13935) );
  NAND3_X1 U12926 ( .A1(n16584), .A2(n16604), .A3(n13659), .ZN(n13660) );
  INV_X1 U12927 ( .A(n11561), .ZN(n11560) );
  NAND3_X1 U12928 ( .A1(n16584), .A2(n16604), .A3(n11563), .ZN(n11562) );
  INV_X1 U12929 ( .A(n15092), .ZN(n22476) );
  NAND2_X1 U12930 ( .A1(n11570), .A2(n15092), .ZN(n11569) );
  NAND2_X1 U12931 ( .A1(n11572), .A2(n11571), .ZN(n15080) );
  INV_X1 U12932 ( .A(n14076), .ZN(n11572) );
  NAND2_X1 U12933 ( .A1(n14532), .A2(n11838), .ZN(n14076) );
  OR2_X2 U12934 ( .A1(n16358), .A2(n11574), .ZN(n16313) );
  NOR2_X2 U12935 ( .A1(n16382), .A2(n11579), .ZN(n16357) );
  AND2_X2 U12936 ( .A1(n15593), .A2(n11282), .ZN(n15850) );
  NAND2_X1 U12937 ( .A1(n12446), .A2(n11590), .ZN(n11593) );
  NAND2_X1 U12938 ( .A1(n12446), .A2(n12447), .ZN(n16290) );
  INV_X1 U12939 ( .A(n11593), .ZN(n16289) );
  XNOR2_X2 U12940 ( .A(n12002), .B(n15118), .ZN(n14569) );
  OR2_X2 U12941 ( .A1(n11963), .A2(n11962), .ZN(n12002) );
  NOR2_X1 U12942 ( .A1(n11597), .A2(n11594), .ZN(n11598) );
  NAND3_X1 U12943 ( .A1(n18111), .A2(n11596), .A3(n11595), .ZN(n11594) );
  NAND2_X1 U12944 ( .A1(n18116), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11606) );
  NAND3_X1 U12945 ( .A1(n18351), .A2(n18341), .A3(n11310), .ZN(n18373) );
  AND2_X2 U12946 ( .A1(n18282), .A2(n11297), .ZN(n18341) );
  NOR2_X2 U12948 ( .A1(n18181), .A2(n11609), .ZN(n18457) );
  AND2_X2 U12949 ( .A1(n11611), .A2(n18416), .ZN(n18181) );
  INV_X2 U12950 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21296) );
  OR2_X1 U12951 ( .A1(n16929), .A2(n16082), .ZN(n11612) );
  NAND2_X1 U12952 ( .A1(n16921), .A2(n16923), .ZN(n16922) );
  NAND2_X1 U12953 ( .A1(n11661), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12853) );
  NAND2_X1 U12954 ( .A1(n16912), .A2(n11613), .ZN(n16904) );
  NAND3_X1 U12955 ( .A1(n11614), .A2(n16897), .A3(n16904), .ZN(n16119) );
  OAI21_X1 U12956 ( .B1(n16091), .B2(n11617), .A(n16905), .ZN(n11616) );
  INV_X1 U12957 ( .A(n16098), .ZN(n11617) );
  NAND2_X1 U12958 ( .A1(n11618), .A2(n16098), .ZN(n16895) );
  NAND2_X1 U12959 ( .A1(n15890), .A2(n11283), .ZN(n16939) );
  NAND4_X1 U12960 ( .A1(n20069), .A2(n12815), .A3(n19967), .A4(n13389), .ZN(
        n12738) );
  INV_X2 U12961 ( .A(n13381), .ZN(n19967) );
  NAND2_X2 U12962 ( .A1(n12734), .A2(n12733), .ZN(n12740) );
  INV_X2 U12963 ( .A(n13389), .ZN(n12745) );
  NAND2_X1 U12964 ( .A1(n13188), .A2(n14153), .ZN(n12826) );
  INV_X1 U12965 ( .A(n12888), .ZN(n11625) );
  INV_X1 U12966 ( .A(n11693), .ZN(n11629) );
  NAND3_X1 U12967 ( .A1(n11632), .A2(n11635), .A3(n15233), .ZN(n13232) );
  INV_X1 U12968 ( .A(n13212), .ZN(n11636) );
  NAND3_X1 U12969 ( .A1(n13561), .A2(n13560), .A3(n11262), .ZN(n11656) );
  XNOR2_X1 U12970 ( .A(n11657), .B(n17097), .ZN(n17238) );
  NAND2_X1 U12971 ( .A1(n12700), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11659) );
  NAND2_X1 U12972 ( .A1(n11661), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12867) );
  NAND2_X1 U12973 ( .A1(n16239), .A2(n11234), .ZN(P2_U2983) );
  CLKBUF_X1 U12974 ( .A(n11670), .Z(n11665) );
  NAND2_X1 U12975 ( .A1(n13559), .A2(n13558), .ZN(n13554) );
  NAND2_X1 U12976 ( .A1(n11676), .A2(n11679), .ZN(n13624) );
  NAND3_X1 U12977 ( .A1(n17152), .A2(n13075), .A3(n13078), .ZN(n11676) );
  NAND2_X1 U12978 ( .A1(n13081), .A2(n11309), .ZN(n13717) );
  NAND2_X1 U12979 ( .A1(n13081), .A2(n11211), .ZN(n17075) );
  NOR2_X1 U12980 ( .A1(n13656), .A2(n11683), .ZN(n13657) );
  NOR2_X2 U12981 ( .A1(n11702), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11711) );
  NOR2_X1 U12982 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11713) );
  NAND2_X1 U12983 ( .A1(n11937), .A2(n11936), .ZN(n11945) );
  NOR2_X1 U12984 ( .A1(n14341), .A2(n20676), .ZN(n14440) );
  NAND2_X1 U12985 ( .A1(n14235), .A2(n14234), .ZN(n14258) );
  NAND2_X1 U12986 ( .A1(n11971), .A2(n11970), .ZN(n14312) );
  CLKBUF_X1 U12987 ( .A(n15497), .Z(n15494) );
  NAND2_X1 U12988 ( .A1(n17038), .A2(n19138), .ZN(n13606) );
  NAND2_X2 U12989 ( .A1(n13060), .A2(n13050), .ZN(n13452) );
  AND2_X4 U12990 ( .A1(n11711), .A2(n16830), .ZN(n11863) );
  NOR2_X1 U12991 ( .A1(n12901), .A2(n12904), .ZN(n12991) );
  NAND2_X1 U12992 ( .A1(n15264), .A2(n11698), .ZN(n15497) );
  NAND2_X1 U12993 ( .A1(n16983), .A2(n16973), .ZN(n16975) );
  INV_X1 U12994 ( .A(n15263), .ZN(n15264) );
  INV_X1 U12995 ( .A(n15326), .ZN(n12075) );
  NAND2_X1 U12996 ( .A1(n15108), .A2(n11696), .ZN(n15263) );
  INV_X1 U12997 ( .A(n13624), .ZN(n13080) );
  NAND2_X1 U12998 ( .A1(n17280), .A2(n17025), .ZN(n17026) );
  CLKBUF_X1 U12999 ( .A(n16357), .Z(n16439) );
  BUF_X1 U13000 ( .A(n16313), .Z(n16326) );
  NAND2_X1 U13001 ( .A1(n15815), .A2(n15816), .ZN(n15889) );
  OAI21_X1 U13002 ( .B1(n12446), .B2(n12447), .A(n16290), .ZN(n16478) );
  NAND2_X1 U13003 ( .A1(n14251), .A2(n14250), .ZN(n14252) );
  INV_X1 U13004 ( .A(n13722), .ZN(n13376) );
  INV_X1 U13005 ( .A(n15889), .ZN(n15890) );
  AND2_X1 U13006 ( .A1(n14253), .A2(n14252), .ZN(n17691) );
  NAND2_X1 U13007 ( .A1(n15619), .A2(n15618), .ZN(n15625) );
  AND2_X1 U13008 ( .A1(n17047), .A2(n19138), .ZN(n11683) );
  OR2_X1 U13009 ( .A1(n19119), .A2(n19052), .ZN(n11684) );
  NAND2_X1 U13010 ( .A1(n16097), .A2(n12824), .ZN(n11686) );
  OR2_X1 U13011 ( .A1(n22215), .A2(n22204), .ZN(n11687) );
  OR2_X1 U13012 ( .A1(n16210), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11689) );
  AND2_X1 U13013 ( .A1(n12815), .A2(n13381), .ZN(n11690) );
  INV_X1 U13014 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18415) );
  OR2_X1 U13015 ( .A1(n11692), .A2(n16233), .ZN(n11691) );
  NOR2_X1 U13016 ( .A1(n13733), .A2(n15225), .ZN(n11692) );
  INV_X1 U13017 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18421) );
  INV_X1 U13018 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15288) );
  INV_X1 U13019 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12584) );
  AND2_X1 U13020 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11693) );
  OR4_X1 U13021 ( .A1(n17184), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13736), .A4(n13735), .ZN(n11694) );
  OR3_X1 U13022 ( .A1(n17184), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13735), .ZN(n11695) );
  INV_X1 U13023 ( .A(n13226), .ZN(n13348) );
  OR2_X1 U13024 ( .A1(n13261), .A2(n13260), .ZN(n11696) );
  OR2_X1 U13025 ( .A1(n15888), .A2(n15887), .ZN(n11697) );
  OR2_X1 U13026 ( .A1(n13274), .A2(n13273), .ZN(n11698) );
  AND2_X1 U13027 ( .A1(n13418), .A2(n16097), .ZN(n11699) );
  INV_X1 U13028 ( .A(n15322), .ZN(n14131) );
  INV_X1 U13029 ( .A(n13195), .ZN(n13363) );
  AND2_X2 U13030 ( .A1(n14191), .A2(n16830), .ZN(n11983) );
  AND4_X1 U13031 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11700) );
  INV_X1 U13032 ( .A(n11184), .ZN(n12388) );
  AND4_X1 U13033 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11701) );
  NAND2_X1 U13034 ( .A1(n11945), .A2(n11944), .ZN(n11973) );
  NAND2_X1 U13035 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12834) );
  OR2_X1 U13036 ( .A1(n12036), .A2(n12035), .ZN(n12498) );
  AND2_X1 U13037 ( .A1(n15376), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12562) );
  OR2_X1 U13038 ( .A1(n12012), .A2(n12011), .ZN(n12488) );
  OR2_X1 U13039 ( .A1(n11892), .A2(n12549), .ZN(n11877) );
  AOI22_X1 U13040 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12753), .B1(
        n12756), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U13041 ( .A1(n12856), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12866) );
  AND2_X1 U13042 ( .A1(n16781), .A2(n21975), .ZN(n12532) );
  OR2_X1 U13043 ( .A1(n12059), .A2(n12058), .ZN(n12508) );
  OR2_X1 U13044 ( .A1(n12578), .A2(n12577), .ZN(n13802) );
  NAND2_X1 U13045 ( .A1(n11938), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11854) );
  NAND2_X1 U13046 ( .A1(n11849), .A2(n11848), .ZN(n11851) );
  NAND2_X1 U13047 ( .A1(n13389), .A2(n15211), .ZN(n12825) );
  NAND2_X1 U13048 ( .A1(n12640), .A2(n12639), .ZN(n12638) );
  NAND2_X1 U13049 ( .A1(n11244), .A2(n17191), .ZN(n13583) );
  NAND2_X1 U13050 ( .A1(n13218), .A2(n16097), .ZN(n12912) );
  NAND2_X1 U13051 ( .A1(n15322), .A2(n14215), .ZN(n14161) );
  NAND2_X2 U13052 ( .A1(n21333), .A2(n21772), .ZN(n14338) );
  OR2_X1 U13053 ( .A1(n21399), .A2(n18147), .ZN(n18165) );
  INV_X1 U13054 ( .A(n14565), .ZN(n13838) );
  OR2_X1 U13055 ( .A1(n12423), .A2(n16577), .ZN(n12424) );
  NOR2_X1 U13056 ( .A1(n12229), .A2(n16458), .ZN(n12230) );
  NAND2_X1 U13057 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11993) );
  AND2_X1 U13058 ( .A1(n13828), .A2(n11861), .ZN(n14062) );
  NOR2_X1 U13059 ( .A1(n15284), .A2(n11832), .ZN(n11833) );
  OR2_X1 U13060 ( .A1(n11908), .A2(n11907), .ZN(n12455) );
  INV_X1 U13061 ( .A(n11910), .ZN(n11911) );
  INV_X1 U13062 ( .A(n12831), .ZN(n15203) );
  NAND2_X1 U13063 ( .A1(n14225), .A2(n19733), .ZN(n14219) );
  AND2_X1 U13064 ( .A1(n17628), .A2(n17629), .ZN(n13612) );
  OR2_X1 U13065 ( .A1(n12950), .A2(n12949), .ZN(n13428) );
  OR2_X1 U13066 ( .A1(n13204), .A2(n13203), .ZN(n13208) );
  NOR2_X1 U13067 ( .A1(n12901), .A2(n12902), .ZN(n12990) );
  INV_X1 U13068 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18094) );
  AND2_X1 U13069 ( .A1(n21151), .A2(n18193), .ZN(n18191) );
  INV_X1 U13070 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12123) );
  OAI21_X1 U13071 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11935), .A(
        n11934), .ZN(n11936) );
  OR2_X1 U13072 ( .A1(n14043), .A2(n22153), .ZN(n13685) );
  OR2_X1 U13073 ( .A1(n15286), .A2(n15285), .ZN(n15287) );
  OR2_X1 U13074 ( .A1(n12424), .A2(n16318), .ZN(n13664) );
  AND2_X1 U13075 ( .A1(n12299), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12318) );
  AND2_X1 U13076 ( .A1(n12214), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12199) );
  INV_X1 U13077 ( .A(n12182), .ZN(n12226) );
  AND3_X1 U13078 ( .A1(n11833), .A2(n11919), .A3(n14077), .ZN(n14053) );
  OR2_X1 U13079 ( .A1(n12790), .A2(n12652), .ZN(n12653) );
  INV_X1 U13080 ( .A(n15626), .ZN(n15627) );
  OR2_X1 U13081 ( .A1(n13070), .A2(n13069), .ZN(n13455) );
  NAND2_X1 U13082 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  NOR2_X1 U13083 ( .A1(n18996), .A2(n13507), .ZN(n17053) );
  OR2_X1 U13084 ( .A1(n13591), .A2(n13590), .ZN(n17087) );
  OR2_X1 U13085 ( .A1(n17381), .A2(n17365), .ZN(n13399) );
  NOR2_X1 U13086 ( .A1(n17345), .A2(n13609), .ZN(n17132) );
  INV_X1 U13087 ( .A(n19109), .ZN(n17365) );
  NOR2_X1 U13088 ( .A1(n19140), .A2(n19141), .ZN(n17367) );
  INV_X1 U13089 ( .A(n14137), .ZN(n13213) );
  NAND2_X1 U13090 ( .A1(n12806), .A2(n20177), .ZN(n12818) );
  NOR2_X1 U13091 ( .A1(n12905), .A2(n12898), .ZN(n12981) );
  AND2_X2 U13093 ( .A1(n12637), .A2(n12636), .ZN(n15241) );
  NOR2_X1 U13094 ( .A1(n21263), .A2(n19407), .ZN(n18052) );
  NOR2_X1 U13095 ( .A1(n21138), .A2(n18169), .ZN(n18144) );
  NOR2_X1 U13096 ( .A1(n18492), .A2(n18526), .ZN(n18490) );
  INV_X1 U13097 ( .A(n22096), .ZN(n22125) );
  NOR2_X1 U13098 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  AND2_X1 U13099 ( .A1(n16557), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15300) );
  NAND2_X1 U13100 ( .A1(n11943), .A2(n11942), .ZN(n11944) );
  INV_X1 U13101 ( .A(n16206), .ZN(n16209) );
  XNOR2_X1 U13102 ( .A(n15287), .B(n16285), .ZN(n16557) );
  NAND2_X1 U13103 ( .A1(n12370), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12423) );
  OR2_X1 U13104 ( .A1(n12593), .A2(n13808), .ZN(n12594) );
  AND2_X1 U13105 ( .A1(n21971), .A2(n16616), .ZN(n20511) );
  OR2_X1 U13106 ( .A1(n15529), .A2(n15531), .ZN(n15527) );
  AND2_X1 U13107 ( .A1(n15175), .A2(n15174), .ZN(n22263) );
  NOR2_X1 U13108 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22253) );
  NOR2_X1 U13109 ( .A1(n15697), .A2(n22479), .ZN(n22278) );
  INV_X1 U13110 ( .A(n22292), .ZN(n22266) );
  OR3_X1 U13111 ( .A1(n22280), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14531), 
        .ZN(n22477) );
  INV_X1 U13112 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12293) );
  MUX2_X1 U13113 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12653), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12677) );
  OR2_X1 U13114 ( .A1(n18717), .A2(n15238), .ZN(n19041) );
  NAND2_X1 U13115 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19041), .ZN(n19036) );
  AND3_X1 U13116 ( .A1(n13334), .A2(n13333), .A3(n13332), .ZN(n18827) );
  AND3_X1 U13117 ( .A1(n13225), .A2(n13224), .A3(n13223), .ZN(n15201) );
  INV_X1 U13118 ( .A(n18945), .ZN(n17101) );
  INV_X1 U13119 ( .A(n15272), .ZN(n15491) );
  AOI21_X1 U13120 ( .B1(n16894), .B2(n19103), .A(n11691), .ZN(n13734) );
  AND2_X1 U13121 ( .A1(n17197), .A2(n13400), .ZN(n17189) );
  INV_X1 U13122 ( .A(n13405), .ZN(n13079) );
  AND3_X1 U13123 ( .A1(n13277), .A2(n13276), .A3(n13275), .ZN(n18793) );
  AND2_X1 U13124 ( .A1(n13379), .A2(n13378), .ZN(n14632) );
  NAND2_X1 U13125 ( .A1(n19795), .A2(n20060), .ZN(n19766) );
  INV_X1 U13126 ( .A(n19719), .ZN(n19720) );
  INV_X1 U13127 ( .A(n19788), .ZN(n19838) );
  AOI21_X1 U13128 ( .B1(n17462), .B2(n18047), .A(n17461), .ZN(n21795) );
  OR2_X2 U13129 ( .A1(n20811), .A2(n20812), .ZN(n20823) );
  NAND2_X1 U13130 ( .A1(n20666), .A2(n20670), .ZN(n20674) );
  AOI211_X1 U13131 ( .C1(n18067), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14347), .B(n14346), .ZN(n14348) );
  NOR2_X1 U13132 ( .A1(n18092), .A2(n18091), .ZN(n18188) );
  NAND2_X1 U13133 ( .A1(n18364), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18368) );
  INV_X1 U13134 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20826) );
  NAND2_X1 U13135 ( .A1(n18144), .A2(n18183), .ZN(n21637) );
  INV_X1 U13136 ( .A(n21679), .ZN(n21700) );
  INV_X1 U13137 ( .A(n21753), .ZN(n21707) );
  NAND2_X1 U13138 ( .A1(n20604), .A2(n18050), .ZN(n21601) );
  INV_X1 U13139 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21784) );
  INV_X1 U13140 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20664) );
  AND2_X1 U13141 ( .A1(n15842), .A2(n15289), .ZN(n22137) );
  INV_X1 U13142 ( .A(n22059), .ZN(n22136) );
  INV_X1 U13143 ( .A(n16453), .ZN(n16463) );
  OR2_X2 U13144 ( .A1(n13976), .A2(n13975), .ZN(n14028) );
  OR2_X1 U13145 ( .A1(n12320), .A2(n12319), .ZN(n12369) );
  NAND2_X1 U13146 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n12264), .ZN(
        n12298) );
  AND2_X1 U13147 ( .A1(n15828), .A2(n15827), .ZN(n15833) );
  NAND2_X1 U13148 ( .A1(n12060), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12070) );
  INV_X1 U13149 ( .A(n22141), .ZN(n20518) );
  AND2_X1 U13150 ( .A1(n14066), .A2(n15088), .ZN(n21952) );
  AND2_X1 U13151 ( .A1(n14066), .A2(n14056), .ZN(n22017) );
  OAI22_X1 U13152 ( .A1(n22245), .A2(n22244), .B1(n22274), .B2(n22255), .ZN(
        n22481) );
  INV_X1 U13153 ( .A(n22493), .ZN(n22487) );
  AND2_X1 U13154 ( .A1(n15342), .A2(n15353), .ZN(n22509) );
  INV_X1 U13155 ( .A(n22521), .ZN(n22396) );
  NOR2_X1 U13156 ( .A1(n16820), .A2(n14687), .ZN(n15382) );
  NOR2_X1 U13157 ( .A1(n12463), .A2(n15118), .ZN(n15354) );
  AND2_X1 U13158 ( .A1(n15354), .A2(n15353), .ZN(n22537) );
  NOR2_X1 U13159 ( .A1(n16820), .A2(n14520), .ZN(n15386) );
  AND2_X1 U13160 ( .A1(n16820), .A2(n14687), .ZN(n15352) );
  INV_X1 U13161 ( .A(n22567), .ZN(n22411) );
  NOR2_X1 U13162 ( .A1(n14549), .A2(n22479), .ZN(n22291) );
  INV_X1 U13163 ( .A(n22442), .ZN(n22456) );
  NOR2_X1 U13164 ( .A1(n15388), .A2(n15383), .ZN(n22577) );
  INV_X1 U13165 ( .A(n22235), .ZN(n22587) );
  INV_X1 U13166 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20527) );
  NAND2_X1 U13167 ( .A1(n12677), .A2(n12655), .ZN(n14646) );
  NAND2_X1 U13168 ( .A1(n18911), .A2(n17412), .ZN(n18912) );
  INV_X1 U13169 ( .A(n17412), .ZN(n18778) );
  INV_X1 U13170 ( .A(n19036), .ZN(n19012) );
  AND2_X1 U13171 ( .A1(n18717), .A2(n15231), .ZN(n19014) );
  OR2_X1 U13172 ( .A1(n13299), .A2(n13298), .ZN(n15499) );
  OR2_X1 U13173 ( .A1(n15216), .A2(n19955), .ZN(n19643) );
  INV_X1 U13174 ( .A(n17608), .ZN(n17671) );
  INV_X1 U13175 ( .A(n17633), .ZN(n17670) );
  INV_X1 U13176 ( .A(n14126), .ZN(n19106) );
  BUF_X1 U13177 ( .A(n13624), .Z(n19113) );
  AND2_X1 U13178 ( .A1(n13605), .A2(n13184), .ZN(n19103) );
  INV_X1 U13179 ( .A(n18892), .ZN(n19139) );
  AND2_X1 U13180 ( .A1(n13605), .A2(n14635), .ZN(n19108) );
  NAND2_X1 U13181 ( .A1(n13605), .A2(n13187), .ZN(n19119) );
  INV_X1 U13182 ( .A(n19846), .ZN(n20174) );
  OAI21_X1 U13183 ( .B1(n20280), .B2(n19847), .A(n19846), .ZN(n20286) );
  AND2_X1 U13184 ( .A1(n19825), .A2(n19809), .ZN(n20276) );
  AND2_X1 U13185 ( .A1(n19825), .A2(n19792), .ZN(n20258) );
  AND2_X1 U13186 ( .A1(n19825), .A2(n17424), .ZN(n20259) );
  NOR2_X2 U13187 ( .A1(n19766), .A2(n19718), .ZN(n20251) );
  OAI21_X1 U13188 ( .B1(n20224), .B2(n19736), .A(n19846), .ZN(n20227) );
  NOR2_X1 U13189 ( .A1(n19766), .A2(n19729), .ZN(n20233) );
  INV_X1 U13190 ( .A(n19755), .ZN(n19809) );
  INV_X1 U13191 ( .A(n19750), .ZN(n19792) );
  NOR2_X1 U13192 ( .A1(n19720), .A2(n19729), .ZN(n20208) );
  NOR2_X1 U13193 ( .A1(n19691), .A2(n19718), .ZN(n20200) );
  NOR2_X2 U13194 ( .A1(n19691), .A2(n19755), .ZN(n20193) );
  INV_X1 U13195 ( .A(n20153), .ZN(n20156) );
  INV_X1 U13196 ( .A(n19666), .ZN(n19836) );
  INV_X1 U13197 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22205) );
  INV_X1 U13198 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n17492) );
  NOR2_X1 U13199 ( .A1(n21025), .A2(n21024), .ZN(n21066) );
  NOR2_X1 U13200 ( .A1(n20951), .A2(n20950), .ZN(n20986) );
  INV_X1 U13201 ( .A(n21050), .ZN(n21093) );
  INV_X1 U13202 ( .A(n21090), .ZN(n21056) );
  INV_X1 U13203 ( .A(n21815), .ZN(n21069) );
  NOR2_X1 U13204 ( .A1(n21180), .A2(n21185), .ZN(n21179) );
  INV_X1 U13205 ( .A(n19535), .ZN(n20666) );
  INV_X1 U13206 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20742) );
  AOI21_X1 U13207 ( .B1(n21479), .B2(n21500), .A(n21747), .ZN(n21763) );
  INV_X1 U13208 ( .A(n21807), .ZN(n21832) );
  INV_X1 U13209 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n17477) );
  INV_X1 U13210 ( .A(n18711), .ZN(n18709) );
  OAI21_X1 U13211 ( .B1(n13775), .B2(n13774), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13918) );
  NAND2_X1 U13212 ( .A1(n15302), .A2(n15299), .ZN(n22059) );
  INV_X1 U13213 ( .A(n22137), .ZN(n22114) );
  OR2_X1 U13214 ( .A1(n15833), .A2(n15829), .ZN(n22083) );
  INV_X1 U13215 ( .A(n20356), .ZN(n20384) );
  OR2_X2 U13216 ( .A1(n13976), .A2(n15294), .ZN(n14035) );
  OAI21_X1 U13217 ( .B1(n11584), .B2(n11578), .A(n11190), .ZN(n16637) );
  OAI21_X1 U13218 ( .B1(n15833), .B2(n15832), .A(n11585), .ZN(n16675) );
  INV_X1 U13219 ( .A(n20505), .ZN(n20522) );
  AND2_X1 U13220 ( .A1(n16221), .A2(n16220), .ZN(n22022) );
  INV_X1 U13221 ( .A(n21906), .ZN(n22001) );
  INV_X1 U13222 ( .A(n22017), .ZN(n22014) );
  NAND2_X1 U13223 ( .A1(n14066), .A2(n14052), .ZN(n22004) );
  NAND2_X1 U13224 ( .A1(n15342), .A2(n15386), .ZN(n22491) );
  INV_X1 U13225 ( .A(n22495), .ZN(n15543) );
  NAND2_X1 U13226 ( .A1(n15342), .A2(n15352), .ZN(n22500) );
  INV_X1 U13227 ( .A(n22509), .ZN(n22506) );
  NAND2_X1 U13228 ( .A1(n15354), .A2(n15386), .ZN(n22513) );
  NAND2_X1 U13229 ( .A1(n15354), .A2(n15382), .ZN(n22521) );
  NAND2_X1 U13230 ( .A1(n15354), .A2(n15352), .ZN(n22527) );
  INV_X1 U13231 ( .A(n22537), .ZN(n22534) );
  AND2_X1 U13232 ( .A1(n14564), .A2(n14563), .ZN(n22342) );
  NAND2_X1 U13233 ( .A1(n14688), .A2(n15386), .ZN(n22546) );
  AND2_X1 U13234 ( .A1(n14557), .A2(n14556), .ZN(n22371) );
  INV_X1 U13235 ( .A(n22291), .ZN(n16865) );
  INV_X1 U13236 ( .A(n22469), .ZN(n16892) );
  OR2_X1 U13237 ( .A1(n15388), .A2(n15387), .ZN(n22573) );
  OR2_X1 U13238 ( .A1(n15388), .A2(n14528), .ZN(n22591) );
  INV_X1 U13239 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22153) );
  NOR2_X1 U13240 ( .A1(n14649), .A2(n19171), .ZN(n18717) );
  INV_X1 U13241 ( .A(n19014), .ZN(n19051) );
  AND2_X2 U13242 ( .A1(n14102), .A2(n19160), .ZN(n16952) );
  NAND2_X1 U13243 ( .A1(n20162), .A2(n15212), .ZN(n20164) );
  NAND2_X2 U13244 ( .A1(n15210), .A2(n15209), .ZN(n20162) );
  NOR2_X1 U13245 ( .A1(n20167), .A2(n20112), .ZN(n19910) );
  INV_X1 U13246 ( .A(n19643), .ZN(n20173) );
  INV_X1 U13247 ( .A(n17709), .ZN(n17735) );
  OR2_X1 U13248 ( .A1(n13927), .A2(n13860), .ZN(n13880) );
  NOR3_X1 U13249 ( .A1(n13637), .A2(n13636), .A3(n13635), .ZN(n13638) );
  INV_X1 U13250 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17614) );
  INV_X1 U13251 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18801) );
  AND2_X1 U13252 ( .A1(n13737), .A2(n11694), .ZN(n13754) );
  OR3_X1 U13253 ( .A1(n13487), .A2(n19128), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19115) );
  INV_X1 U13254 ( .A(n19108), .ZN(n19134) );
  AND2_X1 U13255 ( .A1(n14126), .A2(n17319), .ZN(n19109) );
  INV_X1 U13256 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19065) );
  INV_X1 U13257 ( .A(n20282), .ZN(n20279) );
  INV_X1 U13258 ( .A(n20258), .ZN(n20271) );
  AND2_X1 U13259 ( .A1(n19791), .A2(n19790), .ZN(n20264) );
  AOI22_X1 U13260 ( .A1(n17429), .A2(n17433), .B1(n17428), .B2(n17427), .ZN(
        n20256) );
  AND2_X1 U13261 ( .A1(n19774), .A2(n19773), .ZN(n20039) );
  INV_X1 U13262 ( .A(n20138), .ZN(n20243) );
  INV_X1 U13263 ( .A(n20233), .ZN(n20230) );
  INV_X1 U13264 ( .A(n20225), .ZN(n20137) );
  NAND2_X1 U13265 ( .A1(n19719), .A2(n19809), .ZN(n20223) );
  NAND2_X1 U13266 ( .A1(n19719), .A2(n19792), .ZN(n20217) );
  INV_X1 U13267 ( .A(n20208), .ZN(n20204) );
  INV_X1 U13268 ( .A(n20200), .ZN(n20197) );
  INV_X1 U13269 ( .A(n20193), .ZN(n19920) );
  OAI22_X1 U13270 ( .A1(n19685), .A2(n19681), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19680), .ZN(n20190) );
  INV_X1 U13271 ( .A(n19999), .ZN(n20008) );
  NAND2_X1 U13272 ( .A1(n20915), .A2(n20914), .ZN(n20951) );
  NAND2_X1 U13273 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n20810), .ZN(n21090) );
  NOR2_X1 U13274 ( .A1(n20988), .A2(n17953), .ZN(n17958) );
  AND2_X1 U13275 ( .A1(n18039), .A2(n21197), .ZN(n18037) );
  INV_X1 U13276 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17812) );
  NOR2_X1 U13277 ( .A1(n21156), .A2(n21122), .ZN(n21126) );
  NOR2_X1 U13278 ( .A1(n18081), .A2(n18080), .ZN(n21138) );
  NOR2_X1 U13279 ( .A1(n21770), .A2(n18672), .ZN(n18685) );
  INV_X1 U13280 ( .A(n18672), .ZN(n18671) );
  INV_X1 U13281 ( .A(n20617), .ZN(n20659) );
  INV_X1 U13282 ( .A(n18535), .ZN(n18508) );
  INV_X1 U13283 ( .A(n18613), .ZN(n18605) );
  INV_X1 U13284 ( .A(n21757), .ZN(n21747) );
  INV_X1 U13285 ( .A(n21765), .ZN(n21750) );
  INV_X1 U13286 ( .A(n21730), .ZN(n21712) );
  INV_X1 U13287 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21774) );
  INV_X2 U13288 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21333) );
  INV_X1 U13289 ( .A(n19340), .ZN(n19363) );
  INV_X1 U13290 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21830) );
  INV_X1 U13291 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21818) );
  OR2_X1 U13292 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n17477), .ZN(n22225) );
  INV_X1 U13293 ( .A(n18709), .ZN(n18708) );
  INV_X1 U13294 ( .A(n18706), .ZN(n18712) );
  INV_X1 U13295 ( .A(n20352), .ZN(n20341) );
  NAND2_X1 U13296 ( .A1(n11688), .A2(n12606), .ZN(P1_U2971) );
  NAND2_X1 U13297 ( .A1(n11682), .A2(n13638), .ZN(P2_U2994) );
  OAI21_X1 U13298 ( .B1(n11216), .B2(n19134), .A(n13657), .ZN(P2_U3017) );
  NAND2_X1 U13299 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11706) );
  NAND2_X1 U13300 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U13301 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11704) );
  NAND2_X1 U13302 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11703) );
  NAND2_X1 U13303 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11710) );
  NAND2_X1 U13304 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11709) );
  NAND2_X1 U13305 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11708) );
  NAND2_X1 U13306 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11707) );
  NAND2_X1 U13307 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11717) );
  NAND2_X1 U13308 ( .A1(n12053), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11716) );
  BUF_X4 U13309 ( .A(n12237), .Z(n13693) );
  NAND2_X1 U13310 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11715) );
  NAND2_X1 U13311 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11714) );
  AND2_X4 U13312 ( .A1(n11718), .A2(n13935), .ZN(n12338) );
  NAND2_X1 U13313 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U13314 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U13315 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11722) );
  NAND2_X1 U13316 ( .A1(n11983), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U13317 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U13318 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U13319 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11730) );
  NAND2_X1 U13320 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U13321 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11736) );
  NAND2_X1 U13322 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11735) );
  NAND2_X1 U13323 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11734) );
  NAND2_X1 U13324 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11733) );
  NAND2_X1 U13325 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11740) );
  NAND2_X1 U13326 ( .A1(n12053), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U13327 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11738) );
  NAND2_X1 U13328 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11737) );
  NAND2_X1 U13329 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11744) );
  NAND2_X1 U13330 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U13331 ( .A1(n12030), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U13332 ( .A1(n11983), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11741) );
  NAND4_X4 U13333 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11832) );
  NAND2_X1 U13334 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11752) );
  NAND2_X1 U13335 ( .A1(n12078), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11751) );
  NAND2_X1 U13336 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11750) );
  NAND2_X1 U13337 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U13338 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11756) );
  NAND2_X1 U13339 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U13340 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U13341 ( .A1(n12030), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11753) );
  NAND2_X1 U13342 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11760) );
  NAND2_X1 U13343 ( .A1(n12053), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U13344 ( .A1(n11983), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U13345 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11757) );
  NAND2_X1 U13346 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U13347 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U13348 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11762) );
  NAND2_X1 U13349 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11761) );
  AOI22_X1 U13350 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11803), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U13351 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U13352 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U13353 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U13354 ( .A1(n12053), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11181), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U13355 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U13356 ( .A1(n12030), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U13357 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11864), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U13358 ( .A1(n12053), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U13359 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U13360 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U13361 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11778) );
  NAND4_X1 U13362 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11787) );
  AOI22_X1 U13363 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11803), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U13364 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U13365 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11864), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U13366 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11782) );
  NAND4_X1 U13367 ( .A1(n11785), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n11786) );
  AOI22_X1 U13368 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12053), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U13369 ( .A1(n12078), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U13370 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U13371 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11788) );
  NAND4_X1 U13372 ( .A1(n11791), .A2(n11790), .A3(n11789), .A4(n11788), .ZN(
        n11797) );
  AOI22_X1 U13373 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U13374 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U13375 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U13376 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11864), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11792) );
  NAND4_X1 U13377 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11796) );
  AOI22_X1 U13378 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11949), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U13379 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11883), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U13380 ( .A1(n12078), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U13381 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11864), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U13382 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11869), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U13383 ( .A1(n12053), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U13384 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12030), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U13385 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U13386 ( .A1(n11954), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11811) );
  NAND2_X1 U13387 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U13388 ( .A1(n11949), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U13389 ( .A1(n11883), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U13390 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U13391 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U13392 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11813) );
  NAND2_X1 U13393 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11812) );
  AND4_X2 U13394 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11826) );
  NAND2_X1 U13395 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U13396 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U13397 ( .A1(n12030), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U13398 ( .A1(n11864), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U13399 ( .A1(n12053), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11823) );
  NAND2_X1 U13400 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11822) );
  NAND2_X1 U13401 ( .A1(n11870), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U13402 ( .A1(n11983), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11820) );
  NAND4_X4 U13403 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n15294) );
  NAND2_X1 U13404 ( .A1(n17546), .A2(n16206), .ZN(n11830) );
  INV_X1 U13405 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20528) );
  NAND2_X1 U13406 ( .A1(n20528), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22180) );
  INV_X1 U13407 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n22184) );
  NAND2_X1 U13408 ( .A1(n22184), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U13409 ( .A1(n22180), .A2(n11831), .ZN(n13831) );
  INV_X1 U13410 ( .A(n16272), .ZN(n11919) );
  AOI21_X1 U13411 ( .B1(n13809), .B2(n13831), .A(n14053), .ZN(n11834) );
  NAND2_X1 U13412 ( .A1(n14050), .A2(n11834), .ZN(n11835) );
  NAND2_X1 U13413 ( .A1(n11835), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U13414 ( .A1(n14532), .A2(n11836), .ZN(n11837) );
  AOI21_X1 U13415 ( .B1(n13820), .B2(n14043), .A(n14077), .ZN(n11845) );
  NAND2_X1 U13416 ( .A1(n11840), .A2(n11828), .ZN(n11841) );
  NAND2_X1 U13417 ( .A1(n11841), .A2(n14565), .ZN(n11844) );
  NAND2_X1 U13418 ( .A1(n13823), .A2(n15657), .ZN(n11842) );
  INV_X1 U13419 ( .A(n13801), .ZN(n11846) );
  NAND2_X1 U13420 ( .A1(n11938), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11849) );
  NAND2_X1 U13421 ( .A1(n15288), .A2(n22280), .ZN(n20525) );
  XNOR2_X1 U13422 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22240) );
  OR2_X1 U13423 ( .A1(n17549), .A2(n17517), .ZN(n11933) );
  OAI21_X1 U13424 ( .B1(n12602), .B2(n22240), .A(n11933), .ZN(n11847) );
  INV_X1 U13425 ( .A(n11847), .ZN(n11848) );
  INV_X1 U13426 ( .A(n17549), .ZN(n22150) );
  INV_X1 U13427 ( .A(n12602), .ZN(n11976) );
  MUX2_X1 U13428 ( .A(n22150), .B(n11976), .S(n15376), .Z(n11852) );
  INV_X1 U13429 ( .A(n11852), .ZN(n11853) );
  INV_X1 U13430 ( .A(n11855), .ZN(n11859) );
  NAND3_X1 U13431 ( .A1(n13820), .A2(n14043), .A3(n15294), .ZN(n11857) );
  INV_X1 U13432 ( .A(n20525), .ZN(n22146) );
  INV_X1 U13433 ( .A(n12449), .ZN(n14558) );
  OAI21_X1 U13434 ( .B1(n14558), .B2(n14098), .A(n13818), .ZN(n11856) );
  NAND4_X1 U13435 ( .A1(n11857), .A2(n22146), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n11856), .ZN(n11858) );
  NOR2_X1 U13436 ( .A1(n11859), .A2(n11858), .ZN(n11862) );
  NAND2_X1 U13437 ( .A1(n14077), .A2(n11571), .ZN(n11861) );
  AOI22_X1 U13438 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U13439 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U13440 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U13441 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11865) );
  NAND4_X1 U13442 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n11876) );
  AOI22_X1 U13443 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U13444 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11873) );
  INV_X1 U13445 ( .A(n11870), .ZN(n12390) );
  AOI22_X1 U13446 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U13447 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11871) );
  NAND4_X1 U13448 ( .A1(n11874), .A2(n11873), .A3(n11872), .A4(n11871), .ZN(
        n11875) );
  OAI21_X2 U13449 ( .B1(n15410), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11877), 
        .ZN(n12453) );
  AOI22_X1 U13450 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U13451 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11180), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U13452 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11880) );
  BUF_X1 U13453 ( .A(n11983), .Z(n11878) );
  AOI22_X1 U13454 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U13455 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11889) );
  AOI22_X1 U13456 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U13457 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U13458 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U13459 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11884) );
  NAND4_X1 U13460 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n11888) );
  OR2_X1 U13461 ( .A1(n12549), .A2(n12521), .ZN(n11897) );
  NAND2_X1 U13462 ( .A1(n12546), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11891) );
  OAI211_X1 U13463 ( .C1(n11948), .C2(n11892), .A(n11897), .B(n11891), .ZN(
        n11893) );
  INV_X1 U13464 ( .A(n12521), .ZN(n11896) );
  INV_X1 U13465 ( .A(n11897), .ZN(n11909) );
  AOI22_X1 U13466 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12108), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U13467 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U13468 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U13469 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U13470 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11908) );
  AOI22_X1 U13471 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U13472 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U13473 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U13474 ( .A1(n11181), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11903) );
  NAND4_X1 U13475 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11907) );
  MUX2_X1 U13476 ( .A(n12515), .B(n11909), .S(n12455), .Z(n11910) );
  INV_X1 U13477 ( .A(n12455), .ZN(n11914) );
  NAND2_X1 U13478 ( .A1(n12546), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11913) );
  AOI21_X1 U13479 ( .B1(n11838), .B2(n12521), .A(n22153), .ZN(n11912) );
  OAI211_X1 U13480 ( .C1(n11914), .C2(n14245), .A(n11913), .B(n11912), .ZN(
        n11924) );
  INV_X1 U13481 ( .A(n11915), .ZN(n11916) );
  NAND2_X1 U13482 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  NAND2_X1 U13483 ( .A1(n11571), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U13484 ( .A1(n16820), .A2(n12226), .ZN(n11923) );
  AND2_X1 U13485 ( .A1(n11919), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11999) );
  INV_X1 U13486 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11920) );
  INV_X1 U13487 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14168) );
  OAI22_X1 U13488 ( .A1(n12442), .A2(n11920), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14168), .ZN(n11921) );
  AOI21_X1 U13489 ( .B1(n11999), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11921), .ZN(n11922) );
  NAND2_X1 U13490 ( .A1(n14687), .A2(n11571), .ZN(n11926) );
  NAND2_X1 U13491 ( .A1(n11926), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13961) );
  INV_X1 U13492 ( .A(n14523), .ZN(n15432) );
  INV_X1 U13493 ( .A(n11999), .ZN(n12016) );
  NAND2_X1 U13494 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n12293), .ZN(
        n11928) );
  NAND2_X1 U13495 ( .A1(n16281), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11927) );
  OAI211_X1 U13496 ( .C1(n12016), .C2(n11419), .A(n11928), .B(n11927), .ZN(
        n11929) );
  AOI21_X1 U13497 ( .B1(n15432), .B2(n12226), .A(n11929), .ZN(n13962) );
  OR2_X1 U13498 ( .A1(n13961), .A2(n13962), .ZN(n13959) );
  NAND2_X1 U13499 ( .A1(n13962), .A2(n13710), .ZN(n11930) );
  NAND2_X1 U13500 ( .A1(n13959), .A2(n11930), .ZN(n14144) );
  NAND2_X1 U13501 ( .A1(n14145), .A2(n14144), .ZN(n14314) );
  INV_X1 U13502 ( .A(n11933), .ZN(n11935) );
  NAND2_X1 U13503 ( .A1(n11938), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11943) );
  NAND2_X1 U13504 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U13505 ( .A1(n17523), .A2(n11939), .ZN(n11940) );
  NOR2_X1 U13506 ( .A1(n17523), .A2(n17517), .ZN(n15347) );
  NAND2_X1 U13507 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15347), .ZN(
        n11974) );
  NAND2_X1 U13508 ( .A1(n11940), .A2(n11974), .ZN(n15528) );
  OAI22_X1 U13509 ( .A1(n12602), .A2(n15528), .B1(n17549), .B2(n17523), .ZN(
        n11941) );
  INV_X1 U13510 ( .A(n11941), .ZN(n11942) );
  AOI22_X1 U13511 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U13512 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U13513 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U13514 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11950) );
  NAND4_X1 U13515 ( .A1(n11953), .A2(n11952), .A3(n11951), .A4(n11950), .ZN(
        n11960) );
  AOI22_X1 U13516 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13517 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U13518 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U13519 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11955) );
  NAND4_X1 U13520 ( .A1(n11958), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11959) );
  AOI22_X1 U13521 ( .A1(n12582), .A2(n12464), .B1(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12546), .ZN(n11961) );
  NAND2_X1 U13522 ( .A1(n11963), .A2(n11962), .ZN(n11964) );
  NAND2_X1 U13523 ( .A1(n12002), .A2(n11964), .ZN(n12463) );
  INV_X1 U13524 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11966) );
  XNOR2_X1 U13525 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15301) );
  AOI21_X1 U13526 ( .B1(n13710), .B2(n15301), .A(n16280), .ZN(n11965) );
  OAI21_X1 U13527 ( .B1(n12442), .B2(n11966), .A(n11965), .ZN(n11967) );
  AOI21_X1 U13528 ( .B1(n11999), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11967), .ZN(n11968) );
  NAND2_X1 U13529 ( .A1(n16280), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11972) );
  NAND2_X1 U13530 ( .A1(n11969), .A2(n11972), .ZN(n14315) );
  INV_X1 U13531 ( .A(n14315), .ZN(n11970) );
  NAND2_X1 U13532 ( .A1(n11938), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11978) );
  INV_X1 U13533 ( .A(n11974), .ZN(n14524) );
  INV_X1 U13534 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17526) );
  NAND2_X1 U13535 ( .A1(n14524), .A2(n17526), .ZN(n15364) );
  NAND2_X1 U13536 ( .A1(n11974), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11975) );
  NAND2_X1 U13537 ( .A1(n15364), .A2(n11975), .ZN(n16853) );
  AOI22_X1 U13538 ( .A1(n11976), .A2(n16853), .B1(n22150), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11977) );
  XNOR2_X2 U13539 ( .A(n11973), .B(n15165), .ZN(n15419) );
  AOI22_X1 U13540 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U13541 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U13542 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U13543 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11979) );
  NAND4_X1 U13544 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n11989) );
  AOI22_X1 U13545 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U13546 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U13547 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U13548 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11984) );
  NAND4_X1 U13549 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n11988) );
  AOI22_X1 U13550 ( .A1(n12582), .A2(n12480), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12546), .ZN(n11990) );
  NAND2_X1 U13551 ( .A1(n14569), .A2(n12226), .ZN(n12001) );
  INV_X1 U13552 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11997) );
  INV_X1 U13553 ( .A(n11993), .ZN(n11992) );
  INV_X1 U13554 ( .A(n12018), .ZN(n12019) );
  INV_X1 U13555 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U13556 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  NAND2_X1 U13557 ( .A1(n12019), .A2(n11995), .ZN(n15423) );
  AOI22_X1 U13558 ( .A1(n15423), .A2(n13710), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11996) );
  OAI21_X1 U13559 ( .B1(n12442), .B2(n11997), .A(n11996), .ZN(n11998) );
  AOI21_X1 U13560 ( .B1(n11999), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11998), .ZN(n12000) );
  NAND2_X1 U13561 ( .A1(n12001), .A2(n12000), .ZN(n14265) );
  NAND2_X1 U13562 ( .A1(n14266), .A2(n14265), .ZN(n15106) );
  AOI22_X1 U13563 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U13564 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11182), .B1(
        n11180), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U13565 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11184), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U13566 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12307), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12003) );
  NAND4_X1 U13567 ( .A1(n12006), .A2(n12005), .A3(n12004), .A4(n12003), .ZN(
        n12012) );
  AOI22_X1 U13568 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11769), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U13569 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U13570 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U13571 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12007) );
  NAND4_X1 U13572 ( .A1(n12010), .A2(n12009), .A3(n12008), .A4(n12007), .ZN(
        n12011) );
  NAND2_X1 U13573 ( .A1(n12582), .A2(n12488), .ZN(n12014) );
  NAND2_X1 U13574 ( .A1(n12546), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12013) );
  NAND2_X1 U13575 ( .A1(n12014), .A2(n12013), .ZN(n12025) );
  XNOR2_X1 U13576 ( .A(n12024), .B(n12025), .ZN(n12479) );
  AOI22_X1 U13577 ( .A1(n16281), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12293), .ZN(n12015) );
  OAI21_X1 U13578 ( .B1(n12016), .B2(n12584), .A(n12015), .ZN(n12017) );
  NAND2_X1 U13579 ( .A1(n12017), .A2(n13688), .ZN(n12022) );
  INV_X1 U13580 ( .A(n12042), .ZN(n12044) );
  INV_X1 U13581 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15582) );
  NAND2_X1 U13582 ( .A1(n12019), .A2(n15582), .ZN(n12020) );
  NAND2_X1 U13583 ( .A1(n12044), .A2(n12020), .ZN(n20474) );
  NAND2_X1 U13584 ( .A1(n20474), .A2(n13710), .ZN(n12021) );
  NAND2_X1 U13585 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  INV_X1 U13586 ( .A(n12040), .ZN(n12038) );
  AOI22_X1 U13587 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U13588 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U13589 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U13590 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U13591 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12036) );
  AOI22_X1 U13592 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U13593 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U13594 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U13595 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12031) );
  NAND4_X1 U13596 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n12035) );
  AOI22_X1 U13597 ( .A1(n12582), .A2(n12498), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n12546), .ZN(n12039) );
  NAND2_X1 U13598 ( .A1(n12040), .A2(n12039), .ZN(n12041) );
  NAND2_X1 U13599 ( .A1(n12065), .A2(n12041), .ZN(n12487) );
  INV_X1 U13600 ( .A(n12060), .ZN(n12046) );
  INV_X1 U13601 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U13602 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  NAND2_X1 U13603 ( .A1(n12046), .A2(n12045), .ZN(n22034) );
  AOI22_X1 U13604 ( .A1(n22034), .A2(n13710), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U13605 ( .A1(n16281), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n12047) );
  OAI211_X1 U13606 ( .C1(n12487), .C2(n12182), .A(n12048), .B(n12047), .ZN(
        n14670) );
  NAND2_X1 U13607 ( .A1(n14671), .A2(n14670), .ZN(n14669) );
  INV_X1 U13608 ( .A(n14669), .ZN(n12064) );
  AOI22_X1 U13609 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U13610 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U13611 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U13612 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12049) );
  NAND4_X1 U13613 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n12059) );
  AOI22_X1 U13614 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U13615 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U13616 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U13617 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12054) );
  NAND4_X1 U13618 ( .A1(n12057), .A2(n12056), .A3(n12055), .A4(n12054), .ZN(
        n12058) );
  AOI22_X1 U13619 ( .A1(n12582), .A2(n12508), .B1(n12546), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12066) );
  NAND2_X1 U13620 ( .A1(n12065), .A2(n12066), .ZN(n12496) );
  INV_X1 U13621 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n15270) );
  OAI21_X1 U13622 ( .B1(n12060), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n12070), .ZN(n22045) );
  AOI22_X1 U13623 ( .A1(n22045), .A2(n13710), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12061) );
  OAI21_X1 U13624 ( .B1(n12442), .B2(n15270), .A(n12061), .ZN(n12062) );
  INV_X1 U13625 ( .A(n15220), .ZN(n12063) );
  NAND2_X1 U13626 ( .A1(n12064), .A2(n12063), .ZN(n15327) );
  INV_X1 U13627 ( .A(n15327), .ZN(n12076) );
  NAND2_X1 U13628 ( .A1(n12582), .A2(n12521), .ZN(n12068) );
  NAND2_X1 U13629 ( .A1(n12546), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12067) );
  NAND2_X1 U13630 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  INV_X1 U13631 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12073) );
  OAI21_X1 U13632 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12071), .A(
        n12094), .ZN(n22056) );
  AOI22_X1 U13633 ( .A1(n13710), .A2(n22056), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12072) );
  OAI21_X1 U13634 ( .B1(n12442), .B2(n12073), .A(n12072), .ZN(n12074) );
  AOI21_X1 U13635 ( .B1(n12505), .B2(n12226), .A(n12074), .ZN(n15326) );
  NAND2_X1 U13636 ( .A1(n12076), .A2(n12075), .ZN(n15325) );
  NAND2_X1 U13637 ( .A1(n16281), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12092) );
  INV_X1 U13638 ( .A(n12094), .ZN(n12077) );
  XNOR2_X1 U13639 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12077), .ZN(
        n15611) );
  AOI22_X1 U13640 ( .A1(n13710), .A2(n15611), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U13641 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11182), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U13642 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11863), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U13643 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U13644 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12079) );
  NAND4_X1 U13645 ( .A1(n12082), .A2(n12081), .A3(n12080), .A4(n12079), .ZN(
        n12088) );
  AOI22_X1 U13646 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U13647 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U13648 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U13649 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12083) );
  NAND4_X1 U13650 ( .A1(n12086), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n12087) );
  NOR2_X1 U13651 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  OR2_X1 U13652 ( .A1(n12182), .A2(n12089), .ZN(n12090) );
  XOR2_X1 U13653 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12119), .Z(n15777) );
  AOI22_X1 U13654 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U13655 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11863), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U13656 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U13657 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U13658 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12104) );
  AOI22_X1 U13659 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U13660 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U13661 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13662 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U13663 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  OR2_X1 U13664 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  AOI22_X1 U13665 ( .A1(n12226), .A2(n12105), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U13666 ( .A1(n16281), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12106) );
  OAI211_X1 U13667 ( .C1(n15777), .C2(n13688), .A(n12107), .B(n12106), .ZN(
        n15595) );
  AND2_X2 U13668 ( .A1(n15442), .A2(n15595), .ZN(n15593) );
  AOI22_X1 U13669 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U13670 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U13671 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U13672 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12109) );
  NAND4_X1 U13673 ( .A1(n12112), .A2(n12111), .A3(n12110), .A4(n12109), .ZN(
        n12118) );
  AOI22_X1 U13674 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U13675 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U13676 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U13677 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U13678 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12117) );
  NOR2_X1 U13679 ( .A1(n12118), .A2(n12117), .ZN(n12122) );
  XNOR2_X1 U13680 ( .A(n12124), .B(n12123), .ZN(n16678) );
  NAND2_X1 U13681 ( .A1(n16678), .A2(n13710), .ZN(n12121) );
  AOI22_X1 U13682 ( .A1(n16281), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n16280), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12120) );
  OAI211_X1 U13683 ( .C1(n12122), .C2(n12182), .A(n12121), .B(n12120), .ZN(
        n15656) );
  OR2_X1 U13684 ( .A1(n12125), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12126) );
  NAND2_X1 U13685 ( .A1(n12126), .A2(n12164), .ZN(n22069) );
  NAND2_X1 U13686 ( .A1(n22069), .A2(n13710), .ZN(n12128) );
  AOI22_X1 U13687 ( .A1(n16281), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n16280), 
        .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U13688 ( .A1(n12128), .A2(n12127), .ZN(n15762) );
  AOI22_X1 U13689 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U13690 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U13691 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U13692 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12129) );
  NAND4_X1 U13693 ( .A1(n12132), .A2(n12131), .A3(n12130), .A4(n12129), .ZN(
        n12138) );
  AOI22_X1 U13694 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11180), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U13695 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U13696 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U13697 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12133) );
  NAND4_X1 U13698 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(
        n12137) );
  NOR2_X1 U13699 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  NOR2_X1 U13700 ( .A1(n12182), .A2(n12139), .ZN(n15824) );
  XOR2_X1 U13701 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12179), .Z(
        n16672) );
  AOI22_X1 U13702 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11863), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U13703 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U13704 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U13705 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12141) );
  NAND4_X1 U13706 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .ZN(
        n12150) );
  AOI22_X1 U13707 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11182), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U13708 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U13709 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U13710 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12145) );
  NAND4_X1 U13711 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12149) );
  OR2_X1 U13712 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  AOI22_X1 U13713 ( .A1(n12226), .A2(n12151), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12153) );
  NAND2_X1 U13714 ( .A1(n16281), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12152) );
  OAI211_X1 U13715 ( .C1(n16672), .C2(n13688), .A(n12153), .B(n12152), .ZN(
        n15832) );
  AOI22_X1 U13716 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U13717 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11182), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U13718 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U13719 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12154) );
  NAND4_X1 U13720 ( .A1(n12157), .A2(n12156), .A3(n12155), .A4(n12154), .ZN(
        n12163) );
  AOI22_X1 U13721 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11184), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U13722 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12394), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U13723 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U13724 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12158) );
  NAND4_X1 U13725 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12162) );
  NOR2_X1 U13726 ( .A1(n12163), .A2(n12162), .ZN(n12168) );
  NAND2_X1 U13727 ( .A1(n16281), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12167) );
  XNOR2_X1 U13728 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12164), .ZN(
        n22080) );
  INV_X1 U13729 ( .A(n22080), .ZN(n12165) );
  AOI22_X1 U13730 ( .A1(n16280), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13710), .B2(n12165), .ZN(n12166) );
  OAI211_X1 U13731 ( .C1(n12182), .C2(n12168), .A(n12167), .B(n12166), .ZN(
        n15827) );
  AOI22_X1 U13732 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U13733 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U13734 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U13735 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12169) );
  NAND4_X1 U13736 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12178) );
  AOI22_X1 U13737 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U13738 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U13739 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U13740 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12173) );
  NAND4_X1 U13741 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12177) );
  NOR2_X1 U13742 ( .A1(n12178), .A2(n12177), .ZN(n12183) );
  XNOR2_X1 U13743 ( .A(n12184), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16657) );
  NAND2_X1 U13744 ( .A1(n16657), .A2(n13710), .ZN(n12181) );
  AOI22_X1 U13745 ( .A1(n16281), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n16280), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12180) );
  OAI211_X1 U13746 ( .C1(n12183), .C2(n12182), .A(n12181), .B(n12180), .ZN(
        n15851) );
  XNOR2_X1 U13747 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12232), .ZN(
        n20504) );
  INV_X1 U13748 ( .A(n20504), .ZN(n12198) );
  AOI22_X1 U13749 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U13750 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U13751 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U13752 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12185) );
  NAND4_X1 U13753 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n12194) );
  AOI22_X1 U13754 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U13755 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U13756 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U13757 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12189) );
  NAND4_X1 U13758 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12189), .ZN(
        n12193) );
  NOR2_X1 U13759 ( .A1(n12194), .A2(n12193), .ZN(n12196) );
  AOI22_X1 U13760 ( .A1(n16281), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n16280), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12195) );
  OAI21_X1 U13761 ( .B1(n13685), .B2(n12196), .A(n12195), .ZN(n12197) );
  AOI21_X1 U13762 ( .B1(n12198), .B2(n13710), .A(n12197), .ZN(n16391) );
  XNOR2_X1 U13763 ( .A(n12199), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16646) );
  AOI22_X1 U13764 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11184), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U13765 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U13766 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U13767 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U13768 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12209) );
  AOI22_X1 U13769 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U13770 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U13771 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U13772 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U13773 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12208) );
  NOR2_X1 U13774 ( .A1(n12209), .A2(n12208), .ZN(n12211) );
  AOI22_X1 U13775 ( .A1(n16281), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12293), .ZN(n12210) );
  OAI21_X1 U13776 ( .B1(n13685), .B2(n12211), .A(n12210), .ZN(n12212) );
  AND2_X1 U13777 ( .A1(n12212), .A2(n13688), .ZN(n12213) );
  AOI21_X1 U13778 ( .B1(n16646), .B2(n13710), .A(n12213), .ZN(n16405) );
  OR2_X1 U13779 ( .A1(n16391), .A2(n16405), .ZN(n12229) );
  XOR2_X1 U13780 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12214), .Z(
        n22089) );
  AOI22_X1 U13781 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U13782 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U13783 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U13784 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U13785 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12224) );
  AOI22_X1 U13786 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U13787 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U13788 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U13789 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U13790 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12223) );
  OR2_X1 U13791 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  AOI22_X1 U13792 ( .A1(n12226), .A2(n12225), .B1(n16280), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U13793 ( .A1(n16281), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12227) );
  OAI211_X1 U13794 ( .C1(n22089), .C2(n13688), .A(n12228), .B(n12227), .ZN(
        n16454) );
  NAND2_X1 U13795 ( .A1(n15850), .A2(n12230), .ZN(n16382) );
  INV_X1 U13796 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12231) );
  INV_X1 U13797 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16630) );
  XNOR2_X1 U13798 ( .A(n12263), .B(n16630), .ZN(n16632) );
  NAND2_X1 U13799 ( .A1(n16632), .A2(n13710), .ZN(n12248) );
  AOI22_X1 U13800 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U13801 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U13802 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U13803 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12233) );
  NAND4_X1 U13804 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12243) );
  AOI22_X1 U13805 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U13806 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U13807 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U13808 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U13809 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12242) );
  NOR2_X1 U13810 ( .A1(n12243), .A2(n12242), .ZN(n12246) );
  AOI21_X1 U13811 ( .B1(n16630), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12244) );
  AOI21_X1 U13812 ( .B1(n16281), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12244), .ZN(
        n12245) );
  OAI21_X1 U13813 ( .B1(n13685), .B2(n12246), .A(n12245), .ZN(n12247) );
  NAND2_X1 U13814 ( .A1(n12248), .A2(n12247), .ZN(n16381) );
  AOI22_X1 U13815 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11182), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U13816 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U13817 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U13818 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12249) );
  NAND4_X1 U13819 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(
        n12258) );
  AOI22_X1 U13820 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U13821 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U13822 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U13823 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12253) );
  NAND4_X1 U13824 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(
        n12257) );
  NOR2_X1 U13825 ( .A1(n12258), .A2(n12257), .ZN(n12262) );
  NAND2_X1 U13826 ( .A1(n12293), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12259) );
  NAND2_X1 U13827 ( .A1(n13688), .A2(n12259), .ZN(n12260) );
  AOI21_X1 U13828 ( .B1(n16281), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12260), .ZN(
        n12261) );
  OAI21_X1 U13829 ( .B1(n13685), .B2(n12262), .A(n12261), .ZN(n12266) );
  OAI21_X1 U13830 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12264), .A(
        n12298), .ZN(n22097) );
  OR2_X1 U13831 ( .A1(n22097), .A2(n13688), .ZN(n12265) );
  AOI22_X1 U13832 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U13833 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11184), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U13834 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U13835 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11863), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U13836 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12276) );
  AOI22_X1 U13837 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U13838 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U13839 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U13840 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U13841 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12275) );
  NOR2_X1 U13842 ( .A1(n12276), .A2(n12275), .ZN(n12279) );
  INV_X1 U13843 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16624) );
  AOI21_X1 U13844 ( .B1(n16624), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12277) );
  AOI21_X1 U13845 ( .B1(n16281), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12277), .ZN(
        n12278) );
  OAI21_X1 U13846 ( .B1(n13685), .B2(n12279), .A(n12278), .ZN(n12281) );
  XNOR2_X1 U13847 ( .A(n12298), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16628) );
  NAND2_X1 U13848 ( .A1(n16628), .A2(n13710), .ZN(n12280) );
  AOI22_X1 U13849 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U13850 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U13851 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U13852 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12283) );
  NAND4_X1 U13853 ( .A1(n12286), .A2(n12285), .A3(n12284), .A4(n12283), .ZN(
        n12292) );
  AOI22_X1 U13854 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11863), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U13855 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U13856 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U13857 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12287) );
  NAND4_X1 U13858 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12291) );
  NOR2_X1 U13859 ( .A1(n12292), .A2(n12291), .ZN(n12297) );
  NAND2_X1 U13860 ( .A1(n12293), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12294) );
  NAND2_X1 U13861 ( .A1(n13688), .A2(n12294), .ZN(n12295) );
  AOI21_X1 U13862 ( .B1(n16281), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12295), .ZN(
        n12296) );
  OAI21_X1 U13863 ( .B1(n13685), .B2(n12297), .A(n12296), .ZN(n12302) );
  NOR2_X1 U13864 ( .A1(n12299), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12300) );
  OR2_X1 U13865 ( .A1(n12318), .A2(n12300), .ZN(n16613) );
  NAND2_X1 U13866 ( .A1(n22109), .A2(n13710), .ZN(n12301) );
  NAND2_X1 U13867 ( .A1(n12302), .A2(n12301), .ZN(n16437) );
  AOI22_X1 U13868 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U13869 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U13870 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U13871 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U13872 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12313) );
  AOI22_X1 U13873 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U13874 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U13875 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U13876 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12308) );
  NAND4_X1 U13877 ( .A1(n12311), .A2(n12310), .A3(n12309), .A4(n12308), .ZN(
        n12312) );
  OAI21_X1 U13878 ( .B1(n12313), .B2(n12312), .A(n13707), .ZN(n12317) );
  INV_X1 U13879 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12314) );
  AOI21_X1 U13880 ( .B1(n12314), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12315) );
  AOI21_X1 U13881 ( .B1(n16281), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12315), .ZN(
        n12316) );
  XOR2_X1 U13882 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12318), .Z(
        n16360) );
  AOI22_X1 U13883 ( .A1(n12317), .A2(n12316), .B1(n13710), .B2(n16360), .ZN(
        n16359) );
  NAND2_X1 U13884 ( .A1(n16357), .A2(n16359), .ZN(n16358) );
  INV_X1 U13885 ( .A(n12320), .ZN(n12321) );
  INV_X1 U13886 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12319) );
  OAI21_X1 U13887 ( .B1(n12321), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n12369), .ZN(n22129) );
  AOI22_X1 U13888 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U13889 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U13890 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U13891 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12322) );
  NAND4_X1 U13892 ( .A1(n12325), .A2(n12324), .A3(n12323), .A4(n12322), .ZN(
        n12332) );
  AOI22_X1 U13893 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U13894 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U13895 ( .A1(n12326), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U13896 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12327) );
  NAND4_X1 U13897 ( .A1(n12330), .A2(n12329), .A3(n12328), .A4(n12327), .ZN(
        n12331) );
  NOR2_X1 U13898 ( .A1(n12332), .A2(n12331), .ZN(n12363) );
  AOI22_X1 U13899 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11182), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U13900 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U13901 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U13902 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12334) );
  NAND4_X1 U13903 ( .A1(n12337), .A2(n12336), .A3(n12335), .A4(n12334), .ZN(
        n12344) );
  AOI22_X1 U13904 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12338), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U13905 ( .A1(n11180), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U13906 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U13907 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12339) );
  NAND4_X1 U13908 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12343) );
  NOR2_X1 U13909 ( .A1(n12344), .A2(n12343), .ZN(n12364) );
  XNOR2_X1 U13910 ( .A(n12363), .B(n12364), .ZN(n12347) );
  AOI21_X1 U13911 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n12293), .A(
        n13710), .ZN(n12346) );
  NAND2_X1 U13912 ( .A1(n16281), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n12345) );
  OAI211_X1 U13913 ( .C1(n12347), .C2(n13685), .A(n12346), .B(n12345), .ZN(
        n12348) );
  OAI21_X1 U13914 ( .B1(n13688), .B2(n22129), .A(n12348), .ZN(n16430) );
  INV_X1 U13915 ( .A(n12369), .ZN(n12349) );
  XOR2_X1 U13916 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12349), .Z(
        n16601) );
  INV_X1 U13917 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12350) );
  NOR2_X1 U13918 ( .A1(n12388), .A2(n12350), .ZN(n12354) );
  INV_X1 U13919 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12352) );
  INV_X1 U13920 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12351) );
  OAI22_X1 U13921 ( .A1(n11171), .A2(n12352), .B1(n12390), .B2(n12351), .ZN(
        n12353) );
  AOI211_X1 U13922 ( .C1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .C2(n13691), .A(
        n12354), .B(n12353), .ZN(n12362) );
  AOI22_X1 U13923 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U13924 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U13925 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U13926 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12355) );
  AND4_X1 U13927 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12361) );
  AOI22_X1 U13928 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U13929 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12359) );
  NAND4_X1 U13930 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12371) );
  NOR2_X1 U13931 ( .A1(n12364), .A2(n12363), .ZN(n12372) );
  XOR2_X1 U13932 ( .A(n12371), .B(n12372), .Z(n12367) );
  INV_X1 U13933 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n16499) );
  INV_X1 U13934 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22256) );
  NOR2_X1 U13935 ( .A1(n22256), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12365) );
  OAI22_X1 U13936 ( .A1(n12442), .A2(n16499), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12365), .ZN(n12366) );
  AOI21_X1 U13937 ( .B1(n12367), .B2(n13707), .A(n12366), .ZN(n12368) );
  AOI21_X1 U13938 ( .B1(n13710), .B2(n16601), .A(n12368), .ZN(n16347) );
  INV_X1 U13939 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16597) );
  OAI21_X1 U13940 ( .B1(n12370), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n12423), .ZN(n16589) );
  NAND2_X1 U13941 ( .A1(n12372), .A2(n12371), .ZN(n12403) );
  AOI22_X1 U13942 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U13943 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U13944 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U13945 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U13946 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12382) );
  AOI22_X1 U13947 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U13948 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U13949 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U13950 ( .A1(n11878), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12377) );
  NAND4_X1 U13951 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12381) );
  NOR2_X1 U13952 ( .A1(n12382), .A2(n12381), .ZN(n12404) );
  XNOR2_X1 U13953 ( .A(n12403), .B(n12404), .ZN(n12385) );
  AOI21_X1 U13954 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12293), .A(
        n13710), .ZN(n12384) );
  NAND2_X1 U13955 ( .A1(n16281), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n12383) );
  OAI211_X1 U13956 ( .C1(n12385), .C2(n13685), .A(n12384), .B(n12383), .ZN(
        n12386) );
  OAI21_X1 U13957 ( .B1(n13688), .B2(n16589), .A(n12386), .ZN(n16336) );
  XNOR2_X1 U13958 ( .A(n12423), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16581) );
  INV_X1 U13959 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12387) );
  NOR2_X1 U13960 ( .A1(n12388), .A2(n12387), .ZN(n12393) );
  INV_X1 U13961 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12391) );
  INV_X1 U13962 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12389) );
  OAI22_X1 U13963 ( .A1(n11171), .A2(n12391), .B1(n12390), .B2(n12389), .ZN(
        n12392) );
  AOI211_X1 U13964 ( .C1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .C2(n13691), .A(
        n12393), .B(n12392), .ZN(n12402) );
  AOI22_X1 U13965 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U13966 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12326), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U13967 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U13968 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12395) );
  AND4_X1 U13969 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12401) );
  AOI22_X1 U13970 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U13971 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12399) );
  NAND4_X1 U13972 ( .A1(n12402), .A2(n12401), .A3(n12400), .A4(n12399), .ZN(
        n12419) );
  NOR2_X1 U13973 ( .A1(n12404), .A2(n12403), .ZN(n12420) );
  XOR2_X1 U13974 ( .A(n12419), .B(n12420), .Z(n12407) );
  INV_X1 U13975 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n16486) );
  NOR2_X1 U13976 ( .A1(n22256), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12405) );
  OAI22_X1 U13977 ( .A1(n12442), .A2(n16486), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12405), .ZN(n12406) );
  AOI21_X1 U13978 ( .B1(n12407), .B2(n13707), .A(n12406), .ZN(n12408) );
  AOI21_X1 U13979 ( .B1(n13710), .B2(n16581), .A(n12408), .ZN(n16327) );
  AOI22_X1 U13980 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12237), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U13981 ( .A1(n11183), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U13982 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11863), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U13983 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12409) );
  NAND4_X1 U13984 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(
        n12418) );
  AOI22_X1 U13985 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U13986 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11184), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U13987 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U13988 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12413) );
  NAND4_X1 U13989 ( .A1(n12416), .A2(n12415), .A3(n12414), .A4(n12413), .ZN(
        n12417) );
  NOR2_X1 U13990 ( .A1(n12418), .A2(n12417), .ZN(n12440) );
  NAND2_X1 U13991 ( .A1(n12420), .A2(n12419), .ZN(n12439) );
  XNOR2_X1 U13992 ( .A(n12440), .B(n12439), .ZN(n12421) );
  NOR2_X1 U13993 ( .A1(n12421), .A2(n13685), .ZN(n12427) );
  INV_X1 U13994 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n16479) );
  NOR2_X1 U13995 ( .A1(n22256), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12422) );
  OAI22_X1 U13996 ( .A1(n12442), .A2(n16479), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12422), .ZN(n12426) );
  INV_X1 U13997 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16577) );
  INV_X1 U13998 ( .A(n12424), .ZN(n12425) );
  INV_X1 U13999 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16318) );
  OAI21_X1 U14000 ( .B1(n12425), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n13664), .ZN(n16572) );
  OAI22_X1 U14001 ( .A1(n12427), .A2(n12426), .B1(n13688), .B2(n16572), .ZN(
        n16314) );
  INV_X1 U14002 ( .A(n13664), .ZN(n12428) );
  XOR2_X1 U14003 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n12428), .Z(
        n16306) );
  AOI22_X1 U14004 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U14005 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U14006 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U14007 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12429) );
  NAND4_X1 U14008 ( .A1(n12432), .A2(n12431), .A3(n12430), .A4(n12429), .ZN(
        n12438) );
  AOI22_X1 U14009 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U14010 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U14011 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U14012 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12433) );
  NAND4_X1 U14013 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12433), .ZN(
        n12437) );
  OR2_X1 U14014 ( .A1(n12438), .A2(n12437), .ZN(n13671) );
  NOR2_X1 U14015 ( .A1(n12440), .A2(n12439), .ZN(n13672) );
  XOR2_X1 U14016 ( .A(n13671), .B(n13672), .Z(n12444) );
  INV_X1 U14017 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n16472) );
  NOR2_X1 U14018 ( .A1(n22256), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12441) );
  OAI22_X1 U14019 ( .A1(n12442), .A2(n16472), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12441), .ZN(n12443) );
  AOI21_X1 U14020 ( .B1(n12444), .B2(n13707), .A(n12443), .ZN(n12445) );
  AOI21_X1 U14021 ( .B1(n13710), .B2(n16306), .A(n12445), .ZN(n12447) );
  NAND3_X1 U14022 ( .A1(n22153), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17553) );
  INV_X1 U14023 ( .A(n17553), .ZN(n12448) );
  NAND2_X1 U14024 ( .A1(n14520), .A2(n12557), .ZN(n12452) );
  AND2_X1 U14025 ( .A1(n11828), .A2(n14245), .ZN(n17545) );
  INV_X1 U14026 ( .A(n17545), .ZN(n21844) );
  NAND2_X1 U14027 ( .A1(n11829), .A2(n12449), .ZN(n12465) );
  OAI21_X1 U14028 ( .B1(n21844), .B2(n12455), .A(n12465), .ZN(n12450) );
  INV_X1 U14029 ( .A(n12450), .ZN(n12451) );
  NAND2_X1 U14030 ( .A1(n12452), .A2(n12451), .ZN(n13958) );
  OR2_X1 U14031 ( .A1(n12453), .A2(n11828), .ZN(n12459) );
  NAND2_X1 U14032 ( .A1(n12455), .A2(n12454), .ZN(n12472) );
  OAI21_X1 U14033 ( .B1(n12455), .B2(n12454), .A(n12472), .ZN(n12456) );
  OAI211_X1 U14034 ( .C1(n12456), .C2(n21844), .A(n11570), .B(n11832), .ZN(
        n12457) );
  INV_X1 U14035 ( .A(n12457), .ZN(n12458) );
  NAND2_X1 U14036 ( .A1(n12459), .A2(n12458), .ZN(n12460) );
  INV_X1 U14037 ( .A(n12460), .ZN(n12461) );
  OR2_X1 U14038 ( .A1(n13957), .A2(n12461), .ZN(n12462) );
  INV_X1 U14039 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21893) );
  XNOR2_X1 U14040 ( .A(n12469), .B(n21893), .ZN(n14311) );
  INV_X1 U14041 ( .A(n12557), .ZN(n12516) );
  INV_X1 U14042 ( .A(n12464), .ZN(n12471) );
  XNOR2_X1 U14043 ( .A(n12472), .B(n12471), .ZN(n12467) );
  INV_X1 U14044 ( .A(n12465), .ZN(n12466) );
  AOI21_X1 U14045 ( .B1(n12467), .B2(n17545), .A(n12466), .ZN(n12468) );
  OAI21_X1 U14046 ( .B1(n12463), .B2(n12516), .A(n12468), .ZN(n14310) );
  NAND2_X1 U14047 ( .A1(n12469), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12470) );
  NAND2_X1 U14048 ( .A1(n14569), .A2(n12557), .ZN(n12476) );
  NAND2_X1 U14049 ( .A1(n12472), .A2(n12471), .ZN(n12481) );
  INV_X1 U14050 ( .A(n12480), .ZN(n12473) );
  XNOR2_X1 U14051 ( .A(n12481), .B(n12473), .ZN(n12474) );
  NAND2_X1 U14052 ( .A1(n12474), .A2(n17545), .ZN(n12475) );
  INV_X1 U14053 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21909) );
  NAND2_X1 U14054 ( .A1(n12477), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12478) );
  NAND2_X1 U14055 ( .A1(n12479), .A2(n12557), .ZN(n12484) );
  NAND2_X1 U14056 ( .A1(n12481), .A2(n12480), .ZN(n12490) );
  XNOR2_X1 U14057 ( .A(n12490), .B(n12488), .ZN(n12482) );
  NAND2_X1 U14058 ( .A1(n12482), .A2(n17545), .ZN(n12483) );
  NAND2_X1 U14059 ( .A1(n12484), .A2(n12483), .ZN(n12485) );
  INV_X1 U14060 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21896) );
  XNOR2_X1 U14061 ( .A(n12485), .B(n21896), .ZN(n20468) );
  NAND2_X1 U14062 ( .A1(n20469), .A2(n20468), .ZN(n20467) );
  NAND2_X1 U14063 ( .A1(n12485), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12486) );
  NAND2_X1 U14064 ( .A1(n20467), .A2(n12486), .ZN(n20477) );
  INV_X1 U14065 ( .A(n12488), .ZN(n12489) );
  OR2_X1 U14066 ( .A1(n12490), .A2(n12489), .ZN(n12497) );
  XNOR2_X1 U14067 ( .A(n12497), .B(n12498), .ZN(n12491) );
  NAND2_X1 U14068 ( .A1(n12491), .A2(n17545), .ZN(n12492) );
  NAND2_X1 U14069 ( .A1(n12493), .A2(n12492), .ZN(n12494) );
  INV_X1 U14070 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21911) );
  XNOR2_X1 U14071 ( .A(n12494), .B(n21911), .ZN(n20476) );
  NAND2_X1 U14072 ( .A1(n20477), .A2(n20476), .ZN(n20475) );
  NAND2_X1 U14073 ( .A1(n12494), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12495) );
  NAND3_X1 U14074 ( .A1(n12519), .A2(n12557), .A3(n12496), .ZN(n12502) );
  INV_X1 U14075 ( .A(n12497), .ZN(n12499) );
  NAND2_X1 U14076 ( .A1(n12499), .A2(n12498), .ZN(n12507) );
  XNOR2_X1 U14077 ( .A(n12507), .B(n12508), .ZN(n12500) );
  NAND2_X1 U14078 ( .A1(n12500), .A2(n17545), .ZN(n12501) );
  NAND2_X1 U14079 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  INV_X1 U14080 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21922) );
  XNOR2_X1 U14081 ( .A(n12503), .B(n21922), .ZN(n20482) );
  NAND2_X1 U14082 ( .A1(n12503), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12504) );
  INV_X1 U14083 ( .A(n12505), .ZN(n12506) );
  INV_X1 U14084 ( .A(n12507), .ZN(n12509) );
  NAND2_X1 U14085 ( .A1(n12509), .A2(n12508), .ZN(n12523) );
  XNOR2_X1 U14086 ( .A(n12523), .B(n12521), .ZN(n12510) );
  NAND2_X1 U14087 ( .A1(n12510), .A2(n17545), .ZN(n12511) );
  NAND2_X1 U14088 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  INV_X1 U14089 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21939) );
  XNOR2_X1 U14090 ( .A(n12513), .B(n21939), .ZN(n20488) );
  NAND2_X1 U14091 ( .A1(n12513), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12514) );
  INV_X1 U14092 ( .A(n12515), .ZN(n12517) );
  NOR2_X1 U14093 ( .A1(n12517), .A2(n12516), .ZN(n12518) );
  NAND2_X1 U14094 ( .A1(n17545), .A2(n12521), .ZN(n12522) );
  OR2_X1 U14095 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  NAND2_X1 U14096 ( .A1(n12520), .A2(n12524), .ZN(n12525) );
  INV_X1 U14097 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21943) );
  XNOR2_X1 U14098 ( .A(n12525), .B(n21943), .ZN(n15608) );
  NAND2_X1 U14099 ( .A1(n12525), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12526) );
  INV_X2 U14100 ( .A(n16779), .ZN(n20516) );
  XNOR2_X1 U14101 ( .A(n16778), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15771) );
  INV_X1 U14102 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21960) );
  INV_X1 U14103 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21873) );
  NAND2_X1 U14104 ( .A1(n12520), .A2(n21873), .ZN(n12528) );
  NAND2_X1 U14105 ( .A1(n16653), .A2(n12528), .ZN(n16668) );
  INV_X1 U14106 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16803) );
  NAND2_X1 U14107 ( .A1(n12520), .A2(n16803), .ZN(n16666) );
  NAND2_X1 U14108 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U14109 ( .A1(n12520), .A2(n12529), .ZN(n16664) );
  NAND2_X1 U14110 ( .A1(n16666), .A2(n16664), .ZN(n12530) );
  NOR2_X1 U14111 ( .A1(n16668), .A2(n12530), .ZN(n16651) );
  INV_X1 U14112 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21867) );
  NAND2_X1 U14113 ( .A1(n16778), .A2(n21867), .ZN(n12531) );
  NAND2_X1 U14114 ( .A1(n16651), .A2(n12531), .ZN(n16640) );
  AND2_X1 U14115 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21984) );
  NAND2_X1 U14116 ( .A1(n21984), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n21975) );
  NOR2_X1 U14117 ( .A1(n16640), .A2(n12532), .ZN(n12533) );
  INV_X1 U14118 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16796) );
  INV_X1 U14119 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16170) );
  NAND2_X1 U14120 ( .A1(n16796), .A2(n16170), .ZN(n21982) );
  NOR2_X1 U14121 ( .A1(n21982), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12536) );
  NOR2_X1 U14122 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12534) );
  OR2_X1 U14123 ( .A1(n12520), .A2(n12534), .ZN(n16662) );
  OR2_X1 U14124 ( .A1(n12520), .A2(n16803), .ZN(n16665) );
  OR2_X1 U14125 ( .A1(n12520), .A2(n21867), .ZN(n12535) );
  NAND3_X1 U14126 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16218) );
  INV_X1 U14127 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16615) );
  NOR2_X1 U14128 ( .A1(n16218), .A2(n16615), .ZN(n12538) );
  INV_X1 U14129 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21995) );
  INV_X1 U14130 ( .A(n13658), .ZN(n16593) );
  AND2_X1 U14131 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16735) );
  NAND2_X1 U14132 ( .A1(n16735), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16726) );
  INV_X1 U14133 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16721) );
  NOR3_X1 U14134 ( .A1(n16593), .A2(n16726), .A3(n16721), .ZN(n12541) );
  INV_X1 U14135 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20515) );
  INV_X1 U14136 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16583) );
  NAND2_X1 U14137 ( .A1(n20515), .A2(n16583), .ZN(n16743) );
  NOR4_X1 U14138 ( .A1(n13658), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n16743), .ZN(n12540) );
  MUX2_X1 U14139 ( .A(n16721), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n20516), .Z(n12539) );
  OAI21_X1 U14140 ( .B1(n12541), .B2(n12540), .A(n12539), .ZN(n12542) );
  INV_X1 U14141 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16201) );
  XNOR2_X1 U14142 ( .A(n12542), .B(n16201), .ZN(n16713) );
  XNOR2_X1 U14143 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12561) );
  INV_X1 U14144 ( .A(n12561), .ZN(n12543) );
  XNOR2_X1 U14145 ( .A(n12543), .B(n12562), .ZN(n13803) );
  OAI22_X1 U14146 ( .A1(n12579), .A2(n13803), .B1(n22153), .B2(n11832), .ZN(
        n12556) );
  INV_X1 U14147 ( .A(n13803), .ZN(n12544) );
  NAND2_X1 U14148 ( .A1(n11828), .A2(n12544), .ZN(n12555) );
  AND2_X1 U14149 ( .A1(n11419), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12545) );
  NOR2_X1 U14150 ( .A1(n12562), .A2(n12545), .ZN(n12548) );
  NAND2_X1 U14151 ( .A1(n12582), .A2(n12548), .ZN(n12547) );
  NAND2_X1 U14152 ( .A1(n12547), .A2(n12593), .ZN(n12554) );
  NAND2_X1 U14153 ( .A1(n12549), .A2(n12548), .ZN(n12550) );
  NAND3_X1 U14154 ( .A1(n12550), .A2(n14245), .A3(n14076), .ZN(n12552) );
  NAND2_X1 U14155 ( .A1(n14532), .A2(n14245), .ZN(n12551) );
  NAND2_X1 U14156 ( .A1(n12551), .A2(n11828), .ZN(n12568) );
  NAND2_X1 U14157 ( .A1(n12552), .A2(n12568), .ZN(n12553) );
  OAI211_X1 U14158 ( .C1(n12556), .C2(n12555), .A(n12554), .B(n12553), .ZN(
        n12560) );
  OAI21_X1 U14159 ( .B1(n12557), .B2(n13803), .A(n12556), .ZN(n12559) );
  NAND3_X1 U14160 ( .A1(n12582), .A2(n15294), .A3(n13803), .ZN(n12558) );
  NAND3_X1 U14161 ( .A1(n12560), .A2(n12559), .A3(n12558), .ZN(n12567) );
  NAND2_X1 U14162 ( .A1(n12562), .A2(n12561), .ZN(n12564) );
  NAND2_X1 U14163 ( .A1(n17517), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12563) );
  NAND2_X1 U14164 ( .A1(n12564), .A2(n12563), .ZN(n12571) );
  XNOR2_X1 U14165 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12570) );
  INV_X1 U14166 ( .A(n12570), .ZN(n12565) );
  XNOR2_X1 U14167 ( .A(n12571), .B(n12565), .ZN(n13804) );
  NAND2_X1 U14168 ( .A1(n12582), .A2(n13804), .ZN(n12569) );
  OAI211_X1 U14169 ( .C1(n13804), .C2(n12579), .A(n12569), .B(n12568), .ZN(
        n12566) );
  NAND2_X1 U14170 ( .A1(n12567), .A2(n12566), .ZN(n12581) );
  OR2_X1 U14171 ( .A1(n12569), .A2(n12568), .ZN(n12580) );
  NAND2_X1 U14172 ( .A1(n12571), .A2(n12570), .ZN(n12573) );
  NAND2_X1 U14173 ( .A1(n17523), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12572) );
  NAND2_X1 U14174 ( .A1(n12573), .A2(n12572), .ZN(n12576) );
  XNOR2_X1 U14175 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12575) );
  XNOR2_X1 U14176 ( .A(n12576), .B(n12575), .ZN(n12578) );
  NOR2_X1 U14177 ( .A1(n11702), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12574) );
  AOI21_X1 U14178 ( .B1(n12576), .B2(n12575), .A(n12574), .ZN(n12585) );
  AND2_X1 U14179 ( .A1(n12585), .A2(n12584), .ZN(n12583) );
  AND2_X1 U14180 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12583), .ZN(
        n12577) );
  INV_X1 U14181 ( .A(n12582), .ZN(n12591) );
  INV_X1 U14182 ( .A(n12583), .ZN(n12587) );
  OAI21_X1 U14183 ( .B1(n12585), .B2(n12584), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U14184 ( .A1(n12587), .A2(n12586), .ZN(n13808) );
  INV_X1 U14185 ( .A(n12593), .ZN(n12588) );
  NAND2_X1 U14186 ( .A1(n12588), .A2(n13802), .ZN(n12590) );
  NAND2_X1 U14187 ( .A1(n22153), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12589) );
  OAI211_X1 U14188 ( .C1(n12591), .C2(n13808), .A(n12590), .B(n12589), .ZN(
        n12592) );
  OR2_X1 U14189 ( .A1(n14043), .A2(n13821), .ZN(n13842) );
  OR2_X1 U14190 ( .A1(n13821), .A2(n11829), .ZN(n15079) );
  NAND2_X1 U14191 ( .A1(n13842), .A2(n15079), .ZN(n12596) );
  NAND2_X1 U14192 ( .A1(n14098), .A2(n11838), .ZN(n12595) );
  NAND2_X1 U14193 ( .A1(n13834), .A2(n13823), .ZN(n17539) );
  NAND2_X1 U14194 ( .A1(n17549), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22162) );
  NOR2_X1 U14195 ( .A1(n17539), .A2(n22162), .ZN(n12597) );
  NAND2_X1 U14196 ( .A1(n22290), .A2(n12602), .ZN(n21840) );
  NAND2_X1 U14197 ( .A1(n21840), .A2(n22153), .ZN(n12598) );
  NOR2_X1 U14198 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12293), .ZN(n17548) );
  INV_X1 U14199 ( .A(n17548), .ZN(n12600) );
  NAND2_X1 U14200 ( .A1(n22256), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12599) );
  AND2_X1 U14201 ( .A1(n12600), .A2(n12599), .ZN(n13963) );
  INV_X1 U14202 ( .A(n13963), .ZN(n12601) );
  INV_X1 U14203 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13663) );
  NOR2_X1 U14204 ( .A1(n12602), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21906) );
  NAND2_X1 U14205 ( .A1(n21906), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16707) );
  OAI21_X1 U14206 ( .B1(n16670), .B2(n13663), .A(n16707), .ZN(n12603) );
  AOI21_X1 U14207 ( .B1(n16306), .B2(n20505), .A(n12603), .ZN(n12604) );
  INV_X1 U14208 ( .A(n12605), .ZN(n12606) );
  MUX2_X1 U14209 ( .A(n19807), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12644) );
  NAND2_X1 U14210 ( .A1(n12644), .A2(n12643), .ZN(n12608) );
  NAND2_X1 U14211 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19807), .ZN(
        n12607) );
  MUX2_X1 U14212 ( .A(n19787), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n17422), .Z(n12639) );
  NAND2_X1 U14213 ( .A1(n17422), .A2(n19787), .ZN(n12609) );
  INV_X1 U14214 ( .A(n12615), .ZN(n12610) );
  INV_X1 U14215 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17497) );
  NOR2_X1 U14216 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17497), .ZN(
        n12612) );
  NAND3_X1 U14217 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12613), .A3(
        n19065), .ZN(n12769) );
  XNOR2_X1 U14218 ( .A(n12615), .B(n12614), .ZN(n12786) );
  NAND2_X1 U14219 ( .A1(n12769), .A2(n12786), .ZN(n12679) );
  AND2_X4 U14220 ( .A1(n14598), .A2(n14282), .ZN(n15970) );
  AOI22_X1 U14221 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U14222 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U14223 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12617) );
  INV_X2 U14224 ( .A(n16131), .ZN(n12755) );
  AOI22_X1 U14225 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12755), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12616) );
  NAND4_X1 U14226 ( .A1(n12619), .A2(n12618), .A3(n12617), .A4(n12616), .ZN(
        n12625) );
  AOI22_X1 U14227 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U14228 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U14229 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U14230 ( .A1(n11185), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12755), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12620) );
  NAND4_X1 U14231 ( .A1(n12623), .A2(n12622), .A3(n12621), .A4(n12620), .ZN(
        n12624) );
  AOI22_X1 U14232 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U14233 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U14234 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12626) );
  INV_X2 U14235 ( .A(n16124), .ZN(n14587) );
  AOI22_X1 U14236 ( .A1(n11185), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12755), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12627) );
  NAND4_X1 U14237 ( .A1(n12630), .A2(n12629), .A3(n12628), .A4(n12627), .ZN(
        n12637) );
  AOI22_X1 U14238 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U14239 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U14240 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12634) );
  INV_X2 U14241 ( .A(n16131), .ZN(n12727) );
  AOI22_X1 U14242 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12633) );
  NAND3_X1 U14243 ( .A1(n12635), .A2(n12634), .A3(n12633), .ZN(n12636) );
  NAND2_X2 U14244 ( .A1(n13189), .A2(n15241), .ZN(n13603) );
  OAI21_X1 U14245 ( .B1(n12640), .B2(n12639), .A(n12638), .ZN(n12680) );
  INV_X1 U14246 ( .A(n12680), .ZN(n12641) );
  NAND2_X1 U14247 ( .A1(n15241), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12654) );
  AOI21_X1 U14248 ( .B1(n12654), .B2(n19060), .A(n12641), .ZN(n12649) );
  INV_X4 U14249 ( .A(n13189), .ZN(n16097) );
  INV_X2 U14250 ( .A(n15241), .ZN(n20177) );
  OAI21_X1 U14251 ( .B1(n19819), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12642), .ZN(n12770) );
  INV_X1 U14252 ( .A(n12644), .ZN(n12771) );
  OAI21_X1 U14253 ( .B1(n12770), .B2(n12771), .A(n15234), .ZN(n12647) );
  INV_X1 U14254 ( .A(n12770), .ZN(n13429) );
  XNOR2_X1 U14255 ( .A(n12644), .B(n12643), .ZN(n12681) );
  INV_X1 U14256 ( .A(n12681), .ZN(n12645) );
  OAI211_X1 U14257 ( .C1(n19060), .C2(n13429), .A(n20177), .B(n12645), .ZN(
        n12646) );
  OAI211_X1 U14258 ( .C1(n12823), .C2(n12680), .A(n12647), .B(n12646), .ZN(
        n12648) );
  OAI21_X1 U14259 ( .B1(n13411), .B2(n12649), .A(n12648), .ZN(n12651) );
  NAND2_X1 U14260 ( .A1(n12679), .A2(n15234), .ZN(n12650) );
  OAI21_X1 U14261 ( .B1(n12679), .B2(n12651), .A(n12650), .ZN(n12652) );
  NAND2_X1 U14262 ( .A1(n12790), .A2(n13865), .ZN(n12655) );
  NAND2_X1 U14263 ( .A1(n14646), .A2(n19060), .ZN(n14304) );
  AOI22_X1 U14264 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12660) );
  CLKBUF_X3 U14265 ( .A(n12656), .Z(n16135) );
  AOI22_X1 U14266 ( .A1(n16135), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U14267 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U14268 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U14269 ( .A1(n16135), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U14270 ( .A1(n11166), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U14271 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U14272 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19164) );
  INV_X1 U14273 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n17736) );
  NAND2_X1 U14274 ( .A1(n17492), .A2(n17736), .ZN(n22199) );
  OAI21_X1 U14275 ( .B1(n22205), .B2(n22199), .A(n17745), .ZN(n18722) );
  NAND2_X1 U14276 ( .A1(n19164), .A2(n18722), .ZN(n14663) );
  INV_X1 U14277 ( .A(n14663), .ZN(n14647) );
  NAND2_X1 U14278 ( .A1(n12793), .A2(n14647), .ZN(n12800) );
  AOI22_X1 U14279 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U14280 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U14281 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12665) );
  NAND4_X1 U14282 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12669) );
  NAND2_X1 U14283 ( .A1(n12669), .A2(n14603), .ZN(n12676) );
  AOI22_X1 U14284 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U14285 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U14286 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12755), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12670) );
  NAND4_X1 U14287 ( .A1(n12673), .A2(n12672), .A3(n12671), .A4(n12670), .ZN(
        n12674) );
  AOI21_X1 U14288 ( .B1(n12677), .B2(n20177), .A(n19967), .ZN(n12678) );
  NAND2_X1 U14289 ( .A1(n14304), .A2(n12678), .ZN(n12799) );
  OR2_X1 U14290 ( .A1(n12680), .A2(n12679), .ZN(n12684) );
  NOR2_X1 U14291 ( .A1(n12681), .A2(n12684), .ZN(n12682) );
  OR2_X1 U14292 ( .A1(n12790), .A2(n12682), .ZN(n14638) );
  INV_X1 U14293 ( .A(n14638), .ZN(n12683) );
  OAI21_X1 U14294 ( .B1(n12770), .B2(n12684), .A(n12683), .ZN(n12685) );
  INV_X1 U14295 ( .A(n12685), .ZN(n12686) );
  NAND2_X1 U14296 ( .A1(n12686), .A2(n15237), .ZN(n12691) );
  NAND2_X1 U14297 ( .A1(n12687), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U14298 ( .A1(n12688), .A2(n19065), .ZN(n19059) );
  INV_X1 U14299 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12689) );
  OAI21_X1 U14300 ( .B1(n13303), .B2(n19059), .A(n12689), .ZN(n12690) );
  NAND2_X1 U14301 ( .A1(n12690), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17683) );
  NAND2_X1 U14302 ( .A1(n12691), .A2(n17683), .ZN(n19156) );
  AOI22_X1 U14303 ( .A1(n16135), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U14304 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U14305 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U14306 ( .A1(n11185), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12692) );
  NAND4_X1 U14307 ( .A1(n12695), .A2(n12694), .A3(n12693), .A4(n12692), .ZN(
        n12701) );
  AOI22_X1 U14308 ( .A1(n16135), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U14309 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U14310 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U14311 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12696) );
  NAND4_X1 U14312 ( .A1(n12699), .A2(n12698), .A3(n12697), .A4(n12696), .ZN(
        n12700) );
  AOI22_X1 U14313 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U14314 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U14315 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U14316 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U14317 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12711) );
  AOI22_X1 U14318 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U14319 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U14320 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U14321 ( .A1(n11185), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12755), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12706) );
  NAND4_X1 U14322 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n12710) );
  MUX2_X2 U14323 ( .A(n12711), .B(n12710), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12815) );
  INV_X1 U14324 ( .A(n12738), .ZN(n12736) );
  AOI22_X1 U14325 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U14326 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U14327 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12753), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U14328 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12712) );
  NAND4_X1 U14329 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n12712), .ZN(
        n12716) );
  NAND2_X1 U14330 ( .A1(n12716), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12723) );
  AOI22_X1 U14331 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U14332 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U14333 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12717) );
  NAND4_X1 U14334 ( .A1(n12720), .A2(n12719), .A3(n12718), .A4(n12717), .ZN(
        n12721) );
  NAND2_X1 U14335 ( .A1(n12721), .A2(n14603), .ZN(n12722) );
  INV_X2 U14336 ( .A(n14153), .ZN(n15649) );
  AOI22_X1 U14337 ( .A1(n12756), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11186), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U14338 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16134), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U14339 ( .A1(n11167), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U14340 ( .A1(n14587), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12727), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12728) );
  NAND4_X1 U14341 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12732) );
  NAND2_X1 U14342 ( .A1(n12732), .A2(n14603), .ZN(n12733) );
  NAND2_X1 U14343 ( .A1(n15649), .A2(n12740), .ZN(n12807) );
  INV_X1 U14344 ( .A(n12807), .ZN(n12735) );
  INV_X1 U14345 ( .A(n13604), .ZN(n12737) );
  NAND3_X1 U14346 ( .A1(n19156), .A2(n12737), .A3(n19060), .ZN(n12797) );
  NAND2_X1 U14347 ( .A1(n14665), .A2(n14647), .ZN(n12739) );
  OR2_X1 U14348 ( .A1(n14638), .A2(n12739), .ZN(n12752) );
  NAND2_X2 U14349 ( .A1(n12740), .A2(n14153), .ZN(n12824) );
  NAND2_X1 U14350 ( .A1(n12824), .A2(n13389), .ZN(n12742) );
  NAND2_X1 U14351 ( .A1(n14153), .A2(n19967), .ZN(n12741) );
  NAND3_X1 U14352 ( .A1(n12742), .A2(n12815), .A3(n12741), .ZN(n12809) );
  NAND3_X1 U14353 ( .A1(n19967), .A2(n12740), .A3(n12793), .ZN(n12743) );
  NAND2_X1 U14354 ( .A1(n12824), .A2(n13381), .ZN(n12802) );
  NAND2_X1 U14355 ( .A1(n12802), .A2(n20069), .ZN(n12744) );
  NAND2_X1 U14356 ( .A1(n19062), .A2(n12744), .ZN(n12751) );
  NAND2_X1 U14357 ( .A1(n16097), .A2(n13381), .ZN(n13377) );
  INV_X2 U14358 ( .A(n12815), .ZN(n15212) );
  AOI21_X1 U14359 ( .B1(n13377), .B2(n20177), .A(n15212), .ZN(n12746) );
  NAND2_X1 U14360 ( .A1(n12747), .A2(n19967), .ZN(n12804) );
  OAI211_X1 U14361 ( .C1(n12746), .C2(n12793), .A(n12804), .B(n12832), .ZN(
        n12749) );
  INV_X1 U14362 ( .A(n12747), .ZN(n12748) );
  NAND2_X1 U14363 ( .A1(n16097), .A2(n15241), .ZN(n18721) );
  AOI21_X1 U14364 ( .B1(n12748), .B2(n12815), .A(n18721), .ZN(n13387) );
  NOR2_X1 U14365 ( .A1(n12749), .A2(n13387), .ZN(n12750) );
  AND2_X1 U14366 ( .A1(n12752), .A2(n13379), .ZN(n14297) );
  INV_X1 U14367 ( .A(n12753), .ZN(n15925) );
  AND2_X2 U14368 ( .A1(n12754), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13304) );
  AOI22_X1 U14369 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U14370 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12759) );
  AND2_X1 U14371 ( .A1(n15970), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12774) );
  AOI22_X1 U14372 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12758) );
  AND2_X1 U14373 ( .A1(n12756), .A2(n14603), .ZN(n12939) );
  AOI22_X1 U14374 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12757) );
  NAND4_X1 U14375 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12768) );
  AND2_X1 U14376 ( .A1(n16134), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12779) );
  AOI22_X1 U14377 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12766) );
  AND2_X2 U14378 ( .A1(n11186), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14285) );
  AOI22_X1 U14379 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U14380 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n16060), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12764) );
  AND2_X2 U14381 ( .A1(n14608), .A2(n15926), .ZN(n16062) );
  AND2_X1 U14382 ( .A1(n12762), .A2(n15926), .ZN(n12932) );
  AOI22_X1 U14383 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12763) );
  NAND4_X1 U14384 ( .A1(n12766), .A2(n12765), .A3(n12764), .A4(n12763), .ZN(
        n12767) );
  MUX2_X1 U14385 ( .A(n12769), .B(n13222), .S(n15234), .Z(n13408) );
  INV_X1 U14386 ( .A(n13408), .ZN(n12789) );
  NOR2_X1 U14387 ( .A1(n12771), .A2(n12770), .ZN(n12787) );
  AOI22_X1 U14388 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U14389 ( .A1(n13303), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12773), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U14390 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U14391 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12952), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12775) );
  NAND4_X1 U14392 ( .A1(n12778), .A2(n12777), .A3(n12776), .A4(n12775), .ZN(
        n12785) );
  AOI22_X1 U14393 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U14394 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U14395 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12932), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12781) );
  AOI22_X1 U14396 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n16062), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12780) );
  NAND4_X1 U14397 ( .A1(n12783), .A2(n12782), .A3(n12781), .A4(n12780), .ZN(
        n12784) );
  OAI21_X1 U14398 ( .B1(n13411), .B2(n12787), .A(n13417), .ZN(n12788) );
  NOR2_X1 U14399 ( .A1(n12789), .A2(n12788), .ZN(n12791) );
  OR2_X1 U14400 ( .A1(n12791), .A2(n12790), .ZN(n14636) );
  INV_X1 U14401 ( .A(n14636), .ZN(n12792) );
  NOR2_X1 U14402 ( .A1(n13604), .A2(n18721), .ZN(n14635) );
  NAND2_X1 U14403 ( .A1(n12792), .A2(n14635), .ZN(n13622) );
  MUX2_X1 U14404 ( .A(n14665), .B(n12793), .S(n16097), .Z(n12794) );
  NAND2_X1 U14405 ( .A1(n12794), .A2(n19164), .ZN(n12795) );
  OR2_X1 U14406 ( .A1(n14638), .A2(n12795), .ZN(n12796) );
  OAI211_X1 U14407 ( .C1(n14304), .C2(n12800), .A(n12799), .B(n12798), .ZN(
        n12801) );
  NAND3_X1 U14408 ( .A1(n15237), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19171) );
  AND2_X1 U14409 ( .A1(n12802), .A2(n12815), .ZN(n12803) );
  NAND2_X1 U14410 ( .A1(n12807), .A2(n20069), .ZN(n12808) );
  OAI21_X1 U14411 ( .B1(n12809), .B2(n12808), .A(n20177), .ZN(n12810) );
  NAND2_X1 U14412 ( .A1(n11686), .A2(n20177), .ZN(n12811) );
  AND2_X1 U14413 ( .A1(n20069), .A2(n19060), .ZN(n12812) );
  NAND2_X1 U14414 ( .A1(n13604), .A2(n12812), .ZN(n13185) );
  INV_X1 U14415 ( .A(n12820), .ZN(n12829) );
  NAND3_X1 U14416 ( .A1(n13185), .A2(n13865), .A3(n12829), .ZN(n12848) );
  NAND2_X1 U14417 ( .A1(n12876), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12822) );
  INV_X1 U14418 ( .A(n12823), .ZN(n12814) );
  AND2_X1 U14419 ( .A1(n12815), .A2(n15649), .ZN(n15214) );
  INV_X1 U14420 ( .A(n15214), .ZN(n12816) );
  NOR2_X1 U14421 ( .A1(n12816), .A2(n12740), .ZN(n12817) );
  NAND2_X1 U14422 ( .A1(n15204), .A2(n12817), .ZN(n12819) );
  NOR2_X1 U14423 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12877) );
  NAND2_X1 U14424 ( .A1(n12822), .A2(n12821), .ZN(n12841) );
  INV_X1 U14425 ( .A(n12841), .ZN(n12840) );
  NAND2_X1 U14426 ( .A1(n13603), .A2(n12745), .ZN(n12827) );
  INV_X1 U14427 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15227) );
  NOR2_X1 U14428 ( .A1(n12832), .A2(n13603), .ZN(n12833) );
  AND2_X2 U14429 ( .A1(n15203), .A2(n12833), .ZN(n13394) );
  AND2_X4 U14430 ( .A1(n13394), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12856) );
  NOR2_X1 U14431 ( .A1(n12837), .A2(n12836), .ZN(n12838) );
  OAI21_X2 U14432 ( .B1(n12872), .B2(n15227), .A(n12838), .ZN(n12842) );
  INV_X1 U14433 ( .A(n12842), .ZN(n12839) );
  NAND2_X1 U14434 ( .A1(n12840), .A2(n12839), .ZN(n12862) );
  NAND2_X1 U14435 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  NAND2_X1 U14436 ( .A1(n12844), .A2(n11686), .ZN(n12845) );
  INV_X1 U14437 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12850) );
  INV_X1 U14438 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15368) );
  INV_X1 U14439 ( .A(n12877), .ZN(n19147) );
  OAI21_X1 U14440 ( .B1(n15237), .B2(n15368), .A(n19147), .ZN(n12847) );
  AOI21_X1 U14441 ( .B1(n12856), .B2(P2_EBX_REG_0__SCAN_IN), .A(n12847), .ZN(
        n12849) );
  OAI211_X1 U14442 ( .C1(n12864), .C2(n12850), .A(n12849), .B(n12848), .ZN(
        n12851) );
  INV_X1 U14443 ( .A(n12851), .ZN(n12852) );
  OAI211_X2 U14444 ( .C1(n12854), .C2(n15635), .A(n12853), .B(n12852), .ZN(
        n12888) );
  NAND2_X1 U14445 ( .A1(n15234), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12855) );
  NOR2_X1 U14446 ( .A1(n12855), .A2(n12832), .ZN(n12857) );
  OAI22_X1 U14447 ( .A1(n12876), .A2(n12857), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12856), .ZN(n12861) );
  NAND2_X1 U14448 ( .A1(n12877), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12858) );
  AND2_X1 U14449 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  NAND2_X1 U14450 ( .A1(n12861), .A2(n12860), .ZN(n12889) );
  AOI21_X1 U14451 ( .B1(n15635), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12863) );
  INV_X1 U14452 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n12868) );
  INV_X1 U14453 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12865) );
  NAND2_X1 U14454 ( .A1(n12870), .A2(n12869), .ZN(n12871) );
  INV_X1 U14455 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n15481) );
  NAND2_X1 U14456 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12873) );
  OAI211_X1 U14457 ( .C1(n13097), .C2(n15481), .A(n12874), .B(n12873), .ZN(
        n12875) );
  AOI21_X2 U14458 ( .B1(n13727), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12875), .ZN(n13091) );
  NAND2_X1 U14459 ( .A1(n12876), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12879) );
  NAND2_X1 U14460 ( .A1(n12877), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12878) );
  XNOR2_X2 U14461 ( .A(n13091), .B(n13090), .ZN(n13088) );
  XNOR2_X2 U14462 ( .A(n13089), .B(n13088), .ZN(n14254) );
  INV_X1 U14463 ( .A(n12880), .ZN(n12883) );
  INV_X1 U14464 ( .A(n12881), .ZN(n12882) );
  NAND2_X1 U14465 ( .A1(n12883), .A2(n12882), .ZN(n12884) );
  NAND2_X1 U14466 ( .A1(n12886), .A2(n11220), .ZN(n12887) );
  NAND2_X1 U14467 ( .A1(n14605), .A2(n14615), .ZN(n12904) );
  INV_X1 U14468 ( .A(n12904), .ZN(n12893) );
  AOI22_X1 U14470 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12983), .B1(
        n19682), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12897) );
  OR2_X2 U14471 ( .A1(n14254), .A2(n15322), .ZN(n12905) );
  AOI22_X1 U14472 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12992), .B1(
        n15644), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12896) );
  INV_X1 U14473 ( .A(n12885), .ZN(n12892) );
  AOI22_X1 U14474 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12981), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12895) );
  NOR2_X2 U14475 ( .A1(n12905), .A2(n12902), .ZN(n12982) );
  AND2_X2 U14476 ( .A1(n12903), .A2(n12893), .ZN(n12995) );
  AOI22_X1 U14477 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12982), .B1(
        n12995), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12894) );
  NOR2_X2 U14478 ( .A1(n12901), .A2(n12898), .ZN(n19745) );
  AND2_X2 U14479 ( .A1(n12907), .A2(n12899), .ZN(n19668) );
  AOI22_X1 U14480 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19745), .B1(
        n19668), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U14481 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12990), .B1(
        n12991), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12910) );
  NOR2_X2 U14482 ( .A1(n12901), .A2(n12900), .ZN(n12984) );
  AOI22_X1 U14483 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12984), .B1(
        n12985), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12909) );
  AND2_X2 U14484 ( .A1(n12907), .A2(n12906), .ZN(n12994) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12992), .B1(
        n19682), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U14486 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n15644), .B1(
        n12985), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U14487 ( .A1(n12915), .A2(n12914), .ZN(n12916) );
  NOR2_X1 U14488 ( .A1(n12917), .A2(n12916), .ZN(n12927) );
  INV_X1 U14489 ( .A(n12982), .ZN(n19824) );
  INV_X1 U14490 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12919) );
  NAND2_X1 U14491 ( .A1(n12991), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12918) );
  INV_X1 U14492 ( .A(n12920), .ZN(n12926) );
  AOI22_X1 U14493 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12983), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U14494 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19745), .B1(
        n12995), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U14495 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12990), .B1(
        n19668), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U14496 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12981), .B1(
        n12994), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U14497 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12773), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U14498 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U14499 ( .A1(n13303), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U14500 ( .A1(n12944), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12928) );
  NAND4_X1 U14501 ( .A1(n12931), .A2(n12930), .A3(n12929), .A4(n12928), .ZN(
        n12938) );
  AOI22_X1 U14502 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16060), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U14503 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U14504 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U14505 ( .A1(n12779), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12933) );
  NAND4_X1 U14506 ( .A1(n12936), .A2(n12935), .A3(n12934), .A4(n12933), .ZN(
        n12937) );
  AOI22_X1 U14507 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U14508 ( .A1(n13303), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U14509 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U14510 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12940) );
  NAND4_X1 U14511 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        n12950) );
  AOI22_X1 U14512 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U14513 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12773), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U14514 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n16062), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U14515 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12932), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12945) );
  NAND4_X1 U14516 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12949) );
  AND2_X1 U14517 ( .A1(n16097), .A2(n13428), .ZN(n13950) );
  NAND2_X1 U14518 ( .A1(n13410), .A2(n13950), .ZN(n12968) );
  AOI22_X1 U14519 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U14520 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U14521 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U14522 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12953) );
  NAND4_X1 U14523 ( .A1(n12956), .A2(n12955), .A3(n12954), .A4(n12953), .ZN(
        n12962) );
  AOI22_X1 U14524 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U14525 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n16059), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U14526 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n16060), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U14527 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12957) );
  NAND4_X1 U14528 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        n12961) );
  OR2_X2 U14529 ( .A1(n12962), .A2(n12961), .ZN(n13412) );
  INV_X1 U14530 ( .A(n13412), .ZN(n12963) );
  NAND2_X1 U14531 ( .A1(n12968), .A2(n12963), .ZN(n12964) );
  INV_X1 U14532 ( .A(n13428), .ZN(n12965) );
  XNOR2_X1 U14533 ( .A(n13410), .B(n12965), .ZN(n12966) );
  INV_X1 U14534 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19073) );
  NOR2_X1 U14535 ( .A1(n13950), .A2(n19073), .ZN(n13952) );
  NAND2_X1 U14536 ( .A1(n12966), .A2(n13952), .ZN(n12967) );
  XOR2_X1 U14537 ( .A(n12966), .B(n13952), .Z(n13785) );
  NAND2_X1 U14538 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13785), .ZN(
        n13784) );
  NAND2_X1 U14539 ( .A1(n12967), .A2(n13784), .ZN(n12969) );
  XOR2_X1 U14540 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12969), .Z(
        n13872) );
  XOR2_X1 U14541 ( .A(n13412), .B(n12968), .Z(n13871) );
  NAND2_X1 U14542 ( .A1(n13872), .A2(n13871), .ZN(n13870) );
  NAND2_X1 U14543 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12969), .ZN(
        n12970) );
  NAND2_X1 U14544 ( .A1(n13870), .A2(n12970), .ZN(n12971) );
  INV_X1 U14545 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15516) );
  XNOR2_X1 U14546 ( .A(n12971), .B(n15516), .ZN(n15465) );
  NAND2_X1 U14547 ( .A1(n15466), .A2(n15465), .ZN(n12973) );
  NAND2_X1 U14548 ( .A1(n12971), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12972) );
  NAND2_X1 U14549 ( .A1(n12973), .A2(n12972), .ZN(n12976) );
  XNOR2_X1 U14550 ( .A(n11222), .B(n12980), .ZN(n12977) );
  XNOR2_X1 U14551 ( .A(n12976), .B(n12977), .ZN(n15509) );
  INV_X1 U14552 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15686) );
  NAND2_X1 U14553 ( .A1(n15509), .A2(n15686), .ZN(n15508) );
  INV_X1 U14554 ( .A(n12976), .ZN(n12978) );
  NAND2_X1 U14555 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  INV_X1 U14556 ( .A(n13222), .ZN(n12980) );
  AOI22_X1 U14557 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19798), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U14558 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n12983), .B1(
        n19682), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U14559 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19745), .B1(
        n15644), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U14560 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n12984), .B1(
        n12985), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12986) );
  NAND4_X1 U14561 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n12986), .ZN(
        n13004) );
  AOI22_X1 U14562 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19777), .B1(
        n19759), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U14563 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12992), .B1(
        n19668), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U14564 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n12993), .B1(
        n12994), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13000) );
  INV_X1 U14565 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12997) );
  INV_X1 U14566 ( .A(n12995), .ZN(n12996) );
  INV_X1 U14567 ( .A(n13027), .ZN(n19702) );
  INV_X1 U14568 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13305) );
  OAI22_X1 U14569 ( .A1(n12997), .A2(n12996), .B1(n19702), .B2(n13305), .ZN(
        n12998) );
  INV_X1 U14570 ( .A(n12998), .ZN(n12999) );
  NAND4_X1 U14571 ( .A1(n13002), .A2(n13001), .A3(n13000), .A4(n12999), .ZN(
        n13003) );
  NOR2_X1 U14572 ( .A1(n13004), .A2(n13003), .ZN(n13015) );
  AOI22_X1 U14573 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U14574 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U14575 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U14576 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U14577 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13014) );
  AOI22_X1 U14578 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U14579 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U14580 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n16060), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13010) );
  AOI22_X1 U14581 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13009) );
  NAND4_X1 U14582 ( .A1(n13012), .A2(n13011), .A3(n13010), .A4(n13009), .ZN(
        n13013) );
  NOR2_X1 U14583 ( .A1(n13014), .A2(n13013), .ZN(n13418) );
  INV_X1 U14584 ( .A(n13017), .ZN(n13016) );
  NAND2_X1 U14585 ( .A1(n11347), .A2(n13016), .ZN(n13019) );
  NAND2_X1 U14586 ( .A1(n13018), .A2(n13017), .ZN(n13049) );
  INV_X1 U14587 ( .A(n13053), .ZN(n13021) );
  NAND2_X1 U14588 ( .A1(n13021), .A2(n13020), .ZN(n13022) );
  INV_X1 U14589 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15685) );
  AOI22_X1 U14590 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12982), .B1(
        n12983), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U14591 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19745), .B1(
        n15644), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U14592 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12993), .B1(
        n12985), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U14593 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19759), .B1(
        n12994), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13023) );
  NAND4_X1 U14594 ( .A1(n13026), .A2(n13025), .A3(n13024), .A4(n13023), .ZN(
        n13033) );
  AOI22_X1 U14595 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12984), .B1(
        n19777), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U14596 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12995), .B1(
        n19682), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U14597 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19798), .B1(
        n13027), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13029) );
  AOI22_X1 U14598 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12992), .B1(
        n19668), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13028) );
  NAND4_X1 U14599 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13032) );
  AOI22_X1 U14600 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U14601 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U14602 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U14603 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13034) );
  NAND4_X1 U14604 ( .A1(n13037), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        n13043) );
  AOI22_X1 U14605 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U14606 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U14607 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U14608 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13038) );
  NAND4_X1 U14609 ( .A1(n13041), .A2(n13040), .A3(n13039), .A4(n13038), .ZN(
        n13042) );
  INV_X1 U14610 ( .A(n13449), .ZN(n13044) );
  NAND2_X1 U14611 ( .A1(n13044), .A2(n16097), .ZN(n13045) );
  NOR2_X1 U14612 ( .A1(n13049), .A2(n13048), .ZN(n13047) );
  INV_X1 U14613 ( .A(n13047), .ZN(n13060) );
  NAND2_X1 U14614 ( .A1(n13049), .A2(n13048), .ZN(n13050) );
  INV_X1 U14615 ( .A(n13452), .ZN(n13058) );
  AND2_X1 U14616 ( .A1(n13051), .A2(n15685), .ZN(n13052) );
  OR2_X1 U14617 ( .A1(n13053), .A2(n13052), .ZN(n13055) );
  NAND3_X1 U14618 ( .A1(n13020), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n13048), .ZN(n13054) );
  NAND2_X1 U14619 ( .A1(n13059), .A2(n13058), .ZN(n17151) );
  AOI22_X1 U14620 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U14621 ( .A1(n13303), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U14622 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12773), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U14623 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13061) );
  NAND4_X1 U14624 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13070) );
  AOI22_X1 U14625 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U14626 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U14627 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16060), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U14628 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13065) );
  NAND4_X1 U14629 ( .A1(n13068), .A2(n13067), .A3(n13066), .A4(n13065), .ZN(
        n13069) );
  INV_X1 U14630 ( .A(n13073), .ZN(n13071) );
  NAND2_X1 U14631 ( .A1(n13071), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13072) );
  AND2_X1 U14632 ( .A1(n17151), .A2(n13072), .ZN(n13075) );
  INV_X1 U14633 ( .A(n13072), .ZN(n13074) );
  XNOR2_X1 U14634 ( .A(n13073), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17153) );
  NAND2_X1 U14635 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13077) );
  INV_X1 U14636 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17368) );
  NAND2_X1 U14637 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17364) );
  NOR2_X1 U14638 ( .A1(n17368), .A2(n17364), .ZN(n17334) );
  NAND4_X1 U14639 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n17334), .ZN(n17271) );
  INV_X1 U14640 ( .A(n17271), .ZN(n17265) );
  INV_X1 U14641 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13522) );
  NAND3_X1 U14642 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17267) );
  NOR2_X1 U14643 ( .A1(n13522), .A2(n17267), .ZN(n17273) );
  AND2_X1 U14644 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17273), .ZN(
        n17275) );
  NAND2_X1 U14645 ( .A1(n17275), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13405) );
  INV_X1 U14646 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17258) );
  AND2_X1 U14647 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17231) );
  INV_X1 U14648 ( .A(n17231), .ZN(n13406) );
  NAND2_X1 U14649 ( .A1(n17099), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17216) );
  INV_X1 U14650 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13590) );
  INV_X1 U14651 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13570) );
  AND2_X1 U14652 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13640) );
  NAND2_X1 U14653 ( .A1(n13640), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13735) );
  XNOR2_X1 U14654 ( .A(n13716), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17040) );
  NAND2_X1 U14655 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13087) );
  INV_X1 U14656 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17217) );
  NAND2_X1 U14657 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13083) );
  OAI211_X1 U14658 ( .C1(n13730), .C2(n17217), .A(n13084), .B(n13083), .ZN(
        n13085) );
  INV_X1 U14659 ( .A(n13085), .ZN(n13086) );
  NAND2_X1 U14660 ( .A1(n13087), .A2(n13086), .ZN(n16934) );
  INV_X1 U14661 ( .A(n13090), .ZN(n13092) );
  NAND2_X1 U14662 ( .A1(n13092), .A2(n13091), .ZN(n13093) );
  NAND2_X1 U14663 ( .A1(n13094), .A2(n13093), .ZN(n14237) );
  INV_X1 U14664 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n13221) );
  NAND2_X1 U14665 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13095) );
  OAI211_X1 U14666 ( .C1(n13097), .C2(n13221), .A(n13096), .B(n13095), .ZN(
        n13098) );
  AOI21_X1 U14667 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13098), .ZN(n14236) );
  INV_X1 U14668 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13230) );
  NAND2_X1 U14669 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13100) );
  OAI211_X1 U14670 ( .C1(n13730), .C2(n13230), .A(n13101), .B(n13100), .ZN(
        n13102) );
  AOI21_X1 U14671 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13102), .ZN(n14230) );
  INV_X1 U14672 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U14673 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13104) );
  AOI22_X1 U14674 ( .A1(n12856), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13103) );
  OAI211_X1 U14675 ( .C1(n13730), .C2(n13105), .A(n13104), .B(n13103), .ZN(
        n14260) );
  INV_X1 U14676 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n17160) );
  NAND2_X1 U14677 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13106) );
  OAI211_X1 U14678 ( .C1(n13730), .C2(n17160), .A(n13107), .B(n13106), .ZN(
        n13108) );
  AOI21_X1 U14679 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13108), .ZN(n14276) );
  INV_X1 U14680 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U14681 ( .A1(n12856), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13111) );
  NAND2_X1 U14682 ( .A1(n13109), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n13110) );
  OAI211_X1 U14683 ( .C1(n13112), .C2(n13465), .A(n13111), .B(n13110), .ZN(
        n14320) );
  INV_X1 U14684 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n17147) );
  NAND2_X1 U14685 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13113) );
  OAI211_X1 U14686 ( .C1(n13730), .C2(n17147), .A(n13114), .B(n13113), .ZN(
        n13115) );
  AOI21_X1 U14687 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n13115), .ZN(n15110) );
  NAND2_X1 U14688 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13120) );
  INV_X1 U14689 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U14690 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13116) );
  OAI211_X1 U14691 ( .C1(n13730), .C2(n13264), .A(n13117), .B(n13116), .ZN(
        n13118) );
  INV_X1 U14692 ( .A(n13118), .ZN(n13119) );
  NAND2_X1 U14693 ( .A1(n13120), .A2(n13119), .ZN(n15265) );
  INV_X1 U14694 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U14695 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13121) );
  OAI211_X1 U14696 ( .C1(n13730), .C2(n13123), .A(n13122), .B(n13121), .ZN(
        n13124) );
  AOI21_X1 U14697 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n13124), .ZN(n15273) );
  INV_X1 U14698 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n13301) );
  NAND2_X1 U14699 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13125) );
  OAI211_X1 U14700 ( .C1(n13730), .C2(n13301), .A(n13126), .B(n13125), .ZN(
        n13127) );
  AOI21_X1 U14701 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n13127), .ZN(n15490) );
  INV_X1 U14702 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U14703 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13129) );
  OAI211_X1 U14704 ( .C1(n13730), .C2(n13131), .A(n13130), .B(n13129), .ZN(
        n13132) );
  AOI21_X1 U14705 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n13132), .ZN(n15544) );
  INV_X1 U14706 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U14707 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13134) );
  AOI22_X1 U14708 ( .A1(n12856), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n13133) );
  OAI211_X1 U14709 ( .C1(n13730), .C2(n13320), .A(n13134), .B(n13133), .ZN(
        n15616) );
  INV_X1 U14710 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n18839) );
  NAND2_X1 U14711 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13136) );
  AOI22_X1 U14712 ( .A1(n12856), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n13135) );
  OAI211_X1 U14713 ( .C1(n13730), .C2(n18839), .A(n13136), .B(n13135), .ZN(
        n15629) );
  INV_X1 U14714 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n13139) );
  NAND2_X1 U14715 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13138) );
  AOI22_X1 U14716 ( .A1(n12856), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n13137) );
  OAI211_X1 U14717 ( .C1(n13139), .C2(n13730), .A(n13138), .B(n13137), .ZN(
        n15730) );
  NAND2_X1 U14718 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13145) );
  INV_X1 U14719 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U14720 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13140) );
  OAI211_X1 U14721 ( .C1(n13730), .C2(n13142), .A(n13141), .B(n13140), .ZN(
        n13143) );
  INV_X1 U14722 ( .A(n13143), .ZN(n13144) );
  NAND2_X1 U14723 ( .A1(n13145), .A2(n13144), .ZN(n15792) );
  INV_X1 U14724 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U14725 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13146) );
  OAI211_X1 U14726 ( .C1(n13730), .C2(n13351), .A(n13147), .B(n13146), .ZN(
        n13148) );
  AOI21_X1 U14727 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n13148), .ZN(n15853) );
  INV_X1 U14728 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n18894) );
  NAND2_X1 U14729 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13149) );
  OAI211_X1 U14730 ( .C1(n13730), .C2(n18894), .A(n13150), .B(n13149), .ZN(
        n13151) );
  AOI21_X1 U14731 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n13151), .ZN(n15898) );
  INV_X1 U14732 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n18905) );
  NAND2_X1 U14733 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13152) );
  OAI211_X1 U14734 ( .C1(n13730), .C2(n18905), .A(n13153), .B(n13152), .ZN(
        n13154) );
  AOI21_X1 U14735 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n13154), .ZN(n13632) );
  INV_X1 U14736 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n18917) );
  NAND2_X1 U14737 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13156) );
  AOI22_X1 U14738 ( .A1(n12856), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n13155) );
  OAI211_X1 U14739 ( .C1(n13730), .C2(n18917), .A(n13156), .B(n13155), .ZN(
        n16958) );
  INV_X1 U14740 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U14741 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13158) );
  AOI22_X1 U14742 ( .A1(n12856), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n13157) );
  OAI211_X1 U14743 ( .C1(n13730), .C2(n13360), .A(n13158), .B(n13157), .ZN(
        n16949) );
  INV_X1 U14744 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U14745 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13159) );
  OAI211_X1 U14746 ( .C1(n13730), .C2(n13161), .A(n13160), .B(n13159), .ZN(
        n13162) );
  AOI21_X1 U14747 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n13162), .ZN(n16941) );
  INV_X1 U14748 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17740) );
  NAND2_X1 U14749 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13163) );
  OAI211_X1 U14750 ( .C1(n13730), .C2(n17740), .A(n13164), .B(n13163), .ZN(
        n13165) );
  AOI21_X1 U14751 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n13165), .ZN(n16924) );
  INV_X1 U14752 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17742) );
  NAND2_X1 U14753 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13166) );
  OAI211_X1 U14754 ( .C1(n13730), .C2(n17742), .A(n13167), .B(n13166), .ZN(
        n13168) );
  AOI21_X1 U14755 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13168), .ZN(n16907) );
  INV_X1 U14756 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17741) );
  NAND2_X1 U14757 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13169) );
  OAI211_X1 U14758 ( .C1(n13730), .C2(n17741), .A(n13170), .B(n13169), .ZN(
        n13171) );
  AOI21_X1 U14759 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13171), .ZN(n16916) );
  OR2_X1 U14760 ( .A1(n16907), .A2(n16916), .ZN(n13172) );
  INV_X1 U14761 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17058) );
  NAND2_X1 U14762 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13174) );
  AOI22_X1 U14763 ( .A1(n12856), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n13173) );
  OAI211_X1 U14764 ( .C1(n13730), .C2(n17058), .A(n13174), .B(n13173), .ZN(
        n16899) );
  NAND2_X1 U14765 ( .A1(n16908), .A2(n16899), .ZN(n16901) );
  INV_X1 U14766 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17743) );
  NAND2_X1 U14767 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13175) );
  OAI211_X1 U14768 ( .C1(n13730), .C2(n17743), .A(n13176), .B(n13175), .ZN(
        n13177) );
  AOI21_X1 U14769 ( .B1(n11165), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13177), .ZN(n13642) );
  INV_X1 U14770 ( .A(n13726), .ZN(n13644) );
  INV_X1 U14771 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19023) );
  NAND2_X1 U14772 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13179) );
  AOI22_X1 U14773 ( .A1(n12856), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13178) );
  OAI211_X1 U14774 ( .C1(n13730), .C2(n19023), .A(n13179), .B(n13178), .ZN(
        n13725) );
  NAND2_X1 U14775 ( .A1(n13180), .A2(n16097), .ZN(n13183) );
  INV_X1 U14776 ( .A(n13181), .ZN(n13182) );
  NAND2_X1 U14777 ( .A1(n13183), .A2(n13182), .ZN(n13184) );
  AND2_X1 U14778 ( .A1(n13797), .A2(n19062), .ZN(n14634) );
  NOR2_X1 U14779 ( .A1(n14606), .A2(n13185), .ZN(n14642) );
  INV_X1 U14780 ( .A(n14642), .ZN(n13186) );
  OAI21_X1 U14781 ( .B1(n14634), .B2(n16097), .A(n13186), .ZN(n13187) );
  AND2_X2 U14782 ( .A1(n13192), .A2(n13448), .ZN(n13331) );
  NAND2_X1 U14783 ( .A1(n13331), .A2(n13428), .ZN(n13191) );
  MUX2_X1 U14784 ( .A(n12815), .B(n19819), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13190) );
  AND2_X1 U14785 ( .A1(n13189), .A2(n19733), .ZN(n13215) );
  NAND2_X1 U14786 ( .A1(n15211), .A2(n13215), .ZN(n13205) );
  NAND3_X1 U14787 ( .A1(n13191), .A2(n13190), .A3(n13205), .ZN(n15193) );
  INV_X1 U14788 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n20161) );
  OAI21_X1 U14789 ( .B1(n12815), .B2(n20161), .A(n19733), .ZN(n13193) );
  AOI21_X1 U14790 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13215), .A(
        n13193), .ZN(n13194) );
  INV_X1 U14791 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17738) );
  OR2_X1 U14792 ( .A1(n13722), .A2(n17738), .ZN(n13197) );
  NOR2_X1 U14793 ( .A1(n12815), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U14794 ( .A1(n13195), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13215), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13196) );
  NAND2_X1 U14795 ( .A1(n13197), .A2(n13196), .ZN(n13203) );
  INV_X1 U14796 ( .A(n13203), .ZN(n13198) );
  NAND2_X1 U14797 ( .A1(n13410), .A2(n13331), .ZN(n13201) );
  NAND2_X1 U14798 ( .A1(n12824), .A2(n12815), .ZN(n13199) );
  MUX2_X1 U14799 ( .A(n13199), .B(n19807), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13200) );
  NAND2_X1 U14800 ( .A1(n13201), .A2(n13200), .ZN(n13780) );
  INV_X1 U14801 ( .A(n13780), .ZN(n13202) );
  NAND2_X1 U14802 ( .A1(n13779), .A2(n13202), .ZN(n13783) );
  NAND2_X1 U14803 ( .A1(n13331), .A2(n13412), .ZN(n13206) );
  OAI211_X1 U14804 ( .C1(n19733), .C2(n19787), .A(n13206), .B(n13205), .ZN(
        n13207) );
  AND3_X1 U14805 ( .A1(n13783), .A2(n13208), .A3(n13207), .ZN(n13209) );
  INV_X1 U14806 ( .A(n14136), .ZN(n13214) );
  OR2_X1 U14807 ( .A1(n13722), .A2(n12868), .ZN(n13211) );
  INV_X2 U14808 ( .A(n13363), .ZN(n13720) );
  INV_X1 U14809 ( .A(n13215), .ZN(n13226) );
  AOI22_X1 U14810 ( .A1(n13720), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13215), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U14811 ( .A1(n13211), .A2(n13210), .ZN(n14137) );
  AOI22_X1 U14812 ( .A1(n13348), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13217) );
  NAND2_X1 U14813 ( .A1(n13720), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n13216) );
  AND2_X1 U14814 ( .A1(n13217), .A2(n13216), .ZN(n13220) );
  NAND2_X1 U14815 ( .A1(n13331), .A2(n13218), .ZN(n13219) );
  OAI211_X1 U14816 ( .C1(n13722), .C2(n15481), .A(n13220), .B(n13219), .ZN(
        n15197) );
  OR2_X1 U14817 ( .A1(n13722), .A2(n13221), .ZN(n13225) );
  NAND2_X1 U14818 ( .A1(n13331), .A2(n13222), .ZN(n13224) );
  AOI22_X1 U14819 ( .A1(n13720), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13215), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U14820 ( .A1(n13720), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13348), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13229) );
  INV_X1 U14821 ( .A(n13418), .ZN(n13227) );
  NAND2_X1 U14822 ( .A1(n13331), .A2(n13227), .ZN(n13228) );
  OAI211_X1 U14823 ( .C1(n13722), .C2(n13230), .A(n13229), .B(n13228), .ZN(
        n15233) );
  NAND2_X1 U14824 ( .A1(n13331), .A2(n13449), .ZN(n13231) );
  OR2_X1 U14825 ( .A1(n13722), .A2(n13105), .ZN(n13234) );
  AOI22_X1 U14826 ( .A1(n13720), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13348), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13233) );
  NAND2_X1 U14827 ( .A1(n13234), .A2(n13233), .ZN(n17404) );
  NAND2_X1 U14828 ( .A1(n17403), .A2(n17404), .ZN(n13236) );
  NAND2_X1 U14829 ( .A1(n13331), .A2(n13455), .ZN(n13235) );
  OR2_X1 U14830 ( .A1(n13722), .A2(n17160), .ZN(n13238) );
  AOI22_X1 U14831 ( .A1(n13720), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13348), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U14832 ( .A1(n13238), .A2(n13237), .ZN(n17390) );
  INV_X1 U14833 ( .A(n13331), .ZN(n13347) );
  AOI22_X1 U14834 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U14835 ( .A1(n12772), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U14836 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12773), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U14837 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12952), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13239) );
  NAND4_X1 U14838 ( .A1(n13242), .A2(n13241), .A3(n13240), .A4(n13239), .ZN(
        n13248) );
  AOI22_X1 U14839 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U14840 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U14841 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12932), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U14842 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n16062), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13243) );
  NAND4_X1 U14843 ( .A1(n13246), .A2(n13245), .A3(n13244), .A4(n13243), .ZN(
        n13247) );
  INV_X1 U14844 ( .A(n14324), .ZN(n13250) );
  AOI22_X1 U14845 ( .A1(n13720), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13348), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13249) );
  OAI21_X1 U14846 ( .B1(n13347), .B2(n13250), .A(n13249), .ZN(n13251) );
  AOI21_X1 U14847 ( .B1(n13376), .B2(P2_REIP_REG_8__SCAN_IN), .A(n13251), .ZN(
        n18773) );
  AOI22_X1 U14848 ( .A1(n13720), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13348), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U14849 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U14850 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U14851 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13253) );
  AOI22_X1 U14852 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13252) );
  NAND4_X1 U14853 ( .A1(n13255), .A2(n13254), .A3(n13253), .A4(n13252), .ZN(
        n13261) );
  AOI22_X1 U14854 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13259) );
  AOI22_X1 U14855 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U14856 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U14857 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13256) );
  NAND4_X1 U14858 ( .A1(n13259), .A2(n13258), .A3(n13257), .A4(n13256), .ZN(
        n13260) );
  NAND2_X1 U14859 ( .A1(n13331), .A2(n11696), .ZN(n13262) );
  OAI211_X1 U14860 ( .C1(n13722), .C2(n17147), .A(n13263), .B(n13262), .ZN(
        n17377) );
  OR2_X1 U14861 ( .A1(n13722), .A2(n13264), .ZN(n13277) );
  AOI22_X1 U14862 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12951), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U14863 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U14864 ( .A1(n12772), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U14865 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12773), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13265) );
  NAND4_X1 U14866 ( .A1(n13268), .A2(n13267), .A3(n13266), .A4(n13265), .ZN(
        n13274) );
  AOI22_X1 U14867 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U14868 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12952), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13271) );
  AOI22_X1 U14869 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U14870 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13269) );
  NAND4_X1 U14871 ( .A1(n13272), .A2(n13271), .A3(n13270), .A4(n13269), .ZN(
        n13273) );
  NAND2_X1 U14872 ( .A1(n13331), .A2(n11698), .ZN(n13276) );
  AOI22_X1 U14873 ( .A1(n13720), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13275) );
  AOI22_X1 U14874 ( .A1(n13376), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n13348), .ZN(n13289) );
  AOI22_X1 U14875 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U14876 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U14877 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U14878 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13278) );
  NAND4_X1 U14879 ( .A1(n13281), .A2(n13280), .A3(n13279), .A4(n13278), .ZN(
        n13287) );
  AOI22_X1 U14880 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13285) );
  AOI22_X1 U14881 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13284) );
  AOI22_X1 U14882 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U14883 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13282) );
  NAND4_X1 U14884 ( .A1(n13285), .A2(n13284), .A3(n13283), .A4(n13282), .ZN(
        n13286) );
  OR2_X1 U14885 ( .A1(n13287), .A2(n13286), .ZN(n15495) );
  AOI22_X1 U14886 ( .A1(n13331), .A2(n15495), .B1(n13720), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n13288) );
  NAND2_X1 U14887 ( .A1(n13289), .A2(n13288), .ZN(n17363) );
  AOI22_X1 U14888 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U14889 ( .A1(n12772), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13292) );
  AOI22_X1 U14890 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12773), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13291) );
  AOI22_X1 U14891 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12952), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13290) );
  NAND4_X1 U14892 ( .A1(n13293), .A2(n13292), .A3(n13291), .A4(n13290), .ZN(
        n13299) );
  AOI22_X1 U14893 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U14894 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13296) );
  AOI22_X1 U14895 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12932), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U14896 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n16062), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13294) );
  NAND4_X1 U14897 ( .A1(n13297), .A2(n13296), .A3(n13295), .A4(n13294), .ZN(
        n13298) );
  AOI22_X1 U14898 ( .A1(n13720), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13300) );
  OAI21_X1 U14899 ( .B1(n13722), .B2(n13301), .A(n13300), .ZN(n13302) );
  AOI21_X1 U14900 ( .B1(n13331), .B2(n15499), .A(n13302), .ZN(n17350) );
  AOI22_X1 U14901 ( .A1(n13376), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n13720), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13319) );
  INV_X1 U14902 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13306) );
  INV_X1 U14903 ( .A(n13303), .ZN(n15913) );
  INV_X1 U14904 ( .A(n13304), .ZN(n15912) );
  OAI22_X1 U14905 ( .A1(n13306), .A2(n15913), .B1(n15912), .B2(n13305), .ZN(
        n13307) );
  INV_X1 U14906 ( .A(n13307), .ZN(n13311) );
  AOI22_X1 U14907 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U14908 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U14909 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13308) );
  NAND4_X1 U14910 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13317) );
  AOI22_X1 U14911 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U14912 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U14913 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U14914 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13312) );
  NAND4_X1 U14915 ( .A1(n13315), .A2(n13314), .A3(n13313), .A4(n13312), .ZN(
        n13316) );
  AOI22_X1 U14916 ( .A1(n13331), .A2(n15621), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13348), .ZN(n13318) );
  NAND2_X1 U14917 ( .A1(n13319), .A2(n13318), .ZN(n15561) );
  OR2_X1 U14918 ( .A1(n13722), .A2(n13320), .ZN(n13334) );
  AOI22_X1 U14919 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U14920 ( .A1(n13303), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12773), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U14921 ( .A1(n13304), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13322) );
  AOI22_X1 U14922 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12952), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13321) );
  NAND4_X1 U14923 ( .A1(n13324), .A2(n13323), .A3(n13322), .A4(n13321), .ZN(
        n13330) );
  AOI22_X1 U14924 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U14925 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14285), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13327) );
  AOI22_X1 U14926 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12932), .B1(
        n16061), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13326) );
  AOI22_X1 U14927 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n16062), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13325) );
  NAND4_X1 U14928 ( .A1(n13328), .A2(n13327), .A3(n13326), .A4(n13325), .ZN(
        n13329) );
  OR2_X1 U14929 ( .A1(n13330), .A2(n13329), .ZN(n15620) );
  NAND2_X1 U14930 ( .A1(n13331), .A2(n15620), .ZN(n13333) );
  AOI22_X1 U14931 ( .A1(n13720), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U14932 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n13304), .B1(
        n13303), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U14933 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U14934 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13336) );
  AOI22_X1 U14935 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13335) );
  NAND4_X1 U14936 ( .A1(n13338), .A2(n13337), .A3(n13336), .A4(n13335), .ZN(
        n13344) );
  AOI22_X1 U14937 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U14938 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U14939 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13340) );
  AOI22_X1 U14940 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13339) );
  NAND4_X1 U14941 ( .A1(n13342), .A2(n13341), .A3(n13340), .A4(n13339), .ZN(
        n13343) );
  NOR2_X1 U14942 ( .A1(n13344), .A2(n13343), .ZN(n15626) );
  OR2_X1 U14943 ( .A1(n13722), .A2(n18839), .ZN(n13346) );
  AOI22_X1 U14944 ( .A1(n13720), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13345) );
  OAI211_X1 U14945 ( .C1(n15626), .C2(n13347), .A(n13346), .B(n13345), .ZN(
        n17313) );
  AOI222_X1 U14946 ( .A1(n13376), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n13215), .C1(n13720), .C2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n15749) );
  OR2_X1 U14947 ( .A1(n13722), .A2(n13142), .ZN(n13350) );
  AOI22_X1 U14948 ( .A1(n13720), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13349) );
  NAND2_X1 U14949 ( .A1(n13350), .A2(n13349), .ZN(n15797) );
  OR2_X1 U14950 ( .A1(n13722), .A2(n13351), .ZN(n13353) );
  AOI22_X1 U14951 ( .A1(n13720), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U14952 ( .A1(n13353), .A2(n13352), .ZN(n15818) );
  OR2_X1 U14953 ( .A1(n13722), .A2(n18894), .ZN(n13355) );
  AOI22_X1 U14954 ( .A1(n13720), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13354) );
  OR2_X1 U14955 ( .A1(n13722), .A2(n18905), .ZN(n13357) );
  AOI22_X1 U14956 ( .A1(n13720), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13215), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U14957 ( .A1(n13357), .A2(n13356), .ZN(n17277) );
  OR2_X1 U14958 ( .A1(n13722), .A2(n18917), .ZN(n13359) );
  AOI22_X1 U14959 ( .A1(n13720), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13358) );
  NAND2_X1 U14960 ( .A1(n13359), .A2(n13358), .ZN(n17025) );
  OR2_X1 U14961 ( .A1(n13722), .A2(n13360), .ZN(n13362) );
  AOI22_X1 U14962 ( .A1(n13720), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13215), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13361) );
  AND2_X1 U14963 ( .A1(n13362), .A2(n13361), .ZN(n17239) );
  INV_X1 U14964 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17232) );
  INV_X1 U14965 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n17019) );
  OAI222_X1 U14966 ( .A1(n13226), .A2(n17232), .B1(n13363), .B2(n17019), .C1(
        n13722), .C2(n13161), .ZN(n17018) );
  OR2_X1 U14967 ( .A1(n13722), .A2(n17217), .ZN(n13365) );
  AOI22_X1 U14968 ( .A1(n13720), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13364) );
  OR2_X1 U14969 ( .A1(n13722), .A2(n17740), .ZN(n13367) );
  AOI22_X1 U14970 ( .A1(n13720), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13366) );
  AND2_X1 U14971 ( .A1(n13367), .A2(n13366), .ZN(n16999) );
  OR2_X1 U14972 ( .A1(n13722), .A2(n17741), .ZN(n13369) );
  AOI22_X1 U14973 ( .A1(n13720), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13215), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13368) );
  NAND2_X1 U14974 ( .A1(n13369), .A2(n13368), .ZN(n16990) );
  OR2_X1 U14975 ( .A1(n13722), .A2(n17742), .ZN(n13371) );
  AOI22_X1 U14976 ( .A1(n13720), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U14977 ( .A1(n13371), .A2(n13370), .ZN(n16981) );
  OR2_X1 U14978 ( .A1(n13722), .A2(n17058), .ZN(n13373) );
  AOI22_X1 U14979 ( .A1(n13720), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13215), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13372) );
  NAND2_X1 U14980 ( .A1(n13373), .A2(n13372), .ZN(n16973) );
  OR2_X1 U14981 ( .A1(n13722), .A2(n17743), .ZN(n13375) );
  AOI22_X1 U14982 ( .A1(n13720), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13374) );
  AND2_X1 U14983 ( .A1(n13375), .A2(n13374), .ZN(n13645) );
  AOI222_X1 U14984 ( .A1(n13376), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13348), .C1(n13720), .C2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n13718) );
  NOR2_X2 U14985 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19788) );
  NAND2_X1 U14986 ( .A1(n19788), .A2(n15237), .ZN(n17559) );
  OR2_X1 U14987 ( .A1(n17559), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18892) );
  INV_X1 U14988 ( .A(n19139), .ZN(n18813) );
  OR2_X1 U14989 ( .A1(n18813), .A2(n19023), .ZN(n17034) );
  INV_X1 U14990 ( .A(n13377), .ZN(n13378) );
  NAND2_X1 U14991 ( .A1(n13605), .A2(n14632), .ZN(n14126) );
  NAND3_X1 U14992 ( .A1(n12844), .A2(n13380), .A3(n11686), .ZN(n13393) );
  INV_X1 U14993 ( .A(n14296), .ZN(n13813) );
  OAI21_X1 U14994 ( .B1(n13380), .B2(n13381), .A(n13813), .ZN(n13382) );
  OAI21_X1 U14995 ( .B1(n20177), .B2(n20069), .A(n13382), .ZN(n13383) );
  INV_X1 U14996 ( .A(n13383), .ZN(n13384) );
  AND2_X1 U14997 ( .A1(n13385), .A2(n13384), .ZN(n13392) );
  NAND2_X1 U14998 ( .A1(n13386), .A2(n19060), .ZN(n14607) );
  INV_X1 U14999 ( .A(n13387), .ZN(n13388) );
  NAND2_X1 U15000 ( .A1(n14607), .A2(n13388), .ZN(n13390) );
  NAND2_X1 U15001 ( .A1(n13390), .A2(n13389), .ZN(n13391) );
  AND3_X1 U15002 ( .A1(n13393), .A2(n13392), .A3(n13391), .ZN(n14614) );
  INV_X1 U15003 ( .A(n13394), .ZN(n14589) );
  NAND2_X1 U15004 ( .A1(n14614), .A2(n14589), .ZN(n13395) );
  NAND2_X1 U15005 ( .A1(n13605), .A2(n13395), .ZN(n17319) );
  INV_X1 U15006 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17401) );
  NAND3_X1 U15007 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13403) );
  NOR2_X1 U15008 ( .A1(n17401), .A2(n13403), .ZN(n17389) );
  NAND3_X1 U15009 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n17389), .ZN(n13396) );
  NAND2_X1 U15010 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14129) );
  NAND2_X1 U15011 ( .A1(n12865), .A2(n14129), .ZN(n14127) );
  INV_X1 U15012 ( .A(n18892), .ZN(n19095) );
  OR2_X1 U15013 ( .A1(n13605), .A2(n19095), .ZN(n19074) );
  OAI21_X1 U15014 ( .B1(n14126), .B2(n14127), .A(n19074), .ZN(n15468) );
  AOI21_X1 U15015 ( .B1(n19106), .B2(n13396), .A(n15468), .ZN(n17269) );
  NOR2_X1 U15016 ( .A1(n12865), .A2(n14129), .ZN(n15470) );
  INV_X1 U15017 ( .A(n15470), .ZN(n14128) );
  NOR2_X1 U15018 ( .A1(n14128), .A2(n13396), .ZN(n17266) );
  OR2_X1 U15019 ( .A1(n17319), .A2(n17266), .ZN(n13397) );
  NAND2_X1 U15020 ( .A1(n17269), .A2(n13397), .ZN(n17381) );
  NAND3_X1 U15021 ( .A1(n17265), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n13079), .ZN(n13398) );
  OAI21_X1 U15022 ( .B1(n17381), .B2(n13398), .A(n13399), .ZN(n17257) );
  OAI211_X1 U15023 ( .C1(n17231), .C2(n19109), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17257), .ZN(n17219) );
  NAND2_X1 U15024 ( .A1(n17219), .A2(n13399), .ZN(n17197) );
  NAND2_X1 U15025 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13407) );
  NAND2_X1 U15026 ( .A1(n13399), .A2(n13407), .ZN(n13400) );
  INV_X1 U15027 ( .A(n13735), .ZN(n13401) );
  NAND2_X1 U15028 ( .A1(n17189), .A2(n13401), .ZN(n13641) );
  INV_X1 U15029 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13736) );
  INV_X1 U15030 ( .A(n17189), .ZN(n17176) );
  OAI22_X1 U15031 ( .A1(n13641), .A2(n13736), .B1(n17365), .B2(n17176), .ZN(
        n13733) );
  OR2_X1 U15032 ( .A1(n13733), .A2(n13736), .ZN(n13402) );
  INV_X1 U15033 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13404) );
  INV_X1 U15034 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17348) );
  INV_X1 U15035 ( .A(n17319), .ZN(n17268) );
  AOI21_X1 U15036 ( .B1(n17268), .B2(n15470), .A(n15469), .ZN(n15515) );
  NOR2_X1 U15037 ( .A1(n15515), .A2(n13403), .ZN(n17402) );
  NAND2_X1 U15038 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17402), .ZN(
        n19140) );
  NAND2_X1 U15039 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19141) );
  NAND2_X1 U15040 ( .A1(n17334), .A2(n17367), .ZN(n17349) );
  NOR3_X1 U15041 ( .A1(n13404), .A2(n17348), .A3(n17349), .ZN(n19087) );
  NAND2_X1 U15042 ( .A1(n19087), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n19112) );
  NOR2_X1 U15043 ( .A1(n19112), .A2(n13405), .ZN(n17251) );
  NAND2_X1 U15044 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17251), .ZN(
        n17245) );
  NOR2_X1 U15045 ( .A1(n13406), .A2(n17245), .ZN(n17220) );
  NAND2_X1 U15046 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17220), .ZN(
        n17210) );
  INV_X1 U15047 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14240) );
  MUX2_X1 U15048 ( .A(n13408), .B(n14240), .S(n13479), .Z(n13425) );
  NOR2_X1 U15049 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n13409) );
  MUX2_X1 U15050 ( .A(n13410), .B(n13409), .S(n13479), .Z(n13435) );
  INV_X1 U15051 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13416) );
  INV_X1 U15052 ( .A(n13411), .ZN(n13414) );
  NAND2_X1 U15053 ( .A1(n15234), .A2(n13412), .ZN(n13413) );
  NAND2_X1 U15054 ( .A1(n13414), .A2(n13413), .ZN(n13415) );
  MUX2_X1 U15055 ( .A(n13416), .B(n13415), .S(n13448), .Z(n13434) );
  NAND2_X1 U15056 ( .A1(n13435), .A2(n13434), .ZN(n13437) );
  MUX2_X1 U15057 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n13418), .S(n13448), .Z(
        n13419) );
  INV_X1 U15058 ( .A(n13451), .ZN(n13421) );
  NAND2_X1 U15059 ( .A1(n13423), .A2(n13419), .ZN(n13420) );
  NAND2_X1 U15060 ( .A1(n13421), .A2(n13420), .ZN(n15247) );
  NAND2_X1 U15061 ( .A1(n13422), .A2(n15247), .ZN(n13445) );
  XNOR2_X1 U15062 ( .A(n13445), .B(n15685), .ZN(n15682) );
  OAI21_X1 U15063 ( .B1(n13425), .B2(n13424), .A(n13423), .ZN(n18734) );
  NAND2_X1 U15064 ( .A1(n15466), .A2(n13507), .ZN(n13427) );
  XNOR2_X1 U15065 ( .A(n13437), .B(n13426), .ZN(n15256) );
  NAND2_X1 U15066 ( .A1(n13427), .A2(n15256), .ZN(n15503) );
  MUX2_X1 U15067 ( .A(n13429), .B(n13428), .S(n15234), .Z(n13430) );
  MUX2_X1 U15068 ( .A(n13430), .B(P2_EBX_REG_0__SCAN_IN), .S(n13479), .Z(
        n15370) );
  INV_X1 U15069 ( .A(n15370), .ZN(n13431) );
  NOR2_X1 U15070 ( .A1(n13431), .A2(n19073), .ZN(n13433) );
  INV_X1 U15071 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14107) );
  INV_X1 U15072 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15574) );
  NOR3_X1 U15073 ( .A1(n13448), .A2(n14107), .A3(n15574), .ZN(n13432) );
  NOR2_X1 U15074 ( .A1(n13435), .A2(n13432), .ZN(n15578) );
  NOR2_X1 U15075 ( .A1(n13433), .A2(n15578), .ZN(n13791) );
  AND2_X1 U15076 ( .A1(n13433), .A2(n15578), .ZN(n13790) );
  NOR2_X1 U15077 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13790), .ZN(
        n13789) );
  NOR2_X1 U15078 ( .A1(n13791), .A2(n13789), .ZN(n13869) );
  OR2_X1 U15079 ( .A1(n13435), .A2(n13434), .ZN(n13436) );
  NAND2_X1 U15080 ( .A1(n13437), .A2(n13436), .ZN(n15314) );
  XNOR2_X1 U15081 ( .A(n15314), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13868) );
  NOR2_X1 U15082 ( .A1(n15314), .A2(n12865), .ZN(n13438) );
  AOI21_X1 U15083 ( .B1(n13869), .B2(n13868), .A(n13438), .ZN(n13441) );
  NAND2_X1 U15084 ( .A1(n18734), .A2(n15686), .ZN(n13442) );
  INV_X1 U15085 ( .A(n13442), .ZN(n13439) );
  AOI21_X1 U15086 ( .B1(n13441), .B2(n15516), .A(n13439), .ZN(n13440) );
  NAND2_X1 U15087 ( .A1(n15503), .A2(n13440), .ZN(n13444) );
  INV_X1 U15088 ( .A(n13441), .ZN(n15504) );
  NAND3_X1 U15089 ( .A1(n15504), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n13442), .ZN(n13443) );
  OAI211_X1 U15090 ( .C1(n18734), .C2(n15686), .A(n13444), .B(n13443), .ZN(
        n15683) );
  NAND2_X1 U15091 ( .A1(n15682), .A2(n15683), .ZN(n13447) );
  NAND2_X1 U15092 ( .A1(n13445), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13446) );
  NAND2_X1 U15093 ( .A1(n13447), .A2(n13446), .ZN(n17164) );
  INV_X1 U15094 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18744) );
  MUX2_X1 U15095 ( .A(n18744), .B(n13449), .S(n13448), .Z(n13450) );
  OAI21_X1 U15096 ( .B1(n13451), .B2(n13450), .A(n13460), .ZN(n18745) );
  OAI21_X2 U15097 ( .B1(n13452), .B2(n13455), .A(n18745), .ZN(n13453) );
  XNOR2_X1 U15098 ( .A(n13453), .B(n17401), .ZN(n17165) );
  NAND2_X1 U15099 ( .A1(n13453), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13454) );
  MUX2_X1 U15100 ( .A(n13507), .B(P2_EBX_REG_7__SCAN_IN), .S(n13479), .Z(
        n13459) );
  INV_X1 U15101 ( .A(n13459), .ZN(n13456) );
  XNOR2_X1 U15102 ( .A(n13460), .B(n13456), .ZN(n18758) );
  AND2_X1 U15103 ( .A1(n18758), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17155) );
  INV_X1 U15104 ( .A(n18758), .ZN(n13458) );
  INV_X1 U15105 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13457) );
  NAND2_X1 U15106 ( .A1(n13458), .A2(n13457), .ZN(n13463) );
  NAND2_X1 U15107 ( .A1(n13479), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13461) );
  NOR2_X1 U15108 ( .A1(n11253), .A2(n13461), .ZN(n13462) );
  OR2_X1 U15109 ( .A1(n13746), .A2(n13462), .ZN(n18766) );
  NOR2_X1 U15110 ( .A1(n18766), .A2(n13507), .ZN(n13464) );
  NAND2_X1 U15111 ( .A1(n13464), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17570) );
  INV_X1 U15112 ( .A(n13463), .ZN(n17156) );
  INV_X1 U15113 ( .A(n13464), .ZN(n13466) );
  NAND2_X1 U15114 ( .A1(n13479), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13470) );
  INV_X1 U15115 ( .A(n13470), .ZN(n13468) );
  XNOR2_X1 U15116 ( .A(n13746), .B(n13468), .ZN(n18781) );
  NAND2_X1 U15117 ( .A1(n18781), .A2(n13749), .ZN(n13469) );
  INV_X1 U15118 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17366) );
  NAND2_X1 U15119 ( .A1(n13469), .A2(n17366), .ZN(n17144) );
  INV_X1 U15120 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n15269) );
  NOR2_X1 U15121 ( .A1(n13448), .A2(n15269), .ZN(n13471) );
  NAND2_X1 U15122 ( .A1(n13472), .A2(n13471), .ZN(n13473) );
  NAND2_X1 U15123 ( .A1(n13513), .A2(n13473), .ZN(n18789) );
  INV_X1 U15124 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U15125 ( .A1(n13540), .A2(n13474), .ZN(n17585) );
  INV_X1 U15126 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13475) );
  NOR2_X2 U15127 ( .A1(n13513), .A2(n13511), .ZN(n13501) );
  NAND2_X1 U15128 ( .A1(n13479), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13499) );
  AND2_X2 U15129 ( .A1(n13501), .A2(n13499), .ZN(n13504) );
  NAND2_X1 U15130 ( .A1(n13479), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13503) );
  INV_X1 U15131 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13476) );
  NOR2_X1 U15132 ( .A1(n13448), .A2(n13476), .ZN(n13494) );
  INV_X1 U15133 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13477) );
  NOR2_X1 U15134 ( .A1(n13448), .A2(n13477), .ZN(n13490) );
  INV_X1 U15135 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13478) );
  NOR2_X1 U15136 ( .A1(n13448), .A2(n13478), .ZN(n13484) );
  NAND2_X1 U15137 ( .A1(n13479), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13515) );
  INV_X1 U15138 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15856) );
  NOR2_X1 U15139 ( .A1(n13448), .A2(n15856), .ZN(n13519) );
  INV_X1 U15140 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n15897) );
  NOR2_X1 U15141 ( .A1(n13448), .A2(n15897), .ZN(n13527) );
  NOR2_X2 U15142 ( .A1(n13529), .A2(n13527), .ZN(n13481) );
  NAND2_X1 U15143 ( .A1(n13479), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13480) );
  AND2_X2 U15144 ( .A1(n13481), .A2(n13480), .ZN(n13525) );
  NOR2_X1 U15145 ( .A1(n13481), .A2(n13480), .ZN(n13482) );
  OR2_X1 U15146 ( .A1(n13525), .A2(n13482), .ZN(n18907) );
  INV_X1 U15147 ( .A(n18907), .ZN(n13483) );
  NAND2_X1 U15148 ( .A1(n13483), .A2(n13749), .ZN(n13618) );
  INV_X1 U15149 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17274) );
  AND2_X1 U15150 ( .A1(n13492), .A2(n13484), .ZN(n13485) );
  OR2_X1 U15151 ( .A1(n13485), .A2(n13516), .ZN(n18856) );
  NOR2_X1 U15152 ( .A1(n18856), .A2(n13507), .ZN(n13486) );
  NAND2_X1 U15153 ( .A1(n13486), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13613) );
  INV_X1 U15154 ( .A(n13486), .ZN(n13488) );
  INV_X1 U15155 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13487) );
  NAND2_X1 U15156 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  AND2_X1 U15157 ( .A1(n13613), .A2(n13489), .ZN(n17628) );
  NAND2_X1 U15158 ( .A1(n13496), .A2(n13490), .ZN(n13491) );
  NAND2_X1 U15159 ( .A1(n13492), .A2(n13491), .ZN(n18841) );
  INV_X1 U15160 ( .A(n18841), .ZN(n13493) );
  NAND2_X1 U15161 ( .A1(n13493), .A2(n13749), .ZN(n17137) );
  INV_X1 U15162 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17316) );
  NAND2_X1 U15163 ( .A1(n17137), .A2(n17316), .ZN(n13510) );
  NAND2_X1 U15164 ( .A1(n13506), .A2(n13494), .ZN(n13495) );
  NAND2_X1 U15165 ( .A1(n13496), .A2(n13495), .ZN(n18825) );
  OR2_X1 U15166 ( .A1(n18825), .A2(n13507), .ZN(n13498) );
  INV_X1 U15167 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13497) );
  NAND2_X1 U15168 ( .A1(n13498), .A2(n13497), .ZN(n17136) );
  INV_X1 U15169 ( .A(n13499), .ZN(n13500) );
  XNOR2_X1 U15170 ( .A(n13501), .B(n13500), .ZN(n18812) );
  NAND2_X1 U15171 ( .A1(n18812), .A2(n13749), .ZN(n13502) );
  NAND2_X1 U15172 ( .A1(n13502), .A2(n17348), .ZN(n17343) );
  OR2_X1 U15173 ( .A1(n13504), .A2(n13503), .ZN(n13505) );
  NAND2_X1 U15174 ( .A1(n13506), .A2(n13505), .ZN(n15565) );
  OR2_X1 U15175 ( .A1(n15565), .A2(n13507), .ZN(n13508) );
  NAND2_X1 U15176 ( .A1(n13508), .A2(n13404), .ZN(n17134) );
  AND3_X1 U15177 ( .A1(n17136), .A2(n17343), .A3(n17134), .ZN(n13509) );
  INV_X1 U15178 ( .A(n13511), .ZN(n13512) );
  XNOR2_X1 U15179 ( .A(n13513), .B(n13512), .ZN(n18803) );
  NAND2_X1 U15180 ( .A1(n18803), .A2(n13749), .ZN(n13514) );
  NAND2_X1 U15181 ( .A1(n13514), .A2(n17368), .ZN(n13607) );
  OR2_X1 U15182 ( .A1(n13516), .A2(n13515), .ZN(n13517) );
  NAND2_X1 U15183 ( .A1(n13521), .A2(n13517), .ZN(n18868) );
  INV_X1 U15184 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13625) );
  OAI21_X1 U15185 ( .B1(n18868), .B2(n13507), .A(n13625), .ZN(n17642) );
  NAND4_X1 U15186 ( .A1(n17628), .A2(n17629), .A3(n13607), .A4(n17642), .ZN(
        n13518) );
  AOI21_X1 U15187 ( .B1(n13618), .B2(n17274), .A(n13518), .ZN(n13531) );
  INV_X1 U15188 ( .A(n13519), .ZN(n13520) );
  XNOR2_X1 U15189 ( .A(n13521), .B(n13520), .ZN(n18881) );
  NAND2_X1 U15190 ( .A1(n18881), .A2(n13749), .ZN(n13523) );
  NAND2_X1 U15191 ( .A1(n13523), .A2(n13522), .ZN(n17302) );
  NAND2_X1 U15192 ( .A1(n13479), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n13524) );
  OR2_X1 U15193 ( .A1(n13525), .A2(n13524), .ZN(n13526) );
  NAND2_X1 U15194 ( .A1(n13563), .A2(n13526), .ZN(n18920) );
  OAI21_X1 U15195 ( .B1(n18920), .B2(n13507), .A(n17258), .ZN(n17109) );
  INV_X1 U15196 ( .A(n13527), .ZN(n13528) );
  XNOR2_X1 U15197 ( .A(n13529), .B(n13528), .ZN(n18891) );
  NAND2_X1 U15198 ( .A1(n18891), .A2(n13749), .ZN(n13530) );
  INV_X1 U15199 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17293) );
  NAND2_X1 U15200 ( .A1(n13530), .A2(n17293), .ZN(n17123) );
  AND4_X1 U15201 ( .A1(n13531), .A2(n17302), .A3(n17109), .A4(n17123), .ZN(
        n13532) );
  INV_X1 U15202 ( .A(n13618), .ZN(n13533) );
  NAND2_X1 U15203 ( .A1(n13533), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13553) );
  AND2_X1 U15204 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13534) );
  NAND2_X1 U15205 ( .A1(n18881), .A2(n13534), .ZN(n17301) );
  INV_X1 U15206 ( .A(n17137), .ZN(n13535) );
  NAND2_X1 U15207 ( .A1(n13535), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13539) );
  NAND2_X1 U15208 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13536) );
  OR2_X1 U15209 ( .A1(n18825), .A2(n13536), .ZN(n17135) );
  NAND2_X1 U15210 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13537) );
  OR2_X1 U15211 ( .A1(n15565), .A2(n13537), .ZN(n17133) );
  AND2_X1 U15212 ( .A1(n17135), .A2(n17133), .ZN(n13538) );
  NAND2_X1 U15213 ( .A1(n13539), .A2(n13538), .ZN(n13610) );
  INV_X1 U15214 ( .A(n13540), .ZN(n13541) );
  NAND2_X1 U15215 ( .A1(n13541), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17586) );
  AND2_X1 U15216 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13542) );
  NAND2_X1 U15217 ( .A1(n18781), .A2(n13542), .ZN(n17582) );
  NAND2_X1 U15218 ( .A1(n17586), .A2(n17582), .ZN(n17359) );
  AND2_X1 U15219 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13543) );
  AND2_X1 U15220 ( .A1(n18803), .A2(n13543), .ZN(n17357) );
  NOR2_X1 U15221 ( .A1(n17359), .A2(n17357), .ZN(n13608) );
  INV_X1 U15222 ( .A(n18812), .ZN(n13544) );
  NAND2_X1 U15223 ( .A1(n13608), .A2(n17342), .ZN(n13545) );
  NOR2_X1 U15224 ( .A1(n13610), .A2(n13545), .ZN(n13548) );
  INV_X1 U15225 ( .A(n18868), .ZN(n13547) );
  AND2_X1 U15226 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13546) );
  NAND2_X1 U15227 ( .A1(n13547), .A2(n13546), .ZN(n17641) );
  AND4_X1 U15228 ( .A1(n17301), .A2(n13548), .A3(n13613), .A4(n17641), .ZN(
        n13552) );
  INV_X1 U15229 ( .A(n18920), .ZN(n13550) );
  AND2_X1 U15230 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13549) );
  NAND2_X1 U15231 ( .A1(n13550), .A2(n13549), .ZN(n17108) );
  AND2_X1 U15232 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13551) );
  NAND2_X1 U15233 ( .A1(n18891), .A2(n13551), .ZN(n17122) );
  NAND2_X1 U15234 ( .A1(n13554), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13557) );
  INV_X1 U15235 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n13555) );
  NOR2_X1 U15236 ( .A1(n13448), .A2(n13555), .ZN(n13562) );
  INV_X1 U15237 ( .A(n13562), .ZN(n13556) );
  XNOR2_X1 U15238 ( .A(n13563), .B(n13556), .ZN(n18931) );
  NAND2_X1 U15239 ( .A1(n18931), .A2(n13749), .ZN(n17241) );
  NAND2_X1 U15240 ( .A1(n13557), .A2(n17241), .ZN(n13561) );
  INV_X1 U15241 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17244) );
  NAND2_X1 U15242 ( .A1(n17240), .A2(n17244), .ZN(n13560) );
  NAND2_X1 U15243 ( .A1(n13479), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n13564) );
  OR2_X1 U15244 ( .A1(n11236), .A2(n13564), .ZN(n13565) );
  NAND2_X1 U15245 ( .A1(n13567), .A2(n13565), .ZN(n18942) );
  OR2_X1 U15246 ( .A1(n18942), .A2(n13507), .ZN(n13566) );
  INV_X1 U15247 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16932) );
  XNOR2_X1 U15248 ( .A(n13567), .B(n11287), .ZN(n18953) );
  NAND2_X1 U15249 ( .A1(n18953), .A2(n13749), .ZN(n17225) );
  INV_X1 U15250 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n13568) );
  NOR2_X1 U15251 ( .A1(n13448), .A2(n13568), .ZN(n13574) );
  INV_X1 U15252 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16915) );
  NOR2_X1 U15253 ( .A1(n13448), .A2(n16915), .ZN(n13578) );
  INV_X1 U15254 ( .A(n13578), .ZN(n13569) );
  XNOR2_X1 U15255 ( .A(n13579), .B(n13569), .ZN(n18974) );
  NAND2_X1 U15256 ( .A1(n18974), .A2(n13749), .ZN(n13571) );
  NAND2_X1 U15257 ( .A1(n13571), .A2(n13570), .ZN(n13573) );
  AND2_X1 U15258 ( .A1(n13749), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13572) );
  NAND2_X1 U15259 ( .A1(n18974), .A2(n13572), .ZN(n13592) );
  NAND2_X1 U15260 ( .A1(n13573), .A2(n13592), .ZN(n17078) );
  INV_X1 U15261 ( .A(n13574), .ZN(n13575) );
  XNOR2_X1 U15262 ( .A(n13576), .B(n13575), .ZN(n18962) );
  NAND2_X1 U15263 ( .A1(n18962), .A2(n13749), .ZN(n13591) );
  NAND2_X1 U15264 ( .A1(n13479), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13580) );
  OR2_X1 U15265 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  NAND2_X1 U15266 ( .A1(n13586), .A2(n13582), .ZN(n18985) );
  INV_X1 U15267 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n13584) );
  NOR2_X1 U15268 ( .A1(n13448), .A2(n13584), .ZN(n13585) );
  NAND2_X1 U15269 ( .A1(n13586), .A2(n13585), .ZN(n13587) );
  NAND2_X1 U15270 ( .A1(n13598), .A2(n13587), .ZN(n18996) );
  OAI21_X1 U15271 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n17053), .ZN(n13588) );
  INV_X1 U15272 ( .A(n17053), .ZN(n13589) );
  INV_X1 U15273 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17052) );
  NAND2_X1 U15274 ( .A1(n13589), .A2(n17052), .ZN(n13593) );
  NAND2_X1 U15275 ( .A1(n13592), .A2(n17087), .ZN(n17049) );
  INV_X1 U15276 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n13594) );
  XNOR2_X1 U15277 ( .A(n13598), .B(n11295), .ZN(n19010) );
  NAND2_X1 U15278 ( .A1(n19010), .A2(n13749), .ZN(n13596) );
  INV_X1 U15279 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13595) );
  AND2_X1 U15280 ( .A1(n13596), .A2(n13595), .ZN(n13653) );
  INV_X1 U15281 ( .A(n13596), .ZN(n13597) );
  NOR2_X1 U15282 ( .A1(n13744), .A2(n13739), .ZN(n13602) );
  INV_X1 U15283 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n19026) );
  NOR2_X1 U15284 ( .A1(n13448), .A2(n19026), .ZN(n13599) );
  XNOR2_X1 U15285 ( .A(n13745), .B(n13599), .ZN(n19024) );
  NOR3_X1 U15286 ( .A1(n19024), .A2(n13507), .A3(n13736), .ZN(n13738) );
  OAI21_X1 U15287 ( .B1(n19024), .B2(n13507), .A(n13736), .ZN(n13743) );
  INV_X1 U15288 ( .A(n13743), .ZN(n13600) );
  NOR2_X1 U15289 ( .A1(n13738), .A2(n13600), .ZN(n13601) );
  XNOR2_X1 U15290 ( .A(n13602), .B(n13601), .ZN(n17038) );
  NOR2_X1 U15291 ( .A1(n13604), .A2(n13603), .ZN(n14633) );
  OAI211_X1 U15292 ( .C1(n19134), .C2(n17040), .A(n11685), .B(n13606), .ZN(
        P2_U3016) );
  INV_X1 U15293 ( .A(n13607), .ZN(n17358) );
  INV_X1 U15294 ( .A(n17342), .ZN(n13609) );
  INV_X1 U15295 ( .A(n13610), .ZN(n13611) );
  NAND2_X1 U15296 ( .A1(n13614), .A2(n17641), .ZN(n13615) );
  AND2_X1 U15297 ( .A1(n17123), .A2(n17302), .ZN(n13616) );
  NAND2_X1 U15298 ( .A1(n13617), .A2(n13616), .ZN(n13619) );
  NAND2_X1 U15299 ( .A1(n13619), .A2(n13618), .ZN(n13620) );
  NAND2_X1 U15300 ( .A1(n19156), .A2(n14633), .ZN(n13623) );
  NAND2_X1 U15301 ( .A1(n13623), .A2(n13622), .ZN(n14650) );
  NAND2_X1 U15302 ( .A1(n17645), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17300) );
  NAND2_X1 U15303 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n15636) );
  INV_X1 U15304 ( .A(n15636), .ZN(n13626) );
  NOR2_X1 U15305 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13626), .ZN(n17682) );
  NAND2_X1 U15306 ( .A1(n17682), .A2(n15635), .ZN(n13627) );
  NOR2_X1 U15307 ( .A1(n18813), .A2(n18905), .ZN(n17281) );
  AOI21_X1 U15308 ( .B1(n17670), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17281), .ZN(n13631) );
  INV_X1 U15309 ( .A(n14215), .ZN(n14661) );
  INV_X1 U15310 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22169) );
  NAND2_X1 U15311 ( .A1(n22169), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13628) );
  NAND2_X1 U15312 ( .A1(n14661), .A2(n13628), .ZN(n13954) );
  NAND2_X1 U15313 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n15229), .ZN(
        n15228) );
  NOR2_X2 U15314 ( .A1(n15228), .A2(n15510), .ZN(n15226) );
  INV_X1 U15315 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17130) );
  INV_X1 U15316 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18864) );
  INV_X1 U15317 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17120) );
  OAI21_X1 U15318 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11245), .A(
        n17114), .ZN(n18913) );
  INV_X1 U15319 ( .A(n18913), .ZN(n13629) );
  NAND2_X1 U15320 ( .A1(n17640), .A2(n13629), .ZN(n13630) );
  NAND2_X1 U15321 ( .A1(n13631), .A2(n13630), .ZN(n13636) );
  AND2_X1 U15322 ( .A1(n15901), .A2(n13632), .ZN(n13633) );
  OR2_X1 U15323 ( .A1(n13633), .A2(n16959), .ZN(n18916) );
  INV_X1 U15324 ( .A(n18916), .ZN(n13634) );
  AND2_X1 U15325 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17494) );
  AND2_X1 U15326 ( .A1(n13634), .A2(n17673), .ZN(n13635) );
  INV_X1 U15327 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17191) );
  AOI21_X1 U15328 ( .B1(n17072), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13639) );
  AOI22_X1 U15329 ( .A1(n13641), .A2(n13640), .B1(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n13735), .ZN(n13652) );
  NAND2_X1 U15330 ( .A1(n16901), .A2(n13642), .ZN(n13643) );
  NOR2_X1 U15331 ( .A1(n18892), .A2(n17743), .ZN(n17043) );
  NAND2_X1 U15332 ( .A1(n16975), .A2(n13645), .ZN(n13646) );
  OR2_X1 U15333 ( .A1(n16247), .A2(n19119), .ZN(n13648) );
  NAND2_X1 U15334 ( .A1(n17176), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13647) );
  OAI21_X1 U15335 ( .B1(n17184), .B2(n13652), .A(n13651), .ZN(n13656) );
  NOR2_X1 U15336 ( .A1(n13739), .A2(n13653), .ZN(n13654) );
  XNOR2_X1 U15337 ( .A(n13655), .B(n13654), .ZN(n17047) );
  NOR2_X1 U15338 ( .A1(n16743), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13659) );
  NAND2_X1 U15339 ( .A1(n13660), .A2(n16779), .ZN(n13661) );
  NOR2_X1 U15340 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16706) );
  XNOR2_X1 U15341 ( .A(n20516), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16562) );
  AND2_X1 U15342 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16705) );
  INV_X1 U15343 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16688) );
  XNOR2_X1 U15344 ( .A(n13662), .B(n16688), .ZN(n16694) );
  OR2_X2 U15345 ( .A1(n16694), .A2(n22141), .ZN(n13667) );
  NAND2_X1 U15346 ( .A1(n13668), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15286) );
  XNOR2_X1 U15347 ( .A(n15286), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16257) );
  INV_X1 U15348 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U15349 ( .A1(n21906), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16685) );
  OAI21_X1 U15350 ( .B1(n16670), .B2(n15285), .A(n16685), .ZN(n13665) );
  AOI21_X1 U15351 ( .B1(n16257), .B2(n20505), .A(n13665), .ZN(n13666) );
  INV_X1 U15352 ( .A(n13668), .ZN(n13669) );
  INV_X1 U15353 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16292) );
  NAND2_X1 U15354 ( .A1(n13669), .A2(n16292), .ZN(n13670) );
  NAND2_X1 U15355 ( .A1(n15286), .A2(n13670), .ZN(n16565) );
  NAND2_X1 U15356 ( .A1(n13672), .A2(n13671), .ZN(n13689) );
  AOI22_X1 U15357 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U15358 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11769), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13675) );
  AOI22_X1 U15359 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U15360 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11878), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13673) );
  NAND4_X1 U15361 ( .A1(n13676), .A2(n13675), .A3(n13674), .A4(n13673), .ZN(
        n13682) );
  AOI22_X1 U15362 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U15363 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U15364 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12030), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U15365 ( .A1(n12108), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13677) );
  NAND4_X1 U15366 ( .A1(n13680), .A2(n13679), .A3(n13678), .A4(n13677), .ZN(
        n13681) );
  NOR2_X1 U15367 ( .A1(n13682), .A2(n13681), .ZN(n13690) );
  XNOR2_X1 U15368 ( .A(n13689), .B(n13690), .ZN(n13686) );
  AOI21_X1 U15369 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n12293), .A(
        n13710), .ZN(n13684) );
  NAND2_X1 U15370 ( .A1(n16281), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13683) );
  OAI211_X1 U15371 ( .C1(n13686), .C2(n13685), .A(n13684), .B(n13683), .ZN(
        n13687) );
  OAI21_X1 U15372 ( .B1(n13688), .B2(n16565), .A(n13687), .ZN(n16291) );
  NOR2_X1 U15373 ( .A1(n13690), .A2(n13689), .ZN(n13706) );
  AOI22_X1 U15374 ( .A1(n11184), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U15375 ( .A1(n11182), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U15376 ( .A1(n11863), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11870), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U15377 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13694) );
  NAND4_X1 U15378 ( .A1(n13697), .A2(n13696), .A3(n13695), .A4(n13694), .ZN(
        n13704) );
  AOI22_X1 U15379 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U15380 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11183), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U15381 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12030), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U15382 ( .A1(n12338), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11983), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U15383 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13703) );
  NOR2_X1 U15384 ( .A1(n13704), .A2(n13703), .ZN(n13705) );
  XNOR2_X1 U15385 ( .A(n13706), .B(n13705), .ZN(n13708) );
  NAND2_X1 U15386 ( .A1(n13708), .A2(n13707), .ZN(n13713) );
  AOI21_X1 U15387 ( .B1(n15285), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13709) );
  AOI21_X1 U15388 ( .B1(n16281), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13709), .ZN(
        n13712) );
  AOI21_X1 U15389 ( .B1(n13713), .B2(n13712), .A(n13711), .ZN(n16279) );
  NAND2_X1 U15390 ( .A1(n13715), .A2(n13714), .ZN(P1_U2969) );
  XOR2_X1 U15391 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13717), .Z(
        n16240) );
  INV_X1 U15392 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19042) );
  AOI22_X1 U15393 ( .A1(n13720), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n13348), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13721) );
  OAI21_X1 U15394 ( .B1(n13722), .B2(n19042), .A(n13721), .ZN(n13723) );
  NAND2_X1 U15395 ( .A1(n13726), .A2(n13725), .ZN(n13732) );
  NAND2_X1 U15396 ( .A1(n11165), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13729) );
  AOI22_X1 U15397 ( .A1(n12856), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13728) );
  OAI211_X1 U15398 ( .C1(n13730), .C2(n19042), .A(n13729), .B(n13728), .ZN(
        n13731) );
  INV_X1 U15399 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15225) );
  NOR2_X1 U15400 ( .A1(n18892), .A2(n19042), .ZN(n16233) );
  AND2_X1 U15401 ( .A1(n11684), .A2(n13734), .ZN(n13737) );
  INV_X1 U15402 ( .A(n13739), .ZN(n13740) );
  AOI21_X1 U15403 ( .B1(n13744), .B2(n13743), .A(n13742), .ZN(n13752) );
  NOR2_X1 U15404 ( .A1(n13745), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13748) );
  INV_X1 U15405 ( .A(n13746), .ZN(n13747) );
  MUX2_X1 U15406 ( .A(n13748), .B(n13747), .S(n13448), .Z(n19035) );
  NAND2_X1 U15407 ( .A1(n19035), .A2(n13749), .ZN(n13750) );
  XNOR2_X1 U15408 ( .A(n13750), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13751) );
  XNOR2_X1 U15409 ( .A(n13752), .B(n13751), .ZN(n16238) );
  NAND2_X1 U15410 ( .A1(n16238), .A2(n19138), .ZN(n13753) );
  OAI211_X1 U15411 ( .C1(n16240), .C2(n19134), .A(n13754), .B(n13753), .ZN(
        P2_U3015) );
  NOR4_X1 U15412 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13758) );
  NOR4_X1 U15413 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13757) );
  NOR4_X1 U15414 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13756) );
  NOR4_X1 U15415 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13755) );
  AND4_X1 U15416 ( .A1(n13758), .A2(n13757), .A3(n13756), .A4(n13755), .ZN(
        n13763) );
  NOR4_X1 U15417 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13761) );
  NOR4_X1 U15418 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13760) );
  NOR4_X1 U15419 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13759) );
  INV_X1 U15420 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20386) );
  AND4_X1 U15421 ( .A1(n13761), .A2(n13760), .A3(n13759), .A4(n20386), .ZN(
        n13762) );
  NAND2_X1 U15422 ( .A1(n13763), .A2(n13762), .ZN(n13764) );
  AND2_X2 U15423 ( .A1(n13764), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n16270)
         );
  INV_X1 U15424 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22594) );
  INV_X1 U15425 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20599) );
  NOR4_X1 U15426 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n22594), .A4(n20599), .ZN(n13766) );
  NOR4_X1 U15427 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13765) );
  NAND3_X1 U15428 ( .A1(n16270), .A2(n13766), .A3(n13765), .ZN(U214) );
  NOR4_X1 U15429 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13770) );
  NOR4_X1 U15430 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13769) );
  NOR4_X1 U15431 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13768) );
  NOR4_X1 U15432 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13767) );
  NAND4_X1 U15433 ( .A1(n13770), .A2(n13769), .A3(n13768), .A4(n13767), .ZN(
        n13775) );
  NOR4_X1 U15434 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13773) );
  NOR4_X1 U15435 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13772) );
  NOR4_X1 U15436 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13771) );
  INV_X1 U15437 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20293) );
  NAND4_X1 U15438 ( .A1(n13773), .A2(n13772), .A3(n13771), .A4(n20293), .ZN(
        n13774) );
  NOR2_X1 U15439 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n13777) );
  NOR4_X1 U15440 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13776) );
  NAND4_X1 U15441 ( .A1(n13777), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n13776), .ZN(n13778) );
  OR2_X1 U15442 ( .A1(n13918), .A2(n13778), .ZN(n20531) );
  INV_X2 U15443 ( .A(U214), .ZN(n20584) );
  NOR2_X1 U15444 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13778), .ZN(n19529)
         );
  INV_X1 U15445 ( .A(n14605), .ZN(n15575) );
  OAI22_X1 U15446 ( .A1(n19133), .A2(n15575), .B1(n15227), .B2(n19074), .ZN(
        n13796) );
  INV_X1 U15447 ( .A(n13779), .ZN(n13781) );
  NAND2_X1 U15448 ( .A1(n13781), .A2(n13780), .ZN(n13782) );
  NAND2_X1 U15449 ( .A1(n13783), .A2(n13782), .ZN(n20111) );
  INV_X1 U15450 ( .A(n20111), .ZN(n15194) );
  OAI21_X1 U15451 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13785), .A(
        n13784), .ZN(n13970) );
  INV_X1 U15452 ( .A(n13970), .ZN(n13786) );
  NAND2_X1 U15453 ( .A1(n19108), .A2(n13786), .ZN(n13787) );
  OR2_X1 U15454 ( .A1(n18813), .A2(n17738), .ZN(n13968) );
  OAI211_X1 U15455 ( .C1(n15194), .C2(n19119), .A(n13787), .B(n13968), .ZN(
        n13795) );
  INV_X1 U15456 ( .A(n13791), .ZN(n13788) );
  AOI222_X1 U15457 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13791), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13790), .C1(n13789), .C2(
        n13788), .ZN(n13974) );
  NOR2_X1 U15458 ( .A1(n13974), .A2(n19091), .ZN(n13794) );
  OAI21_X1 U15459 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n14129), .ZN(n13792) );
  NOR2_X1 U15460 ( .A1(n19109), .A2(n13792), .ZN(n13793) );
  OR4_X1 U15461 ( .A1(n13796), .A2(n13795), .A3(n13794), .A4(n13793), .ZN(
        P2_U3045) );
  OR2_X1 U15462 ( .A1(n19062), .A2(n19171), .ZN(n13863) );
  OR2_X1 U15463 ( .A1(n14638), .A2(n13863), .ZN(n15581) );
  INV_X1 U15464 ( .A(n15581), .ZN(n18736) );
  INV_X1 U15465 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n17706) );
  OR2_X1 U15466 ( .A1(n13797), .A2(n19171), .ZN(n13798) );
  INV_X1 U15467 ( .A(n13859), .ZN(n13799) );
  OAI211_X1 U15468 ( .C1(n18736), .C2(n17706), .A(n13799), .B(n17559), .ZN(
        P2_U2814) );
  AND2_X1 U15469 ( .A1(n13823), .A2(n11829), .ZN(n13800) );
  AND2_X1 U15470 ( .A1(n13801), .A2(n13800), .ZN(n15087) );
  INV_X1 U15471 ( .A(n13802), .ZN(n13806) );
  AND2_X1 U15472 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  NAND2_X1 U15473 ( .A1(n13806), .A2(n13805), .ZN(n13807) );
  NAND2_X1 U15474 ( .A1(n15087), .A2(n15085), .ZN(n15097) );
  NOR2_X1 U15475 ( .A1(n15097), .A2(n22162), .ZN(n13812) );
  INV_X1 U15476 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22595) );
  AND2_X1 U15477 ( .A1(n13809), .A2(n14093), .ZN(n13810) );
  AND2_X1 U15478 ( .A1(n15381), .A2(n15288), .ZN(n15446) );
  INV_X1 U15479 ( .A(n15446), .ZN(n13811) );
  OAI211_X1 U15480 ( .C1(n13812), .C2(n22595), .A(n13976), .B(n13811), .ZN(
        P1_U2801) );
  OR2_X1 U15481 ( .A1(n14638), .A2(n14634), .ZN(n14649) );
  NOR2_X1 U15482 ( .A1(n18717), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13814)
         );
  AOI22_X1 U15483 ( .A1(n13814), .A2(n17559), .B1(n13813), .B2(n18717), .ZN(
        P2_U3612) );
  AND2_X1 U15484 ( .A1(n15087), .A2(n15294), .ZN(n16833) );
  NAND3_X1 U15485 ( .A1(n15095), .A2(n14093), .A3(n16833), .ZN(n14242) );
  INV_X1 U15486 ( .A(n13815), .ZN(n22145) );
  NAND3_X1 U15487 ( .A1(n22145), .A2(n14093), .A3(n15085), .ZN(n13816) );
  OAI21_X1 U15488 ( .B1(n15446), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n21838), 
        .ZN(n13817) );
  OAI21_X1 U15489 ( .B1(n13818), .B2(n21838), .A(n13817), .ZN(P1_U3487) );
  AOI21_X1 U15490 ( .B1(n14098), .B2(n15294), .A(n11829), .ZN(n13819) );
  NAND2_X1 U15491 ( .A1(n13820), .A2(n13819), .ZN(n13833) );
  NAND2_X1 U15492 ( .A1(n13821), .A2(n14245), .ZN(n13822) );
  OAI21_X1 U15493 ( .B1(n13823), .B2(n15283), .A(n13822), .ZN(n13824) );
  INV_X1 U15494 ( .A(n13824), .ZN(n13827) );
  OR2_X1 U15495 ( .A1(n13825), .A2(n14558), .ZN(n13826) );
  AND3_X1 U15496 ( .A1(n13833), .A2(n13827), .A3(n13826), .ZN(n14061) );
  NAND4_X1 U15497 ( .A1(n14061), .A2(n11832), .A3(n13815), .A4(n13828), .ZN(
        n13932) );
  INV_X1 U15498 ( .A(n13932), .ZN(n16829) );
  OAI22_X1 U15499 ( .A1(n14523), .A2(n16829), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14043), .ZN(n17514) );
  INV_X1 U15500 ( .A(n22156), .ZN(n16849) );
  OAI22_X1 U15501 ( .A1(n16849), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15288), .ZN(n13830) );
  AOI21_X1 U15502 ( .B1(n17514), .B2(n22146), .A(n13830), .ZN(n13856) );
  NAND2_X1 U15503 ( .A1(n13831), .A2(n20527), .ZN(n22189) );
  NAND2_X1 U15504 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21842) );
  INV_X1 U15505 ( .A(n21842), .ZN(n22181) );
  NOR2_X1 U15506 ( .A1(n22189), .A2(n22181), .ZN(n13832) );
  OAI211_X1 U15507 ( .C1(n16833), .C2(n17546), .A(n13832), .B(n15095), .ZN(
        n13841) );
  INV_X1 U15508 ( .A(n15087), .ZN(n13836) );
  NAND2_X1 U15509 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  NAND2_X1 U15510 ( .A1(n13836), .A2(n13835), .ZN(n14045) );
  NOR2_X1 U15511 ( .A1(n15079), .A2(n11828), .ZN(n13837) );
  INV_X1 U15512 ( .A(n14043), .ZN(n16831) );
  INV_X1 U15513 ( .A(n15088), .ZN(n13934) );
  OR2_X1 U15514 ( .A1(n15095), .A2(n13934), .ZN(n13840) );
  OR2_X1 U15515 ( .A1(n15283), .A2(n13838), .ZN(n13839) );
  AND4_X1 U15516 ( .A1(n13841), .A2(n14045), .A3(n13840), .A4(n13839), .ZN(
        n13848) );
  NAND2_X1 U15517 ( .A1(n17546), .A2(n21842), .ZN(n14039) );
  INV_X1 U15518 ( .A(n13842), .ZN(n13843) );
  NAND2_X1 U15519 ( .A1(n13843), .A2(n15094), .ZN(n14049) );
  OAI21_X1 U15520 ( .B1(n14039), .B2(n16209), .A(n14049), .ZN(n13844) );
  NAND2_X1 U15521 ( .A1(n15095), .A2(n13844), .ZN(n13846) );
  NAND3_X1 U15522 ( .A1(n22145), .A2(n15085), .A3(n21842), .ZN(n13845) );
  NAND2_X1 U15523 ( .A1(n13846), .A2(n13845), .ZN(n14094) );
  INV_X1 U15524 ( .A(n14094), .ZN(n13847) );
  NAND2_X1 U15525 ( .A1(n13848), .A2(n13847), .ZN(n17515) );
  NAND2_X1 U15526 ( .A1(n17515), .A2(n14093), .ZN(n13852) );
  INV_X1 U15527 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22142) );
  NAND2_X1 U15528 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22152) );
  NOR3_X1 U15529 ( .A1(n22142), .A2(n22153), .A3(n22152), .ZN(n13850) );
  NOR2_X1 U15530 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22280), .ZN(n13849) );
  NOR2_X1 U15531 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  NAND2_X1 U15532 ( .A1(n13852), .A2(n13851), .ZN(n22149) );
  INV_X1 U15533 ( .A(n22149), .ZN(n13855) );
  NAND2_X1 U15534 ( .A1(n16833), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17512) );
  INV_X1 U15535 ( .A(n17512), .ZN(n13853) );
  AOI22_X1 U15536 ( .A1(n13855), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n22146), .B2(n13853), .ZN(n13854) );
  OAI21_X1 U15537 ( .B1(n13856), .B2(n13855), .A(n13854), .ZN(P1_U3474) );
  AND2_X1 U15538 ( .A1(n13859), .A2(n19164), .ZN(n13860) );
  INV_X1 U15539 ( .A(n13860), .ZN(n13857) );
  INV_X1 U15540 ( .A(n13858), .ZN(n13862) );
  AOI22_X1 U15541 ( .A1(n15753), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15750), .ZN(n19634) );
  NAND2_X1 U15542 ( .A1(n13859), .A2(n16097), .ZN(n13883) );
  INV_X2 U15543 ( .A(n13883), .ZN(n13927) );
  INV_X1 U15544 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13861) );
  INV_X1 U15545 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19635) );
  OAI222_X1 U15546 ( .A1(n13862), .A2(n19634), .B1(n13880), .B2(n13861), .C1(
        n13883), .C2(n19635), .ZN(P2_U2982) );
  INV_X1 U15547 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n16146) );
  OAI21_X1 U15548 ( .B1(n14304), .B2(n13863), .A(n13883), .ZN(n13864) );
  NAND2_X1 U15549 ( .A1(n17709), .A2(n13865), .ZN(n14125) );
  NOR2_X1 U15550 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15636), .ZN(n17725) );
  AOI22_X1 U15551 ( .A1(n17725), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13866) );
  OAI21_X1 U15552 ( .B1(n16146), .B2(n14125), .A(n13866), .ZN(P2_U2921) );
  INV_X1 U15553 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15798) );
  AOI22_X1 U15554 ( .A1(n17725), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13867) );
  OAI21_X1 U15555 ( .B1(n15798), .B2(n14125), .A(n13867), .ZN(P2_U2934) );
  XNOR2_X1 U15556 ( .A(n13869), .B(n13868), .ZN(n14141) );
  OAI21_X1 U15557 ( .B1(n13872), .B2(n13871), .A(n13870), .ZN(n14132) );
  NOR2_X1 U15558 ( .A1(n18892), .A2(n12868), .ZN(n14138) );
  AOI21_X1 U15559 ( .B1(n17670), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14138), .ZN(n13874) );
  AOI21_X1 U15560 ( .B1(n13967), .B2(n15315), .A(n15229), .ZN(n15312) );
  NAND2_X1 U15561 ( .A1(n17640), .A2(n15312), .ZN(n13873) );
  OAI211_X1 U15562 ( .C1(n14132), .C2(n17676), .A(n13874), .B(n13873), .ZN(
        n13875) );
  AOI21_X1 U15563 ( .B1(n17673), .B2(n15322), .A(n13875), .ZN(n13876) );
  OAI21_X1 U15564 ( .B1(n17608), .B2(n14141), .A(n13876), .ZN(P2_U3012) );
  INV_X1 U15565 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17729) );
  INV_X2 U15566 ( .A(n13880), .ZN(n13924) );
  NAND2_X1 U15567 ( .A1(n13924), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U15568 ( .A1(n15750), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13878) );
  INV_X1 U15569 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20557) );
  OR2_X1 U15570 ( .A1(n15750), .A2(n20557), .ZN(n13877) );
  NAND2_X1 U15571 ( .A1(n13878), .A2(n13877), .ZN(n19644) );
  NAND2_X1 U15572 ( .A1(n13858), .A2(n19644), .ZN(n13881) );
  OAI211_X1 U15573 ( .C1(n17729), .C2(n13883), .A(n13879), .B(n13881), .ZN(
        P2_U2979) );
  INV_X1 U15574 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14112) );
  NAND2_X1 U15575 ( .A1(n13924), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13882) );
  OAI211_X1 U15576 ( .C1(n14112), .C2(n13883), .A(n13882), .B(n13881), .ZN(
        P2_U2964) );
  AOI22_X1 U15577 ( .A1(n13924), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U15578 ( .A1(n15753), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13918), .ZN(n20016) );
  INV_X1 U15579 ( .A(n20016), .ZN(n15894) );
  NAND2_X1 U15580 ( .A1(n13858), .A2(n15894), .ZN(n13913) );
  NAND2_X1 U15581 ( .A1(n13884), .A2(n13913), .ZN(P2_U2955) );
  AOI22_X1 U15582 ( .A1(n13924), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n13927), .ZN(n13886) );
  AOI22_X1 U15583 ( .A1(n15753), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13918), .ZN(n20175) );
  INV_X1 U15584 ( .A(n20175), .ZN(n13885) );
  NAND2_X1 U15585 ( .A1(n13858), .A2(n13885), .ZN(n13892) );
  NAND2_X1 U15586 ( .A1(n13886), .A2(n13892), .ZN(P2_U2952) );
  AOI22_X1 U15587 ( .A1(n13924), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13927), .ZN(n13887) );
  AOI22_X1 U15588 ( .A1(n15753), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n15750), .ZN(n19647) );
  INV_X1 U15589 ( .A(n19647), .ZN(n16986) );
  NAND2_X1 U15590 ( .A1(n13858), .A2(n16986), .ZN(n13907) );
  NAND2_X1 U15591 ( .A1(n13887), .A2(n13907), .ZN(P2_U2963) );
  AOI22_X1 U15592 ( .A1(n13924), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n13927), .ZN(n13889) );
  INV_X1 U15593 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20561) );
  NOR2_X1 U15594 ( .A1(n15750), .A2(n20561), .ZN(n13888) );
  AOI21_X1 U15595 ( .B1(n15750), .B2(BUF2_REG_14__SCAN_IN), .A(n13888), .ZN(
        n19637) );
  INV_X1 U15596 ( .A(n19637), .ZN(n16148) );
  NAND2_X1 U15597 ( .A1(n13858), .A2(n16148), .ZN(n13925) );
  NAND2_X1 U15598 ( .A1(n13889), .A2(n13925), .ZN(P2_U2966) );
  AOI22_X1 U15599 ( .A1(n13924), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13927), .ZN(n13890) );
  AOI22_X1 U15600 ( .A1(n15753), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13918), .ZN(n20068) );
  INV_X1 U15601 ( .A(n20068), .ZN(n15821) );
  NAND2_X1 U15602 ( .A1(n13858), .A2(n15821), .ZN(n13930) );
  NAND2_X1 U15603 ( .A1(n13890), .A2(n13930), .ZN(P2_U2954) );
  AOI22_X1 U15604 ( .A1(n13924), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n13927), .ZN(n13891) );
  INV_X1 U15605 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20541) );
  INV_X1 U15606 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19367) );
  AOI22_X1 U15607 ( .A1(n15753), .A2(n20541), .B1(n19367), .B2(n13918), .ZN(
        n19965) );
  NAND2_X1 U15608 ( .A1(n13858), .A2(n19965), .ZN(n13902) );
  NAND2_X1 U15609 ( .A1(n13891), .A2(n13902), .ZN(P2_U2971) );
  AOI22_X1 U15610 ( .A1(n13924), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n13927), .ZN(n13893) );
  NAND2_X1 U15611 ( .A1(n13893), .A2(n13892), .ZN(P2_U2967) );
  AOI22_X1 U15612 ( .A1(n13924), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U15613 ( .A1(n15753), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13918), .ZN(n19661) );
  INV_X1 U15614 ( .A(n19661), .ZN(n17021) );
  NAND2_X1 U15615 ( .A1(n13858), .A2(n17021), .ZN(n13900) );
  NAND2_X1 U15616 ( .A1(n13894), .A2(n13900), .ZN(P2_U2959) );
  AOI22_X1 U15617 ( .A1(n13924), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n13927), .ZN(n13896) );
  INV_X1 U15618 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20553) );
  NOR2_X1 U15619 ( .A1(n15750), .A2(n20553), .ZN(n13895) );
  AOI21_X1 U15620 ( .B1(n15750), .B2(BUF2_REG_10__SCAN_IN), .A(n13895), .ZN(
        n19651) );
  INV_X1 U15621 ( .A(n19651), .ZN(n16995) );
  NAND2_X1 U15622 ( .A1(n13858), .A2(n16995), .ZN(n13905) );
  NAND2_X1 U15623 ( .A1(n13896), .A2(n13905), .ZN(P2_U2962) );
  AOI22_X1 U15624 ( .A1(n13924), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U15625 ( .A1(n15753), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13918), .ZN(n20119) );
  INV_X1 U15626 ( .A(n20119), .ZN(n15801) );
  NAND2_X1 U15627 ( .A1(n13858), .A2(n15801), .ZN(n13909) );
  NAND2_X1 U15628 ( .A1(n13897), .A2(n13909), .ZN(P2_U2953) );
  AOI22_X1 U15629 ( .A1(n13924), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U15630 ( .A1(n15753), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n15750), .ZN(n19654) );
  INV_X1 U15631 ( .A(n19654), .ZN(n17004) );
  NAND2_X1 U15632 ( .A1(n13858), .A2(n17004), .ZN(n13928) );
  NAND2_X1 U15633 ( .A1(n13898), .A2(n13928), .ZN(P2_U2961) );
  AOI22_X1 U15634 ( .A1(n13924), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13899) );
  INV_X1 U15635 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20545) );
  INV_X1 U15636 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21136) );
  AOI22_X1 U15637 ( .A1(n15753), .A2(n20545), .B1(n21136), .B2(n13918), .ZN(
        n19854) );
  NAND2_X1 U15638 ( .A1(n13858), .A2(n19854), .ZN(n13911) );
  NAND2_X1 U15639 ( .A1(n13899), .A2(n13911), .ZN(P2_U2973) );
  AOI22_X1 U15640 ( .A1(n13924), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13901) );
  NAND2_X1 U15641 ( .A1(n13901), .A2(n13900), .ZN(P2_U2974) );
  AOI22_X1 U15642 ( .A1(n13924), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13927), .ZN(n13903) );
  NAND2_X1 U15643 ( .A1(n13903), .A2(n13902), .ZN(P2_U2956) );
  AOI22_X1 U15644 ( .A1(n13924), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13927), .ZN(n13904) );
  AOI22_X1 U15645 ( .A1(n15753), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n15750), .ZN(n19640) );
  INV_X1 U15646 ( .A(n19640), .ZN(n16249) );
  NAND2_X1 U15647 ( .A1(n13858), .A2(n16249), .ZN(n13915) );
  NAND2_X1 U15648 ( .A1(n13904), .A2(n13915), .ZN(P2_U2965) );
  AOI22_X1 U15649 ( .A1(n13924), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n13927), .ZN(n13906) );
  NAND2_X1 U15650 ( .A1(n13906), .A2(n13905), .ZN(P2_U2977) );
  AOI22_X1 U15651 ( .A1(n13924), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13908) );
  NAND2_X1 U15652 ( .A1(n13908), .A2(n13907), .ZN(P2_U2978) );
  AOI22_X1 U15653 ( .A1(n13924), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13910) );
  NAND2_X1 U15654 ( .A1(n13910), .A2(n13909), .ZN(P2_U2968) );
  AOI22_X1 U15655 ( .A1(n13924), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13927), .ZN(n13912) );
  NAND2_X1 U15656 ( .A1(n13912), .A2(n13911), .ZN(P2_U2958) );
  AOI22_X1 U15657 ( .A1(n13924), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n13927), .ZN(n13914) );
  NAND2_X1 U15658 ( .A1(n13914), .A2(n13913), .ZN(P2_U2970) );
  AOI22_X1 U15659 ( .A1(n13924), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13916) );
  NAND2_X1 U15660 ( .A1(n13916), .A2(n13915), .ZN(P2_U2980) );
  AOI22_X1 U15661 ( .A1(n13924), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n13927), .ZN(n13917) );
  AOI22_X1 U15662 ( .A1(n15753), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15750), .ZN(n19658) );
  INV_X1 U15663 ( .A(n19658), .ZN(n17012) );
  NAND2_X1 U15664 ( .A1(n13858), .A2(n17012), .ZN(n13920) );
  NAND2_X1 U15665 ( .A1(n13917), .A2(n13920), .ZN(P2_U2960) );
  AOI22_X1 U15666 ( .A1(n13924), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n13927), .ZN(n13919) );
  AOI22_X1 U15667 ( .A1(n15753), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13918), .ZN(n19911) );
  INV_X1 U15668 ( .A(n19911), .ZN(n17030) );
  NAND2_X1 U15669 ( .A1(n13858), .A2(n17030), .ZN(n13922) );
  NAND2_X1 U15670 ( .A1(n13919), .A2(n13922), .ZN(P2_U2972) );
  AOI22_X1 U15671 ( .A1(n13924), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n13927), .ZN(n13921) );
  NAND2_X1 U15672 ( .A1(n13921), .A2(n13920), .ZN(P2_U2975) );
  AOI22_X1 U15673 ( .A1(n13924), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13923) );
  NAND2_X1 U15674 ( .A1(n13923), .A2(n13922), .ZN(P2_U2957) );
  AOI22_X1 U15675 ( .A1(n13924), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n13927), .ZN(n13926) );
  NAND2_X1 U15676 ( .A1(n13926), .A2(n13925), .ZN(P2_U2981) );
  AOI22_X1 U15677 ( .A1(n13924), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13927), .ZN(n13929) );
  NAND2_X1 U15678 ( .A1(n13929), .A2(n13928), .ZN(P2_U2976) );
  AOI22_X1 U15679 ( .A1(n13924), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n13927), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13931) );
  NAND2_X1 U15680 ( .A1(n13931), .A2(n13930), .ZN(P2_U2969) );
  NAND2_X1 U15681 ( .A1(n15419), .A2(n13932), .ZN(n13946) );
  XNOR2_X1 U15682 ( .A(n11702), .B(n13933), .ZN(n13944) );
  NAND2_X1 U15683 ( .A1(n13934), .A2(n14049), .ZN(n14177) );
  MUX2_X1 U15684 ( .A(n13935), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16830), .Z(n13936) );
  NOR2_X1 U15685 ( .A1(n13936), .A2(n14191), .ZN(n13937) );
  NAND2_X1 U15686 ( .A1(n14177), .A2(n13937), .ZN(n13942) );
  NAND2_X1 U15687 ( .A1(n14077), .A2(n15094), .ZN(n13938) );
  NOR2_X1 U15688 ( .A1(n14043), .A2(n13938), .ZN(n14174) );
  INV_X1 U15689 ( .A(n16830), .ZN(n13939) );
  AOI21_X1 U15690 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13939), .A(
        n11711), .ZN(n13940) );
  NAND2_X1 U15691 ( .A1(n11179), .A2(n13940), .ZN(n13947) );
  NAND2_X1 U15692 ( .A1(n14174), .A2(n13947), .ZN(n13941) );
  NAND2_X1 U15693 ( .A1(n13942), .A2(n13941), .ZN(n13943) );
  AOI21_X1 U15694 ( .B1(n16833), .B2(n13944), .A(n13943), .ZN(n13945) );
  NAND2_X1 U15695 ( .A1(n13946), .A2(n13945), .ZN(n14173) );
  AOI22_X1 U15696 ( .A1(n14173), .A2(n22146), .B1(n22156), .B2(n13947), .ZN(
        n13948) );
  MUX2_X1 U15697 ( .A(n11702), .B(n13948), .S(n22149), .Z(n13949) );
  INV_X1 U15698 ( .A(n13949), .ZN(P1_U3469) );
  AND2_X1 U15699 ( .A1(n13950), .A2(n19073), .ZN(n13951) );
  NOR2_X1 U15700 ( .A1(n13952), .A2(n13951), .ZN(n19070) );
  NOR2_X1 U15701 ( .A1(n18892), .A2(n12850), .ZN(n19068) );
  XNOR2_X1 U15702 ( .A(n15370), .B(n19073), .ZN(n19067) );
  AND2_X1 U15703 ( .A1(n17671), .A2(n19067), .ZN(n13953) );
  AOI211_X1 U15704 ( .C1(n17664), .C2(n19070), .A(n19068), .B(n13953), .ZN(
        n13956) );
  OAI21_X1 U15705 ( .B1(n17670), .B2(n13954), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13955) );
  OAI211_X1 U15706 ( .C1(n17657), .C2(n14615), .A(n13956), .B(n13955), .ZN(
        P2_U3014) );
  OAI21_X1 U15707 ( .B1(n13958), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13957), .ZN(n14089) );
  INV_X1 U15708 ( .A(n13959), .ZN(n13960) );
  AOI21_X1 U15709 ( .B1(n13962), .B2(n13961), .A(n13960), .ZN(n14081) );
  NAND2_X1 U15710 ( .A1(n14081), .A2(n20519), .ZN(n13966) );
  NAND2_X1 U15711 ( .A1(n13963), .A2(n16670), .ZN(n13964) );
  INV_X2 U15712 ( .A(n22001), .ZN(n22016) );
  AND2_X1 U15713 ( .A1(n22016), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14086) );
  AOI21_X1 U15714 ( .B1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13964), .A(
        n14086), .ZN(n13965) );
  OAI211_X1 U15715 ( .C1(n22141), .C2(n14089), .A(n13966), .B(n13965), .ZN(
        P1_U2999) );
  OR2_X1 U15716 ( .A1(n17633), .A2(n13967), .ZN(n13969) );
  OAI211_X1 U15717 ( .C1(n17676), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        n13972) );
  NOR2_X1 U15718 ( .A1(n17657), .A2(n15575), .ZN(n13971) );
  AOI211_X1 U15719 ( .C1(n17640), .C2(n13967), .A(n13972), .B(n13971), .ZN(
        n13973) );
  OAI21_X1 U15720 ( .B1(n13974), .B2(n17608), .A(n13973), .ZN(P2_U3013) );
  NOR2_X1 U15721 ( .A1(n17545), .A2(n21842), .ZN(n13975) );
  INV_X1 U15722 ( .A(DATAI_8_), .ZN(n13977) );
  INV_X1 U15723 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20549) );
  MUX2_X1 U15724 ( .A(n13977), .B(n20549), .S(n16270), .Z(n16501) );
  INV_X1 U15725 ( .A(n16501), .ZN(n13978) );
  NAND2_X1 U15726 ( .A1(n11272), .A2(n13978), .ZN(n13981) );
  NAND2_X1 U15727 ( .A1(n14028), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13979) );
  OAI211_X1 U15728 ( .C1(n15479), .C2(n14035), .A(n13981), .B(n13979), .ZN(
        P1_U2960) );
  NAND2_X1 U15729 ( .A1(n14028), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13980) );
  OAI211_X1 U15730 ( .C1(n14035), .C2(n16499), .A(n13981), .B(n13980), .ZN(
        P1_U2945) );
  INV_X1 U15731 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n16492) );
  MUX2_X1 U15732 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n16270), .Z(
        n16495) );
  NAND2_X1 U15733 ( .A1(n11272), .A2(n16495), .ZN(n13998) );
  NAND2_X1 U15734 ( .A1(n14028), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13982) );
  OAI211_X1 U15735 ( .C1(n14035), .C2(n16492), .A(n13998), .B(n13982), .ZN(
        P1_U2946) );
  MUX2_X1 U15736 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n16270), .Z(
        n16489) );
  NAND2_X1 U15737 ( .A1(n11272), .A2(n16489), .ZN(n14001) );
  NAND2_X1 U15738 ( .A1(n14028), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13983) );
  OAI211_X1 U15739 ( .C1(n14035), .C2(n16486), .A(n14001), .B(n13983), .ZN(
        P1_U2947) );
  INV_X1 U15740 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15157) );
  MUX2_X1 U15741 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n16270), .Z(
        n16274) );
  NAND2_X1 U15742 ( .A1(n11272), .A2(n16274), .ZN(n13992) );
  NAND2_X1 U15743 ( .A1(n14028), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13984) );
  OAI211_X1 U15744 ( .C1(n14035), .C2(n15157), .A(n13992), .B(n13984), .ZN(
        P1_U2951) );
  INV_X1 U15745 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20375) );
  MUX2_X1 U15746 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n16270), .Z(
        n16482) );
  NAND2_X1 U15747 ( .A1(n11272), .A2(n16482), .ZN(n13996) );
  NAND2_X1 U15748 ( .A1(n14028), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13985) );
  OAI211_X1 U15749 ( .C1(n20375), .C2(n14035), .A(n13996), .B(n13985), .ZN(
        P1_U2963) );
  NAND2_X1 U15750 ( .A1(n16270), .A2(n20545), .ZN(n13986) );
  OAI21_X1 U15751 ( .B1(n16270), .B2(DATAI_6_), .A(n13986), .ZN(n16513) );
  INV_X1 U15752 ( .A(n16513), .ZN(n14542) );
  NAND2_X1 U15753 ( .A1(n11272), .A2(n14542), .ZN(n13990) );
  NAND2_X1 U15754 ( .A1(n14028), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n13987) );
  OAI211_X1 U15755 ( .C1(n15270), .C2(n14035), .A(n13990), .B(n13987), .ZN(
        P1_U2958) );
  INV_X1 U15756 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15149) );
  MUX2_X1 U15757 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n16270), .Z(
        n16468) );
  NAND2_X1 U15758 ( .A1(n11272), .A2(n16468), .ZN(n13994) );
  NAND2_X1 U15759 ( .A1(n14028), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13988) );
  OAI211_X1 U15760 ( .C1(n14035), .C2(n15149), .A(n13994), .B(n13988), .ZN(
        P1_U2950) );
  INV_X1 U15761 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n16511) );
  NAND2_X1 U15762 ( .A1(n14028), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13989) );
  OAI211_X1 U15763 ( .C1(n14035), .C2(n16511), .A(n13990), .B(n13989), .ZN(
        P1_U2943) );
  INV_X1 U15764 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20382) );
  NAND2_X1 U15765 ( .A1(n14028), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13991) );
  OAI211_X1 U15766 ( .C1(n20382), .C2(n14035), .A(n13992), .B(n13991), .ZN(
        P1_U2966) );
  INV_X1 U15767 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20380) );
  NAND2_X1 U15768 ( .A1(n14028), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n13993) );
  OAI211_X1 U15769 ( .C1(n20380), .C2(n14035), .A(n13994), .B(n13993), .ZN(
        P1_U2965) );
  NAND2_X1 U15770 ( .A1(n14028), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13995) );
  OAI211_X1 U15771 ( .C1(n14035), .C2(n16479), .A(n13996), .B(n13995), .ZN(
        P1_U2948) );
  INV_X1 U15772 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20370) );
  NAND2_X1 U15773 ( .A1(n14028), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n13997) );
  OAI211_X1 U15774 ( .C1(n20370), .C2(n14035), .A(n13998), .B(n13997), .ZN(
        P1_U2961) );
  MUX2_X1 U15775 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n16270), .Z(
        n16475) );
  NAND2_X1 U15776 ( .A1(n11272), .A2(n16475), .ZN(n14003) );
  NAND2_X1 U15777 ( .A1(n14028), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13999) );
  OAI211_X1 U15778 ( .C1(n14035), .C2(n16472), .A(n14003), .B(n13999), .ZN(
        P1_U2949) );
  INV_X1 U15779 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20373) );
  NAND2_X1 U15780 ( .A1(n14028), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14000) );
  OAI211_X1 U15781 ( .C1(n20373), .C2(n14035), .A(n14001), .B(n14000), .ZN(
        P1_U2962) );
  INV_X1 U15782 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20378) );
  NAND2_X1 U15783 ( .A1(n14028), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n14002) );
  OAI211_X1 U15784 ( .C1(n20378), .C2(n14035), .A(n14003), .B(n14002), .ZN(
        P1_U2964) );
  INV_X1 U15785 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20539) );
  NAND2_X1 U15786 ( .A1(n16270), .A2(n20539), .ZN(n14004) );
  OAI21_X1 U15787 ( .B1(n16270), .B2(DATAI_3_), .A(n14004), .ZN(n14555) );
  INV_X1 U15788 ( .A(n14555), .ZN(n16531) );
  NAND2_X1 U15789 ( .A1(n11272), .A2(n16531), .ZN(n14007) );
  NAND2_X1 U15790 ( .A1(n14028), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n14005) );
  OAI211_X1 U15791 ( .C1(n11997), .C2(n14035), .A(n14007), .B(n14005), .ZN(
        P1_U2955) );
  INV_X1 U15792 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15163) );
  NAND2_X1 U15793 ( .A1(n14028), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14006) );
  OAI211_X1 U15794 ( .C1(n15163), .C2(n14035), .A(n14007), .B(n14006), .ZN(
        P1_U2940) );
  INV_X1 U15795 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15147) );
  INV_X1 U15796 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20533) );
  NAND2_X1 U15797 ( .A1(n16270), .A2(n20533), .ZN(n14008) );
  OAI21_X1 U15798 ( .B1(n16270), .B2(DATAI_0_), .A(n14008), .ZN(n14549) );
  INV_X1 U15799 ( .A(n14549), .ZN(n16544) );
  NAND2_X1 U15800 ( .A1(n11272), .A2(n16544), .ZN(n14011) );
  NAND2_X1 U15801 ( .A1(n14028), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14009) );
  OAI211_X1 U15802 ( .C1(n15147), .C2(n14035), .A(n14011), .B(n14009), .ZN(
        P1_U2937) );
  INV_X1 U15803 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20358) );
  NAND2_X1 U15804 ( .A1(n14028), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14010) );
  OAI211_X1 U15805 ( .C1(n20358), .C2(n14035), .A(n14011), .B(n14010), .ZN(
        P1_U2952) );
  INV_X1 U15806 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14247) );
  INV_X1 U15807 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20535) );
  NAND2_X1 U15808 ( .A1(n16270), .A2(n20535), .ZN(n14012) );
  OAI21_X1 U15809 ( .B1(n16270), .B2(DATAI_1_), .A(n14012), .ZN(n14536) );
  INV_X1 U15810 ( .A(n14536), .ZN(n16538) );
  NAND2_X1 U15811 ( .A1(n11272), .A2(n16538), .ZN(n14015) );
  NAND2_X1 U15812 ( .A1(n14028), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14013) );
  OAI211_X1 U15813 ( .C1(n14247), .C2(n14035), .A(n14015), .B(n14013), .ZN(
        P1_U2938) );
  NAND2_X1 U15814 ( .A1(n14028), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n14014) );
  OAI211_X1 U15815 ( .C1(n11920), .C2(n14035), .A(n14015), .B(n14014), .ZN(
        P1_U2953) );
  INV_X1 U15816 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20537) );
  NAND2_X1 U15817 ( .A1(n16270), .A2(n20537), .ZN(n14016) );
  OAI21_X1 U15818 ( .B1(n16270), .B2(DATAI_2_), .A(n14016), .ZN(n14562) );
  INV_X1 U15819 ( .A(n14562), .ZN(n16535) );
  NAND2_X1 U15820 ( .A1(n11272), .A2(n16535), .ZN(n14019) );
  NAND2_X1 U15821 ( .A1(n14028), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n14017) );
  OAI211_X1 U15822 ( .C1(n11966), .C2(n14035), .A(n14019), .B(n14017), .ZN(
        P1_U2954) );
  INV_X1 U15823 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14249) );
  NAND2_X1 U15824 ( .A1(n14028), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14018) );
  OAI211_X1 U15825 ( .C1(n14249), .C2(n14035), .A(n14019), .B(n14018), .ZN(
        P1_U2939) );
  INV_X1 U15826 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20363) );
  NAND2_X1 U15827 ( .A1(n16270), .A2(n20541), .ZN(n14020) );
  OAI21_X1 U15828 ( .B1(n16270), .B2(DATAI_4_), .A(n14020), .ZN(n22383) );
  INV_X1 U15829 ( .A(n22383), .ZN(n14021) );
  NAND2_X1 U15830 ( .A1(n11272), .A2(n14021), .ZN(n14024) );
  NAND2_X1 U15831 ( .A1(n14028), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n14022) );
  OAI211_X1 U15832 ( .C1(n20363), .C2(n14035), .A(n14024), .B(n14022), .ZN(
        P1_U2956) );
  INV_X1 U15833 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n16524) );
  NAND2_X1 U15834 ( .A1(n14028), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14023) );
  OAI211_X1 U15835 ( .C1(n14035), .C2(n16524), .A(n14024), .B(n14023), .ZN(
        P1_U2941) );
  INV_X1 U15836 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n16505) );
  INV_X1 U15837 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20547) );
  NAND2_X1 U15838 ( .A1(n16270), .A2(n20547), .ZN(n14025) );
  OAI21_X1 U15839 ( .B1(n16270), .B2(DATAI_7_), .A(n14025), .ZN(n22480) );
  INV_X1 U15840 ( .A(n22480), .ZN(n14026) );
  NAND2_X1 U15841 ( .A1(n11272), .A2(n14026), .ZN(n14030) );
  NAND2_X1 U15842 ( .A1(n14028), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14027) );
  OAI211_X1 U15843 ( .C1(n14035), .C2(n16505), .A(n14030), .B(n14027), .ZN(
        P1_U2944) );
  NAND2_X1 U15844 ( .A1(n14028), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n14029) );
  OAI211_X1 U15845 ( .C1(n12073), .C2(n14035), .A(n14030), .B(n14029), .ZN(
        P1_U2959) );
  INV_X1 U15846 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20365) );
  INV_X1 U15847 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20543) );
  NOR2_X1 U15848 ( .A1(n16270), .A2(DATAI_5_), .ZN(n14031) );
  AOI21_X1 U15849 ( .B1(n16270), .B2(n20543), .A(n14031), .ZN(n16520) );
  NAND2_X1 U15850 ( .A1(n11272), .A2(n16520), .ZN(n14034) );
  NAND2_X1 U15851 ( .A1(n14028), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n14032) );
  OAI211_X1 U15852 ( .C1(n20365), .C2(n14035), .A(n14034), .B(n14032), .ZN(
        P1_U2957) );
  INV_X1 U15853 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n16517) );
  NAND2_X1 U15854 ( .A1(n14028), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14033) );
  OAI211_X1 U15855 ( .C1(n14035), .C2(n16517), .A(n14034), .B(n14033), .ZN(
        P1_U2942) );
  OR2_X1 U15856 ( .A1(n14036), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14170) );
  AOI21_X1 U15857 ( .B1(n15294), .B2(n22189), .A(n22181), .ZN(n14037) );
  NAND2_X1 U15858 ( .A1(n15085), .A2(n14037), .ZN(n14042) );
  NAND2_X1 U15859 ( .A1(n11828), .A2(n22189), .ZN(n15293) );
  INV_X1 U15860 ( .A(n15293), .ZN(n14038) );
  OAI211_X1 U15861 ( .C1(n14039), .C2(n14038), .A(n14245), .B(n16272), .ZN(
        n14040) );
  NAND2_X1 U15862 ( .A1(n15095), .A2(n14040), .ZN(n14041) );
  MUX2_X1 U15863 ( .A(n14042), .B(n14041), .S(n14565), .Z(n14048) );
  OR2_X1 U15864 ( .A1(n14043), .A2(n11828), .ZN(n14044) );
  OR2_X1 U15865 ( .A1(n15095), .A2(n14044), .ZN(n14046) );
  INV_X1 U15866 ( .A(n14053), .ZN(n14051) );
  AND2_X1 U15867 ( .A1(n17539), .A2(n14049), .ZN(n15084) );
  OAI211_X1 U15868 ( .C1(n11838), .C2(n14051), .A(n14050), .B(n15084), .ZN(
        n14052) );
  NAND3_X1 U15869 ( .A1(n14170), .A2(n14169), .A3(n22018), .ZN(n14071) );
  NAND2_X1 U15870 ( .A1(n13809), .A2(n11828), .ZN(n14055) );
  NAND2_X1 U15871 ( .A1(n14053), .A2(n11838), .ZN(n14054) );
  NAND2_X1 U15872 ( .A1(n14055), .A2(n14054), .ZN(n14056) );
  NAND2_X1 U15873 ( .A1(n14558), .A2(n14245), .ZN(n14072) );
  INV_X1 U15874 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14147) );
  INV_X1 U15875 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21879) );
  NAND2_X1 U15876 ( .A1(n14072), .A2(n21879), .ZN(n14058) );
  NAND2_X1 U15877 ( .A1(n16206), .A2(n14147), .ZN(n14057) );
  NAND3_X1 U15878 ( .A1(n14058), .A2(n16261), .A3(n14057), .ZN(n14059) );
  XNOR2_X1 U15879 ( .A(n14074), .B(n14267), .ZN(n15413) );
  NAND2_X1 U15880 ( .A1(n15413), .A2(n16206), .ZN(n14268) );
  OAI21_X1 U15881 ( .B1(n15413), .B2(n16206), .A(n14268), .ZN(n14146) );
  INV_X1 U15882 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21878) );
  NAND2_X1 U15883 ( .A1(n14062), .A2(n14061), .ZN(n14063) );
  NAND2_X1 U15884 ( .A1(n14066), .A2(n14063), .ZN(n21855) );
  OR2_X1 U15885 ( .A1(n21855), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14065) );
  OR2_X1 U15886 ( .A1(n14066), .A2(n22016), .ZN(n14064) );
  INV_X1 U15887 ( .A(n21880), .ZN(n21934) );
  AOI21_X1 U15888 ( .B1(n21952), .B2(n21878), .A(n21934), .ZN(n14084) );
  NAND2_X1 U15889 ( .A1(n22016), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14166) );
  OAI21_X1 U15890 ( .B1(n14084), .B2(n21879), .A(n14166), .ZN(n14069) );
  NAND2_X1 U15891 ( .A1(n14066), .A2(n16833), .ZN(n21850) );
  INV_X1 U15892 ( .A(n21952), .ZN(n21884) );
  AND2_X1 U15893 ( .A1(n21932), .A2(n21884), .ZN(n16785) );
  INV_X1 U15894 ( .A(n21850), .ZN(n14067) );
  NOR2_X1 U15895 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14067), .ZN(
        n16215) );
  NOR3_X1 U15896 ( .A1(n16785), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n16215), .ZN(n14068) );
  AOI211_X1 U15897 ( .C1(n22017), .C2(n14146), .A(n14069), .B(n14068), .ZN(
        n14070) );
  NAND2_X1 U15898 ( .A1(n14071), .A2(n14070), .ZN(P1_U3030) );
  OR2_X1 U15899 ( .A1(n16210), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14073) );
  NAND2_X1 U15900 ( .A1(n14074), .A2(n14073), .ZN(n15436) );
  NAND2_X1 U15901 ( .A1(n15088), .A2(n14093), .ZN(n14075) );
  OR2_X1 U15902 ( .A1(n15095), .A2(n14075), .ZN(n14080) );
  NOR3_X1 U15903 ( .A1(n11571), .A2(n15092), .A3(n22162), .ZN(n14078) );
  NAND3_X1 U15904 ( .A1(n11572), .A2(n14078), .A3(n14077), .ZN(n14095) );
  OR2_X1 U15905 ( .A1(n14095), .A2(n16209), .ZN(n14079) );
  NAND2_X2 U15906 ( .A1(n16451), .A2(n22476), .ZN(n16453) );
  INV_X1 U15907 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14082) );
  INV_X1 U15908 ( .A(n14081), .ZN(n15438) );
  OAI222_X1 U15909 ( .A1(n15436), .A2(n16453), .B1(n14082), .B2(n16451), .C1(
        n16425), .C2(n15438), .ZN(P1_U2872) );
  INV_X1 U15910 ( .A(n15436), .ZN(n14087) );
  INV_X1 U15911 ( .A(n21855), .ZN(n21852) );
  NOR2_X1 U15912 ( .A1(n21852), .A2(n21952), .ZN(n14083) );
  AOI22_X1 U15913 ( .A1(n14084), .A2(n21850), .B1(n14083), .B2(n21878), .ZN(
        n14085) );
  AOI211_X1 U15914 ( .C1(n22017), .C2(n14087), .A(n14086), .B(n14085), .ZN(
        n14088) );
  OAI21_X1 U15915 ( .B1(n14089), .B2(n22004), .A(n14088), .ZN(P1_U3031) );
  INV_X1 U15916 ( .A(DATAI_15_), .ZN(n14917) );
  NAND2_X1 U15917 ( .A1(n16270), .A2(BUF1_REG_15__SCAN_IN), .ZN(n14090) );
  OAI21_X1 U15918 ( .B1(n16270), .B2(n14917), .A(n14090), .ZN(n16550) );
  AOI222_X1 U15919 ( .A1(n16550), .A2(n11272), .B1(P1_EAX_REG_15__SCAN_IN), 
        .B2(n14091), .C1(n14028), .C2(P1_LWORD_REG_15__SCAN_IN), .ZN(n14092)
         );
  INV_X1 U15920 ( .A(n14092), .ZN(P1_U2967) );
  NAND2_X1 U15921 ( .A1(n14094), .A2(n14093), .ZN(n14097) );
  OR2_X1 U15922 ( .A1(n14095), .A2(n15284), .ZN(n14096) );
  INV_X1 U15923 ( .A(n14098), .ZN(n14099) );
  NAND2_X1 U15924 ( .A1(n14099), .A2(n15092), .ZN(n14100) );
  INV_X1 U15925 ( .A(n16551), .ZN(n15478) );
  OAI222_X1 U15926 ( .A1(n15478), .A2(n14549), .B1(n16523), .B2(n20358), .C1(
        n16553), .C2(n15438), .ZN(P1_U2904) );
  INV_X1 U15927 ( .A(n14646), .ZN(n14101) );
  NAND2_X1 U15928 ( .A1(n14101), .A2(n14642), .ZN(n14301) );
  NAND2_X1 U15929 ( .A1(n14301), .A2(n14589), .ZN(n14102) );
  NAND2_X1 U15930 ( .A1(n15649), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14225) );
  NOR2_X1 U15931 ( .A1(n19838), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14103) );
  AOI21_X1 U15932 ( .B1(n14219), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14103), .ZN(n14104) );
  NAND2_X1 U15933 ( .A1(n19060), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14105) );
  AND4_X1 U15934 ( .A1(n14153), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14105), 
        .A4(n19733), .ZN(n14106) );
  MUX2_X1 U15935 ( .A(n14107), .B(n14615), .S(n16952), .Z(n14108) );
  OAI21_X1 U15936 ( .B1(n16968), .B2(n19674), .A(n14108), .ZN(P2_U2887) );
  INV_X1 U15937 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15751) );
  AOI22_X1 U15938 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n17733), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17732), .ZN(n14109) );
  OAI21_X1 U15939 ( .B1(n15751), .B2(n14125), .A(n14109), .ZN(P2_U2935) );
  INV_X1 U15940 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U15941 ( .A1(n17733), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14110) );
  OAI21_X1 U15942 ( .B1(n16993), .B2(n14125), .A(n14110), .ZN(P2_U2925) );
  AOI22_X1 U15943 ( .A1(n17733), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14111) );
  OAI21_X1 U15944 ( .B1(n14112), .B2(n14125), .A(n14111), .ZN(P2_U2923) );
  INV_X1 U15945 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U15946 ( .A1(n17733), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14113) );
  OAI21_X1 U15947 ( .B1(n17010), .B2(n14125), .A(n14113), .ZN(P2_U2927) );
  INV_X1 U15948 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U15949 ( .A1(n17733), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14114) );
  OAI21_X1 U15950 ( .B1(n17002), .B2(n14125), .A(n14114), .ZN(P2_U2926) );
  INV_X1 U15951 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16246) );
  AOI22_X1 U15952 ( .A1(n17733), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14115) );
  OAI21_X1 U15953 ( .B1(n16246), .B2(n14125), .A(n14115), .ZN(P2_U2922) );
  INV_X1 U15954 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U15955 ( .A1(n17733), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14116) );
  OAI21_X1 U15956 ( .B1(n14117), .B2(n14125), .A(n14116), .ZN(P2_U2931) );
  INV_X1 U15957 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14119) );
  AOI22_X1 U15958 ( .A1(n17733), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14118) );
  OAI21_X1 U15959 ( .B1(n14119), .B2(n14125), .A(n14118), .ZN(P2_U2929) );
  AOI22_X1 U15960 ( .A1(n17733), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14120) );
  OAI21_X1 U15961 ( .B1(n17019), .B2(n14125), .A(n14120), .ZN(P2_U2928) );
  INV_X1 U15962 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U15963 ( .A1(n17733), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14121) );
  OAI21_X1 U15964 ( .B1(n16984), .B2(n14125), .A(n14121), .ZN(P2_U2924) );
  INV_X1 U15965 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U15966 ( .A1(n17733), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14122) );
  OAI21_X1 U15967 ( .B1(n17028), .B2(n14125), .A(n14122), .ZN(P2_U2930) );
  INV_X1 U15968 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15819) );
  AOI22_X1 U15969 ( .A1(n17725), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14123) );
  OAI21_X1 U15970 ( .B1(n15819), .B2(n14125), .A(n14123), .ZN(P2_U2933) );
  INV_X1 U15971 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15891) );
  AOI22_X1 U15972 ( .A1(n17725), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14124) );
  OAI21_X1 U15973 ( .B1(n15891), .B2(n14125), .A(n14124), .ZN(P2_U2932) );
  AOI21_X1 U15974 ( .B1(n14128), .B2(n14127), .A(n14126), .ZN(n14143) );
  INV_X1 U15975 ( .A(n14129), .ZN(n14130) );
  OAI22_X1 U15976 ( .A1(n12865), .A2(n14130), .B1(n14129), .B2(n15470), .ZN(
        n14135) );
  NOR2_X1 U15977 ( .A1(n19133), .A2(n14131), .ZN(n14134) );
  OAI22_X1 U15978 ( .A1(n19134), .A2(n14132), .B1(n19074), .B2(n12865), .ZN(
        n14133) );
  AOI211_X1 U15979 ( .C1(n17268), .C2(n14135), .A(n14134), .B(n14133), .ZN(
        n14140) );
  XNOR2_X1 U15980 ( .A(n14136), .B(n14137), .ZN(n20059) );
  AOI21_X1 U15981 ( .B1(n19129), .B2(n20059), .A(n14138), .ZN(n14139) );
  OAI211_X1 U15982 ( .C1(n19091), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        n14142) );
  OR2_X1 U15983 ( .A1(n14143), .A2(n14142), .ZN(P2_U3044) );
  OAI21_X1 U15984 ( .B1(n14145), .B2(n14144), .A(n14314), .ZN(n15418) );
  INV_X1 U15985 ( .A(n14146), .ZN(n14148) );
  OAI22_X1 U15986 ( .A1(n16453), .A2(n14148), .B1(n14147), .B2(n16451), .ZN(
        n14149) );
  INV_X1 U15987 ( .A(n14149), .ZN(n14150) );
  OAI21_X1 U15988 ( .B1(n15418), .B2(n16425), .A(n14150), .ZN(P1_U2871) );
  NAND2_X1 U15989 ( .A1(n14219), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14151) );
  NAND2_X1 U15990 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19789) );
  NAND2_X1 U15991 ( .A1(n19819), .A2(n19807), .ZN(n19835) );
  AND2_X1 U15992 ( .A1(n19789), .A2(n19835), .ZN(n19754) );
  NAND2_X1 U15993 ( .A1(n19754), .A2(n19788), .ZN(n19810) );
  NAND2_X1 U15994 ( .A1(n14151), .A2(n19810), .ZN(n14152) );
  NAND2_X1 U15995 ( .A1(n16085), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14155) );
  INV_X1 U15996 ( .A(n14154), .ZN(n14156) );
  NAND2_X1 U15997 ( .A1(n14156), .A2(n14155), .ZN(n14157) );
  INV_X1 U15998 ( .A(n19789), .ZN(n14216) );
  NAND2_X1 U15999 ( .A1(n14216), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19664) );
  NAND2_X1 U16000 ( .A1(n19789), .A2(n19787), .ZN(n14158) );
  NAND2_X1 U16001 ( .A1(n19664), .A2(n14158), .ZN(n15633) );
  NOR2_X1 U16002 ( .A1(n15633), .A2(n19838), .ZN(n14159) );
  AOI21_X1 U16003 ( .B1(n14219), .B2(n17422), .A(n14159), .ZN(n14160) );
  NAND2_X1 U16004 ( .A1(n16085), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14210) );
  MUX2_X1 U16005 ( .A(n13416), .B(n14131), .S(n16952), .Z(n14165) );
  OAI21_X1 U16006 ( .B1(n17686), .B2(n16968), .A(n14165), .ZN(P2_U2885) );
  OAI21_X1 U16007 ( .B1(n16670), .B2(n14168), .A(n14166), .ZN(n14167) );
  AOI21_X1 U16008 ( .B1(n20505), .B2(n14168), .A(n14167), .ZN(n14172) );
  NAND3_X1 U16009 ( .A1(n14170), .A2(n14169), .A3(n20518), .ZN(n14171) );
  OAI211_X1 U16010 ( .C1(n15418), .C2(n20496), .A(n14172), .B(n14171), .ZN(
        P1_U2998) );
  OAI222_X1 U16011 ( .A1(n15478), .A2(n14536), .B1(n16523), .B2(n11920), .C1(
        n16553), .C2(n15418), .ZN(P1_U2903) );
  MUX2_X1 U16012 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14173), .S(
        n17515), .Z(n17529) );
  XNOR2_X1 U16013 ( .A(n16830), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16848) );
  INV_X1 U16014 ( .A(n14174), .ZN(n14175) );
  NOR2_X1 U16015 ( .A1(n14175), .A2(n16848), .ZN(n14176) );
  AOI21_X1 U16016 ( .B1(n14177), .B2(n16848), .A(n14176), .ZN(n14180) );
  NAND3_X1 U16017 ( .A1(n16833), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n14178), .ZN(n14179) );
  OAI211_X1 U16018 ( .C1(n16826), .C2(n16829), .A(n14180), .B(n14179), .ZN(
        n16843) );
  INV_X1 U16019 ( .A(n17515), .ZN(n14181) );
  MUX2_X1 U16020 ( .A(n16843), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14181), .Z(n14183) );
  AND2_X1 U16021 ( .A1(n16832), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14182) );
  AND2_X1 U16022 ( .A1(n16833), .A2(n14182), .ZN(n16842) );
  OR2_X1 U16023 ( .A1(n14183), .A2(n16842), .ZN(n17524) );
  NAND3_X1 U16024 ( .A1(n17529), .A2(n17524), .A3(n15288), .ZN(n14194) );
  INV_X1 U16025 ( .A(n15165), .ZN(n14522) );
  OR2_X1 U16026 ( .A1(n11973), .A2(n14522), .ZN(n14184) );
  XNOR2_X1 U16027 ( .A(n14184), .B(n12584), .ZN(n22144) );
  NAND2_X1 U16028 ( .A1(n22145), .A2(n15288), .ZN(n14185) );
  OR2_X1 U16029 ( .A1(n22144), .A2(n14185), .ZN(n14189) );
  NAND2_X1 U16030 ( .A1(n17515), .A2(n15288), .ZN(n14187) );
  NOR2_X1 U16031 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n12584), .ZN(n14186) );
  NAND2_X1 U16032 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  NAND2_X1 U16033 ( .A1(n14189), .A2(n14188), .ZN(n14195) );
  AND2_X1 U16034 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22142), .ZN(n14190) );
  AND2_X1 U16035 ( .A1(n14191), .A2(n14190), .ZN(n14192) );
  NOR2_X1 U16036 ( .A1(n14195), .A2(n14192), .ZN(n14193) );
  NAND2_X1 U16037 ( .A1(n14194), .A2(n14193), .ZN(n17533) );
  INV_X1 U16038 ( .A(n14195), .ZN(n14196) );
  NAND2_X1 U16039 ( .A1(n14196), .A2(n11719), .ZN(n14197) );
  NAND2_X1 U16040 ( .A1(n17533), .A2(n14197), .ZN(n14201) );
  NAND2_X1 U16041 ( .A1(n14201), .A2(n22142), .ZN(n14199) );
  NOR2_X1 U16042 ( .A1(n22153), .A2(n22152), .ZN(n14198) );
  NAND2_X1 U16043 ( .A1(n14199), .A2(n14198), .ZN(n14200) );
  NOR2_X1 U16044 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22157) );
  INV_X1 U16045 ( .A(n22157), .ZN(n15279) );
  NAND2_X1 U16046 ( .A1(n14200), .A2(n22479), .ZN(n17556) );
  INV_X1 U16047 ( .A(n14201), .ZN(n14202) );
  NOR2_X1 U16048 ( .A1(n14202), .A2(n22152), .ZN(n22160) );
  NAND2_X1 U16049 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22280), .ZN(n15123) );
  INV_X1 U16050 ( .A(n15123), .ZN(n16827) );
  OAI22_X1 U16051 ( .A1(n14687), .A2(n22290), .B1(n14523), .B2(n16827), .ZN(
        n14203) );
  OAI21_X1 U16052 ( .B1(n22160), .B2(n14203), .A(n17556), .ZN(n14204) );
  OAI21_X1 U16053 ( .B1(n17556), .B2(n15376), .A(n14204), .ZN(P1_U3478) );
  NAND2_X1 U16054 ( .A1(n19690), .A2(n15746), .ZN(n14209) );
  NAND2_X1 U16055 ( .A1(n16952), .A2(n14605), .ZN(n14208) );
  OAI211_X1 U16056 ( .C1(n16952), .C2(n15574), .A(n14209), .B(n14208), .ZN(
        P2_U2886) );
  INV_X1 U16057 ( .A(n14210), .ZN(n14211) );
  NAND2_X1 U16058 ( .A1(n14212), .A2(n14211), .ZN(n14213) );
  NAND2_X1 U16059 ( .A1(n14254), .A2(n14215), .ZN(n14221) );
  NAND2_X1 U16060 ( .A1(n19664), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14217) );
  NAND2_X1 U16061 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19786), .ZN(
        n19757) );
  INV_X1 U16062 ( .A(n19757), .ZN(n19769) );
  NAND2_X1 U16063 ( .A1(n14216), .A2(n19769), .ZN(n19746) );
  NAND2_X1 U16064 ( .A1(n14217), .A2(n19746), .ZN(n14218) );
  AND2_X1 U16065 ( .A1(n14218), .A2(n19788), .ZN(n15643) );
  AOI21_X1 U16066 ( .B1(n14219), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n15643), .ZN(n14220) );
  NAND2_X1 U16067 ( .A1(n14221), .A2(n14220), .ZN(n14223) );
  INV_X1 U16068 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15992) );
  NOR2_X1 U16069 ( .A1(n16092), .A2(n15992), .ZN(n14222) );
  OR2_X1 U16070 ( .A1(n14223), .A2(n14222), .ZN(n14224) );
  NAND2_X1 U16071 ( .A1(n14223), .A2(n14222), .ZN(n14228) );
  INV_X1 U16072 ( .A(n14225), .ZN(n14226) );
  NAND2_X1 U16073 ( .A1(n14226), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14227) );
  INV_X1 U16074 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16001) );
  NOR2_X1 U16075 ( .A1(n16092), .A2(n16001), .ZN(n14234) );
  XOR2_X1 U16076 ( .A(n14258), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14233)
         );
  AND2_X1 U16077 ( .A1(n14239), .A2(n14230), .ZN(n14231) );
  OR2_X1 U16078 ( .A1(n14231), .A2(n14261), .ZN(n15687) );
  INV_X1 U16079 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n15243) );
  MUX2_X1 U16080 ( .A(n15687), .B(n15243), .S(n16966), .Z(n14232) );
  OAI21_X1 U16081 ( .B1(n14233), .B2(n16968), .A(n14232), .ZN(P2_U2882) );
  OAI21_X1 U16082 ( .B1(n14235), .B2(n14234), .A(n14258), .ZN(n18729) );
  NAND2_X1 U16083 ( .A1(n14237), .A2(n14236), .ZN(n14238) );
  NAND2_X1 U16084 ( .A1(n14239), .A2(n14238), .ZN(n18743) );
  MUX2_X1 U16085 ( .A(n18743), .B(n14240), .S(n16966), .Z(n14241) );
  OAI21_X1 U16086 ( .B1(n18729), .B2(n16968), .A(n14241), .ZN(P2_U2883) );
  NAND2_X1 U16087 ( .A1(n14035), .A2(n14242), .ZN(n14244) );
  INV_X1 U16088 ( .A(n22189), .ZN(n14243) );
  NAND2_X1 U16089 ( .A1(n20356), .A2(n14245), .ZN(n15162) );
  NOR2_X1 U16090 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22152), .ZN(n20376) );
  NOR2_X4 U16091 ( .A1(n20356), .A2(n21841), .ZN(n20371) );
  AOI22_X1 U16092 ( .A1(n21841), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14246) );
  OAI21_X1 U16093 ( .B1(n14247), .B2(n15162), .A(n14246), .ZN(P1_U2919) );
  AOI22_X1 U16094 ( .A1(n21841), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14248) );
  OAI21_X1 U16095 ( .B1(n14249), .B2(n15162), .A(n14248), .ZN(P1_U2918) );
  OR2_X1 U16096 ( .A1(n14250), .A2(n14251), .ZN(n14253) );
  INV_X1 U16097 ( .A(n14255), .ZN(n15473) );
  NOR2_X1 U16098 ( .A1(n15473), .A2(n16966), .ZN(n14256) );
  AOI21_X1 U16099 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16966), .A(n14256), .ZN(
        n14257) );
  OAI21_X1 U16100 ( .B1(n19795), .B2(n16968), .A(n14257), .ZN(P2_U2884) );
  INV_X1 U16101 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16018) );
  NOR2_X1 U16102 ( .A1(n14258), .A2(n16018), .ZN(n14259) );
  OAI211_X1 U16103 ( .C1(n14259), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15746), .B(n14321), .ZN(n14264) );
  OR2_X1 U16104 ( .A1(n14261), .A2(n14260), .ZN(n14262) );
  AND2_X1 U16105 ( .A1(n14262), .A2(n14275), .ZN(n18751) );
  NAND2_X1 U16106 ( .A1(n18751), .A2(n16952), .ZN(n14263) );
  OAI211_X1 U16107 ( .C1(n16952), .C2(n18744), .A(n14264), .B(n14263), .ZN(
        P2_U2881) );
  OAI21_X1 U16108 ( .B1(n14266), .B2(n14265), .A(n15106), .ZN(n14332) );
  INV_X1 U16109 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14329) );
  NAND2_X1 U16110 ( .A1(n14072), .A2(n21893), .ZN(n14270) );
  NAND2_X1 U16111 ( .A1(n16206), .A2(n14329), .ZN(n14269) );
  NAND3_X1 U16112 ( .A1(n14270), .A2(n16261), .A3(n14269), .ZN(n14271) );
  NAND2_X1 U16113 ( .A1(n14272), .A2(n14271), .ZN(n14327) );
  NAND2_X1 U16114 ( .A1(n14328), .A2(n14327), .ZN(n14676) );
  MUX2_X1 U16115 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n14273) );
  OAI21_X1 U16116 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16210), .A(
        n14273), .ZN(n14677) );
  XOR2_X1 U16117 ( .A(n14676), .B(n14677), .Z(n21904) );
  INV_X1 U16118 ( .A(n16451), .ZN(n16462) );
  AOI22_X1 U16119 ( .A1(n16463), .A2(n21904), .B1(n16462), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14274) );
  OAI21_X1 U16120 ( .B1(n14332), .B2(n16425), .A(n14274), .ZN(P1_U2869) );
  XOR2_X1 U16121 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14321), .Z(n14281)
         );
  INV_X1 U16122 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14279) );
  NAND2_X1 U16123 ( .A1(n14276), .A2(n14275), .ZN(n14278) );
  INV_X1 U16124 ( .A(n14319), .ZN(n14277) );
  NAND2_X1 U16125 ( .A1(n14278), .A2(n14277), .ZN(n18760) );
  MUX2_X1 U16126 ( .A(n14279), .B(n18760), .S(n16952), .Z(n14280) );
  OAI21_X1 U16127 ( .B1(n14281), .B2(n16968), .A(n14280), .ZN(P2_U2880) );
  INV_X1 U16128 ( .A(n14614), .ZN(n14604) );
  OR2_X1 U16129 ( .A1(n14632), .A2(n14642), .ZN(n14592) );
  NOR2_X1 U16130 ( .A1(n14282), .A2(n17422), .ZN(n14588) );
  INV_X1 U16131 ( .A(n14588), .ZN(n14288) );
  NAND2_X1 U16132 ( .A1(n14592), .A2(n14288), .ZN(n14293) );
  NAND2_X1 U16133 ( .A1(n16124), .A2(n14603), .ZN(n14283) );
  AOI21_X1 U16134 ( .B1(n13180), .B2(n12687), .A(n14283), .ZN(n14292) );
  INV_X1 U16135 ( .A(n12687), .ZN(n14284) );
  NAND2_X1 U16136 ( .A1(n13180), .A2(n14284), .ZN(n14290) );
  NAND2_X1 U16137 ( .A1(n14589), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14287) );
  INV_X1 U16138 ( .A(n14285), .ZN(n14286) );
  OAI21_X1 U16139 ( .B1(n13181), .B2(n14287), .A(n14286), .ZN(n14289) );
  AND3_X1 U16140 ( .A1(n14290), .A2(n14289), .A3(n14288), .ZN(n14291) );
  AOI21_X1 U16141 ( .B1(n14293), .B2(n14292), .A(n14291), .ZN(n14294) );
  AOI21_X1 U16142 ( .B1(n14255), .B2(n14604), .A(n14294), .ZN(n14602) );
  INV_X1 U16143 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U16144 ( .A1(n15237), .A2(n19733), .ZN(n19148) );
  NOR2_X1 U16145 ( .A1(n14602), .A2(n19148), .ZN(n14295) );
  AOI21_X1 U16146 ( .B1(n17691), .B2(n19162), .A(n14295), .ZN(n14307) );
  OR2_X1 U16147 ( .A1(n19062), .A2(n14663), .ZN(n14303) );
  AND2_X1 U16148 ( .A1(n14296), .A2(n19164), .ZN(n15208) );
  INV_X1 U16149 ( .A(n15208), .ZN(n14298) );
  OAI21_X1 U16150 ( .B1(n14298), .B2(n14649), .A(n14297), .ZN(n14299) );
  INV_X1 U16151 ( .A(n14299), .ZN(n14300) );
  NAND2_X1 U16152 ( .A1(n14646), .A2(n14632), .ZN(n15206) );
  AND2_X1 U16153 ( .A1(n14300), .A2(n15206), .ZN(n14302) );
  OAI211_X1 U16154 ( .C1(n14304), .C2(n14303), .A(n14302), .B(n14301), .ZN(
        n14601) );
  NAND2_X1 U16155 ( .A1(n14601), .A2(n19160), .ZN(n14306) );
  NOR2_X1 U16156 ( .A1(n15635), .A2(n15636), .ZN(n19157) );
  AOI22_X1 U16157 ( .A1(n15635), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19157), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n14305) );
  NAND2_X1 U16158 ( .A1(n14306), .A2(n14305), .ZN(n19066) );
  INV_X1 U16159 ( .A(n19066), .ZN(n19057) );
  MUX2_X1 U16160 ( .A(n14307), .B(n14603), .S(n19057), .Z(n14308) );
  INV_X1 U16161 ( .A(n14308), .ZN(P2_U3596) );
  OAI222_X1 U16162 ( .A1(n15478), .A2(n14555), .B1(n16523), .B2(n11997), .C1(
        n16553), .C2(n14332), .ZN(P1_U2901) );
  OAI21_X1 U16163 ( .B1(n14311), .B2(n14310), .A(n14309), .ZN(n21883) );
  INV_X1 U16164 ( .A(n14312), .ZN(n14313) );
  AOI21_X1 U16165 ( .B1(n14315), .B2(n14314), .A(n14313), .ZN(n15291) );
  AOI22_X1 U16166 ( .A1(n20514), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21906), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14316) );
  OAI21_X1 U16167 ( .B1(n20522), .B2(n15301), .A(n14316), .ZN(n14317) );
  AOI21_X1 U16168 ( .B1(n15291), .B2(n20519), .A(n14317), .ZN(n14318) );
  OAI21_X1 U16169 ( .B1(n22141), .B2(n21883), .A(n14318), .ZN(P1_U2997) );
  OAI21_X1 U16170 ( .B1(n14320), .B2(n14319), .A(n15109), .ZN(n19132) );
  INV_X1 U16171 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16120) );
  INV_X1 U16172 ( .A(n15108), .ZN(n14323) );
  OAI211_X1 U16173 ( .C1(n14322), .C2(n14324), .A(n14323), .B(n15746), .ZN(
        n14326) );
  NAND2_X1 U16174 ( .A1(n16966), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14325) );
  OAI211_X1 U16175 ( .C1(n19132), .C2(n16966), .A(n14326), .B(n14325), .ZN(
        P2_U2879) );
  OAI21_X1 U16176 ( .B1(n14328), .B2(n14327), .A(n14676), .ZN(n21886) );
  INV_X1 U16177 ( .A(n15291), .ZN(n14548) );
  OAI222_X1 U16178 ( .A1(n21886), .A2(n16453), .B1(n14329), .B2(n16451), .C1(
        n14548), .C2(n16425), .ZN(P1_U2870) );
  INV_X1 U16179 ( .A(n14332), .ZN(n15420) );
  AOI22_X1 U16180 ( .A1(n20514), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n21906), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14333) );
  OAI21_X1 U16181 ( .B1(n20522), .B2(n15423), .A(n14333), .ZN(n14334) );
  AOI21_X1 U16182 ( .B1(n15420), .B2(n20519), .A(n14334), .ZN(n14335) );
  OAI21_X1 U16183 ( .B1(n22141), .B2(n21903), .A(n14335), .ZN(P1_U2996) );
  INV_X1 U16184 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n21038) );
  INV_X1 U16185 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21030) );
  NOR2_X1 U16186 ( .A1(n21038), .A2(n21030), .ZN(n14439) );
  INV_X2 U16187 ( .A(n17909), .ZN(n17895) );
  AOI22_X1 U16188 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14350) );
  NOR2_X2 U16189 ( .A1(n14339), .A2(n14337), .ZN(n14388) );
  AOI22_X1 U16190 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18116), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14349) );
  NOR2_X2 U16191 ( .A1(n14340), .A2(n14338), .ZN(n18108) );
  AOI22_X1 U16192 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14336) );
  OAI21_X1 U16193 ( .B1(n11214), .B2(n18060), .A(n14336), .ZN(n14347) );
  NOR2_X2 U16194 ( .A1(n21294), .A2(n14338), .ZN(n14484) );
  AOI22_X1 U16195 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14345) );
  AOI22_X1 U16196 ( .A1(n18156), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14344) );
  OR2_X2 U16197 ( .A1(n21296), .A2(n14341), .ZN(n21316) );
  NOR2_X2 U16198 ( .A1(n21310), .A2(n21316), .ZN(n18106) );
  INV_X2 U16199 ( .A(n20700), .ZN(n18148) );
  AOI22_X1 U16200 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14343) );
  AOI22_X1 U16201 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14342) );
  NAND4_X1 U16202 ( .A1(n14345), .A2(n14344), .A3(n14343), .A4(n14342), .ZN(
        n14346) );
  AOI22_X1 U16203 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11168), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U16204 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14354) );
  AOI22_X1 U16205 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18105), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14353) );
  INV_X2 U16206 ( .A(n20700), .ZN(n17901) );
  AOI22_X1 U16207 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14352) );
  NAND4_X1 U16208 ( .A1(n14355), .A2(n14354), .A3(n14353), .A4(n14352), .ZN(
        n14361) );
  AOI22_X1 U16209 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14359) );
  BUF_X2 U16210 ( .A(n14388), .Z(n18154) );
  AOI22_X1 U16211 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14358) );
  AOI22_X1 U16212 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14357) );
  INV_X2 U16213 ( .A(n11218), .ZN(n18126) );
  AOI22_X1 U16214 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14356) );
  NAND4_X1 U16215 ( .A1(n14359), .A2(n14358), .A3(n14357), .A4(n14356), .ZN(
        n14360) );
  AOI22_X1 U16216 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14362) );
  OAI21_X1 U16217 ( .B1(n11214), .B2(n18107), .A(n14362), .ZN(n14368) );
  AOI22_X1 U16218 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14455), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14366) );
  INV_X2 U16219 ( .A(n17909), .ZN(n18132) );
  AOI22_X1 U16220 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14365) );
  AOI22_X1 U16221 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14364) );
  AOI22_X1 U16222 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14363) );
  NAND4_X1 U16223 ( .A1(n14366), .A2(n14365), .A3(n14364), .A4(n14363), .ZN(
        n14367) );
  OAI22_X1 U16224 ( .A1(n21772), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21791), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U16225 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21784), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21296), .ZN(n17460) );
  OAI22_X1 U16226 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21774), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14373), .ZN(n14379) );
  NOR2_X1 U16227 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21774), .ZN(
        n14374) );
  NAND2_X1 U16228 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14373), .ZN(
        n14378) );
  AOI22_X1 U16229 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14379), .B1(
        n14374), .B2(n14378), .ZN(n14382) );
  AOI21_X1 U16230 ( .B1(n21310), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n17459), .ZN(n18046) );
  AND2_X1 U16231 ( .A1(n17460), .A2(n18046), .ZN(n14381) );
  OAI21_X1 U16232 ( .B1(n14377), .B2(n14376), .A(n14382), .ZN(n14375) );
  INV_X1 U16233 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21798) );
  OAI22_X1 U16234 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21798), .B1(
        n14380), .B2(n14379), .ZN(n17461) );
  AOI211_X1 U16235 ( .C1(n14382), .C2(n14381), .A(n18047), .B(n17461), .ZN(
        n21348) );
  AOI22_X1 U16236 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14386) );
  AOI22_X1 U16237 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U16238 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18129), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U16239 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14383) );
  NAND4_X1 U16240 ( .A1(n14386), .A2(n14385), .A3(n14384), .A4(n14383), .ZN(
        n14394) );
  AOI22_X1 U16241 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U16242 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18116), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U16243 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14390) );
  AOI22_X1 U16244 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14389) );
  NAND4_X1 U16245 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n14393) );
  AOI22_X1 U16246 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U16247 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U16248 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14455), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14395) );
  OAI21_X1 U16249 ( .B1(n11214), .B2(n17812), .A(n14395), .ZN(n14401) );
  AOI22_X1 U16250 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14400) );
  AOI22_X1 U16251 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18116), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U16252 ( .A1(n18156), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14398) );
  AOI22_X1 U16253 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U16254 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U16255 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U16256 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14404) );
  OAI21_X1 U16257 ( .B1(n11214), .B2(n18094), .A(n14404), .ZN(n14410) );
  AOI22_X1 U16258 ( .A1(n14472), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18156), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U16259 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14388), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U16260 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18105), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U16261 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14405) );
  NAND4_X1 U16262 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14409) );
  NOR2_X1 U16263 ( .A1(n19325), .A2(n21338), .ZN(n21344) );
  AOI22_X1 U16264 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U16265 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18126), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U16266 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U16267 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14415) );
  NAND4_X1 U16268 ( .A1(n14418), .A2(n14417), .A3(n14416), .A4(n14415), .ZN(
        n14424) );
  AOI22_X1 U16269 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U16270 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U16271 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U16272 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18116), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14419) );
  NAND4_X1 U16273 ( .A1(n14422), .A2(n14421), .A3(n14420), .A4(n14419), .ZN(
        n14423) );
  AOI22_X1 U16274 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11168), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U16275 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U16276 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U16277 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14425) );
  NAND4_X1 U16278 ( .A1(n14428), .A2(n14427), .A3(n14426), .A4(n14425), .ZN(
        n14434) );
  AOI22_X1 U16279 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U16280 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U16281 ( .A1(n14472), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14430) );
  AOI22_X1 U16282 ( .A1(n18156), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14429) );
  NAND4_X1 U16283 ( .A1(n14432), .A2(n14431), .A3(n14430), .A4(n14429), .ZN(
        n14433) );
  NAND2_X1 U16284 ( .A1(n21342), .A2(n19407), .ZN(n18051) );
  NOR2_X1 U16285 ( .A1(n21197), .A2(n17449), .ZN(n14435) );
  NOR2_X1 U16286 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n21830), .ZN(n21812) );
  NAND2_X1 U16287 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21812), .ZN(n21807) );
  NAND2_X1 U16288 ( .A1(n21263), .A2(n18039), .ZN(n18035) );
  INV_X1 U16289 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20988) );
  INV_X1 U16290 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n20963) );
  INV_X1 U16291 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20926) );
  INV_X1 U16292 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20912) );
  INV_X1 U16293 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20804) );
  INV_X1 U16294 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20780) );
  NAND4_X1 U16295 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .A4(P3_EBX_REG_11__SCAN_IN), .ZN(n14438)
         );
  INV_X1 U16296 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20753) );
  INV_X1 U16297 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n14436) );
  NAND3_X1 U16298 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n17754) );
  NOR3_X1 U16299 ( .A1(n14436), .A2(n20705), .A3(n17754), .ZN(n17753) );
  NAND3_X1 U16300 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17753), .ZN(n17775) );
  NOR2_X1 U16301 ( .A1(n20753), .A2(n17775), .ZN(n17774) );
  NAND4_X1 U16302 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n17774), .ZN(n14437) );
  NOR4_X1 U16303 ( .A1(n20804), .A2(n20780), .A3(n14438), .A4(n14437), .ZN(
        n18029) );
  NAND2_X1 U16304 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18029), .ZN(n18028) );
  NOR2_X1 U16305 ( .A1(n20912), .A2(n18028), .ZN(n18000) );
  NAND2_X1 U16306 ( .A1(n18039), .A2(n18000), .ZN(n18003) );
  NOR2_X1 U16307 ( .A1(n20926), .A2(n18003), .ZN(n18016) );
  NAND2_X1 U16308 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18016), .ZN(n17932) );
  NOR2_X1 U16309 ( .A1(n21197), .A2(n17932), .ZN(n17933) );
  NAND2_X1 U16310 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17933), .ZN(n17977) );
  NOR2_X1 U16311 ( .A1(n20963), .A2(n17977), .ZN(n17959) );
  NAND2_X1 U16312 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17959), .ZN(n17953) );
  NAND3_X1 U16313 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17958), .ZN(n17938) );
  NAND2_X1 U16314 ( .A1(n18034), .A2(n17938), .ZN(n17948) );
  OAI21_X1 U16315 ( .B1(n14439), .B2(n18035), .A(n17948), .ZN(n17942) );
  AOI22_X1 U16316 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14444) );
  AOI22_X1 U16317 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U16318 ( .A1(n18158), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U16319 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14441) );
  NAND4_X1 U16320 ( .A1(n14444), .A2(n14443), .A3(n14442), .A4(n14441), .ZN(
        n14450) );
  AOI22_X1 U16321 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U16322 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14447) );
  AOI22_X1 U16323 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U16324 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14445) );
  NAND4_X1 U16325 ( .A1(n14448), .A2(n14447), .A3(n14446), .A4(n14445), .ZN(
        n14449) );
  NOR2_X1 U16326 ( .A1(n14450), .A2(n14449), .ZN(n14514) );
  AOI22_X1 U16327 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U16328 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18156), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14453) );
  AOI22_X1 U16329 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14452) );
  AOI22_X1 U16330 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14451) );
  NAND4_X1 U16331 ( .A1(n14454), .A2(n14453), .A3(n14452), .A4(n14451), .ZN(
        n14461) );
  AOI22_X1 U16332 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U16333 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14458) );
  AOI22_X1 U16334 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14457) );
  AOI22_X1 U16335 ( .A1(n18116), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14456) );
  NAND4_X1 U16336 ( .A1(n14459), .A2(n14458), .A3(n14457), .A4(n14456), .ZN(
        n14460) );
  NOR2_X1 U16337 ( .A1(n14461), .A2(n14460), .ZN(n17946) );
  AOI22_X1 U16338 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18108), .ZN(n14465) );
  AOI22_X1 U16339 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14464) );
  AOI22_X1 U16340 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n18105), .ZN(n14463) );
  AOI22_X1 U16341 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18148), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n18082), .ZN(n14462) );
  NAND4_X1 U16342 ( .A1(n14465), .A2(n14464), .A3(n14463), .A4(n14462), .ZN(
        n14471) );
  AOI22_X1 U16343 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18127), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14469) );
  AOI22_X1 U16344 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18116), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14468) );
  AOI22_X1 U16345 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11174), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U16346 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18157), .ZN(n14466) );
  NAND4_X1 U16347 ( .A1(n14469), .A2(n14468), .A3(n14467), .A4(n14466), .ZN(
        n14470) );
  NOR2_X1 U16348 ( .A1(n14471), .A2(n14470), .ZN(n17955) );
  AOI22_X1 U16349 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U16350 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14481) );
  INV_X1 U16351 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U16352 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14473) );
  OAI21_X1 U16353 ( .B1(n17909), .B2(n17761), .A(n14473), .ZN(n14479) );
  AOI22_X1 U16354 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U16355 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U16356 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14475) );
  AOI22_X1 U16357 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14474) );
  NAND4_X1 U16358 ( .A1(n14477), .A2(n14476), .A3(n14475), .A4(n14474), .ZN(
        n14478) );
  AOI211_X1 U16359 ( .C1(n11175), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n14479), .B(n14478), .ZN(n14480) );
  NAND3_X1 U16360 ( .A1(n14482), .A2(n14481), .A3(n14480), .ZN(n17961) );
  AOI22_X1 U16361 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14388), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14493) );
  AOI22_X1 U16362 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U16363 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14483) );
  OAI21_X1 U16364 ( .B1(n11218), .B2(n18060), .A(n14483), .ZN(n14490) );
  AOI22_X1 U16365 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U16366 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U16367 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U16368 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14485) );
  NAND4_X1 U16369 ( .A1(n14488), .A2(n14487), .A3(n14486), .A4(n14485), .ZN(
        n14489) );
  AOI211_X1 U16370 ( .C1(n18128), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n14490), .B(n14489), .ZN(n14491) );
  NAND3_X1 U16371 ( .A1(n14493), .A2(n14492), .A3(n14491), .ZN(n17962) );
  NAND2_X1 U16372 ( .A1(n17961), .A2(n17962), .ZN(n17960) );
  NOR2_X1 U16373 ( .A1(n17955), .A2(n17960), .ZN(n17954) );
  AOI22_X1 U16374 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14503) );
  AOI22_X1 U16375 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U16376 ( .A1(n18116), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14494) );
  OAI21_X1 U16377 ( .B1(n17909), .B2(n18094), .A(n14494), .ZN(n14500) );
  AOI22_X1 U16378 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14498) );
  AOI22_X1 U16379 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14497) );
  AOI22_X1 U16380 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U16381 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14495) );
  NAND4_X1 U16382 ( .A1(n14498), .A2(n14497), .A3(n14496), .A4(n14495), .ZN(
        n14499) );
  AOI211_X1 U16383 ( .C1(n11176), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n14500), .B(n14499), .ZN(n14501) );
  NAND3_X1 U16384 ( .A1(n14503), .A2(n14502), .A3(n14501), .ZN(n17950) );
  NAND2_X1 U16385 ( .A1(n17954), .A2(n17950), .ZN(n17949) );
  NOR2_X1 U16386 ( .A1(n17946), .A2(n17949), .ZN(n17945) );
  AOI22_X1 U16387 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14388), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14513) );
  AOI22_X1 U16388 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14512) );
  INV_X1 U16389 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18115) );
  AOI22_X1 U16390 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14504) );
  OAI21_X1 U16391 ( .B1(n17909), .B2(n18115), .A(n14504), .ZN(n14510) );
  AOI22_X1 U16392 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18156), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14508) );
  AOI22_X1 U16393 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14507) );
  AOI22_X1 U16394 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U16395 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14505) );
  NAND4_X1 U16396 ( .A1(n14508), .A2(n14507), .A3(n14506), .A4(n14505), .ZN(
        n14509) );
  AOI211_X1 U16397 ( .C1(n18155), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n14510), .B(n14509), .ZN(n14511) );
  NAND3_X1 U16398 ( .A1(n14513), .A2(n14512), .A3(n14511), .ZN(n17936) );
  NAND2_X1 U16399 ( .A1(n17945), .A2(n17936), .ZN(n17935) );
  NOR2_X1 U16400 ( .A1(n14514), .A2(n17935), .ZN(n17941) );
  AOI21_X1 U16401 ( .B1(n14514), .B2(n17935), .A(n17941), .ZN(n21219) );
  AOI22_X1 U16402 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17942), .B1(n21219), 
        .B2(n18037), .ZN(n14517) );
  INV_X1 U16403 ( .A(n17938), .ZN(n14515) );
  NAND3_X1 U16404 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n21038), .A3(n14515), 
        .ZN(n14516) );
  NAND2_X1 U16405 ( .A1(n14517), .A2(n14516), .ZN(P3_U2675) );
  NAND2_X1 U16406 ( .A1(n15127), .A2(n15118), .ZN(n15388) );
  NAND2_X1 U16407 ( .A1(n16820), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15336) );
  INV_X1 U16408 ( .A(n15336), .ZN(n14518) );
  NAND2_X1 U16409 ( .A1(n14518), .A2(n22253), .ZN(n16823) );
  NOR2_X1 U16410 ( .A1(n15388), .A2(n16823), .ZN(n14519) );
  NAND2_X1 U16411 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15347), .ZN(
        n22285) );
  INV_X1 U16412 ( .A(n22285), .ZN(n14526) );
  OAI21_X1 U16413 ( .B1(n14519), .B2(n14526), .A(n15379), .ZN(n22588) );
  INV_X1 U16414 ( .A(n15353), .ZN(n14521) );
  OR2_X1 U16415 ( .A1(n16826), .A2(n14522), .ZN(n16852) );
  INV_X1 U16416 ( .A(n15349), .ZN(n14525) );
  NAND2_X1 U16417 ( .A1(n14524), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22425) );
  OAI21_X1 U16418 ( .B1(n16852), .B2(n14525), .A(n22425), .ZN(n14527) );
  AOI22_X1 U16419 ( .A1(n14527), .A2(n22253), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14526), .ZN(n22426) );
  AND2_X1 U16420 ( .A1(n16520), .A2(n15699), .ZN(n22454) );
  INV_X1 U16421 ( .A(n22454), .ZN(n16885) );
  OAI22_X1 U16422 ( .A1(n22235), .A2(n22459), .B1(n22426), .B2(n16885), .ZN(
        n14534) );
  INV_X1 U16423 ( .A(n15352), .ZN(n14528) );
  NAND2_X1 U16424 ( .A1(n11152), .A2(DATAI_29_), .ZN(n14530) );
  NAND2_X1 U16425 ( .A1(n22474), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14529) );
  AND2_X1 U16426 ( .A1(n14530), .A2(n14529), .ZN(n22442) );
  NOR2_X1 U16427 ( .A1(n22477), .A2(n14532), .ZN(n22455) );
  INV_X1 U16428 ( .A(n22455), .ZN(n22441) );
  OAI22_X1 U16429 ( .A1(n22591), .A2(n22442), .B1(n22441), .B2(n22425), .ZN(
        n14533) );
  AOI211_X1 U16430 ( .C1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .C2(n22588), .A(
        n14534), .B(n14533), .ZN(n14535) );
  INV_X1 U16431 ( .A(n14535), .ZN(P1_U3158) );
  AOI22_X2 U16432 ( .A1(DATAI_17_), .A2(n11152), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n22474), .ZN(n22330) );
  INV_X1 U16433 ( .A(n22325), .ZN(n16870) );
  OAI22_X1 U16434 ( .A1(n22235), .A2(n22330), .B1(n22426), .B2(n16870), .ZN(
        n14540) );
  NAND2_X1 U16435 ( .A1(n11152), .A2(DATAI_25_), .ZN(n14538) );
  NAND2_X1 U16436 ( .A1(n22474), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U16437 ( .A1(n14538), .A2(n14537), .ZN(n22327) );
  INV_X1 U16438 ( .A(n22327), .ZN(n22309) );
  NOR2_X1 U16439 ( .A1(n22477), .A2(n11828), .ZN(n22326) );
  INV_X1 U16440 ( .A(n22326), .ZN(n22308) );
  OAI22_X1 U16441 ( .A1(n22591), .A2(n22309), .B1(n22425), .B2(n22308), .ZN(
        n14539) );
  AOI211_X1 U16442 ( .C1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n22588), .A(
        n14540), .B(n14539), .ZN(n14541) );
  INV_X1 U16443 ( .A(n14541), .ZN(P1_U3154) );
  AND2_X1 U16444 ( .A1(n15699), .A2(n14542), .ZN(n22469) );
  OAI22_X1 U16445 ( .A1(n22235), .A2(n22473), .B1(n16892), .B2(n22426), .ZN(
        n14546) );
  NAND2_X1 U16446 ( .A1(n11152), .A2(DATAI_30_), .ZN(n14544) );
  NAND2_X1 U16447 ( .A1(n22474), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14543) );
  NAND2_X1 U16448 ( .A1(n14544), .A2(n14543), .ZN(n22470) );
  INV_X1 U16449 ( .A(n22470), .ZN(n15712) );
  NOR2_X1 U16450 ( .A1(n22477), .A2(n11571), .ZN(n22468) );
  INV_X1 U16451 ( .A(n22468), .ZN(n16889) );
  OAI22_X1 U16452 ( .A1(n22591), .A2(n15712), .B1(n22425), .B2(n16889), .ZN(
        n14545) );
  AOI211_X1 U16453 ( .C1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n22588), .A(
        n14546), .B(n14545), .ZN(n14547) );
  INV_X1 U16454 ( .A(n14547), .ZN(P1_U3159) );
  OAI222_X1 U16455 ( .A1(n15478), .A2(n14562), .B1(n16523), .B2(n11966), .C1(
        n16553), .C2(n14548), .ZN(P1_U2902) );
  OAI22_X1 U16456 ( .A1(n22235), .A2(n22302), .B1(n22426), .B2(n16865), .ZN(
        n14553) );
  NAND2_X1 U16457 ( .A1(n11152), .A2(DATAI_24_), .ZN(n14551) );
  NAND2_X1 U16458 ( .A1(n22474), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14550) );
  NAND2_X1 U16459 ( .A1(n14551), .A2(n14550), .ZN(n22299) );
  INV_X1 U16460 ( .A(n22299), .ZN(n22267) );
  NOR2_X1 U16461 ( .A1(n22477), .A2(n11829), .ZN(n22292) );
  OAI22_X1 U16462 ( .A1(n22591), .A2(n22267), .B1(n22425), .B2(n22266), .ZN(
        n14552) );
  AOI211_X1 U16463 ( .C1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .C2(n22588), .A(
        n14553), .B(n14552), .ZN(n14554) );
  INV_X1 U16464 ( .A(n14554), .ZN(P1_U3153) );
  NOR2_X1 U16465 ( .A1(n14555), .A2(n22479), .ZN(n22377) );
  INV_X1 U16466 ( .A(n22377), .ZN(n16880) );
  OAI22_X1 U16467 ( .A1(n22235), .A2(n22382), .B1(n22426), .B2(n16880), .ZN(
        n14560) );
  NAND2_X1 U16468 ( .A1(n11152), .A2(DATAI_27_), .ZN(n14557) );
  NAND2_X1 U16469 ( .A1(n22474), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14556) );
  NOR2_X1 U16470 ( .A1(n22477), .A2(n14558), .ZN(n22378) );
  OAI22_X1 U16471 ( .A1(n22591), .A2(n22371), .B1(n22425), .B2(n22370), .ZN(
        n14559) );
  AOI211_X1 U16472 ( .C1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .C2(n22588), .A(
        n14560), .B(n14559), .ZN(n14561) );
  INV_X1 U16473 ( .A(n14561), .ZN(P1_U3156) );
  INV_X1 U16474 ( .A(n22354), .ZN(n16875) );
  OAI22_X1 U16475 ( .A1(n22235), .A2(n22359), .B1(n22426), .B2(n16875), .ZN(
        n14567) );
  NAND2_X1 U16476 ( .A1(n11152), .A2(DATAI_26_), .ZN(n14564) );
  NAND2_X1 U16477 ( .A1(n22474), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14563) );
  NOR2_X1 U16478 ( .A1(n22477), .A2(n14565), .ZN(n22355) );
  OAI22_X1 U16479 ( .A1(n22591), .A2(n22342), .B1(n22425), .B2(n22341), .ZN(
        n14566) );
  AOI211_X1 U16480 ( .C1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .C2(n22588), .A(
        n14567), .B(n14566), .ZN(n14568) );
  INV_X1 U16481 ( .A(n14568), .ZN(P1_U3155) );
  NAND3_X1 U16482 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n17523), .ZN(n15720) );
  INV_X1 U16483 ( .A(n15720), .ZN(n14572) );
  INV_X1 U16484 ( .A(n14688), .ZN(n15120) );
  NAND2_X1 U16485 ( .A1(n15419), .A2(n16826), .ZN(n15719) );
  INV_X1 U16486 ( .A(n15719), .ZN(n22272) );
  NOR2_X1 U16487 ( .A1(n15376), .A2(n15720), .ZN(n22554) );
  AOI21_X1 U16488 ( .B1(n22272), .B2(n15349), .A(n22554), .ZN(n14571) );
  OAI211_X1 U16489 ( .C1(n15120), .C2(n15336), .A(n15381), .B(n14571), .ZN(
        n14570) );
  OAI211_X1 U16490 ( .C1(n15381), .C2(n14572), .A(n14570), .B(n15379), .ZN(
        n22557) );
  NAND2_X1 U16491 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14576) );
  INV_X1 U16492 ( .A(n22382), .ZN(n16876) );
  INV_X1 U16493 ( .A(n14571), .ZN(n14573) );
  AOI22_X1 U16494 ( .A1(n14573), .A2(n15381), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14572), .ZN(n22322) );
  INV_X1 U16495 ( .A(n22554), .ZN(n14583) );
  OAI22_X1 U16496 ( .A1(n22322), .A2(n16880), .B1(n22370), .B2(n14583), .ZN(
        n14574) );
  AOI21_X1 U16497 ( .B1(n22411), .B2(n16876), .A(n14574), .ZN(n14575) );
  OAI211_X1 U16498 ( .C1(n22371), .C2(n22553), .A(n14576), .B(n14575), .ZN(
        P1_U3124) );
  NAND2_X1 U16499 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14579) );
  INV_X1 U16500 ( .A(n22473), .ZN(n16886) );
  OAI22_X1 U16501 ( .A1(n16892), .A2(n22322), .B1(n16889), .B2(n14583), .ZN(
        n14577) );
  AOI21_X1 U16502 ( .B1(n22411), .B2(n16886), .A(n14577), .ZN(n14578) );
  OAI211_X1 U16503 ( .C1(n15712), .C2(n22553), .A(n14579), .B(n14578), .ZN(
        P1_U3127) );
  NAND2_X1 U16504 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14582) );
  INV_X1 U16505 ( .A(n22459), .ZN(n16881) );
  OAI22_X1 U16506 ( .A1(n22322), .A2(n16885), .B1(n22441), .B2(n14583), .ZN(
        n14580) );
  AOI21_X1 U16507 ( .B1(n22411), .B2(n16881), .A(n14580), .ZN(n14581) );
  OAI211_X1 U16508 ( .C1(n22442), .C2(n22553), .A(n14582), .B(n14581), .ZN(
        P1_U3126) );
  NAND2_X1 U16509 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14586) );
  INV_X1 U16510 ( .A(n22302), .ZN(n16861) );
  OAI22_X1 U16511 ( .A1(n22322), .A2(n16865), .B1(n22266), .B2(n14583), .ZN(
        n14584) );
  AOI21_X1 U16512 ( .B1(n22411), .B2(n16861), .A(n14584), .ZN(n14585) );
  OAI211_X1 U16513 ( .C1(n22267), .C2(n22553), .A(n14586), .B(n14585), .ZN(
        P1_U3121) );
  NOR2_X1 U16514 ( .A1(n14588), .A2(n15953), .ZN(n14591) );
  NAND2_X1 U16515 ( .A1(n14589), .A2(n14591), .ZN(n14590) );
  OAI22_X1 U16516 ( .A1(n14592), .A2(n14591), .B1(n13181), .B2(n14590), .ZN(
        n14596) );
  NOR2_X1 U16517 ( .A1(n14593), .A2(n12687), .ZN(n14594) );
  NAND2_X1 U16518 ( .A1(n13180), .A2(n14594), .ZN(n14595) );
  NAND2_X1 U16519 ( .A1(n14596), .A2(n14595), .ZN(n14597) );
  AOI21_X1 U16520 ( .B1(n15322), .B2(n14604), .A(n14597), .ZN(n17419) );
  NAND2_X1 U16521 ( .A1(n17419), .A2(n14601), .ZN(n14600) );
  INV_X1 U16522 ( .A(n14601), .ZN(n14656) );
  NAND2_X1 U16523 ( .A1(n14656), .A2(n14598), .ZN(n14599) );
  NAND2_X1 U16524 ( .A1(n14600), .A2(n14599), .ZN(n14660) );
  MUX2_X1 U16525 ( .A(n14603), .B(n14602), .S(n14601), .Z(n14659) );
  NAND2_X1 U16526 ( .A1(n14605), .A2(n14604), .ZN(n14613) );
  NAND2_X1 U16527 ( .A1(n14607), .A2(n14606), .ZN(n14616) );
  INV_X1 U16528 ( .A(n14608), .ZN(n14610) );
  INV_X1 U16529 ( .A(n12762), .ZN(n14609) );
  NAND2_X1 U16530 ( .A1(n14610), .A2(n14609), .ZN(n14611) );
  AOI22_X1 U16531 ( .A1(n13180), .A2(n11464), .B1(n14616), .B2(n14611), .ZN(
        n14612) );
  NAND2_X1 U16532 ( .A1(n14613), .A2(n14612), .ZN(n17415) );
  OR2_X1 U16533 ( .A1(n14615), .A2(n14614), .ZN(n14620) );
  INV_X1 U16534 ( .A(n13180), .ZN(n14618) );
  INV_X1 U16535 ( .A(n14616), .ZN(n14617) );
  NAND2_X1 U16536 ( .A1(n14620), .A2(n14619), .ZN(n19053) );
  OAI22_X1 U16537 ( .A1(n17415), .A2(n19807), .B1(n19819), .B2(n19053), .ZN(
        n14622) );
  NAND2_X1 U16538 ( .A1(n17415), .A2(n19807), .ZN(n14621) );
  AOI21_X1 U16539 ( .B1(n14622), .B2(n14621), .A(n14656), .ZN(n14624) );
  NAND2_X1 U16540 ( .A1(n14624), .A2(n19787), .ZN(n14623) );
  NAND2_X1 U16541 ( .A1(n14623), .A2(n14660), .ZN(n14627) );
  INV_X1 U16542 ( .A(n14624), .ZN(n14625) );
  NAND2_X1 U16543 ( .A1(n14625), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14626) );
  NAND2_X1 U16544 ( .A1(n14627), .A2(n14626), .ZN(n14628) );
  NAND2_X1 U16545 ( .A1(n14659), .A2(n14628), .ZN(n14631) );
  OR2_X1 U16546 ( .A1(n14628), .A2(n14659), .ZN(n14629) );
  AOI21_X1 U16547 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14629), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14630) );
  NAND2_X1 U16548 ( .A1(n14631), .A2(n14630), .ZN(n14658) );
  INV_X1 U16549 ( .A(n14632), .ZN(n14645) );
  INV_X1 U16550 ( .A(n14633), .ZN(n14640) );
  INV_X1 U16551 ( .A(n14634), .ZN(n14637) );
  AOI22_X1 U16552 ( .A1(n14638), .A2(n14637), .B1(n14636), .B2(n14635), .ZN(
        n14639) );
  OAI21_X1 U16553 ( .B1(n19156), .B2(n14640), .A(n14639), .ZN(n14641) );
  INV_X1 U16554 ( .A(n14641), .ZN(n14644) );
  NAND2_X1 U16555 ( .A1(n14646), .A2(n14642), .ZN(n14643) );
  OAI211_X1 U16556 ( .C1(n14646), .C2(n14645), .A(n14644), .B(n14643), .ZN(
        n19173) );
  NAND2_X1 U16557 ( .A1(n16097), .A2(n19059), .ZN(n14653) );
  OR2_X1 U16558 ( .A1(n15208), .A2(n14647), .ZN(n14648) );
  NOR2_X1 U16559 ( .A1(n14649), .A2(n14648), .ZN(n19172) );
  OAI21_X1 U16560 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19172), .ZN(n14652) );
  INV_X1 U16561 ( .A(n14650), .ZN(n14651) );
  OAI211_X1 U16562 ( .C1(n19062), .C2(n14653), .A(n14652), .B(n14651), .ZN(
        n14654) );
  OR2_X1 U16563 ( .A1(n19173), .A2(n14654), .ZN(n14655) );
  AOI21_X1 U16564 ( .B1(n14656), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n14655), .ZN(n14657) );
  OAI211_X1 U16565 ( .C1(n14660), .C2(n14659), .A(n14658), .B(n14657), .ZN(
        n19159) );
  NAND2_X1 U16566 ( .A1(n15237), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14662) );
  OAI21_X1 U16567 ( .B1(n19159), .B2(n14662), .A(n14661), .ZN(n14667) );
  NOR2_X1 U16568 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14663), .ZN(n15239) );
  INV_X1 U16569 ( .A(n15239), .ZN(n14664) );
  NOR2_X1 U16570 ( .A1(n18721), .A2(n14664), .ZN(n15231) );
  NAND2_X1 U16571 ( .A1(n14665), .A2(n15231), .ZN(n14666) );
  AND2_X1 U16572 ( .A1(n14667), .A2(n14666), .ZN(n19161) );
  OAI21_X1 U16573 ( .B1(n19161), .B2(n15635), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14668) );
  INV_X1 U16574 ( .A(n19157), .ZN(n17496) );
  NAND2_X1 U16575 ( .A1(n14668), .A2(n17496), .ZN(P2_U3593) );
  OR2_X1 U16576 ( .A1(n14671), .A2(n14670), .ZN(n14672) );
  AND2_X1 U16577 ( .A1(n14669), .A2(n14672), .ZN(n22031) );
  INV_X1 U16578 ( .A(n22031), .ZN(n14684) );
  AOI22_X1 U16579 ( .A1(n16551), .A2(n16520), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n16549), .ZN(n14673) );
  OAI21_X1 U16580 ( .B1(n14684), .B2(n16553), .A(n14673), .ZN(P1_U2899) );
  NAND2_X1 U16581 ( .A1(n16261), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14674) );
  OAI211_X1 U16582 ( .C1(n16209), .C2(P1_EBX_REG_5__SCAN_IN), .A(n14674), .B(
        n14072), .ZN(n14675) );
  OAI21_X1 U16583 ( .B1(n16199), .B2(P1_EBX_REG_5__SCAN_IN), .A(n14675), .ZN(
        n14682) );
  INV_X1 U16584 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n15588) );
  NAND2_X1 U16585 ( .A1(n14072), .A2(n21896), .ZN(n14679) );
  NAND2_X1 U16586 ( .A1(n16206), .A2(n15588), .ZN(n14678) );
  NAND3_X1 U16587 ( .A1(n14679), .A2(n16261), .A3(n14678), .ZN(n14680) );
  NAND2_X1 U16588 ( .A1(n14681), .A2(n14680), .ZN(n15103) );
  AOI21_X1 U16589 ( .B1(n14682), .B2(n15104), .A(n15331), .ZN(n22025) );
  AOI22_X1 U16590 ( .A1(n16463), .A2(n22025), .B1(n16462), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n14683) );
  OAI21_X1 U16591 ( .B1(n14684), .B2(n16425), .A(n14683), .ZN(P1_U2867) );
  NAND3_X1 U16592 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17523), .A3(
        n17517), .ZN(n22271) );
  INV_X1 U16593 ( .A(n22271), .ZN(n14689) );
  OR2_X1 U16594 ( .A1(n16820), .A2(n22256), .ZN(n15164) );
  NOR2_X1 U16595 ( .A1(n15376), .A2(n22271), .ZN(n22541) );
  INV_X1 U16596 ( .A(n22541), .ZN(n14706) );
  OAI21_X1 U16597 ( .B1(n15719), .B2(n15377), .A(n14706), .ZN(n14690) );
  INV_X1 U16598 ( .A(n14690), .ZN(n14685) );
  OAI211_X1 U16599 ( .C1(n15120), .C2(n15164), .A(n15381), .B(n14685), .ZN(
        n14686) );
  OAI211_X1 U16600 ( .C1(n22253), .C2(n14689), .A(n15379), .B(n14686), .ZN(
        n22543) );
  NAND2_X1 U16601 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n14693) );
  INV_X1 U16602 ( .A(n22330), .ZN(n16866) );
  AOI22_X1 U16603 ( .A1(n14690), .A2(n15381), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14689), .ZN(n22406) );
  OAI22_X1 U16604 ( .A1(n22308), .A2(n14706), .B1(n22406), .B2(n16870), .ZN(
        n14691) );
  AOI21_X1 U16605 ( .B1(n22548), .B2(n16866), .A(n14691), .ZN(n14692) );
  OAI211_X1 U16606 ( .C1(n22309), .C2(n22546), .A(n14693), .B(n14692), .ZN(
        P1_U3106) );
  NAND2_X1 U16607 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n14696) );
  OAI22_X1 U16608 ( .A1(n22266), .A2(n14706), .B1(n22406), .B2(n16865), .ZN(
        n14694) );
  AOI21_X1 U16609 ( .B1(n22548), .B2(n16861), .A(n14694), .ZN(n14695) );
  OAI211_X1 U16610 ( .C1(n22267), .C2(n22546), .A(n14696), .B(n14695), .ZN(
        P1_U3105) );
  NAND2_X1 U16611 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14699) );
  INV_X1 U16612 ( .A(n22359), .ZN(n16871) );
  OAI22_X1 U16613 ( .A1(n22341), .A2(n14706), .B1(n22406), .B2(n16875), .ZN(
        n14697) );
  AOI21_X1 U16614 ( .B1(n22548), .B2(n16871), .A(n14697), .ZN(n14698) );
  OAI211_X1 U16615 ( .C1(n22342), .C2(n22546), .A(n14699), .B(n14698), .ZN(
        P1_U3107) );
  NAND2_X1 U16616 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n14702) );
  OAI22_X1 U16617 ( .A1(n22441), .A2(n14706), .B1(n22406), .B2(n16885), .ZN(
        n14700) );
  AOI21_X1 U16618 ( .B1(n22548), .B2(n16881), .A(n14700), .ZN(n14701) );
  OAI211_X1 U16619 ( .C1(n22442), .C2(n22546), .A(n14702), .B(n14701), .ZN(
        P1_U3110) );
  NAND2_X1 U16620 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n14705) );
  OAI22_X1 U16621 ( .A1(n16892), .A2(n22406), .B1(n16889), .B2(n14706), .ZN(
        n14703) );
  AOI21_X1 U16622 ( .B1(n22548), .B2(n16886), .A(n14703), .ZN(n14704) );
  OAI211_X1 U16623 ( .C1(n15712), .C2(n22546), .A(n14705), .B(n14704), .ZN(
        P1_U3111) );
  NAND2_X1 U16624 ( .A1(n22543), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n14709) );
  OAI22_X1 U16625 ( .A1(n22370), .A2(n14706), .B1(n22406), .B2(n16880), .ZN(
        n14707) );
  AOI21_X1 U16626 ( .B1(n22548), .B2(n16876), .A(n14707), .ZN(n14708) );
  OAI211_X1 U16627 ( .C1(n22371), .C2(n22546), .A(n14709), .B(n14708), .ZN(
        P1_U3108) );
  XOR2_X1 U16628 ( .A(keyinput_127), .B(keyinput_255), .Z(n15078) );
  XOR2_X1 U16629 ( .A(DATAI_30_), .B(keyinput_130), .Z(n14713) );
  XOR2_X1 U16630 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_128), .Z(n14712) );
  INV_X1 U16631 ( .A(DATAI_31_), .ZN(n16467) );
  XNOR2_X1 U16632 ( .A(n16467), .B(keyinput_129), .ZN(n14711) );
  XNOR2_X1 U16633 ( .A(DATAI_29_), .B(keyinput_131), .ZN(n14710) );
  NAND4_X1 U16634 ( .A1(n14713), .A2(n14712), .A3(n14711), .A4(n14710), .ZN(
        n14716) );
  INV_X1 U16635 ( .A(DATAI_28_), .ZN(n16473) );
  XNOR2_X1 U16636 ( .A(n16473), .B(keyinput_132), .ZN(n14715) );
  XOR2_X1 U16637 ( .A(DATAI_27_), .B(keyinput_133), .Z(n14714) );
  AOI21_X1 U16638 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(n14724) );
  XOR2_X1 U16639 ( .A(DATAI_23_), .B(keyinput_137), .Z(n14720) );
  INV_X1 U16640 ( .A(DATAI_22_), .ZN(n16512) );
  XNOR2_X1 U16641 ( .A(n16512), .B(keyinput_138), .ZN(n14719) );
  XNOR2_X1 U16642 ( .A(DATAI_26_), .B(keyinput_134), .ZN(n14718) );
  XNOR2_X1 U16643 ( .A(DATAI_21_), .B(keyinput_139), .ZN(n14717) );
  NAND4_X1 U16644 ( .A1(n14720), .A2(n14719), .A3(n14718), .A4(n14717), .ZN(
        n14723) );
  XNOR2_X1 U16645 ( .A(DATAI_25_), .B(keyinput_135), .ZN(n14722) );
  XNOR2_X1 U16646 ( .A(DATAI_24_), .B(keyinput_136), .ZN(n14721) );
  NOR4_X1 U16647 ( .A1(n14724), .A2(n14723), .A3(n14722), .A4(n14721), .ZN(
        n14727) );
  INV_X1 U16648 ( .A(DATAI_20_), .ZN(n16525) );
  XNOR2_X1 U16649 ( .A(n16525), .B(keyinput_140), .ZN(n14726) );
  XNOR2_X1 U16650 ( .A(DATAI_19_), .B(keyinput_141), .ZN(n14725) );
  OAI21_X1 U16651 ( .B1(n14727), .B2(n14726), .A(n14725), .ZN(n14730) );
  XNOR2_X1 U16652 ( .A(DATAI_18_), .B(keyinput_142), .ZN(n14729) );
  XOR2_X1 U16653 ( .A(DATAI_17_), .B(keyinput_143), .Z(n14728) );
  AOI21_X1 U16654 ( .B1(n14730), .B2(n14729), .A(n14728), .ZN(n14736) );
  XNOR2_X1 U16655 ( .A(DATAI_16_), .B(keyinput_144), .ZN(n14735) );
  XNOR2_X1 U16656 ( .A(DATAI_15_), .B(keyinput_145), .ZN(n14733) );
  XNOR2_X1 U16657 ( .A(DATAI_13_), .B(keyinput_147), .ZN(n14732) );
  XNOR2_X1 U16658 ( .A(DATAI_14_), .B(keyinput_146), .ZN(n14731) );
  NOR3_X1 U16659 ( .A1(n14733), .A2(n14732), .A3(n14731), .ZN(n14734) );
  OAI21_X1 U16660 ( .B1(n14736), .B2(n14735), .A(n14734), .ZN(n14746) );
  XOR2_X1 U16661 ( .A(DATAI_12_), .B(keyinput_148), .Z(n14745) );
  INV_X1 U16662 ( .A(DATAI_9_), .ZN(n14738) );
  OAI22_X1 U16663 ( .A1(n14738), .A2(keyinput_151), .B1(DATAI_11_), .B2(
        keyinput_149), .ZN(n14737) );
  AOI221_X1 U16664 ( .B1(n14738), .B2(keyinput_151), .C1(keyinput_149), .C2(
        DATAI_11_), .A(n14737), .ZN(n14743) );
  XNOR2_X1 U16665 ( .A(keyinput_152), .B(DATAI_8_), .ZN(n14742) );
  INV_X1 U16666 ( .A(keyinput_153), .ZN(n14739) );
  XNOR2_X1 U16667 ( .A(n14739), .B(DATAI_7_), .ZN(n14741) );
  XNOR2_X1 U16668 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n14740) );
  NAND4_X1 U16669 ( .A1(n14743), .A2(n14742), .A3(n14741), .A4(n14740), .ZN(
        n14744) );
  AOI21_X1 U16670 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(n14749) );
  XOR2_X1 U16671 ( .A(DATAI_6_), .B(keyinput_154), .Z(n14748) );
  XOR2_X1 U16672 ( .A(DATAI_5_), .B(keyinput_155), .Z(n14747) );
  OAI21_X1 U16673 ( .B1(n14749), .B2(n14748), .A(n14747), .ZN(n14752) );
  XOR2_X1 U16674 ( .A(DATAI_4_), .B(keyinput_156), .Z(n14751) );
  XNOR2_X1 U16675 ( .A(DATAI_3_), .B(keyinput_157), .ZN(n14750) );
  AOI21_X1 U16676 ( .B1(n14752), .B2(n14751), .A(n14750), .ZN(n14755) );
  XOR2_X1 U16677 ( .A(DATAI_2_), .B(keyinput_158), .Z(n14754) );
  XNOR2_X1 U16678 ( .A(keyinput_159), .B(DATAI_1_), .ZN(n14753) );
  OAI21_X1 U16679 ( .B1(n14755), .B2(n14754), .A(n14753), .ZN(n14758) );
  XOR2_X1 U16680 ( .A(keyinput_161), .B(HOLD), .Z(n14757) );
  XOR2_X1 U16681 ( .A(keyinput_160), .B(DATAI_0_), .Z(n14756) );
  NAND3_X1 U16682 ( .A1(n14758), .A2(n14757), .A3(n14756), .ZN(n14761) );
  XNOR2_X1 U16683 ( .A(keyinput_162), .B(NA), .ZN(n14760) );
  XOR2_X1 U16684 ( .A(keyinput_163), .B(BS16), .Z(n14759) );
  AOI21_X1 U16685 ( .B1(n14761), .B2(n14760), .A(n14759), .ZN(n14764) );
  XOR2_X1 U16686 ( .A(READY1), .B(keyinput_164), .Z(n14763) );
  XOR2_X1 U16687 ( .A(READY2), .B(keyinput_165), .Z(n14762) );
  OAI21_X1 U16688 ( .B1(n14764), .B2(n14763), .A(n14762), .ZN(n14770) );
  INV_X1 U16689 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20530) );
  OAI22_X1 U16690 ( .A1(n20530), .A2(keyinput_170), .B1(P1_M_IO_N_REG_SCAN_IN), 
        .B2(keyinput_169), .ZN(n14765) );
  AOI221_X1 U16691 ( .B1(n20530), .B2(keyinput_170), .C1(keyinput_169), .C2(
        P1_M_IO_N_REG_SCAN_IN), .A(n14765), .ZN(n14769) );
  XOR2_X1 U16692 ( .A(keyinput_166), .B(P1_READREQUEST_REG_SCAN_IN), .Z(n14768) );
  INV_X1 U16693 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17557) );
  OAI22_X1 U16694 ( .A1(n17557), .A2(keyinput_167), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_168), .ZN(n14766) );
  AOI221_X1 U16695 ( .B1(n17557), .B2(keyinput_167), .C1(keyinput_168), .C2(
        P1_CODEFETCH_REG_SCAN_IN), .A(n14766), .ZN(n14767) );
  NAND4_X1 U16696 ( .A1(n14770), .A2(n14769), .A3(n14768), .A4(n14767), .ZN(
        n14773) );
  XOR2_X1 U16697 ( .A(keyinput_171), .B(P1_REQUESTPENDING_REG_SCAN_IN), .Z(
        n14772) );
  XNOR2_X1 U16698 ( .A(P1_STATEBS16_REG_SCAN_IN), .B(keyinput_172), .ZN(n14771) );
  AOI21_X1 U16699 ( .B1(n14773), .B2(n14772), .A(n14771), .ZN(n14779) );
  XNOR2_X1 U16700 ( .A(keyinput_175), .B(P1_W_R_N_REG_SCAN_IN), .ZN(n14776) );
  XNOR2_X1 U16701 ( .A(keyinput_174), .B(P1_FLUSH_REG_SCAN_IN), .ZN(n14775) );
  XNOR2_X1 U16702 ( .A(keyinput_173), .B(P1_MORE_REG_SCAN_IN), .ZN(n14774) );
  NAND3_X1 U16703 ( .A1(n14776), .A2(n14775), .A3(n14774), .ZN(n14778) );
  XOR2_X1 U16704 ( .A(keyinput_176), .B(P1_BYTEENABLE_REG_0__SCAN_IN), .Z(
        n14777) );
  OAI21_X1 U16705 ( .B1(n14779), .B2(n14778), .A(n14777), .ZN(n14783) );
  XOR2_X1 U16706 ( .A(keyinput_177), .B(P1_BYTEENABLE_REG_1__SCAN_IN), .Z(
        n14782) );
  XOR2_X1 U16707 ( .A(keyinput_179), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .Z(
        n14781) );
  XNOR2_X1 U16708 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_178), .ZN(
        n14780) );
  AOI211_X1 U16709 ( .C1(n14783), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        n14790) );
  XOR2_X1 U16710 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_183), .Z(n14787)
         );
  XOR2_X1 U16711 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_182), .Z(n14786)
         );
  INV_X1 U16712 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20435) );
  XNOR2_X1 U16713 ( .A(n20435), .B(keyinput_180), .ZN(n14785) );
  XNOR2_X1 U16714 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .ZN(n14784)
         );
  NAND4_X1 U16715 ( .A1(n14787), .A2(n14786), .A3(n14785), .A4(n14784), .ZN(
        n14789) );
  XOR2_X1 U16716 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_184), .Z(n14788)
         );
  OAI21_X1 U16717 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14797) );
  XOR2_X1 U16718 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_186), .Z(n14793)
         );
  XOR2_X1 U16719 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_187), .Z(n14792)
         );
  XNOR2_X1 U16720 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_189), .ZN(n14791)
         );
  NOR3_X1 U16721 ( .A1(n14793), .A2(n14792), .A3(n14791), .ZN(n14796) );
  XNOR2_X1 U16722 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_185), .ZN(n14795)
         );
  XNOR2_X1 U16723 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_188), .ZN(n14794)
         );
  NAND4_X1 U16724 ( .A1(n14797), .A2(n14796), .A3(n14795), .A4(n14794), .ZN(
        n14800) );
  XOR2_X1 U16725 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_191), .Z(n14799)
         );
  INV_X1 U16726 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n22123) );
  XNOR2_X1 U16727 ( .A(n22123), .B(keyinput_190), .ZN(n14798) );
  NAND3_X1 U16728 ( .A1(n14800), .A2(n14799), .A3(n14798), .ZN(n14814) );
  AOI22_X1 U16729 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_195), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(keyinput_193), .ZN(n14813) );
  INV_X1 U16730 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20407) );
  AOI22_X1 U16731 ( .A1(n20407), .A2(keyinput_197), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_194), .ZN(n14812) );
  INV_X1 U16732 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21853) );
  INV_X1 U16733 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n22000) );
  INV_X1 U16734 ( .A(keyinput_192), .ZN(n14806) );
  OAI22_X1 U16735 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_195), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(keyinput_193), .ZN(n14804) );
  OAI22_X1 U16736 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_192), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_194), .ZN(n14803) );
  INV_X1 U16737 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20404) );
  OAI22_X1 U16738 ( .A1(n20404), .A2(keyinput_199), .B1(n20407), .B2(
        keyinput_197), .ZN(n14802) );
  INV_X1 U16739 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20408) );
  OAI22_X1 U16740 ( .A1(n20408), .A2(keyinput_196), .B1(n21853), .B2(
        keyinput_198), .ZN(n14801) );
  NOR4_X1 U16741 ( .A1(n14804), .A2(n14803), .A3(n14802), .A4(n14801), .ZN(
        n14805) );
  OAI21_X1 U16742 ( .B1(n22000), .B2(n14806), .A(n14805), .ZN(n14810) );
  INV_X1 U16743 ( .A(keyinput_199), .ZN(n14808) );
  INV_X1 U16744 ( .A(keyinput_196), .ZN(n14807) );
  OAI22_X1 U16745 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n14808), .B1(n14807), 
        .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14809) );
  AOI211_X1 U16746 ( .C1(keyinput_198), .C2(n21853), .A(n14810), .B(n14809), 
        .ZN(n14811) );
  NAND4_X1 U16747 ( .A1(n14814), .A2(n14813), .A3(n14812), .A4(n14811), .ZN(
        n14818) );
  XOR2_X1 U16748 ( .A(keyinput_200), .B(P1_REIP_REG_11__SCAN_IN), .Z(n14817)
         );
  XOR2_X1 U16749 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_202), .Z(n14816) );
  XNOR2_X1 U16750 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_201), .ZN(n14815)
         );
  AOI211_X1 U16751 ( .C1(n14818), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        n14821) );
  XNOR2_X1 U16752 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_203), .ZN(n14820)
         );
  XOR2_X1 U16753 ( .A(keyinput_204), .B(P1_REIP_REG_7__SCAN_IN), .Z(n14819) );
  OAI21_X1 U16754 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n14824) );
  XNOR2_X1 U16755 ( .A(keyinput_205), .B(P1_REIP_REG_6__SCAN_IN), .ZN(n14823)
         );
  XOR2_X1 U16756 ( .A(keyinput_206), .B(P1_REIP_REG_5__SCAN_IN), .Z(n14822) );
  AOI21_X1 U16757 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n14835) );
  XOR2_X1 U16758 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_211), .Z(n14828) );
  XOR2_X1 U16759 ( .A(keyinput_210), .B(P1_REIP_REG_1__SCAN_IN), .Z(n14827) );
  XNOR2_X1 U16760 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_208), .ZN(n14826)
         );
  XNOR2_X1 U16761 ( .A(keyinput_207), .B(P1_REIP_REG_4__SCAN_IN), .ZN(n14825)
         );
  NOR4_X1 U16762 ( .A1(n14828), .A2(n14827), .A3(n14826), .A4(n14825), .ZN(
        n14831) );
  XOR2_X1 U16763 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .Z(n14830) );
  XOR2_X1 U16764 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_209), .Z(n14829) );
  NAND3_X1 U16765 ( .A1(n14831), .A2(n14830), .A3(n14829), .ZN(n14834) );
  INV_X1 U16766 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16419) );
  XNOR2_X1 U16767 ( .A(n16419), .B(keyinput_214), .ZN(n14833) );
  XNOR2_X1 U16768 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n14832)
         );
  OAI211_X1 U16769 ( .C1(n14835), .C2(n14834), .A(n14833), .B(n14832), .ZN(
        n14839) );
  INV_X1 U16770 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16422) );
  XNOR2_X1 U16771 ( .A(n16422), .B(keyinput_217), .ZN(n14838) );
  XNOR2_X1 U16772 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_216), .ZN(n14837)
         );
  XNOR2_X1 U16773 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_215), .ZN(n14836)
         );
  NAND4_X1 U16774 ( .A1(n14839), .A2(n14838), .A3(n14837), .A4(n14836), .ZN(
        n14841) );
  XOR2_X1 U16775 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_218), .Z(n14840) );
  NAND2_X1 U16776 ( .A1(n14841), .A2(n14840), .ZN(n14845) );
  XOR2_X1 U16777 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_220), .Z(n14844) );
  XNOR2_X1 U16778 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_221), .ZN(n14843)
         );
  XNOR2_X1 U16779 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_219), .ZN(n14842)
         );
  NAND4_X1 U16780 ( .A1(n14845), .A2(n14844), .A3(n14843), .A4(n14842), .ZN(
        n14848) );
  XNOR2_X1 U16781 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_222), .ZN(n14847)
         );
  XNOR2_X1 U16782 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_223), .ZN(n14846)
         );
  AOI21_X1 U16783 ( .B1(n14848), .B2(n14847), .A(n14846), .ZN(n14855) );
  XOR2_X1 U16784 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_226), .Z(n14852) );
  INV_X1 U16785 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16448) );
  XNOR2_X1 U16786 ( .A(n16448), .B(keyinput_225), .ZN(n14851) );
  XNOR2_X1 U16787 ( .A(keyinput_227), .B(P1_EBX_REG_16__SCAN_IN), .ZN(n14850)
         );
  XNOR2_X1 U16788 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_224), .ZN(n14849)
         );
  NAND4_X1 U16789 ( .A1(n14852), .A2(n14851), .A3(n14850), .A4(n14849), .ZN(
        n14854) );
  XOR2_X1 U16790 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_228), .Z(n14853) );
  OAI21_X1 U16791 ( .B1(n14855), .B2(n14854), .A(n14853), .ZN(n14858) );
  XNOR2_X1 U16792 ( .A(keyinput_229), .B(P1_EBX_REG_14__SCAN_IN), .ZN(n14857)
         );
  XOR2_X1 U16793 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_230), .Z(n14856) );
  AOI21_X1 U16794 ( .B1(n14858), .B2(n14857), .A(n14856), .ZN(n14862) );
  XOR2_X1 U16795 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_232), .Z(n14861) );
  INV_X1 U16796 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15695) );
  XNOR2_X1 U16797 ( .A(n15695), .B(keyinput_233), .ZN(n14860) );
  INV_X1 U16798 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n22078) );
  XNOR2_X1 U16799 ( .A(n22078), .B(keyinput_231), .ZN(n14859) );
  NOR4_X1 U16800 ( .A1(n14862), .A2(n14861), .A3(n14860), .A4(n14859), .ZN(
        n14866) );
  XOR2_X1 U16801 ( .A(keyinput_234), .B(P1_EBX_REG_9__SCAN_IN), .Z(n14865) );
  XOR2_X1 U16802 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .Z(n14864) );
  XOR2_X1 U16803 ( .A(keyinput_236), .B(P1_EBX_REG_7__SCAN_IN), .Z(n14863) );
  OAI211_X1 U16804 ( .C1(n14866), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        n14869) );
  XNOR2_X1 U16805 ( .A(keyinput_237), .B(P1_EBX_REG_6__SCAN_IN), .ZN(n14868)
         );
  XNOR2_X1 U16806 ( .A(keyinput_238), .B(P1_EBX_REG_5__SCAN_IN), .ZN(n14867)
         );
  AOI21_X1 U16807 ( .B1(n14869), .B2(n14868), .A(n14867), .ZN(n14873) );
  XOR2_X1 U16808 ( .A(keyinput_241), .B(P1_EBX_REG_2__SCAN_IN), .Z(n14872) );
  XNOR2_X1 U16809 ( .A(keyinput_239), .B(P1_EBX_REG_4__SCAN_IN), .ZN(n14871)
         );
  XNOR2_X1 U16810 ( .A(keyinput_240), .B(P1_EBX_REG_3__SCAN_IN), .ZN(n14870)
         );
  NOR4_X1 U16811 ( .A1(n14873), .A2(n14872), .A3(n14871), .A4(n14870), .ZN(
        n14876) );
  XOR2_X1 U16812 ( .A(keyinput_243), .B(P1_EBX_REG_0__SCAN_IN), .Z(n14875) );
  XNOR2_X1 U16813 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_242), .ZN(n14874)
         );
  NOR3_X1 U16814 ( .A1(n14876), .A2(n14875), .A3(n14874), .ZN(n14879) );
  XNOR2_X1 U16815 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .ZN(n14878)
         );
  XNOR2_X1 U16816 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n14877)
         );
  NOR3_X1 U16817 ( .A1(n14879), .A2(n14878), .A3(n14877), .ZN(n14893) );
  XNOR2_X1 U16818 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .ZN(n14892)
         );
  OAI22_X1 U16819 ( .A1(keyinput_249), .A2(n16486), .B1(n16479), .B2(
        keyinput_248), .ZN(n14890) );
  INV_X1 U16820 ( .A(keyinput_247), .ZN(n14885) );
  AOI22_X1 U16821 ( .A1(n16479), .A2(keyinput_248), .B1(keyinput_252), .B2(
        n16505), .ZN(n14883) );
  AOI22_X1 U16822 ( .A1(n16511), .A2(keyinput_253), .B1(keyinput_249), .B2(
        n16486), .ZN(n14882) );
  AOI22_X1 U16823 ( .A1(keyinput_250), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n16499), .B2(keyinput_251), .ZN(n14881) );
  AOI22_X1 U16824 ( .A1(P1_EAX_REG_28__SCAN_IN), .A2(keyinput_247), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_254), .ZN(n14880) );
  NAND4_X1 U16825 ( .A1(n14883), .A2(n14882), .A3(n14881), .A4(n14880), .ZN(
        n14884) );
  AOI21_X1 U16826 ( .B1(n16472), .B2(n14885), .A(n14884), .ZN(n14886) );
  OAI21_X1 U16827 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput_254), .A(n14886), 
        .ZN(n14889) );
  OAI22_X1 U16828 ( .A1(keyinput_251), .A2(n16499), .B1(n16511), .B2(
        keyinput_253), .ZN(n14888) );
  OAI22_X1 U16829 ( .A1(n16505), .A2(keyinput_252), .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_250), .ZN(n14887) );
  NOR4_X1 U16830 ( .A1(n14890), .A2(n14889), .A3(n14888), .A4(n14887), .ZN(
        n14891) );
  OAI21_X1 U16831 ( .B1(n14893), .B2(n14892), .A(n14891), .ZN(n15077) );
  XOR2_X1 U16832 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_127), .Z(n15076) );
  XOR2_X1 U16833 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_0), .Z(n14897)
         );
  XNOR2_X1 U16834 ( .A(n16467), .B(keyinput_1), .ZN(n14896) );
  XNOR2_X1 U16835 ( .A(DATAI_29_), .B(keyinput_3), .ZN(n14895) );
  XNOR2_X1 U16836 ( .A(DATAI_30_), .B(keyinput_2), .ZN(n14894) );
  NAND4_X1 U16837 ( .A1(n14897), .A2(n14896), .A3(n14895), .A4(n14894), .ZN(
        n14900) );
  XNOR2_X1 U16838 ( .A(n16473), .B(keyinput_4), .ZN(n14899) );
  XOR2_X1 U16839 ( .A(DATAI_27_), .B(keyinput_5), .Z(n14898) );
  AOI21_X1 U16840 ( .B1(n14900), .B2(n14899), .A(n14898), .ZN(n14908) );
  XOR2_X1 U16841 ( .A(DATAI_25_), .B(keyinput_7), .Z(n14907) );
  XNOR2_X1 U16842 ( .A(DATAI_23_), .B(keyinput_9), .ZN(n14906) );
  XNOR2_X1 U16843 ( .A(DATAI_24_), .B(keyinput_8), .ZN(n14904) );
  XNOR2_X1 U16844 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n14903) );
  XNOR2_X1 U16845 ( .A(DATAI_21_), .B(keyinput_11), .ZN(n14902) );
  XNOR2_X1 U16846 ( .A(DATAI_22_), .B(keyinput_10), .ZN(n14901) );
  NAND4_X1 U16847 ( .A1(n14904), .A2(n14903), .A3(n14902), .A4(n14901), .ZN(
        n14905) );
  NOR4_X1 U16848 ( .A1(n14908), .A2(n14907), .A3(n14906), .A4(n14905), .ZN(
        n14911) );
  XNOR2_X1 U16849 ( .A(n16525), .B(keyinput_12), .ZN(n14910) );
  XNOR2_X1 U16850 ( .A(DATAI_19_), .B(keyinput_13), .ZN(n14909) );
  OAI21_X1 U16851 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(n14914) );
  XOR2_X1 U16852 ( .A(DATAI_18_), .B(keyinput_14), .Z(n14913) );
  XNOR2_X1 U16853 ( .A(DATAI_17_), .B(keyinput_15), .ZN(n14912) );
  AOI21_X1 U16854 ( .B1(n14914), .B2(n14913), .A(n14912), .ZN(n14916) );
  XOR2_X1 U16855 ( .A(DATAI_16_), .B(keyinput_16), .Z(n14915) );
  NOR2_X1 U16856 ( .A1(n14916), .A2(n14915), .ZN(n14921) );
  XOR2_X1 U16857 ( .A(DATAI_13_), .B(keyinput_19), .Z(n14920) );
  XOR2_X1 U16858 ( .A(DATAI_14_), .B(keyinput_18), .Z(n14919) );
  XNOR2_X1 U16859 ( .A(n14917), .B(keyinput_17), .ZN(n14918) );
  NOR4_X1 U16860 ( .A1(n14921), .A2(n14920), .A3(n14919), .A4(n14918), .ZN(
        n14930) );
  XOR2_X1 U16861 ( .A(DATAI_12_), .B(keyinput_20), .Z(n14929) );
  XOR2_X1 U16862 ( .A(DATAI_8_), .B(keyinput_24), .Z(n14924) );
  XNOR2_X1 U16863 ( .A(DATAI_11_), .B(keyinput_21), .ZN(n14923) );
  XNOR2_X1 U16864 ( .A(DATAI_7_), .B(keyinput_25), .ZN(n14922) );
  NAND3_X1 U16865 ( .A1(n14924), .A2(n14923), .A3(n14922), .ZN(n14927) );
  XOR2_X1 U16866 ( .A(DATAI_10_), .B(keyinput_22), .Z(n14926) );
  XNOR2_X1 U16867 ( .A(DATAI_9_), .B(keyinput_23), .ZN(n14925) );
  NOR3_X1 U16868 ( .A1(n14927), .A2(n14926), .A3(n14925), .ZN(n14928) );
  OAI21_X1 U16869 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(n14933) );
  XNOR2_X1 U16870 ( .A(DATAI_6_), .B(keyinput_26), .ZN(n14932) );
  XOR2_X1 U16871 ( .A(DATAI_5_), .B(keyinput_27), .Z(n14931) );
  AOI21_X1 U16872 ( .B1(n14933), .B2(n14932), .A(n14931), .ZN(n14936) );
  XNOR2_X1 U16873 ( .A(DATAI_4_), .B(keyinput_28), .ZN(n14935) );
  XOR2_X1 U16874 ( .A(DATAI_3_), .B(keyinput_29), .Z(n14934) );
  OAI21_X1 U16875 ( .B1(n14936), .B2(n14935), .A(n14934), .ZN(n14939) );
  XNOR2_X1 U16876 ( .A(DATAI_2_), .B(keyinput_30), .ZN(n14938) );
  XNOR2_X1 U16877 ( .A(DATAI_1_), .B(keyinput_31), .ZN(n14937) );
  AOI21_X1 U16878 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(n14942) );
  XOR2_X1 U16879 ( .A(DATAI_0_), .B(keyinput_32), .Z(n14941) );
  XOR2_X1 U16880 ( .A(HOLD), .B(keyinput_33), .Z(n14940) );
  NOR3_X1 U16881 ( .A1(n14942), .A2(n14941), .A3(n14940), .ZN(n14945) );
  XNOR2_X1 U16882 ( .A(NA), .B(keyinput_34), .ZN(n14944) );
  XOR2_X1 U16883 ( .A(BS16), .B(keyinput_35), .Z(n14943) );
  OAI21_X1 U16884 ( .B1(n14945), .B2(n14944), .A(n14943), .ZN(n14948) );
  XOR2_X1 U16885 ( .A(READY1), .B(keyinput_36), .Z(n14947) );
  XNOR2_X1 U16886 ( .A(READY2), .B(keyinput_37), .ZN(n14946) );
  AOI21_X1 U16887 ( .B1(n14948), .B2(n14947), .A(n14946), .ZN(n14954) );
  AOI22_X1 U16888 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_42), .B1(n22594), 
        .B2(keyinput_41), .ZN(n14949) );
  OAI221_X1 U16889 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_42), .C1(n22594), 
        .C2(keyinput_41), .A(n14949), .ZN(n14953) );
  AOI22_X1 U16890 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_40), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_38), .ZN(n14950) );
  OAI221_X1 U16891 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_40), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_38), .A(n14950), .ZN(n14952)
         );
  XNOR2_X1 U16892 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_39), .ZN(n14951) );
  NOR4_X1 U16893 ( .A1(n14954), .A2(n14953), .A3(n14952), .A4(n14951), .ZN(
        n14957) );
  XOR2_X1 U16894 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_43), .Z(
        n14956) );
  XNOR2_X1 U16895 ( .A(n22256), .B(keyinput_44), .ZN(n14955) );
  OAI21_X1 U16896 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14963) );
  XOR2_X1 U16897 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_47), .Z(n14960) );
  XNOR2_X1 U16898 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_45), .ZN(n14959) );
  XNOR2_X1 U16899 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_46), .ZN(n14958) );
  NOR3_X1 U16900 ( .A1(n14960), .A2(n14959), .A3(n14958), .ZN(n14962) );
  XNOR2_X1 U16901 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_48), .ZN(
        n14961) );
  AOI21_X1 U16902 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14967) );
  XOR2_X1 U16903 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_49), .Z(
        n14966) );
  XOR2_X1 U16904 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_51), .Z(
        n14965) );
  XOR2_X1 U16905 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_50), .Z(
        n14964) );
  OAI211_X1 U16906 ( .C1(n14967), .C2(n14966), .A(n14965), .B(n14964), .ZN(
        n14974) );
  XOR2_X1 U16907 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_55), .Z(n14971) );
  XOR2_X1 U16908 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_54), .Z(n14970) );
  XNOR2_X1 U16909 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_52), .ZN(n14969)
         );
  XNOR2_X1 U16910 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_53), .ZN(n14968)
         );
  NOR4_X1 U16911 ( .A1(n14971), .A2(n14970), .A3(n14969), .A4(n14968), .ZN(
        n14973) );
  XOR2_X1 U16912 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_56), .Z(n14972) );
  AOI21_X1 U16913 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n14980) );
  INV_X1 U16914 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20422) );
  AOI22_X1 U16915 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_57), .B1(n20422), .B2(keyinput_61), .ZN(n14975) );
  OAI221_X1 U16916 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .C1(
        n20422), .C2(keyinput_61), .A(n14975), .ZN(n14979) );
  INV_X1 U16917 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20425) );
  AOI22_X1 U16918 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_59), .B1(n20425), .B2(keyinput_58), .ZN(n14976) );
  OAI221_X1 U16919 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_59), .C1(
        n20425), .C2(keyinput_58), .A(n14976), .ZN(n14978) );
  XNOR2_X1 U16920 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_60), .ZN(n14977)
         );
  NOR4_X1 U16921 ( .A1(n14980), .A2(n14979), .A3(n14978), .A4(n14977), .ZN(
        n14983) );
  XNOR2_X1 U16922 ( .A(n22123), .B(keyinput_62), .ZN(n14982) );
  XNOR2_X1 U16923 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_63), .ZN(n14981)
         );
  NOR3_X1 U16924 ( .A1(n14983), .A2(n14982), .A3(n14981), .ZN(n14995) );
  INV_X1 U16925 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20414) );
  OAI22_X1 U16926 ( .A1(keyinput_69), .A2(n20407), .B1(n20414), .B2(
        keyinput_65), .ZN(n14994) );
  OAI22_X1 U16927 ( .A1(n20404), .A2(keyinput_71), .B1(P1_REIP_REG_13__SCAN_IN), .B2(keyinput_70), .ZN(n14993) );
  NOR2_X1 U16928 ( .A1(n22000), .A2(keyinput_64), .ZN(n14991) );
  INV_X1 U16929 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20410) );
  INV_X1 U16930 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20413) );
  OAI22_X1 U16931 ( .A1(keyinput_67), .A2(n20410), .B1(n20413), .B2(
        keyinput_66), .ZN(n14990) );
  NOR2_X1 U16932 ( .A1(n20408), .A2(keyinput_68), .ZN(n14989) );
  AOI22_X1 U16933 ( .A1(n20404), .A2(keyinput_71), .B1(keyinput_67), .B2(
        n20410), .ZN(n14987) );
  AOI22_X1 U16934 ( .A1(n20408), .A2(keyinput_68), .B1(keyinput_66), .B2(
        n20413), .ZN(n14986) );
  AOI22_X1 U16935 ( .A1(n22000), .A2(keyinput_64), .B1(n20414), .B2(
        keyinput_65), .ZN(n14985) );
  AOI22_X1 U16936 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(keyinput_70), .B1(n20407), .B2(keyinput_69), .ZN(n14984) );
  NAND4_X1 U16937 ( .A1(n14987), .A2(n14986), .A3(n14985), .A4(n14984), .ZN(
        n14988) );
  OR4_X1 U16938 ( .A1(n14991), .A2(n14990), .A3(n14989), .A4(n14988), .ZN(
        n14992) );
  NOR4_X1 U16939 ( .A1(n14995), .A2(n14994), .A3(n14993), .A4(n14992), .ZN(
        n14999) );
  XNOR2_X1 U16940 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_72), .ZN(n14998)
         );
  XOR2_X1 U16941 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_74), .Z(n14997) );
  XNOR2_X1 U16942 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_73), .ZN(n14996)
         );
  OAI211_X1 U16943 ( .C1(n14999), .C2(n14998), .A(n14997), .B(n14996), .ZN(
        n15002) );
  XOR2_X1 U16944 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_75), .Z(n15001) );
  XOR2_X1 U16945 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_76), .Z(n15000) );
  AOI21_X1 U16946 ( .B1(n15002), .B2(n15001), .A(n15000), .ZN(n15005) );
  XNOR2_X1 U16947 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_77), .ZN(n15004)
         );
  XNOR2_X1 U16948 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_78), .ZN(n15003)
         );
  OAI21_X1 U16949 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(n15013) );
  XOR2_X1 U16950 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_82), .Z(n15012) );
  XOR2_X1 U16951 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_81), .Z(n15011) );
  XOR2_X1 U16952 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_84), .Z(n15009) );
  XOR2_X1 U16953 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_79), .Z(n15008) );
  XOR2_X1 U16954 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_83), .Z(n15007) );
  XNOR2_X1 U16955 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_80), .ZN(n15006)
         );
  NOR4_X1 U16956 ( .A1(n15009), .A2(n15008), .A3(n15007), .A4(n15006), .ZN(
        n15010) );
  NAND4_X1 U16957 ( .A1(n15013), .A2(n15012), .A3(n15011), .A4(n15010), .ZN(
        n15016) );
  XNOR2_X1 U16958 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_85), .ZN(n15015)
         );
  XNOR2_X1 U16959 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_86), .ZN(n15014)
         );
  NAND3_X1 U16960 ( .A1(n15016), .A2(n15015), .A3(n15014), .ZN(n15020) );
  XNOR2_X1 U16961 ( .A(n16422), .B(keyinput_89), .ZN(n15019) );
  XOR2_X1 U16962 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_88), .Z(n15018) );
  XNOR2_X1 U16963 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_87), .ZN(n15017)
         );
  NAND4_X1 U16964 ( .A1(n15020), .A2(n15019), .A3(n15018), .A4(n15017), .ZN(
        n15026) );
  XNOR2_X1 U16965 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .ZN(n15025)
         );
  XOR2_X1 U16966 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_92), .Z(n15023) );
  INV_X1 U16967 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16432) );
  XNOR2_X1 U16968 ( .A(n16432), .B(keyinput_93), .ZN(n15022) );
  INV_X1 U16969 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n16426) );
  XNOR2_X1 U16970 ( .A(n16426), .B(keyinput_91), .ZN(n15021) );
  NAND3_X1 U16971 ( .A1(n15023), .A2(n15022), .A3(n15021), .ZN(n15024) );
  AOI21_X1 U16972 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15029) );
  XNOR2_X1 U16973 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_94), .ZN(n15028)
         );
  INV_X1 U16974 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n16441) );
  XNOR2_X1 U16975 ( .A(n16441), .B(keyinput_95), .ZN(n15027) );
  OAI21_X1 U16976 ( .B1(n15029), .B2(n15028), .A(n15027), .ZN(n15036) );
  XNOR2_X1 U16977 ( .A(n16448), .B(keyinput_97), .ZN(n15033) );
  INV_X1 U16978 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n22098) );
  XNOR2_X1 U16979 ( .A(n22098), .B(keyinput_96), .ZN(n15032) );
  XNOR2_X1 U16980 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_98), .ZN(n15031)
         );
  XNOR2_X1 U16981 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_99), .ZN(n15030)
         );
  NOR4_X1 U16982 ( .A1(n15033), .A2(n15032), .A3(n15031), .A4(n15030), .ZN(
        n15035) );
  XOR2_X1 U16983 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_100), .Z(n15034) );
  AOI21_X1 U16984 ( .B1(n15036), .B2(n15035), .A(n15034), .ZN(n15039) );
  XNOR2_X1 U16985 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n15038)
         );
  XOR2_X1 U16986 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_102), .Z(n15037) );
  OAI21_X1 U16987 ( .B1(n15039), .B2(n15038), .A(n15037), .ZN(n15043) );
  XNOR2_X1 U16988 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_104), .ZN(n15042)
         );
  XNOR2_X1 U16989 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_103), .ZN(n15041)
         );
  XNOR2_X1 U16990 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_105), .ZN(n15040)
         );
  NAND4_X1 U16991 ( .A1(n15043), .A2(n15042), .A3(n15041), .A4(n15040), .ZN(
        n15047) );
  XNOR2_X1 U16992 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n15046)
         );
  XNOR2_X1 U16993 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_108), .ZN(n15045)
         );
  XNOR2_X1 U16994 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_107), .ZN(n15044)
         );
  AOI211_X1 U16995 ( .C1(n15047), .C2(n15046), .A(n15045), .B(n15044), .ZN(
        n15050) );
  XOR2_X1 U16996 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_109), .Z(n15049) );
  XOR2_X1 U16997 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_110), .Z(n15048) );
  OAI21_X1 U16998 ( .B1(n15050), .B2(n15049), .A(n15048), .ZN(n15054) );
  XOR2_X1 U16999 ( .A(P1_EBX_REG_2__SCAN_IN), .B(keyinput_113), .Z(n15053) );
  XNOR2_X1 U17000 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n15052)
         );
  XNOR2_X1 U17001 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_112), .ZN(n15051)
         );
  NAND4_X1 U17002 ( .A1(n15054), .A2(n15053), .A3(n15052), .A4(n15051), .ZN(
        n15057) );
  XOR2_X1 U17003 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_114), .Z(n15056) );
  XNOR2_X1 U17004 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_115), .ZN(n15055)
         );
  NAND3_X1 U17005 ( .A1(n15057), .A2(n15056), .A3(n15055), .ZN(n15060) );
  XNOR2_X1 U17006 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_116), .ZN(n15059)
         );
  XNOR2_X1 U17007 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n15058)
         );
  NAND3_X1 U17008 ( .A1(n15060), .A2(n15059), .A3(n15058), .ZN(n15074) );
  XOR2_X1 U17009 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_118), .Z(n15073) );
  OAI22_X1 U17010 ( .A1(keyinput_122), .A2(n16492), .B1(n16505), .B2(
        keyinput_124), .ZN(n15071) );
  INV_X1 U17011 ( .A(keyinput_119), .ZN(n15066) );
  AOI22_X1 U17012 ( .A1(n16472), .A2(keyinput_119), .B1(n16517), .B2(
        keyinput_126), .ZN(n15064) );
  AOI22_X1 U17013 ( .A1(n16505), .A2(keyinput_124), .B1(keyinput_122), .B2(
        n16492), .ZN(n15063) );
  AOI22_X1 U17014 ( .A1(P1_EAX_REG_26__SCAN_IN), .A2(keyinput_121), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_125), .ZN(n15062) );
  AOI22_X1 U17015 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_123), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(keyinput_120), .ZN(n15061) );
  NAND4_X1 U17016 ( .A1(n15064), .A2(n15063), .A3(n15062), .A4(n15061), .ZN(
        n15065) );
  AOI21_X1 U17017 ( .B1(n15066), .B2(P1_EAX_REG_28__SCAN_IN), .A(n15065), .ZN(
        n15067) );
  OAI21_X1 U17018 ( .B1(keyinput_126), .B2(n16517), .A(n15067), .ZN(n15070) );
  OAI22_X1 U17019 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_120), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_121), .ZN(n15069) );
  OAI22_X1 U17020 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_123), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_125), .ZN(n15068) );
  OR4_X1 U17021 ( .A1(n15071), .A2(n15070), .A3(n15069), .A4(n15068), .ZN(
        n15072) );
  AOI21_X1 U17022 ( .B1(n15074), .B2(n15073), .A(n15072), .ZN(n15075) );
  AOI211_X1 U17023 ( .C1(n15078), .C2(n15077), .A(n15076), .B(n15075), .ZN(
        n15102) );
  INV_X1 U17024 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17534) );
  INV_X1 U17025 ( .A(n15079), .ZN(n15082) );
  INV_X1 U17026 ( .A(n15080), .ZN(n15081) );
  NAND2_X1 U17027 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  AND2_X1 U17028 ( .A1(n15084), .A2(n15083), .ZN(n15091) );
  INV_X1 U17029 ( .A(n15085), .ZN(n15086) );
  NAND2_X1 U17030 ( .A1(n15087), .A2(n15086), .ZN(n15090) );
  NAND2_X1 U17031 ( .A1(n15095), .A2(n15088), .ZN(n15089) );
  OAI211_X1 U17032 ( .C1(n15091), .C2(n15095), .A(n15090), .B(n15089), .ZN(
        n15093) );
  NAND2_X1 U17033 ( .A1(n15093), .A2(n15092), .ZN(n17538) );
  OR2_X1 U17034 ( .A1(n15095), .A2(n15094), .ZN(n15099) );
  INV_X1 U17035 ( .A(n13809), .ZN(n15096) );
  NAND2_X1 U17036 ( .A1(n15097), .A2(n15096), .ZN(n15098) );
  NAND2_X1 U17037 ( .A1(n15099), .A2(n15098), .ZN(n20523) );
  NAND3_X1 U17038 ( .A1(n15284), .A2(n16209), .A3(n22189), .ZN(n15100) );
  AND2_X1 U17039 ( .A1(n15100), .A2(n21842), .ZN(n21843) );
  NOR2_X1 U17040 ( .A1(n20523), .A2(n21843), .ZN(n17536) );
  NOR2_X1 U17041 ( .A1(n17536), .A2(n22162), .ZN(n22143) );
  MUX2_X1 U17042 ( .A(n17534), .B(n17538), .S(n22143), .Z(n15101) );
  XNOR2_X1 U17043 ( .A(n15102), .B(n15101), .ZN(P1_U3484) );
  OR2_X1 U17044 ( .A1(n15103), .A2(n11285), .ZN(n15105) );
  NAND2_X1 U17045 ( .A1(n15105), .A2(n15104), .ZN(n21902) );
  XOR2_X1 U17046 ( .A(n15107), .B(n15106), .Z(n20471) );
  INV_X1 U17047 ( .A(n20471), .ZN(n15117) );
  OAI222_X1 U17048 ( .A1(n21902), .A2(n16453), .B1(n16425), .B2(n15117), .C1(
        n16451), .C2(n15588), .ZN(P1_U2868) );
  INV_X1 U17049 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n15116) );
  OAI211_X1 U17050 ( .C1(n15108), .C2(n11696), .A(n15746), .B(n15263), .ZN(
        n15115) );
  NAND2_X1 U17051 ( .A1(n15110), .A2(n15109), .ZN(n15112) );
  INV_X1 U17052 ( .A(n11263), .ZN(n15111) );
  NAND2_X1 U17053 ( .A1(n15112), .A2(n15111), .ZN(n18783) );
  INV_X1 U17054 ( .A(n18783), .ZN(n15113) );
  NAND2_X1 U17055 ( .A1(n16952), .A2(n15113), .ZN(n15114) );
  OAI211_X1 U17056 ( .C1(n16952), .C2(n15116), .A(n15115), .B(n15114), .ZN(
        P2_U2878) );
  OAI222_X1 U17057 ( .A1(n15478), .A2(n22383), .B1(n16523), .B2(n20363), .C1(
        n16553), .C2(n15117), .ZN(P1_U2900) );
  NOR2_X1 U17058 ( .A1(n15388), .A2(n15164), .ZN(n15378) );
  INV_X1 U17059 ( .A(n15354), .ZN(n15119) );
  NOR2_X1 U17060 ( .A1(n15119), .A2(n15336), .ZN(n15348) );
  AOI21_X1 U17061 ( .B1(n15121), .B2(n15120), .A(n22290), .ZN(n15122) );
  AOI21_X1 U17062 ( .B1(n15123), .B2(n15419), .A(n15122), .ZN(n15126) );
  INV_X1 U17063 ( .A(n17556), .ZN(n15125) );
  NAND2_X1 U17064 ( .A1(n15125), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15124) );
  OAI21_X1 U17065 ( .B1(n15126), .B2(n15125), .A(n15124), .ZN(P1_U3475) );
  NAND3_X1 U17066 ( .A1(n17526), .A2(n17523), .A3(n17517), .ZN(n22234) );
  INV_X1 U17067 ( .A(n22234), .ZN(n15131) );
  INV_X1 U17068 ( .A(n15342), .ZN(n15128) );
  OR2_X1 U17069 ( .A1(n15419), .A2(n11947), .ZN(n22239) );
  INV_X1 U17070 ( .A(n22239), .ZN(n15335) );
  INV_X1 U17071 ( .A(n15377), .ZN(n15166) );
  NOR2_X1 U17072 ( .A1(n15376), .A2(n22234), .ZN(n22485) );
  AOI21_X1 U17073 ( .B1(n15335), .B2(n15166), .A(n22485), .ZN(n15130) );
  OAI211_X1 U17074 ( .C1(n15128), .C2(n15164), .A(n15381), .B(n15130), .ZN(
        n15129) );
  OAI211_X1 U17075 ( .C1(n15381), .C2(n15131), .A(n15129), .B(n15379), .ZN(
        n22488) );
  NAND2_X1 U17076 ( .A1(n22488), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15135) );
  NAND2_X1 U17077 ( .A1(n15342), .A2(n15382), .ZN(n22493) );
  INV_X1 U17078 ( .A(n15130), .ZN(n15132) );
  AOI22_X1 U17079 ( .A1(n15132), .A2(n15381), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15131), .ZN(n22305) );
  INV_X1 U17080 ( .A(n22485), .ZN(n15142) );
  OAI22_X1 U17081 ( .A1(n22305), .A2(n16880), .B1(n22370), .B2(n15142), .ZN(
        n15133) );
  AOI21_X1 U17082 ( .B1(n22487), .B2(n16876), .A(n15133), .ZN(n15134) );
  OAI211_X1 U17083 ( .C1(n22371), .C2(n22491), .A(n15135), .B(n15134), .ZN(
        P1_U3044) );
  NAND2_X1 U17084 ( .A1(n22488), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15138) );
  OAI22_X1 U17085 ( .A1(n22305), .A2(n16865), .B1(n22266), .B2(n15142), .ZN(
        n15136) );
  AOI21_X1 U17086 ( .B1(n22487), .B2(n16861), .A(n15136), .ZN(n15137) );
  OAI211_X1 U17087 ( .C1(n22267), .C2(n22491), .A(n15138), .B(n15137), .ZN(
        P1_U3041) );
  NAND2_X1 U17088 ( .A1(n22488), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n15141) );
  OAI22_X1 U17089 ( .A1(n16892), .A2(n22305), .B1(n16889), .B2(n15142), .ZN(
        n15139) );
  AOI21_X1 U17090 ( .B1(n22487), .B2(n16886), .A(n15139), .ZN(n15140) );
  OAI211_X1 U17091 ( .C1(n15712), .C2(n22491), .A(n15141), .B(n15140), .ZN(
        P1_U3047) );
  NAND2_X1 U17092 ( .A1(n22488), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15145) );
  OAI22_X1 U17093 ( .A1(n22305), .A2(n16875), .B1(n22341), .B2(n15142), .ZN(
        n15143) );
  AOI21_X1 U17094 ( .B1(n22487), .B2(n16871), .A(n15143), .ZN(n15144) );
  OAI211_X1 U17095 ( .C1(n22342), .C2(n22491), .A(n15145), .B(n15144), .ZN(
        P1_U3043) );
  AOI22_X1 U17096 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21841), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20371), .ZN(n15146) );
  OAI21_X1 U17097 ( .B1(n15147), .B2(n15162), .A(n15146), .ZN(P1_U2920) );
  AOI22_X1 U17098 ( .A1(n21841), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15148) );
  OAI21_X1 U17099 ( .B1(n15149), .B2(n15162), .A(n15148), .ZN(P1_U2907) );
  AOI22_X1 U17100 ( .A1(n21841), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15150) );
  OAI21_X1 U17101 ( .B1(n16511), .B2(n15162), .A(n15150), .ZN(P1_U2914) );
  AOI22_X1 U17102 ( .A1(n21841), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15151) );
  OAI21_X1 U17103 ( .B1(n16486), .B2(n15162), .A(n15151), .ZN(P1_U2910) );
  AOI22_X1 U17104 ( .A1(n21841), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15152) );
  OAI21_X1 U17105 ( .B1(n16479), .B2(n15162), .A(n15152), .ZN(P1_U2909) );
  AOI22_X1 U17106 ( .A1(n21841), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15153) );
  OAI21_X1 U17107 ( .B1(n16517), .B2(n15162), .A(n15153), .ZN(P1_U2915) );
  AOI22_X1 U17108 ( .A1(n21841), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15154) );
  OAI21_X1 U17109 ( .B1(n16472), .B2(n15162), .A(n15154), .ZN(P1_U2908) );
  AOI22_X1 U17110 ( .A1(n21841), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15155) );
  OAI21_X1 U17111 ( .B1(n16505), .B2(n15162), .A(n15155), .ZN(P1_U2913) );
  AOI22_X1 U17112 ( .A1(n21841), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15156) );
  OAI21_X1 U17113 ( .B1(n15157), .B2(n15162), .A(n15156), .ZN(P1_U2906) );
  AOI22_X1 U17114 ( .A1(n21841), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15158) );
  OAI21_X1 U17115 ( .B1(n16492), .B2(n15162), .A(n15158), .ZN(P1_U2911) );
  AOI22_X1 U17116 ( .A1(n21841), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15159) );
  OAI21_X1 U17117 ( .B1(n16499), .B2(n15162), .A(n15159), .ZN(P1_U2912) );
  AOI22_X1 U17118 ( .A1(n21841), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15160) );
  OAI21_X1 U17119 ( .B1(n16524), .B2(n15162), .A(n15160), .ZN(P1_U2916) );
  AOI22_X1 U17120 ( .A1(n21841), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15161) );
  OAI21_X1 U17121 ( .B1(n15163), .B2(n15162), .A(n15161), .ZN(P1_U2917) );
  INV_X1 U17122 ( .A(n15164), .ZN(n15168) );
  NOR2_X1 U17123 ( .A1(n16826), .A2(n15165), .ZN(n22258) );
  NAND3_X1 U17124 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17526), .A3(
        n17517), .ZN(n22252) );
  NOR2_X1 U17125 ( .A1(n15376), .A2(n22252), .ZN(n22514) );
  AOI21_X1 U17126 ( .B1(n22258), .B2(n15166), .A(n22514), .ZN(n15172) );
  NAND2_X1 U17127 ( .A1(n15172), .A2(n22253), .ZN(n15167) );
  AOI21_X1 U17128 ( .B1(n15354), .B2(n15168), .A(n15167), .ZN(n15171) );
  INV_X1 U17129 ( .A(n22252), .ZN(n15173) );
  NOR2_X1 U17130 ( .A1(n15381), .A2(n15173), .ZN(n15170) );
  INV_X1 U17131 ( .A(n15379), .ZN(n15169) );
  OR2_X1 U17132 ( .A1(n15172), .A2(n22290), .ZN(n15175) );
  NAND2_X1 U17133 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15173), .ZN(n15174) );
  OAI22_X1 U17134 ( .A1(n22521), .A2(n22359), .B1(n22263), .B2(n16875), .ZN(
        n15177) );
  INV_X1 U17135 ( .A(n22514), .ZN(n15188) );
  OAI22_X1 U17136 ( .A1(n22513), .A2(n22342), .B1(n15188), .B2(n22341), .ZN(
        n15176) );
  AOI211_X1 U17137 ( .C1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .C2(n22517), .A(
        n15177), .B(n15176), .ZN(n15178) );
  INV_X1 U17138 ( .A(n15178), .ZN(P1_U3075) );
  OAI22_X1 U17139 ( .A1(n22521), .A2(n22382), .B1(n22263), .B2(n16880), .ZN(
        n15180) );
  OAI22_X1 U17140 ( .A1(n22513), .A2(n22371), .B1(n15188), .B2(n22370), .ZN(
        n15179) );
  AOI211_X1 U17141 ( .C1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .C2(n22517), .A(
        n15180), .B(n15179), .ZN(n15181) );
  INV_X1 U17142 ( .A(n15181), .ZN(P1_U3076) );
  OAI22_X1 U17143 ( .A1(n22521), .A2(n22459), .B1(n22263), .B2(n16885), .ZN(
        n15183) );
  OAI22_X1 U17144 ( .A1(n22513), .A2(n22442), .B1(n22441), .B2(n15188), .ZN(
        n15182) );
  AOI211_X1 U17145 ( .C1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .C2(n22517), .A(
        n15183), .B(n15182), .ZN(n15184) );
  INV_X1 U17146 ( .A(n15184), .ZN(P1_U3078) );
  OAI22_X1 U17147 ( .A1(n22521), .A2(n22330), .B1(n22263), .B2(n16870), .ZN(
        n15186) );
  OAI22_X1 U17148 ( .A1(n22513), .A2(n22309), .B1(n15188), .B2(n22308), .ZN(
        n15185) );
  AOI211_X1 U17149 ( .C1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n22517), .A(
        n15186), .B(n15185), .ZN(n15187) );
  INV_X1 U17150 ( .A(n15187), .ZN(P1_U3074) );
  OAI22_X1 U17151 ( .A1(n22521), .A2(n22473), .B1(n16892), .B2(n22263), .ZN(
        n15190) );
  OAI22_X1 U17152 ( .A1(n22513), .A2(n15712), .B1(n15188), .B2(n16889), .ZN(
        n15189) );
  AOI211_X1 U17153 ( .C1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .C2(n22517), .A(
        n15190), .B(n15189), .ZN(n15191) );
  INV_X1 U17154 ( .A(n15191), .ZN(P1_U3079) );
  INV_X1 U17155 ( .A(n19690), .ZN(n17690) );
  XNOR2_X1 U17156 ( .A(n19690), .B(n20111), .ZN(n20114) );
  XNOR2_X1 U17157 ( .A(n15193), .B(n15192), .ZN(n20163) );
  NOR2_X1 U17158 ( .A1(n19674), .A2(n20163), .ZN(n20166) );
  NOR2_X1 U17159 ( .A1(n20114), .A2(n20166), .ZN(n20113) );
  AOI21_X1 U17160 ( .B1(n15194), .B2(n17690), .A(n20113), .ZN(n15195) );
  XNOR2_X1 U17161 ( .A(n15195), .B(n20059), .ZN(n20061) );
  NAND2_X1 U17162 ( .A1(n15195), .A2(n20059), .ZN(n15196) );
  OAI21_X1 U17163 ( .B1(n20061), .B2(n17686), .A(n15196), .ZN(n20011) );
  INV_X1 U17164 ( .A(n15197), .ZN(n15198) );
  XNOR2_X1 U17165 ( .A(n15199), .B(n15198), .ZN(n20009) );
  XNOR2_X1 U17166 ( .A(n17691), .B(n20009), .ZN(n20012) );
  NOR2_X1 U17167 ( .A1(n20011), .A2(n20012), .ZN(n20010) );
  NOR2_X1 U17168 ( .A1(n17691), .A2(n20009), .ZN(n15202) );
  XNOR2_X1 U17169 ( .A(n15200), .B(n15201), .ZN(n18730) );
  OAI21_X1 U17170 ( .B1(n20010), .B2(n15202), .A(n18730), .ZN(n19906) );
  XOR2_X1 U17171 ( .A(n18729), .B(n19906), .Z(n15219) );
  NAND2_X1 U17172 ( .A1(n15204), .A2(n15203), .ZN(n15205) );
  NAND2_X1 U17173 ( .A1(n15206), .A2(n15205), .ZN(n15207) );
  NAND2_X1 U17174 ( .A1(n15207), .A2(n19160), .ZN(n15210) );
  NAND2_X1 U17175 ( .A1(n18717), .A2(n15208), .ZN(n15209) );
  NAND2_X1 U17176 ( .A1(n20162), .A2(n15211), .ZN(n20115) );
  INV_X1 U17177 ( .A(n20164), .ZN(n20112) );
  INV_X1 U17178 ( .A(n18730), .ZN(n15213) );
  INV_X1 U17179 ( .A(n20162), .ZN(n20110) );
  AOI22_X1 U17180 ( .A1(n20112), .A2(n15213), .B1(n20110), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U17181 ( .A1(n20162), .A2(n15214), .ZN(n15754) );
  INV_X1 U17182 ( .A(n15754), .ZN(n15216) );
  NAND2_X1 U17183 ( .A1(n19643), .A2(n19965), .ZN(n15217) );
  OAI211_X1 U17184 ( .C1(n15219), .C2(n20115), .A(n15218), .B(n15217), .ZN(
        P2_U2915) );
  XOR2_X1 U17185 ( .A(n14669), .B(n15220), .Z(n22042) );
  INV_X1 U17186 ( .A(n22042), .ZN(n15271) );
  NAND2_X1 U17187 ( .A1(n14072), .A2(n21922), .ZN(n15221) );
  OAI211_X1 U17188 ( .C1(n16209), .C2(P1_EBX_REG_6__SCAN_IN), .A(n16261), .B(
        n15221), .ZN(n15222) );
  OAI21_X1 U17189 ( .B1(n16205), .B2(P1_EBX_REG_6__SCAN_IN), .A(n15222), .ZN(
        n15330) );
  XOR2_X1 U17190 ( .A(n15331), .B(n15330), .Z(n22035) );
  AOI22_X1 U17191 ( .A1(n16463), .A2(n22035), .B1(n16462), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n15223) );
  OAI21_X1 U17192 ( .B1(n15271), .B2(n16425), .A(n15223), .ZN(P1_U2866) );
  OAI21_X1 U17193 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n15226), .A(
        n15551), .ZN(n17567) );
  INV_X1 U17194 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18918) );
  INV_X1 U17195 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18940) );
  INV_X1 U17196 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17092) );
  INV_X1 U17197 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17069) );
  INV_X1 U17198 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15224) );
  AOI21_X1 U17199 ( .B1(n15510), .B2(n15228), .A(n15226), .ZN(n18740) );
  OAI22_X1 U17200 ( .A1(n15635), .A2(n19073), .B1(n15368), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n17413) );
  OAI22_X1 U17201 ( .A1(n15635), .A2(n15227), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15571) );
  OR2_X1 U17202 ( .A1(n17413), .A2(n15571), .ZN(n15311) );
  NOR2_X1 U17203 ( .A1(n15312), .A2(n15311), .ZN(n15253) );
  OAI21_X1 U17204 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n15229), .A(
        n15228), .ZN(n15483) );
  NAND2_X1 U17205 ( .A1(n15253), .A2(n15483), .ZN(n18737) );
  NOR2_X1 U17206 ( .A1(n18740), .A2(n18737), .ZN(n15552) );
  NOR2_X1 U17207 ( .A1(n18778), .A2(n15552), .ZN(n15230) );
  XNOR2_X1 U17208 ( .A(n17567), .B(n15230), .ZN(n15236) );
  INV_X1 U17209 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19734) );
  NAND4_X1 U17210 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15635), .A3(n19734), 
        .A4(n22169), .ZN(n19154) );
  XNOR2_X1 U17211 ( .A(n15233), .B(n15232), .ZN(n19909) );
  AND2_X1 U17212 ( .A1(n18717), .A2(n15234), .ZN(n15246) );
  INV_X1 U17213 ( .A(n19164), .ZN(n22197) );
  NOR2_X1 U17214 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n22197), .ZN(n15244) );
  OAI22_X1 U17215 ( .A1(n19051), .A2(n19909), .B1(n19008), .B2(n15687), .ZN(
        n15235) );
  AOI21_X1 U17216 ( .B1(n15236), .B2(n19003), .A(n15235), .ZN(n15252) );
  NOR2_X1 U17217 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15635), .ZN(n19158) );
  NAND3_X1 U17218 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19158), .A3(n15237), 
        .ZN(n19168) );
  NAND3_X1 U17219 ( .A1(n18892), .A2(n19168), .A3(n19154), .ZN(n15238) );
  OAI22_X1 U17220 ( .A1(n19060), .A2(n15239), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n15244), .ZN(n15240) );
  AND2_X1 U17221 ( .A1(n15241), .A2(n15240), .ZN(n15242) );
  NAND2_X1 U17222 ( .A1(n18717), .A2(n15242), .ZN(n19040) );
  OAI21_X1 U17223 ( .B1(n19040), .B2(n15243), .A(n18813), .ZN(n15250) );
  INV_X1 U17224 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15248) );
  INV_X1 U17225 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n19039) );
  NOR2_X1 U17226 ( .A1(n19039), .A2(n15244), .ZN(n15245) );
  OAI22_X1 U17227 ( .A1(n15248), .A2(n19036), .B1(n15247), .B2(n19037), .ZN(
        n15249) );
  AOI211_X1 U17228 ( .C1(n19011), .C2(P2_REIP_REG_5__SCAN_IN), .A(n15250), .B(
        n15249), .ZN(n15251) );
  NAND2_X1 U17229 ( .A1(n15252), .A2(n15251), .ZN(P2_U2850) );
  NOR2_X1 U17230 ( .A1(n18778), .A2(n15253), .ZN(n15254) );
  XNOR2_X1 U17231 ( .A(n15254), .B(n15483), .ZN(n15255) );
  NAND2_X1 U17232 ( .A1(n15255), .A2(n19003), .ZN(n15262) );
  NOR2_X1 U17233 ( .A1(n19037), .A2(n15256), .ZN(n15258) );
  INV_X1 U17234 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15482) );
  OAI22_X1 U17235 ( .A1(n15482), .A2(n19036), .B1(n15481), .B2(n19041), .ZN(
        n15257) );
  AOI211_X1 U17236 ( .C1(n19013), .C2(P2_EBX_REG_3__SCAN_IN), .A(n15258), .B(
        n15257), .ZN(n15259) );
  OAI21_X1 U17237 ( .B1(n15473), .B2(n19008), .A(n15259), .ZN(n15260) );
  AOI21_X1 U17238 ( .B1(n19014), .B2(n20009), .A(n15260), .ZN(n15261) );
  OAI211_X1 U17239 ( .C1(n15581), .C2(n19795), .A(n15262), .B(n15261), .ZN(
        P2_U2852) );
  OAI211_X1 U17240 ( .C1(n15264), .C2(n11698), .A(n15746), .B(n15494), .ZN(
        n15268) );
  OR2_X1 U17241 ( .A1(n15265), .A2(n11263), .ZN(n15266) );
  NAND2_X1 U17242 ( .A1(n15274), .A2(n15266), .ZN(n18800) );
  INV_X1 U17243 ( .A(n18800), .ZN(n19082) );
  NAND2_X1 U17244 ( .A1(n16952), .A2(n19082), .ZN(n15267) );
  OAI211_X1 U17245 ( .C1(n16952), .C2(n15269), .A(n15268), .B(n15267), .ZN(
        P2_U2877) );
  OAI222_X1 U17246 ( .A1(n15478), .A2(n16513), .B1(n16553), .B2(n15271), .C1(
        n15270), .C2(n16523), .ZN(P1_U2898) );
  INV_X1 U17247 ( .A(n15495), .ZN(n15493) );
  XNOR2_X1 U17248 ( .A(n15494), .B(n15493), .ZN(n15278) );
  NAND2_X1 U17249 ( .A1(n15274), .A2(n15273), .ZN(n15275) );
  AND2_X1 U17250 ( .A1(n15491), .A2(n15275), .ZN(n18807) );
  NOR2_X1 U17251 ( .A1(n16952), .A2(n13475), .ZN(n15276) );
  AOI21_X1 U17252 ( .B1(n18807), .B2(n16952), .A(n15276), .ZN(n15277) );
  OAI21_X1 U17253 ( .B1(n15278), .B2(n16968), .A(n15277), .ZN(P2_U2876) );
  OAI22_X1 U17254 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .B1(n15279), .B2(n22280), .ZN(n15281) );
  OAI211_X1 U17255 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n15288), .A(n20525), 
        .B(n22153), .ZN(n15280) );
  NAND2_X1 U17256 ( .A1(n15281), .A2(n15280), .ZN(n15282) );
  NAND2_X2 U17257 ( .A1(n21838), .A2(n15282), .ZN(n15842) );
  OR2_X1 U17258 ( .A1(n15292), .A2(n15283), .ZN(n15592) );
  NOR2_X1 U17259 ( .A1(n15292), .A2(n15284), .ZN(n15290) );
  INV_X1 U17260 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16285) );
  NOR2_X1 U17261 ( .A1(n16557), .A2(n15288), .ZN(n15289) );
  NAND2_X1 U17262 ( .A1(n15291), .A2(n22030), .ZN(n15310) );
  AND2_X1 U17263 ( .A1(n21842), .A2(n22256), .ZN(n15297) );
  AND2_X1 U17264 ( .A1(n15294), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n15296) );
  NOR2_X1 U17265 ( .A1(n17544), .A2(n15296), .ZN(n15295) );
  INV_X1 U17266 ( .A(n15296), .ZN(n15298) );
  NOR2_X1 U17267 ( .A1(n15298), .A2(n15297), .ZN(n15299) );
  AND2_X1 U17268 ( .A1(n15842), .A2(n15300), .ZN(n22110) );
  INV_X1 U17269 ( .A(n15301), .ZN(n15304) );
  OAI21_X1 U17270 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n22073), .A(n15842), .ZN(
        n15303) );
  AOI22_X1 U17271 ( .A1(n22110), .A2(n15304), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n15303), .ZN(n15306) );
  AND2_X2 U17272 ( .A1(n15842), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22134) );
  NAND2_X1 U17273 ( .A1(n22134), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15305) );
  OAI211_X1 U17274 ( .C1(n22059), .C2(n21886), .A(n15306), .B(n15305), .ZN(
        n15308) );
  INV_X1 U17275 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20387) );
  NOR3_X1 U17276 ( .A1(n22073), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n20387), .ZN(
        n15307) );
  AOI211_X1 U17277 ( .C1(P1_EBX_REG_2__SCAN_IN), .C2(n22118), .A(n15308), .B(
        n15307), .ZN(n15309) );
  OAI211_X1 U17278 ( .C1(n15592), .C2(n16826), .A(n15310), .B(n15309), .ZN(
        P1_U2838) );
  NAND2_X1 U17279 ( .A1(n17412), .A2(n15311), .ZN(n15570) );
  XNOR2_X1 U17280 ( .A(n15312), .B(n15570), .ZN(n15313) );
  NAND2_X1 U17281 ( .A1(n15313), .A2(n19003), .ZN(n15324) );
  INV_X1 U17282 ( .A(n20059), .ZN(n15320) );
  INV_X1 U17283 ( .A(n15314), .ZN(n15318) );
  OAI22_X1 U17284 ( .A1(n15315), .A2(n19036), .B1(n12868), .B2(n19041), .ZN(
        n15317) );
  NOR2_X1 U17285 ( .A1(n19040), .A2(n13416), .ZN(n15316) );
  AOI211_X1 U17286 ( .C1(n19009), .C2(n15318), .A(n15317), .B(n15316), .ZN(
        n15319) );
  OAI21_X1 U17287 ( .B1(n15320), .B2(n19051), .A(n15319), .ZN(n15321) );
  AOI21_X1 U17288 ( .B1(n19045), .B2(n15322), .A(n15321), .ZN(n15323) );
  OAI211_X1 U17289 ( .C1(n15581), .C2(n17686), .A(n15324), .B(n15323), .ZN(
        P2_U2853) );
  NAND2_X1 U17290 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  AND2_X1 U17291 ( .A1(n15325), .A2(n15328), .ZN(n22053) );
  INV_X1 U17292 ( .A(n22053), .ZN(n15409) );
  MUX2_X1 U17293 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n15329) );
  NAND2_X1 U17294 ( .A1(n11689), .A2(n15329), .ZN(n15451) );
  INV_X1 U17295 ( .A(n15452), .ZN(n15332) );
  XNOR2_X1 U17296 ( .A(n15451), .B(n15332), .ZN(n22046) );
  INV_X1 U17297 ( .A(n22046), .ZN(n15334) );
  INV_X1 U17298 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15333) );
  OAI222_X1 U17299 ( .A1(n15409), .A2(n16425), .B1(n16453), .B2(n15334), .C1(
        n16451), .C2(n15333), .ZN(P1_U2865) );
  NAND3_X1 U17300 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17526), .A3(
        n17523), .ZN(n15530) );
  NOR2_X1 U17301 ( .A1(n15376), .A2(n15530), .ZN(n22248) );
  AOI21_X1 U17302 ( .B1(n15335), .B2(n15349), .A(n22248), .ZN(n15340) );
  OR2_X1 U17303 ( .A1(n15342), .A2(n22290), .ZN(n15337) );
  NAND2_X1 U17304 ( .A1(n15336), .A2(n15381), .ZN(n16824) );
  OAI22_X1 U17305 ( .A1(n15340), .A2(n15338), .B1(n12293), .B2(n15530), .ZN(
        n22502) );
  INV_X1 U17306 ( .A(n22502), .ZN(n15346) );
  INV_X1 U17307 ( .A(n15338), .ZN(n15339) );
  AOI22_X1 U17308 ( .A1(n15340), .A2(n15339), .B1(n22290), .B2(n15530), .ZN(
        n15341) );
  NAND2_X1 U17309 ( .A1(n15379), .A2(n15341), .ZN(n22503) );
  AOI22_X1 U17310 ( .A1(n22509), .A2(n16886), .B1(n22248), .B2(n22468), .ZN(
        n15343) );
  OAI21_X1 U17311 ( .B1(n15712), .B2(n22500), .A(n15343), .ZN(n15344) );
  AOI21_X1 U17312 ( .B1(n22503), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n15344), .ZN(n15345) );
  OAI21_X1 U17313 ( .B1(n15346), .B2(n16892), .A(n15345), .ZN(P1_U3063) );
  NAND2_X1 U17314 ( .A1(n15347), .A2(n17526), .ZN(n15701) );
  INV_X1 U17315 ( .A(n15701), .ZN(n15356) );
  INV_X1 U17316 ( .A(n15348), .ZN(n15350) );
  INV_X1 U17317 ( .A(n15364), .ZN(n22528) );
  AOI21_X1 U17318 ( .B1(n22258), .B2(n15349), .A(n22528), .ZN(n15355) );
  NAND3_X1 U17319 ( .A1(n15350), .A2(n15381), .A3(n15355), .ZN(n15351) );
  OAI211_X1 U17320 ( .C1(n15381), .C2(n15356), .A(n15351), .B(n15379), .ZN(
        n22531) );
  OAI22_X1 U17321 ( .A1(n22527), .A2(n22267), .B1(n15364), .B2(n22266), .ZN(
        n15359) );
  INV_X1 U17322 ( .A(n15355), .ZN(n15357) );
  AOI22_X1 U17323 ( .A1(n15357), .A2(n15381), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15356), .ZN(n22315) );
  OAI22_X1 U17324 ( .A1(n22534), .A2(n22302), .B1(n22315), .B2(n16865), .ZN(
        n15358) );
  AOI211_X1 U17325 ( .C1(n22531), .C2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n15359), .B(n15358), .ZN(n15360) );
  INV_X1 U17326 ( .A(n15360), .ZN(P1_U3089) );
  OAI22_X1 U17327 ( .A1(n22527), .A2(n15712), .B1(n15364), .B2(n16889), .ZN(
        n15362) );
  OAI22_X1 U17328 ( .A1(n22534), .A2(n22473), .B1(n22315), .B2(n16892), .ZN(
        n15361) );
  AOI211_X1 U17329 ( .C1(n22531), .C2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n15362), .B(n15361), .ZN(n15363) );
  INV_X1 U17330 ( .A(n15363), .ZN(P1_U3095) );
  OAI22_X1 U17331 ( .A1(n22527), .A2(n22371), .B1(n15364), .B2(n22370), .ZN(
        n15366) );
  OAI22_X1 U17332 ( .A1(n22534), .A2(n22382), .B1(n22315), .B2(n16880), .ZN(
        n15365) );
  AOI211_X1 U17333 ( .C1(n22531), .C2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15366), .B(n15365), .ZN(n15367) );
  INV_X1 U17334 ( .A(n15367), .ZN(P1_U3092) );
  NOR2_X1 U17335 ( .A1(n18778), .A2(n19154), .ZN(n19048) );
  NAND2_X1 U17336 ( .A1(n19003), .A2(n18778), .ZN(n18875) );
  AOI21_X1 U17337 ( .B1(n19036), .B2(n18875), .A(n15368), .ZN(n15369) );
  AOI21_X1 U17338 ( .B1(n19048), .B2(n17413), .A(n15369), .ZN(n15375) );
  AOI22_X1 U17339 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n19011), .B1(n19013), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n15372) );
  NAND2_X1 U17340 ( .A1(n19009), .A2(n15370), .ZN(n15371) );
  OAI211_X1 U17341 ( .C1(n19051), .C2(n20163), .A(n15372), .B(n15371), .ZN(
        n15373) );
  AOI21_X1 U17342 ( .B1(n19069), .B2(n19045), .A(n15373), .ZN(n15374) );
  OAI211_X1 U17343 ( .C1(n19674), .C2(n15581), .A(n15375), .B(n15374), .ZN(
        P2_U2855) );
  NAND3_X1 U17344 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n17517), .ZN(n16855) );
  INV_X1 U17345 ( .A(n16855), .ZN(n15384) );
  NOR2_X1 U17346 ( .A1(n15376), .A2(n16855), .ZN(n22568) );
  INV_X1 U17347 ( .A(n22568), .ZN(n15405) );
  OAI21_X1 U17348 ( .B1(n16852), .B2(n15377), .A(n15405), .ZN(n15385) );
  OR2_X1 U17349 ( .A1(n15378), .A2(n15385), .ZN(n15380) );
  OAI221_X1 U17350 ( .B1(n15381), .B2(n15384), .C1(n22290), .C2(n15380), .A(
        n15379), .ZN(n22570) );
  INV_X1 U17351 ( .A(n15382), .ZN(n15383) );
  INV_X1 U17352 ( .A(n22577), .ZN(n15404) );
  AOI22_X1 U17353 ( .A1(n15385), .A2(n22253), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15384), .ZN(n22418) );
  OAI22_X1 U17354 ( .A1(n15404), .A2(n22302), .B1(n22418), .B2(n16865), .ZN(
        n15390) );
  INV_X1 U17355 ( .A(n15386), .ZN(n15387) );
  OAI22_X1 U17356 ( .A1(n22573), .A2(n22267), .B1(n15405), .B2(n22266), .ZN(
        n15389) );
  AOI211_X1 U17357 ( .C1(n22570), .C2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n15390), .B(n15389), .ZN(n15391) );
  INV_X1 U17358 ( .A(n15391), .ZN(P1_U3137) );
  OAI22_X1 U17359 ( .A1(n15404), .A2(n22459), .B1(n22418), .B2(n16885), .ZN(
        n15393) );
  OAI22_X1 U17360 ( .A1(n22573), .A2(n22442), .B1(n22441), .B2(n15405), .ZN(
        n15392) );
  AOI211_X1 U17361 ( .C1(n22570), .C2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15393), .B(n15392), .ZN(n15394) );
  INV_X1 U17362 ( .A(n15394), .ZN(P1_U3142) );
  OAI22_X1 U17363 ( .A1(n15404), .A2(n22330), .B1(n22418), .B2(n16870), .ZN(
        n15396) );
  OAI22_X1 U17364 ( .A1(n22573), .A2(n22309), .B1(n15405), .B2(n22308), .ZN(
        n15395) );
  AOI211_X1 U17365 ( .C1(n22570), .C2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n15396), .B(n15395), .ZN(n15397) );
  INV_X1 U17366 ( .A(n15397), .ZN(P1_U3138) );
  OAI22_X1 U17367 ( .A1(n15404), .A2(n22473), .B1(n22418), .B2(n16892), .ZN(
        n15399) );
  OAI22_X1 U17368 ( .A1(n22573), .A2(n15712), .B1(n15405), .B2(n16889), .ZN(
        n15398) );
  AOI211_X1 U17369 ( .C1(n22570), .C2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n15399), .B(n15398), .ZN(n15400) );
  INV_X1 U17370 ( .A(n15400), .ZN(P1_U3143) );
  OAI22_X1 U17371 ( .A1(n15404), .A2(n22382), .B1(n22418), .B2(n16880), .ZN(
        n15402) );
  OAI22_X1 U17372 ( .A1(n22573), .A2(n22371), .B1(n15405), .B2(n22370), .ZN(
        n15401) );
  AOI211_X1 U17373 ( .C1(n22570), .C2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n15402), .B(n15401), .ZN(n15403) );
  INV_X1 U17374 ( .A(n15403), .ZN(P1_U3140) );
  OAI22_X1 U17375 ( .A1(n15404), .A2(n22359), .B1(n22418), .B2(n16875), .ZN(
        n15407) );
  OAI22_X1 U17376 ( .A1(n22573), .A2(n22342), .B1(n15405), .B2(n22341), .ZN(
        n15406) );
  AOI211_X1 U17377 ( .C1(n22570), .C2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n15407), .B(n15406), .ZN(n15408) );
  INV_X1 U17378 ( .A(n15408), .ZN(P1_U3139) );
  OAI222_X1 U17379 ( .A1(n15478), .A2(n22480), .B1(n16523), .B2(n12073), .C1(
        n16553), .C2(n15409), .ZN(P1_U2897) );
  INV_X1 U17380 ( .A(n22030), .ZN(n15437) );
  INV_X1 U17381 ( .A(n15410), .ZN(n22286) );
  INV_X1 U17382 ( .A(n15592), .ZN(n15433) );
  NAND2_X1 U17383 ( .A1(n22118), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n15412) );
  INV_X1 U17384 ( .A(n15842), .ZN(n15669) );
  AOI22_X1 U17385 ( .A1(n22134), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15669), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n15411) );
  OAI211_X1 U17386 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n22128), .A(
        n15412), .B(n15411), .ZN(n15416) );
  INV_X1 U17387 ( .A(n15413), .ZN(n15414) );
  OAI22_X1 U17388 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n22073), .B1(n22059), 
        .B2(n15414), .ZN(n15415) );
  AOI211_X1 U17389 ( .C1(n22286), .C2(n15433), .A(n15416), .B(n15415), .ZN(
        n15417) );
  OAI21_X1 U17390 ( .B1(n15418), .B2(n15437), .A(n15417), .ZN(P1_U2839) );
  INV_X1 U17391 ( .A(n15419), .ZN(n15430) );
  NAND2_X1 U17392 ( .A1(n15420), .A2(n22030), .ZN(n15429) );
  NAND2_X1 U17393 ( .A1(n22118), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U17394 ( .A1(n22134), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n15669), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n15421) );
  OAI211_X1 U17395 ( .C1(n22128), .C2(n15423), .A(n15422), .B(n15421), .ZN(
        n15427) );
  NAND2_X1 U17396 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n15425) );
  INV_X1 U17397 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20390) );
  NAND3_X1 U17398 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n15583) );
  INV_X1 U17399 ( .A(n15583), .ZN(n15424) );
  AOI211_X1 U17400 ( .C1(n15425), .C2(n20390), .A(n15424), .B(n22073), .ZN(
        n15426) );
  AOI211_X1 U17401 ( .C1(n22136), .C2(n21904), .A(n15427), .B(n15426), .ZN(
        n15428) );
  OAI211_X1 U17402 ( .C1(n15430), .C2(n15592), .A(n15429), .B(n15428), .ZN(
        P1_U2837) );
  NAND2_X1 U17403 ( .A1(n22073), .A2(n15842), .ZN(n22096) );
  NAND2_X1 U17404 ( .A1(n22118), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n15435) );
  OR2_X1 U17405 ( .A1(n22134), .A2(n22110), .ZN(n15431) );
  AOI22_X1 U17406 ( .A1(n15433), .A2(n15432), .B1(n15431), .B2(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15434) );
  OAI211_X1 U17407 ( .C1(n15436), .C2(n22059), .A(n15435), .B(n15434), .ZN(
        n15440) );
  NOR2_X1 U17408 ( .A1(n15438), .A2(n15437), .ZN(n15439) );
  AOI211_X1 U17409 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n22096), .A(n15440), .B(
        n15439), .ZN(n15441) );
  INV_X1 U17410 ( .A(n15441), .ZN(P1_U2840) );
  AOI21_X1 U17411 ( .B1(n15444), .B2(n15325), .A(n15443), .ZN(n15613) );
  INV_X1 U17412 ( .A(n15613), .ZN(n15480) );
  INV_X1 U17413 ( .A(n15611), .ZN(n15460) );
  INV_X1 U17414 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22050) );
  INV_X1 U17415 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n22039) );
  INV_X1 U17416 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20392) );
  NOR2_X1 U17417 ( .A1(n20392), .A2(n15583), .ZN(n22023) );
  NAND2_X1 U17418 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22023), .ZN(n22040) );
  NOR3_X1 U17419 ( .A1(n22050), .A2(n22039), .A3(n22040), .ZN(n15445) );
  NAND2_X1 U17420 ( .A1(n22024), .A2(n15445), .ZN(n15458) );
  INV_X1 U17421 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20398) );
  NAND2_X1 U17422 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n15445), .ZN(n15667) );
  OAI21_X1 U17423 ( .B1(n15667), .B2(n22073), .A(n22096), .ZN(n15601) );
  INV_X1 U17424 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U17425 ( .A1(n14072), .A2(n21943), .ZN(n15448) );
  NAND2_X1 U17426 ( .A1(n16206), .A2(n15462), .ZN(n15447) );
  NAND3_X1 U17427 ( .A1(n15448), .A2(n16261), .A3(n15447), .ZN(n15449) );
  NAND2_X1 U17428 ( .A1(n15450), .A2(n15449), .ZN(n15453) );
  OR2_X1 U17429 ( .A1(n15453), .A2(n15454), .ZN(n15455) );
  NAND2_X1 U17430 ( .A1(n15455), .A2(n15598), .ZN(n21948) );
  OAI22_X1 U17431 ( .A1(n22131), .A2(n15462), .B1(n22059), .B2(n21948), .ZN(
        n15456) );
  AOI211_X1 U17432 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n22100), .B(n15456), .ZN(n15457) );
  OAI221_X1 U17433 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n15458), .C1(n20398), 
        .C2(n15601), .A(n15457), .ZN(n15459) );
  AOI21_X1 U17434 ( .B1(n22110), .B2(n15460), .A(n15459), .ZN(n15461) );
  OAI21_X1 U17435 ( .B1(n15480), .B2(n22114), .A(n15461), .ZN(P1_U2832) );
  OAI22_X1 U17436 ( .A1(n16453), .A2(n21948), .B1(n15462), .B2(n16451), .ZN(
        n15463) );
  INV_X1 U17437 ( .A(n15463), .ZN(n15464) );
  OAI21_X1 U17438 ( .B1(n15480), .B2(n16425), .A(n15464), .ZN(P1_U2864) );
  XNOR2_X1 U17439 ( .A(n15503), .B(n15516), .ZN(n15505) );
  XNOR2_X1 U17440 ( .A(n15505), .B(n15504), .ZN(n15489) );
  XOR2_X1 U17441 ( .A(n15466), .B(n15465), .Z(n15486) );
  NOR2_X1 U17442 ( .A1(n17319), .A2(n15470), .ZN(n15467) );
  NOR2_X1 U17443 ( .A1(n15468), .A2(n15467), .ZN(n17388) );
  OAI211_X1 U17444 ( .C1(n15470), .C2(n15469), .A(n15516), .B(n17365), .ZN(
        n15472) );
  NAND2_X1 U17445 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19139), .ZN(n15471) );
  OAI211_X1 U17446 ( .C1(n15473), .C2(n19133), .A(n15472), .B(n15471), .ZN(
        n15474) );
  AOI21_X1 U17447 ( .B1(n20009), .B2(n19129), .A(n15474), .ZN(n15475) );
  OAI21_X1 U17448 ( .B1(n17388), .B2(n15516), .A(n15475), .ZN(n15476) );
  AOI21_X1 U17449 ( .B1(n15486), .B2(n19108), .A(n15476), .ZN(n15477) );
  OAI21_X1 U17450 ( .B1(n15489), .B2(n19091), .A(n15477), .ZN(P2_U3043) );
  INV_X1 U17451 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15479) );
  OAI222_X1 U17452 ( .A1(n15480), .A2(n16553), .B1(n16523), .B2(n15479), .C1(
        n16501), .C2(n15478), .ZN(P1_U2896) );
  OAI22_X1 U17453 ( .A1(n17633), .A2(n15482), .B1(n15481), .B2(n18813), .ZN(
        n15485) );
  NOR2_X1 U17454 ( .A1(n17681), .A2(n15483), .ZN(n15484) );
  AOI211_X1 U17455 ( .C1(n17673), .C2(n14255), .A(n15485), .B(n15484), .ZN(
        n15488) );
  NAND2_X1 U17456 ( .A1(n15486), .A2(n17664), .ZN(n15487) );
  OAI211_X1 U17457 ( .C1(n15489), .C2(n17608), .A(n15488), .B(n15487), .ZN(
        P2_U3011) );
  NAND2_X1 U17458 ( .A1(n15491), .A2(n15490), .ZN(n15492) );
  NAND2_X1 U17459 ( .A1(n15545), .A2(n15492), .ZN(n18823) );
  NOR2_X1 U17460 ( .A1(n15494), .A2(n15493), .ZN(n15500) );
  NAND2_X1 U17461 ( .A1(n15495), .A2(n15499), .ZN(n15496) );
  INV_X1 U17462 ( .A(n15619), .ZN(n15498) );
  OAI211_X1 U17463 ( .C1(n15500), .C2(n15499), .A(n15498), .B(n15746), .ZN(
        n15502) );
  NAND2_X1 U17464 ( .A1(n16966), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15501) );
  OAI211_X1 U17465 ( .C1(n18823), .C2(n16966), .A(n15502), .B(n15501), .ZN(
        P2_U2875) );
  AOI22_X1 U17466 ( .A1(n15505), .A2(n15504), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15503), .ZN(n15507) );
  XNOR2_X1 U17467 ( .A(n18734), .B(n15686), .ZN(n15506) );
  XNOR2_X1 U17468 ( .A(n15507), .B(n15506), .ZN(n15523) );
  OAI21_X1 U17469 ( .B1(n15509), .B2(n15686), .A(n15508), .ZN(n15521) );
  OAI22_X1 U17470 ( .A1(n15510), .A2(n17633), .B1(n13221), .B2(n18813), .ZN(
        n15511) );
  AOI21_X1 U17471 ( .B1(n17640), .B2(n18740), .A(n15511), .ZN(n15512) );
  OAI21_X1 U17472 ( .B1(n17657), .B2(n18743), .A(n15512), .ZN(n15513) );
  AOI21_X1 U17473 ( .B1(n15521), .B2(n17664), .A(n15513), .ZN(n15514) );
  OAI21_X1 U17474 ( .B1(n15523), .B2(n17608), .A(n15514), .ZN(P2_U3010) );
  NOR2_X1 U17475 ( .A1(n15516), .A2(n15515), .ZN(n15684) );
  OAI21_X1 U17476 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19109), .A(
        n17388), .ZN(n15688) );
  NOR2_X1 U17477 ( .A1(n13221), .A2(n18813), .ZN(n15517) );
  AOI221_X1 U17478 ( .B1(n15684), .B2(n15686), .C1(n15688), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n15517), .ZN(n15518) );
  INV_X1 U17479 ( .A(n15518), .ZN(n15520) );
  OAI22_X1 U17480 ( .A1(n18743), .A2(n19133), .B1(n19119), .B2(n18730), .ZN(
        n15519) );
  AOI211_X1 U17481 ( .C1(n15521), .C2(n19108), .A(n15520), .B(n15519), .ZN(
        n15522) );
  OAI21_X1 U17482 ( .B1(n15523), .B2(n19091), .A(n15522), .ZN(P2_U3042) );
  NAND2_X1 U17483 ( .A1(n22500), .A2(n22493), .ZN(n15524) );
  NAND2_X1 U17484 ( .A1(n15524), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15525) );
  NAND2_X1 U17485 ( .A1(n15525), .A2(n22253), .ZN(n15529) );
  OR2_X1 U17486 ( .A1(n22239), .A2(n15410), .ZN(n15531) );
  INV_X1 U17487 ( .A(n22240), .ZN(n16854) );
  NAND2_X1 U17488 ( .A1(n16854), .A2(n17526), .ZN(n15698) );
  NAND2_X1 U17489 ( .A1(n15528), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22274) );
  OR2_X1 U17490 ( .A1(n15698), .A2(n22274), .ZN(n15526) );
  NOR2_X1 U17491 ( .A1(n15528), .A2(n12293), .ZN(n15697) );
  INV_X1 U17492 ( .A(n15529), .ZN(n15532) );
  OR2_X1 U17493 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15530), .ZN(
        n22492) );
  AOI22_X1 U17494 ( .A1(n15532), .A2(n15531), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22492), .ZN(n15533) );
  NAND2_X1 U17495 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15698), .ZN(n15704) );
  NAND3_X1 U17496 ( .A1(n22278), .A2(n15533), .A3(n15704), .ZN(n22496) );
  NAND2_X1 U17497 ( .A1(n22496), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n15536) );
  OAI22_X1 U17498 ( .A1(n22500), .A2(n22473), .B1(n22492), .B2(n16889), .ZN(
        n15534) );
  AOI21_X1 U17499 ( .B1(n22487), .B2(n22470), .A(n15534), .ZN(n15535) );
  OAI211_X1 U17500 ( .C1(n15543), .C2(n16892), .A(n15536), .B(n15535), .ZN(
        P1_U3055) );
  NAND2_X1 U17501 ( .A1(n22496), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n15539) );
  OAI22_X1 U17502 ( .A1(n22500), .A2(n22330), .B1(n22492), .B2(n22308), .ZN(
        n15537) );
  AOI21_X1 U17503 ( .B1(n22487), .B2(n22327), .A(n15537), .ZN(n15538) );
  OAI211_X1 U17504 ( .C1(n15543), .C2(n16870), .A(n15539), .B(n15538), .ZN(
        P1_U3050) );
  NAND2_X1 U17505 ( .A1(n22496), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n15542) );
  OAI22_X1 U17506 ( .A1(n22500), .A2(n22302), .B1(n22266), .B2(n22492), .ZN(
        n15540) );
  AOI21_X1 U17507 ( .B1(n22487), .B2(n22299), .A(n15540), .ZN(n15541) );
  OAI211_X1 U17508 ( .C1(n15543), .C2(n16865), .A(n15542), .B(n15541), .ZN(
        P1_U3049) );
  XNOR2_X1 U17509 ( .A(n15619), .B(n15621), .ZN(n15549) );
  INV_X1 U17510 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n15564) );
  AND2_X1 U17511 ( .A1(n15545), .A2(n15544), .ZN(n15547) );
  OR2_X1 U17512 ( .A1(n15547), .A2(n15546), .ZN(n17336) );
  MUX2_X1 U17513 ( .A(n15564), .B(n17336), .S(n16952), .Z(n15548) );
  OAI21_X1 U17514 ( .B1(n15549), .B2(n16968), .A(n15548), .ZN(P2_U2874) );
  AOI21_X1 U17515 ( .B1(n17614), .B2(n15550), .A(n17616), .ZN(n17605) );
  INV_X1 U17516 ( .A(n17605), .ZN(n18832) );
  OAI21_X1 U17517 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15558), .A(
        n15550), .ZN(n17604) );
  INV_X1 U17518 ( .A(n17604), .ZN(n18818) );
  OAI21_X1 U17519 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15555), .A(
        n11255), .ZN(n17592) );
  INV_X1 U17520 ( .A(n17592), .ZN(n18796) );
  AOI21_X1 U17521 ( .B1(n17578), .B2(n15553), .A(n15557), .ZN(n18770) );
  AOI21_X1 U17522 ( .B1(n17167), .B2(n15551), .A(n15554), .ZN(n18750) );
  NAND2_X1 U17523 ( .A1(n15552), .A2(n17567), .ZN(n18748) );
  NOR2_X1 U17524 ( .A1(n18750), .A2(n18748), .ZN(n18755) );
  OAI21_X1 U17525 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n15554), .A(
        n15553), .ZN(n18757) );
  NAND2_X1 U17526 ( .A1(n18755), .A2(n18757), .ZN(n18768) );
  NOR2_X1 U17527 ( .A1(n18770), .A2(n18768), .ZN(n18777) );
  INV_X1 U17528 ( .A(n15555), .ZN(n15556) );
  OAI21_X1 U17529 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n15557), .A(
        n15556), .ZN(n18780) );
  NAND2_X1 U17530 ( .A1(n18777), .A2(n18780), .ZN(n18794) );
  NOR2_X1 U17531 ( .A1(n18796), .A2(n18794), .ZN(n18808) );
  AOI21_X1 U17532 ( .B1(n18801), .B2(n11255), .A(n15558), .ZN(n17593) );
  INV_X1 U17533 ( .A(n17593), .ZN(n18811) );
  NAND2_X1 U17534 ( .A1(n18808), .A2(n18811), .ZN(n18816) );
  NOR2_X1 U17535 ( .A1(n18818), .A2(n18816), .ZN(n18833) );
  NOR2_X1 U17536 ( .A1(n18778), .A2(n18833), .ZN(n15559) );
  XNOR2_X1 U17537 ( .A(n18832), .B(n15559), .ZN(n15563) );
  OAI21_X1 U17538 ( .B1(n15560), .B2(n15561), .A(n18828), .ZN(n19642) );
  OAI22_X1 U17539 ( .A1(n17336), .A2(n19008), .B1(n19642), .B2(n19051), .ZN(
        n15562) );
  AOI21_X1 U17540 ( .B1(n15563), .B2(n19003), .A(n15562), .ZN(n15569) );
  OAI21_X1 U17541 ( .B1(n19040), .B2(n15564), .A(n18892), .ZN(n15567) );
  OAI22_X1 U17542 ( .A1(n17614), .A2(n19036), .B1(n15565), .B2(n19037), .ZN(
        n15566) );
  AOI211_X1 U17543 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n19011), .A(n15567), 
        .B(n15566), .ZN(n15568) );
  NAND2_X1 U17544 ( .A1(n15569), .A2(n15568), .ZN(P2_U2842) );
  AOI21_X1 U17545 ( .B1(n17413), .B2(n15571), .A(n15570), .ZN(n17414) );
  NAND2_X1 U17546 ( .A1(n17414), .A2(n19003), .ZN(n15580) );
  AOI22_X1 U17547 ( .A1(n19011), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n19014), 
        .B2(n20111), .ZN(n15573) );
  MUX2_X1 U17548 ( .A(n18875), .B(n19036), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15572) );
  OAI211_X1 U17549 ( .C1(n19040), .C2(n15574), .A(n15573), .B(n15572), .ZN(
        n15577) );
  NOR2_X1 U17550 ( .A1(n19008), .A2(n15575), .ZN(n15576) );
  AOI211_X1 U17551 ( .C1(n19009), .C2(n15578), .A(n15577), .B(n15576), .ZN(
        n15579) );
  OAI211_X1 U17552 ( .C1(n17690), .C2(n15581), .A(n15580), .B(n15579), .ZN(
        P2_U2854) );
  NAND2_X1 U17553 ( .A1(n20471), .A2(n22030), .ZN(n15591) );
  OAI21_X1 U17554 ( .B1(n22073), .B2(n22023), .A(n15842), .ZN(n22029) );
  NOR2_X1 U17555 ( .A1(n22059), .A2(n21902), .ZN(n15586) );
  OAI22_X1 U17556 ( .A1(n15582), .A2(n22113), .B1(n22128), .B2(n20474), .ZN(
        n15585) );
  NOR3_X1 U17557 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22073), .A3(n15583), .ZN(
        n15584) );
  NOR4_X1 U17558 ( .A1(n15586), .A2(n15585), .A3(n22100), .A4(n15584), .ZN(
        n15587) );
  OAI21_X1 U17559 ( .B1(n22131), .B2(n15588), .A(n15587), .ZN(n15589) );
  AOI21_X1 U17560 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n22029), .A(n15589), .ZN(
        n15590) );
  OAI211_X1 U17561 ( .C1(n22144), .C2(n15592), .A(n15591), .B(n15590), .ZN(
        P1_U2836) );
  INV_X1 U17562 ( .A(n15593), .ZN(n15594) );
  OAI21_X1 U17563 ( .B1(n15443), .B2(n15595), .A(n15594), .ZN(n15774) );
  AOI22_X1 U17564 ( .A1(n16551), .A2(n16495), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16549), .ZN(n15596) );
  OAI21_X1 U17565 ( .B1(n15774), .B2(n16553), .A(n15596), .ZN(P1_U2895) );
  INV_X1 U17566 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20400) );
  MUX2_X1 U17567 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n15597) );
  OAI21_X1 U17568 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16210), .A(
        n15597), .ZN(n15599) );
  AOI21_X1 U17569 ( .B1(n15599), .B2(n15598), .A(n15663), .ZN(n21953) );
  AOI22_X1 U17570 ( .A1(n22136), .A2(n21953), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n22134), .ZN(n15600) );
  OAI21_X1 U17571 ( .B1(n20400), .B2(n15601), .A(n15600), .ZN(n15605) );
  NOR3_X1 U17572 ( .A1(n22073), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n15667), .ZN(
        n15604) );
  INV_X1 U17573 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15654) );
  AOI21_X1 U17574 ( .B1(n15777), .B2(n22110), .A(n22100), .ZN(n15602) );
  OAI21_X1 U17575 ( .B1(n22131), .B2(n15654), .A(n15602), .ZN(n15603) );
  NOR3_X1 U17576 ( .A1(n15605), .A2(n15604), .A3(n15603), .ZN(n15606) );
  OAI21_X1 U17577 ( .B1(n15774), .B2(n22114), .A(n15606), .ZN(P1_U2831) );
  OAI21_X1 U17578 ( .B1(n15609), .B2(n15608), .A(n15607), .ZN(n21940) );
  AOI22_X1 U17579 ( .A1(n20514), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n22016), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15610) );
  OAI21_X1 U17580 ( .B1(n20522), .B2(n15611), .A(n15610), .ZN(n15612) );
  AOI21_X1 U17581 ( .B1(n15613), .B2(n20519), .A(n15612), .ZN(n15614) );
  OAI21_X1 U17582 ( .B1(n21940), .B2(n22141), .A(n15614), .ZN(P1_U2991) );
  NOR2_X1 U17583 ( .A1(n15546), .A2(n15616), .ZN(n15617) );
  OR2_X1 U17584 ( .A1(n15615), .A2(n15617), .ZN(n19090) );
  AND2_X1 U17585 ( .A1(n15621), .A2(n15620), .ZN(n15618) );
  AOI21_X1 U17586 ( .B1(n15619), .B2(n15621), .A(n15620), .ZN(n15622) );
  OR3_X1 U17587 ( .A1(n11623), .A2(n15622), .A3(n16968), .ZN(n15624) );
  NAND2_X1 U17588 ( .A1(n16966), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15623) );
  OAI211_X1 U17589 ( .C1(n19090), .C2(n16966), .A(n15624), .B(n15623), .ZN(
        P2_U2873) );
  OAI211_X1 U17590 ( .C1(n11623), .C2(n15627), .A(n15746), .B(n15743), .ZN(
        n15632) );
  NOR2_X1 U17591 ( .A1(n15615), .A2(n15629), .ZN(n15630) );
  NOR2_X1 U17592 ( .A1(n15628), .A2(n15630), .ZN(n18844) );
  NAND2_X1 U17593 ( .A1(n18844), .A2(n16952), .ZN(n15631) );
  OAI211_X1 U17594 ( .C1(n16952), .C2(n13477), .A(n15632), .B(n15631), .ZN(
        P2_U2872) );
  NOR2_X1 U17595 ( .A1(n15633), .A2(n19754), .ZN(n17426) );
  AOI21_X1 U17596 ( .B1(n20204), .B2(n20197), .A(n22169), .ZN(n15634) );
  AOI21_X1 U17597 ( .B1(n17426), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n15634), .ZN(n15642) );
  NAND3_X1 U17598 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19807), .ZN(n19692) );
  NOR2_X1 U17599 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19692), .ZN(
        n20198) );
  AOI21_X1 U17600 ( .B1(n15237), .B2(n19734), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19165) );
  NAND2_X1 U17601 ( .A1(n15636), .A2(n19165), .ZN(n15638) );
  INV_X1 U17602 ( .A(n19799), .ZN(n19841) );
  INV_X1 U17603 ( .A(n15644), .ZN(n15639) );
  NOR2_X1 U17604 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n15638), .ZN(n19842) );
  INV_X1 U17605 ( .A(n19842), .ZN(n19823) );
  NOR2_X1 U17606 ( .A1(n15639), .A2(n19823), .ZN(n15640) );
  AOI211_X1 U17607 ( .C1(n20198), .C2(n19846), .A(n19841), .B(n15640), .ZN(
        n15641) );
  INV_X1 U17608 ( .A(n20201), .ZN(n15680) );
  INV_X1 U17609 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15653) );
  INV_X1 U17610 ( .A(n15643), .ZN(n15647) );
  INV_X1 U17611 ( .A(n17426), .ZN(n15646) );
  OAI21_X1 U17612 ( .B1(n15644), .B2(n20198), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15645) );
  OAI21_X1 U17613 ( .B1(n15647), .B2(n15646), .A(n15645), .ZN(n20199) );
  INV_X1 U17614 ( .A(n19854), .ZN(n19861) );
  INV_X1 U17615 ( .A(n20176), .ZN(n17431) );
  NAND2_X1 U17616 ( .A1(n15649), .A2(n17431), .ZN(n19864) );
  INV_X1 U17617 ( .A(n20198), .ZN(n15677) );
  AOI22_X1 U17618 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n11151), .ZN(n19902) );
  AOI22_X1 U17619 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n11151), .ZN(n19895) );
  INV_X1 U17620 ( .A(n19895), .ZN(n19899) );
  AOI22_X1 U17621 ( .A1(n20208), .A2(n19892), .B1(n20200), .B2(n19899), .ZN(
        n15650) );
  OAI21_X1 U17622 ( .B1(n19864), .B2(n15677), .A(n15650), .ZN(n15651) );
  AOI21_X1 U17623 ( .B1(n20199), .B2(n15648), .A(n15651), .ZN(n15652) );
  OAI21_X1 U17624 ( .B1(n15680), .B2(n15653), .A(n15652), .ZN(P2_U3150) );
  INV_X1 U17625 ( .A(n21953), .ZN(n15655) );
  OAI222_X1 U17626 ( .A1(n15655), .A2(n16453), .B1(n15654), .B2(n16451), .C1(
        n16425), .C2(n15774), .ZN(P1_U2863) );
  OAI21_X1 U17627 ( .B1(n15593), .B2(n15656), .A(n11586), .ZN(n16683) );
  INV_X1 U17628 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15658) );
  OAI21_X1 U17629 ( .B1(n15657), .B2(n15658), .A(n14072), .ZN(n15659) );
  OAI21_X1 U17630 ( .B1(n16209), .B2(P1_EBX_REG_10__SCAN_IN), .A(n15659), .ZN(
        n15661) );
  NAND2_X1 U17631 ( .A1(n15661), .A2(n15660), .ZN(n15662) );
  OR2_X1 U17632 ( .A1(n15662), .A2(n15663), .ZN(n15664) );
  NAND2_X1 U17633 ( .A1(n15664), .A2(n15768), .ZN(n21962) );
  NOR2_X1 U17634 ( .A1(n22128), .A2(n16678), .ZN(n15665) );
  AOI211_X1 U17635 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n22100), .B(n15665), .ZN(n15666) );
  OAI21_X1 U17636 ( .B1(n22059), .B2(n21962), .A(n15666), .ZN(n15672) );
  INV_X1 U17637 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n22064) );
  NOR2_X1 U17638 ( .A1(n20400), .A2(n15667), .ZN(n15668) );
  NAND2_X1 U17639 ( .A1(n22024), .A2(n15668), .ZN(n22063) );
  NAND2_X1 U17640 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15668), .ZN(n15841) );
  AOI21_X1 U17641 ( .B1(n22024), .B2(n15841), .A(n15669), .ZN(n15670) );
  AOI21_X1 U17642 ( .B1(n22064), .B2(n22063), .A(n15670), .ZN(n15671) );
  AOI211_X1 U17643 ( .C1(P1_EBX_REG_10__SCAN_IN), .C2(n22118), .A(n15672), .B(
        n15671), .ZN(n15673) );
  OAI21_X1 U17644 ( .B1(n16683), .B2(n22114), .A(n15673), .ZN(P1_U2830) );
  AOI22_X1 U17645 ( .A1(n16551), .A2(n16489), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16549), .ZN(n15674) );
  OAI21_X1 U17646 ( .B1(n16683), .B2(n16553), .A(n15674), .ZN(P1_U2894) );
  INV_X1 U17647 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15911) );
  NAND2_X1 U17648 ( .A1(n12815), .A2(n17431), .ZN(n19666) );
  INV_X1 U17649 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20596) );
  INV_X1 U17650 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19200) );
  OAI22_X2 U17651 ( .A1(n20596), .A2(n22599), .B1(n19200), .B2(n20065), .ZN(
        n19837) );
  INV_X1 U17652 ( .A(n19853), .ZN(n19803) );
  AOI22_X1 U17653 ( .A1(n20208), .A2(n19837), .B1(n20200), .B2(n19803), .ZN(
        n15676) );
  OAI21_X1 U17654 ( .B1(n19666), .B2(n15677), .A(n15676), .ZN(n15678) );
  AOI21_X1 U17655 ( .B1(n20199), .B2(n15675), .A(n15678), .ZN(n15679) );
  OAI21_X1 U17656 ( .B1(n15680), .B2(n15911), .A(n15679), .ZN(P2_U3151) );
  XNOR2_X1 U17657 ( .A(n15681), .B(n15685), .ZN(n17562) );
  XNOR2_X1 U17658 ( .A(n15682), .B(n15683), .ZN(n17561) );
  OAI221_X1 U17659 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15686), .C2(n15685), .A(
        n15684), .ZN(n15692) );
  INV_X1 U17660 ( .A(n15687), .ZN(n17564) );
  AOI22_X1 U17661 ( .A1(n19139), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15688), .ZN(n15689) );
  OAI21_X1 U17662 ( .B1(n19119), .B2(n19909), .A(n15689), .ZN(n15690) );
  AOI21_X1 U17663 ( .B1(n17564), .B2(n19103), .A(n15690), .ZN(n15691) );
  OAI211_X1 U17664 ( .C1(n17561), .C2(n19091), .A(n15692), .B(n15691), .ZN(
        n15693) );
  INV_X1 U17665 ( .A(n15693), .ZN(n15694) );
  OAI21_X1 U17666 ( .B1(n19134), .B2(n17562), .A(n15694), .ZN(P2_U3041) );
  OAI222_X1 U17667 ( .A1(n21962), .A2(n16453), .B1(n15695), .B2(n16451), .C1(
        n16683), .C2(n16425), .ZN(P1_U2862) );
  NOR3_X1 U17668 ( .A1(n22396), .A2(n22530), .A3(n22290), .ZN(n15696) );
  NOR2_X1 U17669 ( .A1(n22290), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22236) );
  NOR2_X1 U17670 ( .A1(n15696), .A2(n22236), .ZN(n15700) );
  NAND2_X1 U17671 ( .A1(n22258), .A2(n22286), .ZN(n15702) );
  INV_X1 U17672 ( .A(n15697), .ZN(n22289) );
  OAI22_X1 U17673 ( .A1(n15700), .A2(n15702), .B1(n15698), .B2(n22289), .ZN(
        n22523) );
  INV_X1 U17674 ( .A(n22523), .ZN(n15717) );
  AND2_X1 U17675 ( .A1(n22274), .A2(n15699), .ZN(n22297) );
  INV_X1 U17676 ( .A(n15700), .ZN(n15703) );
  NOR2_X1 U17677 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15701), .ZN(
        n15714) );
  INV_X1 U17678 ( .A(n15714), .ZN(n22520) );
  AOI22_X1 U17679 ( .A1(n15703), .A2(n15702), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22520), .ZN(n15705) );
  NAND3_X1 U17680 ( .A1(n22297), .A2(n15705), .A3(n15704), .ZN(n22524) );
  NAND2_X1 U17681 ( .A1(n22524), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n15708) );
  OAI22_X1 U17682 ( .A1(n22330), .A2(n22527), .B1(n22521), .B2(n22309), .ZN(
        n15706) );
  AOI21_X1 U17683 ( .B1(n22326), .B2(n15714), .A(n15706), .ZN(n15707) );
  OAI211_X1 U17684 ( .C1(n15717), .C2(n16870), .A(n15708), .B(n15707), .ZN(
        P1_U3082) );
  NAND2_X1 U17685 ( .A1(n22524), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n15711) );
  OAI22_X1 U17686 ( .A1(n22459), .A2(n22527), .B1(n22521), .B2(n22442), .ZN(
        n15709) );
  AOI21_X1 U17687 ( .B1(n15714), .B2(n22455), .A(n15709), .ZN(n15710) );
  OAI211_X1 U17688 ( .C1(n15717), .C2(n16885), .A(n15711), .B(n15710), .ZN(
        P1_U3086) );
  NAND2_X1 U17689 ( .A1(n22524), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n15716) );
  OAI22_X1 U17690 ( .A1(n22473), .A2(n22527), .B1(n22521), .B2(n15712), .ZN(
        n15713) );
  AOI21_X1 U17691 ( .B1(n22468), .B2(n15714), .A(n15713), .ZN(n15715) );
  OAI211_X1 U17692 ( .C1(n15717), .C2(n16892), .A(n15716), .B(n15715), .ZN(
        P1_U3087) );
  NOR3_X1 U17693 ( .A1(n22556), .A2(n22548), .A3(n22290), .ZN(n15718) );
  NOR2_X1 U17694 ( .A1(n15718), .A2(n22236), .ZN(n15721) );
  OR2_X1 U17695 ( .A1(n15719), .A2(n15410), .ZN(n15722) );
  NAND2_X1 U17696 ( .A1(n16854), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22288) );
  INV_X1 U17697 ( .A(n22549), .ZN(n15729) );
  INV_X1 U17698 ( .A(n22371), .ZN(n22379) );
  NOR2_X1 U17699 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15720), .ZN(
        n22547) );
  INV_X1 U17700 ( .A(n22547), .ZN(n15724) );
  INV_X1 U17701 ( .A(n15721), .ZN(n15723) );
  AOI22_X1 U17702 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15724), .B1(n15723), 
        .B2(n15722), .ZN(n15725) );
  NAND2_X1 U17703 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22288), .ZN(n22296) );
  NAND3_X1 U17704 ( .A1(n22278), .A2(n15725), .A3(n22296), .ZN(n22550) );
  AOI22_X1 U17705 ( .A1(n22378), .A2(n22547), .B1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n22550), .ZN(n15726) );
  OAI21_X1 U17706 ( .B1(n22553), .B2(n22382), .A(n15726), .ZN(n15727) );
  AOI21_X1 U17707 ( .B1(n22548), .B2(n22379), .A(n15727), .ZN(n15728) );
  OAI21_X1 U17708 ( .B1(n15729), .B2(n16880), .A(n15728), .ZN(P1_U3116) );
  OR2_X1 U17709 ( .A1(n15628), .A2(n15730), .ZN(n15732) );
  INV_X1 U17710 ( .A(n15791), .ZN(n15731) );
  NAND2_X1 U17711 ( .A1(n15732), .A2(n15731), .ZN(n19122) );
  AOI22_X1 U17712 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n13303), .B1(
        n13304), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15736) );
  AOI22_X1 U17713 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15735) );
  AOI22_X1 U17714 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U17715 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15733) );
  NAND4_X1 U17716 ( .A1(n15736), .A2(n15735), .A3(n15734), .A4(n15733), .ZN(
        n15742) );
  AOI22_X1 U17717 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15740) );
  AOI22_X1 U17718 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15739) );
  AOI22_X1 U17719 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15738) );
  AOI22_X1 U17720 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15737) );
  NAND4_X1 U17721 ( .A1(n15740), .A2(n15739), .A3(n15738), .A4(n15737), .ZN(
        n15741) );
  NOR2_X1 U17722 ( .A1(n15742), .A2(n15741), .ZN(n15744) );
  AND2_X1 U17723 ( .A1(n15743), .A2(n15744), .ZN(n15745) );
  NOR2_X1 U17724 ( .A1(n11240), .A2(n15745), .ZN(n15758) );
  NAND2_X1 U17725 ( .A1(n15758), .A2(n15746), .ZN(n15748) );
  NAND2_X1 U17726 ( .A1(n16966), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15747) );
  OAI211_X1 U17727 ( .C1(n19122), .C2(n16966), .A(n15748), .B(n15747), .ZN(
        P2_U2871) );
  XNOR2_X1 U17728 ( .A(n17315), .B(n15749), .ZN(n19120) );
  NOR2_X2 U17729 ( .A1(n15754), .A2(n15750), .ZN(n19957) );
  INV_X1 U17730 ( .A(n19955), .ZN(n15752) );
  OAI22_X1 U17731 ( .A1(n15752), .A2(n20175), .B1(n15751), .B2(n20162), .ZN(
        n15757) );
  NOR2_X2 U17732 ( .A1(n15754), .A2(n15753), .ZN(n19956) );
  INV_X1 U17733 ( .A(n19956), .ZN(n16972) );
  INV_X1 U17734 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n15755) );
  NOR2_X1 U17735 ( .A1(n16972), .A2(n15755), .ZN(n15756) );
  AOI211_X1 U17736 ( .C1(BUF1_REG_16__SCAN_IN), .C2(n19957), .A(n15757), .B(
        n15756), .ZN(n15760) );
  INV_X1 U17737 ( .A(n20115), .ZN(n20167) );
  NAND2_X1 U17738 ( .A1(n15758), .A2(n20167), .ZN(n15759) );
  OAI211_X1 U17739 ( .C1(n19120), .C2(n20164), .A(n15760), .B(n15759), .ZN(
        P2_U2903) );
  OR2_X1 U17740 ( .A1(n15763), .A2(n15762), .ZN(n15764) );
  NAND2_X1 U17741 ( .A1(n15761), .A2(n15764), .ZN(n15826) );
  XNOR2_X1 U17742 ( .A(n15826), .B(n15824), .ZN(n22066) );
  AOI22_X1 U17743 ( .A1(n16551), .A2(n16482), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n16549), .ZN(n15765) );
  OAI21_X1 U17744 ( .B1(n20495), .B2(n16553), .A(n15765), .ZN(P1_U2893) );
  OAI21_X1 U17745 ( .B1(n16209), .B2(P1_EBX_REG_11__SCAN_IN), .A(n14072), .ZN(
        n15767) );
  INV_X1 U17746 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16815) );
  NOR2_X1 U17747 ( .A1(n15657), .A2(n16815), .ZN(n15766) );
  OAI22_X1 U17748 ( .A1(n15767), .A2(n15766), .B1(n16199), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15769) );
  AOI21_X1 U17749 ( .B1(n15769), .B2(n15768), .A(n15874), .ZN(n22057) );
  AOI22_X1 U17750 ( .A1(n16463), .A2(n22057), .B1(n16462), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15770) );
  OAI21_X1 U17751 ( .B1(n20495), .B2(n16425), .A(n15770), .ZN(P1_U2861) );
  OAI21_X1 U17752 ( .B1(n15772), .B2(n15771), .A(n16676), .ZN(n21954) );
  INV_X1 U17753 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15773) );
  OAI22_X1 U17754 ( .A1(n16670), .A2(n15773), .B1(n22001), .B2(n20400), .ZN(
        n15776) );
  NOR2_X1 U17755 ( .A1(n15774), .A2(n20496), .ZN(n15775) );
  AOI211_X1 U17756 ( .C1(n20505), .C2(n15777), .A(n15776), .B(n15775), .ZN(
        n15778) );
  OAI21_X1 U17757 ( .B1(n22141), .B2(n21954), .A(n15778), .ZN(P1_U2990) );
  AOI22_X1 U17758 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13303), .B1(
        n13304), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U17759 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15781) );
  AOI22_X1 U17760 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15780) );
  AOI22_X1 U17761 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15779) );
  NAND4_X1 U17762 ( .A1(n15782), .A2(n15781), .A3(n15780), .A4(n15779), .ZN(
        n15788) );
  AOI22_X1 U17763 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U17764 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15785) );
  AOI22_X1 U17765 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15784) );
  AOI22_X1 U17766 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15783) );
  NAND4_X1 U17767 ( .A1(n15786), .A2(n15785), .A3(n15784), .A4(n15783), .ZN(
        n15787) );
  OR2_X1 U17768 ( .A1(n15788), .A2(n15787), .ZN(n15790) );
  INV_X1 U17769 ( .A(n15815), .ZN(n15789) );
  OAI21_X1 U17770 ( .B1(n11240), .B2(n15790), .A(n15789), .ZN(n15804) );
  OR2_X1 U17771 ( .A1(n15792), .A2(n15791), .ZN(n15793) );
  AND2_X1 U17772 ( .A1(n15854), .A2(n15793), .ZN(n19102) );
  NAND2_X1 U17773 ( .A1(n16952), .A2(n19102), .ZN(n15796) );
  INV_X1 U17774 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n15794) );
  OR2_X1 U17775 ( .A1(n16952), .A2(n15794), .ZN(n15795) );
  OAI211_X1 U17776 ( .C1(n15804), .C2(n16968), .A(n15796), .B(n15795), .ZN(
        P2_U2870) );
  XNOR2_X1 U17777 ( .A(n15797), .B(n11247), .ZN(n19104) );
  INV_X1 U17778 ( .A(n19104), .ZN(n15799) );
  OAI22_X1 U17779 ( .A1(n20164), .A2(n15799), .B1(n15798), .B2(n20162), .ZN(
        n15800) );
  AOI21_X1 U17780 ( .B1(n19955), .B2(n15801), .A(n15800), .ZN(n15803) );
  AOI22_X1 U17781 ( .A1(n19956), .A2(BUF2_REG_17__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15802) );
  OAI211_X1 U17782 ( .C1(n15804), .C2(n20115), .A(n15803), .B(n15802), .ZN(
        P2_U2902) );
  AOI22_X1 U17783 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n13303), .B1(
        n13304), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15808) );
  AOI22_X1 U17784 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15807) );
  AOI22_X1 U17785 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15806) );
  AOI22_X1 U17786 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15805) );
  NAND4_X1 U17787 ( .A1(n15808), .A2(n15807), .A3(n15806), .A4(n15805), .ZN(
        n15814) );
  AOI22_X1 U17788 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U17789 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15811) );
  AOI22_X1 U17790 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15810) );
  AOI22_X1 U17791 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15809) );
  NAND4_X1 U17792 ( .A1(n15812), .A2(n15811), .A3(n15810), .A4(n15809), .ZN(
        n15813) );
  OR2_X1 U17793 ( .A1(n15814), .A2(n15813), .ZN(n15816) );
  OAI21_X1 U17794 ( .B1(n15815), .B2(n15816), .A(n15889), .ZN(n15858) );
  OAI21_X1 U17795 ( .B1(n15818), .B2(n15817), .A(n11271), .ZN(n18883) );
  OAI22_X1 U17796 ( .A1(n20164), .A2(n18883), .B1(n15819), .B2(n20162), .ZN(
        n15820) );
  AOI21_X1 U17797 ( .B1(n19955), .B2(n15821), .A(n15820), .ZN(n15823) );
  AOI22_X1 U17798 ( .A1(n19956), .A2(BUF2_REG_18__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15822) );
  OAI211_X1 U17799 ( .C1(n15858), .C2(n20115), .A(n15823), .B(n15822), .ZN(
        P2_U2901) );
  INV_X1 U17800 ( .A(n15824), .ZN(n15825) );
  OAI21_X1 U17801 ( .B1(n15826), .B2(n15825), .A(n15761), .ZN(n15828) );
  NOR2_X1 U17802 ( .A1(n15828), .A2(n15827), .ZN(n15829) );
  AOI22_X1 U17803 ( .A1(n16551), .A2(n16475), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16549), .ZN(n15830) );
  OAI21_X1 U17804 ( .B1(n22083), .B2(n16553), .A(n15830), .ZN(P1_U2892) );
  MUX2_X1 U17805 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n15834) );
  OAI21_X1 U17806 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16210), .A(
        n15834), .ZN(n15838) );
  OAI21_X1 U17807 ( .B1(n15657), .B2(n16803), .A(n14072), .ZN(n15835) );
  OAI21_X1 U17808 ( .B1(n16209), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15835), .ZN(
        n15837) );
  NAND2_X1 U17809 ( .A1(n15837), .A2(n15836), .ZN(n15875) );
  AOI21_X1 U17810 ( .B1(n15838), .B2(n15876), .A(n15868), .ZN(n21862) );
  AOI22_X1 U17811 ( .A1(n16463), .A2(n21862), .B1(n16462), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15839) );
  OAI21_X1 U17812 ( .B1(n16675), .B2(n16425), .A(n15839), .ZN(P1_U2859) );
  AOI22_X1 U17813 ( .A1(n16551), .A2(n16468), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16549), .ZN(n15840) );
  OAI21_X1 U17814 ( .B1(n16675), .B2(n16553), .A(n15840), .ZN(P1_U2891) );
  INV_X1 U17815 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n22062) );
  NOR2_X1 U17816 ( .A1(n22062), .A2(n15841), .ZN(n22071) );
  OAI21_X1 U17817 ( .B1(n22071), .B2(n22073), .A(n15842), .ZN(n22076) );
  AOI21_X1 U17818 ( .B1(n22024), .B2(n20404), .A(n22076), .ZN(n15847) );
  INV_X1 U17819 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15844) );
  INV_X1 U17820 ( .A(n21862), .ZN(n15843) );
  OAI22_X1 U17821 ( .A1(n22131), .A2(n15844), .B1(n22059), .B2(n15843), .ZN(
        n15845) );
  AOI211_X1 U17822 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n22100), .B(n15845), .ZN(n15846) );
  OAI221_X1 U17823 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15859), .C1(n21853), 
        .C2(n15847), .A(n15846), .ZN(n15848) );
  AOI21_X1 U17824 ( .B1(n16672), .B2(n22110), .A(n15848), .ZN(n15849) );
  OAI21_X1 U17825 ( .B1(n16675), .B2(n22114), .A(n15849), .ZN(P1_U2827) );
  INV_X1 U17826 ( .A(n15850), .ZN(n16457) );
  OAI21_X1 U17827 ( .B1(n15831), .B2(n15851), .A(n16457), .ZN(n16661) );
  AOI22_X1 U17828 ( .A1(n16551), .A2(n16274), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16549), .ZN(n15852) );
  OAI21_X1 U17829 ( .B1(n16661), .B2(n16553), .A(n15852), .ZN(P1_U2890) );
  NAND2_X1 U17830 ( .A1(n15854), .A2(n15853), .ZN(n15855) );
  NAND2_X1 U17831 ( .A1(n15899), .A2(n15855), .ZN(n18884) );
  MUX2_X1 U17832 ( .A(n15856), .B(n18884), .S(n16952), .Z(n15857) );
  OAI21_X1 U17833 ( .B1(n15858), .B2(n16968), .A(n15857), .ZN(P2_U2869) );
  NAND2_X1 U17834 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15861), .ZN(n22087) );
  INV_X1 U17835 ( .A(n22087), .ZN(n15860) );
  NOR2_X1 U17836 ( .A1(n15860), .A2(n22125), .ZN(n22085) );
  OAI21_X1 U17837 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n15861), .A(n22085), 
        .ZN(n15873) );
  AOI21_X1 U17838 ( .B1(n22134), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n22100), .ZN(n15862) );
  OAI21_X1 U17839 ( .B1(n16657), .B2(n22128), .A(n15862), .ZN(n15871) );
  INV_X1 U17840 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15878) );
  NAND2_X1 U17841 ( .A1(n14072), .A2(n21867), .ZN(n15864) );
  NAND2_X1 U17842 ( .A1(n16206), .A2(n15878), .ZN(n15863) );
  NAND3_X1 U17843 ( .A1(n15864), .A2(n16261), .A3(n15863), .ZN(n15865) );
  NAND2_X1 U17844 ( .A1(n15866), .A2(n15865), .ZN(n15867) );
  OR2_X1 U17845 ( .A1(n15867), .A2(n15868), .ZN(n15869) );
  NAND2_X1 U17846 ( .A1(n15869), .A2(n16460), .ZN(n21876) );
  NOR2_X1 U17847 ( .A1(n22059), .A2(n21876), .ZN(n15870) );
  AOI211_X1 U17848 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n22118), .A(n15871), .B(
        n15870), .ZN(n15872) );
  OAI211_X1 U17849 ( .C1(n16661), .C2(n22114), .A(n15873), .B(n15872), .ZN(
        P1_U2826) );
  OR2_X1 U17850 ( .A1(n15875), .A2(n15874), .ZN(n15877) );
  NAND2_X1 U17851 ( .A1(n15877), .A2(n15876), .ZN(n22070) );
  OAI222_X1 U17852 ( .A1(n22070), .A2(n16453), .B1(n22078), .B2(n16451), .C1(
        n16425), .C2(n22083), .ZN(P1_U2860) );
  OAI222_X1 U17853 ( .A1(n21876), .A2(n16453), .B1(n15878), .B2(n16451), .C1(
        n16425), .C2(n16661), .ZN(P1_U2858) );
  AOI22_X1 U17854 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n13303), .B1(
        n13304), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15882) );
  AOI22_X1 U17855 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15881) );
  AOI22_X1 U17856 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15880) );
  AOI22_X1 U17857 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15879) );
  NAND4_X1 U17858 ( .A1(n15882), .A2(n15881), .A3(n15880), .A4(n15879), .ZN(
        n15888) );
  AOI22_X1 U17859 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15886) );
  AOI22_X1 U17860 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15885) );
  AOI22_X1 U17861 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15884) );
  AOI22_X1 U17862 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15883) );
  NAND4_X1 U17863 ( .A1(n15886), .A2(n15885), .A3(n15884), .A4(n15883), .ZN(
        n15887) );
  OAI21_X1 U17864 ( .B1(n15890), .B2(n11697), .A(n16044), .ZN(n15904) );
  XNOR2_X1 U17865 ( .A(n11288), .B(n11271), .ZN(n18896) );
  INV_X1 U17866 ( .A(n18896), .ZN(n15892) );
  OAI22_X1 U17867 ( .A1(n20164), .A2(n15892), .B1(n15891), .B2(n20162), .ZN(
        n15893) );
  AOI21_X1 U17868 ( .B1(n19955), .B2(n15894), .A(n15893), .ZN(n15896) );
  AOI22_X1 U17869 ( .A1(n19956), .A2(BUF2_REG_19__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15895) );
  OAI211_X1 U17870 ( .C1(n15904), .C2(n20115), .A(n15896), .B(n15895), .ZN(
        P2_U2900) );
  OR2_X1 U17871 ( .A1(n16952), .A2(n15897), .ZN(n15903) );
  NAND2_X1 U17872 ( .A1(n15899), .A2(n15898), .ZN(n15900) );
  AND2_X1 U17873 ( .A1(n15901), .A2(n15900), .ZN(n18897) );
  NAND2_X1 U17874 ( .A1(n16952), .A2(n18897), .ZN(n15902) );
  OAI211_X1 U17875 ( .C1(n15904), .C2(n16968), .A(n15903), .B(n15902), .ZN(
        P2_U2868) );
  OAI21_X1 U17876 ( .B1(n15905), .B2(n21296), .A(n21798), .ZN(n17475) );
  NOR2_X1 U17877 ( .A1(n18156), .A2(n17475), .ZN(n18043) );
  INV_X1 U17878 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21810) );
  NOR2_X1 U17879 ( .A1(n20664), .A2(n21810), .ZN(n18042) );
  NAND2_X1 U17880 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18042), .ZN(n21817) );
  NOR2_X1 U17881 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21823) );
  NOR2_X1 U17882 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21818), .ZN(
        n21822) );
  INV_X1 U17883 ( .A(n21822), .ZN(n21309) );
  OAI21_X1 U17884 ( .B1(n21823), .B2(n18042), .A(n21309), .ZN(n19206) );
  NAND2_X1 U17885 ( .A1(n21830), .A2(n19206), .ZN(n19366) );
  INV_X1 U17886 ( .A(n21817), .ZN(n17481) );
  NAND2_X1 U17887 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17481), .ZN(n17473) );
  OAI211_X1 U17888 ( .C1(n18043), .C2(n21817), .A(n19366), .B(n17473), .ZN(
        n17483) );
  INV_X1 U17889 ( .A(n17483), .ZN(n18629) );
  NAND2_X1 U17890 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18528) );
  INV_X1 U17891 ( .A(n18528), .ZN(n18582) );
  NOR2_X1 U17892 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18042), .ZN(n20602) );
  INV_X1 U17893 ( .A(n20602), .ZN(n15906) );
  NOR2_X1 U17894 ( .A1(n18582), .A2(n15906), .ZN(n17440) );
  AOI21_X1 U17895 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n17440), .ZN(n17441) );
  NOR2_X1 U17896 ( .A1(n18629), .A2(n17441), .ZN(n15908) );
  INV_X1 U17897 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n20675) );
  NOR3_X1 U17898 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n20675), .ZN(n19241) );
  INV_X1 U17899 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19234) );
  NAND2_X1 U17900 ( .A1(n19234), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19202) );
  NAND2_X1 U17901 ( .A1(n19202), .A2(n17483), .ZN(n17439) );
  OR2_X1 U17902 ( .A1(n19241), .A2(n17439), .ZN(n15907) );
  MUX2_X1 U17903 ( .A(n15908), .B(n15907), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U17904 ( .A1(n17754), .A2(n18035), .ZN(n17756) );
  INV_X1 U17905 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n21091) );
  INV_X1 U17906 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20682) );
  NOR2_X1 U17907 ( .A1(n21091), .A2(n20682), .ZN(n18032) );
  AOI21_X1 U17908 ( .B1(n18039), .B2(n18032), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n15909) );
  NOR2_X1 U17909 ( .A1(n17756), .A2(n15909), .ZN(n15910) );
  MUX2_X1 U17910 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B(n15910), .S(n18034), 
        .Z(P3_U2701) );
  OAI22_X1 U17911 ( .A1(n16120), .A2(n15913), .B1(n15912), .B2(n15911), .ZN(
        n15914) );
  INV_X1 U17912 ( .A(n15914), .ZN(n15918) );
  AOI22_X1 U17913 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15917) );
  AOI22_X1 U17914 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15916) );
  AOI22_X1 U17915 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15915) );
  NAND4_X1 U17916 ( .A1(n15918), .A2(n15917), .A3(n15916), .A4(n15915), .ZN(
        n15924) );
  AOI22_X1 U17917 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15922) );
  AOI22_X1 U17918 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15921) );
  AOI22_X1 U17919 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15920) );
  AOI22_X1 U17920 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15919) );
  NAND4_X1 U17921 ( .A1(n15922), .A2(n15921), .A3(n15920), .A4(n15919), .ZN(
        n15923) );
  OR2_X1 U17922 ( .A1(n15924), .A2(n15923), .ZN(n16070) );
  AOI22_X1 U17923 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15935) );
  AOI22_X1 U17924 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15933) );
  INV_X1 U17925 ( .A(n16134), .ZN(n16121) );
  INV_X1 U17926 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15930) );
  NAND2_X1 U17927 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n15929) );
  INV_X1 U17928 ( .A(n15926), .ZN(n15928) );
  NAND2_X1 U17929 ( .A1(n17422), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15927) );
  NAND2_X1 U17930 ( .A1(n15928), .A2(n15927), .ZN(n16133) );
  OAI211_X1 U17931 ( .C1(n16121), .C2(n15930), .A(n15929), .B(n16133), .ZN(
        n15931) );
  INV_X1 U17932 ( .A(n15931), .ZN(n15932) );
  NAND4_X1 U17933 ( .A1(n15935), .A2(n15934), .A3(n15933), .A4(n15932), .ZN(
        n15944) );
  AOI22_X1 U17934 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15942) );
  AOI22_X1 U17935 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15940) );
  INV_X1 U17936 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U17937 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n15936) );
  INV_X1 U17938 ( .A(n16133), .ZN(n16102) );
  OAI211_X1 U17939 ( .C1(n16121), .C2(n15937), .A(n15936), .B(n16102), .ZN(
        n15938) );
  INV_X1 U17940 ( .A(n15938), .ZN(n15939) );
  NAND4_X1 U17941 ( .A1(n15942), .A2(n15941), .A3(n15940), .A4(n15939), .ZN(
        n15943) );
  AND2_X1 U17942 ( .A1(n15944), .A2(n15943), .ZN(n16069) );
  AND2_X1 U17943 ( .A1(n16070), .A2(n16069), .ZN(n16071) );
  INV_X1 U17944 ( .A(n16071), .ZN(n16073) );
  AOI22_X1 U17945 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15952) );
  INV_X1 U17946 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15947) );
  INV_X1 U17947 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15945) );
  OR2_X1 U17948 ( .A1(n16121), .A2(n15945), .ZN(n15946) );
  OAI211_X1 U17949 ( .C1(n15947), .C2(n16124), .A(n15946), .B(n16133), .ZN(
        n15948) );
  INV_X1 U17950 ( .A(n15948), .ZN(n15950) );
  AOI22_X1 U17951 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12755), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15949) );
  NAND4_X1 U17952 ( .A1(n15952), .A2(n15951), .A3(n15950), .A4(n15949), .ZN(
        n15962) );
  AOI22_X1 U17953 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15960) );
  AOI22_X1 U17954 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15959) );
  INV_X1 U17955 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15955) );
  NAND2_X1 U17956 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n15954) );
  OAI211_X1 U17957 ( .C1(n16121), .C2(n15955), .A(n15954), .B(n16102), .ZN(
        n15956) );
  INV_X1 U17958 ( .A(n15956), .ZN(n15957) );
  NAND4_X1 U17959 ( .A1(n15960), .A2(n15959), .A3(n15958), .A4(n15957), .ZN(
        n15961) );
  NAND2_X1 U17960 ( .A1(n15962), .A2(n15961), .ZN(n16072) );
  NOR2_X1 U17961 ( .A1(n16073), .A2(n16072), .ZN(n16076) );
  AOI22_X1 U17962 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U17963 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15967) );
  INV_X1 U17964 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15964) );
  NAND2_X1 U17965 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n15963) );
  OAI211_X1 U17966 ( .C1(n16121), .C2(n15964), .A(n15963), .B(n16133), .ZN(
        n15965) );
  INV_X1 U17967 ( .A(n15965), .ZN(n15966) );
  NAND4_X1 U17968 ( .A1(n15969), .A2(n15968), .A3(n15967), .A4(n15966), .ZN(
        n15979) );
  AOI22_X1 U17969 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15977) );
  AOI22_X1 U17970 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15975) );
  INV_X1 U17971 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15972) );
  NAND2_X1 U17972 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n15971) );
  OAI211_X1 U17973 ( .C1(n16121), .C2(n15972), .A(n15971), .B(n16102), .ZN(
        n15973) );
  INV_X1 U17974 ( .A(n15973), .ZN(n15974) );
  NAND4_X1 U17975 ( .A1(n15977), .A2(n15976), .A3(n15975), .A4(n15974), .ZN(
        n15978) );
  AND2_X1 U17976 ( .A1(n15979), .A2(n15978), .ZN(n16077) );
  NAND2_X1 U17977 ( .A1(n16076), .A2(n16077), .ZN(n16084) );
  AOI22_X1 U17978 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15990) );
  INV_X1 U17979 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15982) );
  INV_X1 U17980 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15980) );
  OR2_X1 U17981 ( .A1(n16121), .A2(n15980), .ZN(n15981) );
  OAI211_X1 U17982 ( .C1(n15925), .C2(n15982), .A(n16102), .B(n15981), .ZN(
        n15983) );
  INV_X1 U17983 ( .A(n15983), .ZN(n15989) );
  INV_X1 U17984 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15985) );
  INV_X1 U17985 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15984) );
  OAI22_X1 U17986 ( .A1(n15985), .A2(n16131), .B1(n16124), .B2(n15984), .ZN(
        n15986) );
  INV_X1 U17987 ( .A(n15986), .ZN(n15987) );
  NAND4_X1 U17988 ( .A1(n15990), .A2(n15989), .A3(n15988), .A4(n15987), .ZN(
        n15999) );
  AOI22_X1 U17989 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15997) );
  AOI22_X1 U17990 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U17991 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n15991) );
  OAI211_X1 U17992 ( .C1(n16121), .C2(n15992), .A(n15991), .B(n16133), .ZN(
        n15993) );
  INV_X1 U17993 ( .A(n15993), .ZN(n15994) );
  NAND4_X1 U17994 ( .A1(n15997), .A2(n15996), .A3(n15995), .A4(n15994), .ZN(
        n15998) );
  AND2_X1 U17995 ( .A1(n15999), .A2(n15998), .ZN(n16083) );
  INV_X1 U17996 ( .A(n16083), .ZN(n16087) );
  OR2_X1 U17997 ( .A1(n16084), .A2(n16087), .ZN(n16093) );
  AOI22_X1 U17998 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16006) );
  AOI22_X1 U17999 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16004) );
  NAND2_X1 U18000 ( .A1(n12727), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n16000) );
  OAI211_X1 U18001 ( .C1(n16121), .C2(n16001), .A(n16000), .B(n16133), .ZN(
        n16002) );
  INV_X1 U18002 ( .A(n16002), .ZN(n16003) );
  NAND4_X1 U18003 ( .A1(n16006), .A2(n16005), .A3(n16004), .A4(n16003), .ZN(
        n16016) );
  AOI22_X1 U18004 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16014) );
  AOI22_X1 U18005 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16012) );
  INV_X1 U18006 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16009) );
  NAND2_X1 U18007 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n16008) );
  OAI211_X1 U18008 ( .C1(n16121), .C2(n16009), .A(n16008), .B(n16102), .ZN(
        n16010) );
  INV_X1 U18009 ( .A(n16010), .ZN(n16011) );
  NAND4_X1 U18010 ( .A1(n16014), .A2(n16013), .A3(n16012), .A4(n16011), .ZN(
        n16015) );
  NAND2_X1 U18011 ( .A1(n16016), .A2(n16015), .ZN(n16095) );
  OR2_X1 U18012 ( .A1(n16093), .A2(n16095), .ZN(n16896) );
  AOI22_X1 U18013 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16023) );
  AOI22_X1 U18014 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16021) );
  NAND2_X1 U18015 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n16017) );
  OAI211_X1 U18016 ( .C1(n16121), .C2(n16018), .A(n16017), .B(n16133), .ZN(
        n16019) );
  INV_X1 U18017 ( .A(n16019), .ZN(n16020) );
  NAND4_X1 U18018 ( .A1(n16023), .A2(n16022), .A3(n16021), .A4(n16020), .ZN(
        n16032) );
  AOI22_X1 U18019 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16030) );
  AOI22_X1 U18020 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16028) );
  INV_X1 U18021 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16025) );
  NAND2_X1 U18022 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n16024) );
  OAI211_X1 U18023 ( .C1(n16121), .C2(n16025), .A(n16024), .B(n16102), .ZN(
        n16026) );
  INV_X1 U18024 ( .A(n16026), .ZN(n16027) );
  NAND4_X1 U18025 ( .A1(n16030), .A2(n16029), .A3(n16028), .A4(n16027), .ZN(
        n16031) );
  AND2_X1 U18026 ( .A1(n16032), .A2(n16031), .ZN(n16897) );
  INV_X1 U18027 ( .A(n16897), .ZN(n16033) );
  NOR3_X1 U18028 ( .A1(n16896), .A2(n16097), .A3(n16033), .ZN(n16244) );
  AOI22_X1 U18029 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13303), .B1(
        n13304), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U18030 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U18031 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16035) );
  AOI22_X1 U18032 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16034) );
  NAND4_X1 U18033 ( .A1(n16037), .A2(n16036), .A3(n16035), .A4(n16034), .ZN(
        n16043) );
  AOI22_X1 U18034 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16041) );
  AOI22_X1 U18035 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16040) );
  AOI22_X1 U18036 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16039) );
  AOI22_X1 U18037 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16038) );
  NAND4_X1 U18038 ( .A1(n16041), .A2(n16040), .A3(n16039), .A4(n16038), .ZN(
        n16042) );
  NOR2_X1 U18039 ( .A1(n16043), .A2(n16042), .ZN(n16963) );
  AOI22_X1 U18040 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n13303), .B1(
        n13304), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16048) );
  AOI22_X1 U18041 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16047) );
  AOI22_X1 U18042 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16046) );
  AOI22_X1 U18043 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16045) );
  NAND4_X1 U18044 ( .A1(n16048), .A2(n16047), .A3(n16046), .A4(n16045), .ZN(
        n16054) );
  AOI22_X1 U18045 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16052) );
  AOI22_X1 U18046 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16051) );
  AOI22_X1 U18047 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16050) );
  AOI22_X1 U18048 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16049) );
  NAND4_X1 U18049 ( .A1(n16052), .A2(n16051), .A3(n16050), .A4(n16049), .ZN(
        n16053) );
  OR2_X1 U18050 ( .A1(n16054), .A2(n16053), .ZN(n16957) );
  AOI22_X1 U18051 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n13303), .B1(
        n13304), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16058) );
  AOI22_X1 U18052 ( .A1(n12951), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12772), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16057) );
  AOI22_X1 U18053 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12773), .B1(
        n12774), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16056) );
  AOI22_X1 U18054 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16055) );
  NAND4_X1 U18055 ( .A1(n16058), .A2(n16057), .A3(n16056), .A4(n16055), .ZN(
        n16068) );
  AOI22_X1 U18056 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12944), .B1(
        n12779), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16066) );
  AOI22_X1 U18057 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14285), .B1(
        n16059), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16065) );
  AOI22_X1 U18058 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n16061), .B1(
        n16060), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16064) );
  AOI22_X1 U18059 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n16062), .B1(
        n12932), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16063) );
  NAND4_X1 U18060 ( .A1(n16066), .A2(n16065), .A3(n16064), .A4(n16063), .ZN(
        n16067) );
  OR2_X1 U18061 ( .A1(n16068), .A2(n16067), .ZN(n16947) );
  XNOR2_X1 U18062 ( .A(n16070), .B(n16069), .ZN(n16940) );
  NAND2_X1 U18063 ( .A1(n16076), .A2(n19060), .ZN(n16075) );
  OAI21_X1 U18064 ( .B1(n16092), .B2(n16073), .A(n16072), .ZN(n16074) );
  AND2_X1 U18065 ( .A1(n16075), .A2(n16074), .ZN(n16930) );
  INV_X1 U18066 ( .A(n16076), .ZN(n16078) );
  INV_X1 U18067 ( .A(n16077), .ZN(n16080) );
  NAND2_X1 U18068 ( .A1(n16078), .A2(n16080), .ZN(n16079) );
  AND3_X1 U18069 ( .A1(n16084), .A2(n16085), .A3(n16079), .ZN(n16081) );
  NOR2_X1 U18070 ( .A1(n19060), .A2(n16080), .ZN(n16923) );
  INV_X1 U18071 ( .A(n16081), .ZN(n16082) );
  XNOR2_X1 U18072 ( .A(n16084), .B(n16083), .ZN(n16086) );
  NAND2_X1 U18073 ( .A1(n16086), .A2(n16085), .ZN(n16088) );
  XNOR2_X2 U18074 ( .A(n16090), .B(n16088), .ZN(n16914) );
  NOR2_X1 U18075 ( .A1(n19060), .A2(n16087), .ZN(n16913) );
  NAND2_X2 U18076 ( .A1(n16914), .A2(n16913), .ZN(n16912) );
  INV_X1 U18077 ( .A(n16088), .ZN(n16089) );
  NAND2_X1 U18078 ( .A1(n16090), .A2(n16089), .ZN(n16091) );
  AOI21_X1 U18079 ( .B1(n16093), .B2(n16095), .A(n16092), .ZN(n16094) );
  AND2_X1 U18080 ( .A1(n16896), .A2(n16094), .ZN(n16098) );
  INV_X1 U18081 ( .A(n16095), .ZN(n16096) );
  NAND2_X1 U18082 ( .A1(n16097), .A2(n16096), .ZN(n16905) );
  AOI22_X1 U18083 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16108) );
  INV_X1 U18084 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16103) );
  INV_X1 U18085 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16100) );
  OR2_X1 U18086 ( .A1(n16121), .A2(n16100), .ZN(n16101) );
  OAI211_X1 U18087 ( .C1(n15925), .C2(n16103), .A(n16102), .B(n16101), .ZN(
        n16104) );
  INV_X1 U18088 ( .A(n16104), .ZN(n16107) );
  AOI22_X1 U18089 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n15970), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16105) );
  NAND4_X1 U18090 ( .A1(n16108), .A2(n16107), .A3(n16106), .A4(n16105), .ZN(
        n16117) );
  AOI22_X1 U18091 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16115) );
  AOI22_X1 U18092 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16113) );
  INV_X1 U18093 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16110) );
  NAND2_X1 U18094 ( .A1(n12755), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16109) );
  OAI211_X1 U18095 ( .C1(n16121), .C2(n16110), .A(n16109), .B(n16133), .ZN(
        n16111) );
  INV_X1 U18096 ( .A(n16111), .ZN(n16112) );
  NAND4_X1 U18097 ( .A1(n16115), .A2(n16114), .A3(n16113), .A4(n16112), .ZN(
        n16116) );
  NAND2_X1 U18098 ( .A1(n16117), .A2(n16116), .ZN(n16118) );
  NAND2_X1 U18099 ( .A1(n16119), .A2(n16118), .ZN(n16241) );
  NOR2_X2 U18100 ( .A1(n16119), .A2(n16118), .ZN(n16242) );
  AOI21_X1 U18101 ( .B1(n16244), .B2(n16241), .A(n16242), .ZN(n16143) );
  OAI21_X1 U18102 ( .B1(n16121), .B2(n16120), .A(n16133), .ZN(n16126) );
  INV_X1 U18103 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16123) );
  INV_X1 U18104 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16122) );
  OAI22_X1 U18105 ( .A1(n16124), .A2(n16123), .B1(n16131), .B2(n16122), .ZN(
        n16125) );
  AOI211_X1 U18106 ( .C1(n12754), .C2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n16126), .B(n16125), .ZN(n16129) );
  AOI22_X1 U18107 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16128) );
  NAND3_X1 U18108 ( .A1(n16129), .A2(n16128), .A3(n16127), .ZN(n16141) );
  INV_X1 U18109 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16130) );
  NOR2_X1 U18110 ( .A1(n16131), .A2(n16130), .ZN(n16132) );
  AOI211_X1 U18111 ( .C1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n16134), .A(
        n16133), .B(n16132), .ZN(n16139) );
  AOI22_X1 U18112 ( .A1(n16099), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16135), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16138) );
  AOI22_X1 U18113 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15953), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16136) );
  NAND4_X1 U18114 ( .A1(n16139), .A2(n16138), .A3(n16137), .A4(n16136), .ZN(
        n16140) );
  NAND2_X1 U18115 ( .A1(n16141), .A2(n16140), .ZN(n16142) );
  XNOR2_X1 U18116 ( .A(n16143), .B(n16142), .ZN(n16151) );
  NAND2_X1 U18117 ( .A1(n19029), .A2(n16952), .ZN(n16145) );
  NAND2_X1 U18118 ( .A1(n16966), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16144) );
  OAI211_X1 U18119 ( .C1(n16151), .C2(n16968), .A(n16145), .B(n16144), .ZN(
        P2_U2857) );
  OAI22_X1 U18120 ( .A1(n20164), .A2(n19034), .B1(n16146), .B2(n20162), .ZN(
        n16147) );
  AOI21_X1 U18121 ( .B1(n19955), .B2(n16148), .A(n16147), .ZN(n16150) );
  AOI22_X1 U18122 ( .A1(n19956), .A2(BUF2_REG_30__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n16149) );
  OAI211_X1 U18123 ( .C1(n16151), .C2(n20115), .A(n16150), .B(n16149), .ZN(
        P2_U2889) );
  AND2_X2 U18124 ( .A1(n16153), .A2(n16152), .ZN(n16563) );
  INV_X1 U18125 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16697) );
  NAND2_X1 U18126 ( .A1(n20516), .A2(n16697), .ZN(n16154) );
  NAND2_X1 U18127 ( .A1(n16563), .A2(n16154), .ZN(n16164) );
  INV_X1 U18128 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16836) );
  XNOR2_X1 U18129 ( .A(n20516), .B(n16836), .ZN(n16160) );
  INV_X1 U18130 ( .A(n16160), .ZN(n16155) );
  NAND2_X1 U18131 ( .A1(n16778), .A2(n16688), .ZN(n16157) );
  NAND2_X1 U18132 ( .A1(n16155), .A2(n16157), .ZN(n16163) );
  NOR2_X1 U18133 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16156) );
  OR2_X1 U18134 ( .A1(n16778), .A2(n16156), .ZN(n16159) );
  NAND2_X1 U18135 ( .A1(n16159), .A2(n16157), .ZN(n16158) );
  NAND2_X1 U18136 ( .A1(n16158), .A2(n16836), .ZN(n16162) );
  NAND3_X1 U18137 ( .A1(n16164), .A2(n16160), .A3(n16159), .ZN(n16161) );
  OAI211_X1 U18138 ( .C1(n16164), .C2(n16163), .A(n16162), .B(n16161), .ZN(
        n16561) );
  AOI22_X1 U18139 ( .A1(n16210), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16209), .ZN(n16262) );
  NAND2_X1 U18140 ( .A1(n14072), .A2(n16615), .ZN(n16166) );
  NAND2_X1 U18141 ( .A1(n16206), .A2(n16448), .ZN(n16165) );
  NAND3_X1 U18142 ( .A1(n16166), .A2(n16261), .A3(n16165), .ZN(n16167) );
  NAND2_X1 U18143 ( .A1(n16168), .A2(n16167), .ZN(n16383) );
  MUX2_X1 U18144 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n16169) );
  OAI21_X1 U18145 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16210), .A(
        n16169), .ZN(n16461) );
  INV_X1 U18146 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16452) );
  NAND2_X1 U18147 ( .A1(n14072), .A2(n16170), .ZN(n16172) );
  NAND2_X1 U18148 ( .A1(n16206), .A2(n16452), .ZN(n16171) );
  NAND3_X1 U18149 ( .A1(n16172), .A2(n16261), .A3(n16171), .ZN(n16173) );
  NAND2_X1 U18150 ( .A1(n16174), .A2(n16173), .ZN(n16407) );
  MUX2_X1 U18151 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n16175) );
  NAND2_X1 U18152 ( .A1(n11280), .A2(n16175), .ZN(n16393) );
  OR2_X1 U18153 ( .A1(n16199), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n16178) );
  NAND2_X1 U18154 ( .A1(n16206), .A2(n22098), .ZN(n16176) );
  OAI211_X1 U18155 ( .C1(n15657), .C2(n21995), .A(n16176), .B(n14072), .ZN(
        n16177) );
  NAND2_X1 U18156 ( .A1(n16178), .A2(n16177), .ZN(n16446) );
  INV_X1 U18157 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16179) );
  OAI21_X1 U18158 ( .B1(n15657), .B2(n16179), .A(n14072), .ZN(n16181) );
  NAND2_X1 U18159 ( .A1(n16206), .A2(n16441), .ZN(n16180) );
  NAND2_X1 U18160 ( .A1(n16181), .A2(n16180), .ZN(n16182) );
  OAI21_X1 U18161 ( .B1(n16205), .B2(P1_EBX_REG_20__SCAN_IN), .A(n16182), .ZN(
        n16377) );
  MUX2_X1 U18162 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n16184) );
  OR2_X1 U18163 ( .A1(n16210), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16183) );
  AND2_X1 U18164 ( .A1(n16184), .A2(n16183), .ZN(n16433) );
  INV_X1 U18165 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16605) );
  NAND2_X1 U18166 ( .A1(n14072), .A2(n16605), .ZN(n16186) );
  NAND2_X1 U18167 ( .A1(n16206), .A2(n16432), .ZN(n16185) );
  NAND3_X1 U18168 ( .A1(n16186), .A2(n16261), .A3(n16185), .ZN(n16187) );
  AND2_X1 U18169 ( .A1(n16188), .A2(n16187), .ZN(n16365) );
  MUX2_X1 U18170 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n16190) );
  INV_X1 U18171 ( .A(n16210), .ZN(n16207) );
  NAND2_X1 U18172 ( .A1(n16207), .A2(n20515), .ZN(n16189) );
  NAND2_X1 U18173 ( .A1(n16190), .A2(n16189), .ZN(n16427) );
  OAI21_X1 U18174 ( .B1(n15657), .B2(n16583), .A(n14072), .ZN(n16192) );
  NAND2_X1 U18175 ( .A1(n16206), .A2(n16426), .ZN(n16191) );
  NAND2_X1 U18176 ( .A1(n16192), .A2(n16191), .ZN(n16193) );
  OAI21_X1 U18177 ( .B1(n16205), .B2(P1_EBX_REG_24__SCAN_IN), .A(n16193), .ZN(
        n16350) );
  MUX2_X1 U18178 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n16194) );
  OAI21_X1 U18179 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16210), .A(
        n16194), .ZN(n16339) );
  INV_X1 U18180 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16725) );
  NAND2_X1 U18181 ( .A1(n14072), .A2(n16725), .ZN(n16196) );
  NAND2_X1 U18182 ( .A1(n16206), .A2(n16422), .ZN(n16195) );
  NAND3_X1 U18183 ( .A1(n16196), .A2(n16261), .A3(n16195), .ZN(n16197) );
  AND2_X1 U18184 ( .A1(n16198), .A2(n16197), .ZN(n16328) );
  MUX2_X1 U18185 ( .A(n16199), .B(n16261), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n16200) );
  OAI21_X1 U18186 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16210), .A(
        n16200), .ZN(n16316) );
  NAND2_X1 U18187 ( .A1(n14072), .A2(n16201), .ZN(n16203) );
  INV_X1 U18188 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16420) );
  NAND2_X1 U18189 ( .A1(n16206), .A2(n16420), .ZN(n16202) );
  NAND3_X1 U18190 ( .A1(n16203), .A2(n16261), .A3(n16202), .ZN(n16204) );
  OAI21_X1 U18191 ( .B1(n16205), .B2(P1_EBX_REG_28__SCAN_IN), .A(n16204), .ZN(
        n16303) );
  AND2_X1 U18192 ( .A1(n16206), .A2(n16419), .ZN(n16208) );
  AOI21_X1 U18193 ( .B1(n16207), .B2(n16697), .A(n16208), .ZN(n16259) );
  MUX2_X1 U18194 ( .A(n16208), .B(n16259), .S(n16261), .Z(n16293) );
  MUX2_X1 U18195 ( .A(n16261), .B(n16262), .S(n16295), .Z(n16212) );
  OAI22_X1 U18196 ( .A1(n16210), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n16209), .ZN(n16211) );
  INV_X1 U18197 ( .A(n16418), .ZN(n16225) );
  NOR2_X1 U18198 ( .A1(n22001), .A2(n20435), .ZN(n16555) );
  NAND2_X1 U18199 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21974) );
  NOR3_X1 U18200 ( .A1(n16615), .A2(n21975), .A3(n21974), .ZN(n16217) );
  NAND2_X1 U18201 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21965) );
  NAND2_X1 U18202 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21956) );
  NOR2_X1 U18203 ( .A1(n21922), .A2(n21956), .ZN(n16216) );
  AOI21_X1 U18204 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21895) );
  NOR2_X1 U18205 ( .A1(n21896), .A2(n21909), .ZN(n21915) );
  NAND2_X1 U18206 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21915), .ZN(
        n21918) );
  NOR2_X1 U18207 ( .A1(n21895), .A2(n21918), .ZN(n21931) );
  NAND2_X1 U18208 ( .A1(n16216), .A2(n21931), .ZN(n21951) );
  NOR2_X1 U18209 ( .A1(n21965), .A2(n21951), .ZN(n16760) );
  NAND2_X1 U18210 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16760), .ZN(
        n16807) );
  NOR2_X1 U18211 ( .A1(n16803), .A2(n16807), .ZN(n21856) );
  NAND2_X1 U18212 ( .A1(n16217), .A2(n21856), .ZN(n16770) );
  NAND2_X1 U18213 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16213) );
  NOR2_X1 U18214 ( .A1(n16770), .A2(n16213), .ZN(n16764) );
  AND2_X1 U18215 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16214) );
  AND2_X1 U18216 ( .A1(n16764), .A2(n16214), .ZN(n16228) );
  NAND2_X1 U18217 ( .A1(n21952), .A2(n16228), .ZN(n16221) );
  NOR3_X1 U18218 ( .A1(n21893), .A2(n21879), .A3(n21918), .ZN(n21933) );
  NAND2_X1 U18219 ( .A1(n21933), .A2(n16216), .ZN(n16805) );
  NOR2_X1 U18220 ( .A1(n16805), .A2(n21965), .ZN(n16761) );
  NAND3_X1 U18221 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16761), .ZN(n21854) );
  INV_X1 U18222 ( .A(n21854), .ZN(n21861) );
  AND2_X1 U18223 ( .A1(n21861), .A2(n16217), .ZN(n16752) );
  NOR2_X1 U18224 ( .A1(n16605), .A2(n16218), .ZN(n16219) );
  AND2_X1 U18225 ( .A1(n16752), .A2(n16219), .ZN(n16226) );
  NAND2_X1 U18226 ( .A1(n21877), .A2(n16226), .ZN(n16220) );
  INV_X1 U18227 ( .A(n16726), .ZN(n16222) );
  NAND2_X1 U18228 ( .A1(n16222), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16223) );
  NOR2_X1 U18229 ( .A1(n22022), .A2(n16223), .ZN(n16722) );
  NAND3_X1 U18230 ( .A1(n16722), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16705), .ZN(n16686) );
  NOR3_X1 U18231 ( .A1(n16686), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16688), .ZN(n16224) );
  OR2_X1 U18232 ( .A1(n21932), .A2(n16226), .ZN(n16227) );
  OAI211_X1 U18233 ( .C1(n21884), .C2(n16228), .A(n21880), .B(n16227), .ZN(
        n22015) );
  INV_X1 U18234 ( .A(n16785), .ZN(n21936) );
  OR2_X1 U18235 ( .A1(n22015), .A2(n21936), .ZN(n16716) );
  OR2_X1 U18236 ( .A1(n22015), .A2(n16726), .ZN(n16229) );
  NAND2_X1 U18237 ( .A1(n16716), .A2(n16229), .ZN(n16734) );
  AND2_X1 U18238 ( .A1(n16734), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16718) );
  NAND2_X1 U18239 ( .A1(n16718), .A2(n16705), .ZN(n16687) );
  NAND2_X1 U18240 ( .A1(n21936), .A2(n16697), .ZN(n16689) );
  NAND2_X1 U18241 ( .A1(n16689), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16230) );
  OAI211_X1 U18242 ( .C1(n16687), .C2(n16230), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16716), .ZN(n16231) );
  OAI211_X1 U18243 ( .C1(n16561), .C2(n22004), .A(n16232), .B(n16231), .ZN(
        P1_U3000) );
  AOI21_X1 U18244 ( .B1(n17670), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16233), .ZN(n16235) );
  NAND2_X1 U18245 ( .A1(n16894), .A2(n17673), .ZN(n16234) );
  OAI211_X1 U18246 ( .C1(n16236), .C2(n17681), .A(n16235), .B(n16234), .ZN(
        n16237) );
  AOI21_X1 U18247 ( .B1(n16238), .B2(n17671), .A(n16237), .ZN(n16239) );
  INV_X1 U18248 ( .A(n16241), .ZN(n16243) );
  NOR2_X2 U18249 ( .A1(n16243), .A2(n16242), .ZN(n16245) );
  XNOR2_X1 U18250 ( .A(n16245), .B(n16244), .ZN(n16255) );
  OAI22_X1 U18251 ( .A1(n20164), .A2(n16247), .B1(n16246), .B2(n20162), .ZN(
        n16248) );
  AOI21_X1 U18252 ( .B1(n19955), .B2(n16249), .A(n16248), .ZN(n16251) );
  AOI22_X1 U18253 ( .A1(n19956), .A2(BUF2_REG_29__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16250) );
  OAI211_X1 U18254 ( .C1(n16255), .C2(n20115), .A(n16251), .B(n16250), .ZN(
        P2_U2890) );
  NAND2_X1 U18255 ( .A1(n16966), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16254) );
  NAND2_X1 U18256 ( .A1(n16252), .A2(n16952), .ZN(n16253) );
  OAI211_X1 U18257 ( .C1(n16255), .C2(n16968), .A(n16254), .B(n16253), .ZN(
        P2_U2858) );
  NAND2_X1 U18258 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n16413), .ZN(n16412) );
  NAND2_X1 U18259 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n16362), .ZN(n22126) );
  INV_X1 U18260 ( .A(n22126), .ZN(n16256) );
  INV_X1 U18261 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20430) );
  INV_X1 U18262 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20431) );
  XNOR2_X1 U18263 ( .A(n16298), .B(P1_REIP_REG_30__SCAN_IN), .ZN(n16267) );
  INV_X1 U18264 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16277) );
  AOI22_X1 U18265 ( .A1(n16257), .A2(n22110), .B1(n22134), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16258) );
  OAI21_X1 U18266 ( .B1(n22131), .B2(n16277), .A(n16258), .ZN(n16266) );
  NAND2_X1 U18267 ( .A1(n16305), .A2(n16259), .ZN(n16260) );
  OAI21_X1 U18268 ( .B1(n16295), .B2(n16261), .A(n16260), .ZN(n16264) );
  INV_X1 U18269 ( .A(n16262), .ZN(n16263) );
  NOR2_X1 U18270 ( .A1(n16684), .A2(n22059), .ZN(n16265) );
  AOI211_X1 U18271 ( .C1(n16267), .C2(n22096), .A(n16266), .B(n16265), .ZN(
        n16268) );
  OAI21_X1 U18272 ( .B1(n16278), .B2(n22114), .A(n16268), .ZN(P1_U2810) );
  NOR2_X1 U18273 ( .A1(n16272), .A2(n16270), .ZN(n16269) );
  NAND2_X1 U18274 ( .A1(n16523), .A2(n16269), .ZN(n16526) );
  INV_X1 U18275 ( .A(n16526), .ZN(n16542) );
  AOI22_X1 U18276 ( .A1(n16542), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16549), .ZN(n16276) );
  INV_X1 U18277 ( .A(n16270), .ZN(n16271) );
  NOR3_X1 U18278 ( .A1(n16549), .A2(n16272), .A3(n16271), .ZN(n16273) );
  AOI22_X1 U18279 ( .A1(n11159), .A2(n16274), .B1(n16543), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n16275) );
  OAI211_X1 U18280 ( .C1(n16278), .C2(n16553), .A(n16276), .B(n16275), .ZN(
        P1_U2874) );
  OAI222_X1 U18281 ( .A1(n16425), .A2(n16278), .B1(n16451), .B2(n16277), .C1(
        n16684), .C2(n16453), .ZN(P1_U2842) );
  NAND2_X1 U18282 ( .A1(n16289), .A2(n16279), .ZN(n16284) );
  AOI22_X1 U18283 ( .A1(n16281), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n16280), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16282) );
  INV_X1 U18284 ( .A(n16282), .ZN(n16283) );
  XNOR2_X2 U18285 ( .A(n16284), .B(n16283), .ZN(n16559) );
  NAND2_X1 U18286 ( .A1(n16559), .A2(n22137), .ZN(n16288) );
  INV_X1 U18287 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20437) );
  OAI22_X1 U18288 ( .A1(n22113), .A2(n16285), .B1(P1_REIP_REG_31__SCAN_IN), 
        .B2(n11379), .ZN(n16286) );
  OAI211_X1 U18289 ( .C1(n16418), .C2(n22059), .A(n16288), .B(n16287), .ZN(
        P1_U2809) );
  AOI21_X1 U18290 ( .B1(n16291), .B2(n16290), .A(n16289), .ZN(n16567) );
  INV_X1 U18291 ( .A(n16567), .ZN(n16471) );
  OAI22_X1 U18292 ( .A1(n16292), .A2(n22113), .B1(n22128), .B2(n16565), .ZN(
        n16297) );
  NOR2_X1 U18293 ( .A1(n16305), .A2(n16293), .ZN(n16294) );
  NOR2_X1 U18294 ( .A1(n16700), .A2(n22059), .ZN(n16296) );
  AOI211_X1 U18295 ( .C1(n22118), .C2(P1_EBX_REG_29__SCAN_IN), .A(n16297), .B(
        n16296), .ZN(n16301) );
  INV_X1 U18296 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20433) );
  NOR2_X1 U18297 ( .A1(n22125), .A2(n20433), .ZN(n16299) );
  OAI21_X1 U18298 ( .B1(n16299), .B2(n16302), .A(n16298), .ZN(n16300) );
  OAI211_X1 U18299 ( .C1(n16471), .C2(n22114), .A(n16301), .B(n16300), .ZN(
        P1_U2811) );
  INV_X1 U18300 ( .A(n16302), .ZN(n16311) );
  OAI21_X1 U18301 ( .B1(n22125), .B2(n20431), .A(n16323), .ZN(n16310) );
  NOR2_X1 U18302 ( .A1(n16315), .A2(n16303), .ZN(n16304) );
  OR2_X1 U18303 ( .A1(n16305), .A2(n16304), .ZN(n16708) );
  AOI22_X1 U18304 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n22134), .B1(
        n22110), .B2(n16306), .ZN(n16308) );
  NAND2_X1 U18305 ( .A1(n22118), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n16307) );
  OAI211_X1 U18306 ( .C1(n16708), .C2(n22059), .A(n16308), .B(n16307), .ZN(
        n16309) );
  AOI21_X1 U18307 ( .B1(n16311), .B2(n16310), .A(n16309), .ZN(n16312) );
  OAI21_X1 U18308 ( .B1(n16478), .B2(n22114), .A(n16312), .ZN(P1_U2812) );
  AOI21_X1 U18309 ( .B1(n16314), .B2(n16326), .A(n12446), .ZN(n16574) );
  INV_X1 U18310 ( .A(n16574), .ZN(n16485) );
  OAI21_X1 U18311 ( .B1(n22125), .B2(n20430), .A(n16333), .ZN(n16322) );
  AOI21_X1 U18312 ( .B1(n16316), .B2(n11256), .A(n16315), .ZN(n16317) );
  INV_X1 U18313 ( .A(n16317), .ZN(n16715) );
  OAI22_X1 U18314 ( .A1(n16318), .A2(n22113), .B1(n22128), .B2(n16572), .ZN(
        n16319) );
  AOI21_X1 U18315 ( .B1(n22118), .B2(P1_EBX_REG_27__SCAN_IN), .A(n16319), .ZN(
        n16320) );
  OAI21_X1 U18316 ( .B1(n16715), .B2(n22059), .A(n16320), .ZN(n16321) );
  AOI21_X1 U18317 ( .B1(n16323), .B2(n16322), .A(n16321), .ZN(n16324) );
  OAI21_X1 U18318 ( .B1(n16485), .B2(n22114), .A(n16324), .ZN(P1_U2813) );
  OAI21_X1 U18319 ( .B1(n16325), .B2(n16327), .A(n16326), .ZN(n16578) );
  INV_X1 U18320 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20428) );
  OAI21_X1 U18321 ( .B1(n22125), .B2(n20428), .A(n11243), .ZN(n16334) );
  NAND2_X1 U18322 ( .A1(n16337), .A2(n16328), .ZN(n16329) );
  NAND2_X1 U18323 ( .A1(n11256), .A2(n16329), .ZN(n16728) );
  NAND2_X1 U18324 ( .A1(n22118), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n16331) );
  AOI22_X1 U18325 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n22134), .B1(
        n22110), .B2(n16581), .ZN(n16330) );
  OAI211_X1 U18326 ( .C1(n16728), .C2(n22059), .A(n16331), .B(n16330), .ZN(
        n16332) );
  AOI21_X1 U18327 ( .B1(n16334), .B2(n16333), .A(n16332), .ZN(n16335) );
  OAI21_X1 U18328 ( .B1(n16578), .B2(n22114), .A(n16335), .ZN(P1_U2814) );
  AOI21_X1 U18329 ( .B1(n16336), .B2(n11198), .A(n16325), .ZN(n16591) );
  INV_X1 U18330 ( .A(n16591), .ZN(n16498) );
  OAI21_X1 U18331 ( .B1(n22125), .B2(n20425), .A(n16354), .ZN(n16344) );
  INV_X1 U18332 ( .A(n16337), .ZN(n16338) );
  AOI21_X1 U18333 ( .B1(n16339), .B2(n16349), .A(n16338), .ZN(n16423) );
  INV_X1 U18334 ( .A(n16423), .ZN(n16737) );
  INV_X1 U18335 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16340) );
  OAI22_X1 U18336 ( .A1(n16340), .A2(n22113), .B1(n22128), .B2(n16589), .ZN(
        n16341) );
  AOI21_X1 U18337 ( .B1(n22118), .B2(P1_EBX_REG_25__SCAN_IN), .A(n16341), .ZN(
        n16342) );
  OAI21_X1 U18338 ( .B1(n22059), .B2(n16737), .A(n16342), .ZN(n16343) );
  AOI21_X1 U18339 ( .B1(n11243), .B2(n16344), .A(n16343), .ZN(n16345) );
  OAI21_X1 U18340 ( .B1(n16498), .B2(n22114), .A(n16345), .ZN(P1_U2815) );
  OAI21_X1 U18341 ( .B1(n16346), .B2(n16347), .A(n11198), .ZN(n16598) );
  INV_X1 U18342 ( .A(n22124), .ZN(n16348) );
  OAI21_X1 U18343 ( .B1(n22125), .B2(n11382), .A(n16348), .ZN(n16355) );
  OAI21_X1 U18344 ( .B1(n11241), .B2(n16350), .A(n16349), .ZN(n16748) );
  NAND2_X1 U18345 ( .A1(n22118), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n16352) );
  AOI22_X1 U18346 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n22134), .B1(
        n22110), .B2(n16601), .ZN(n16351) );
  OAI211_X1 U18347 ( .C1(n16748), .C2(n22059), .A(n16352), .B(n16351), .ZN(
        n16353) );
  AOI21_X1 U18348 ( .B1(n16355), .B2(n16354), .A(n16353), .ZN(n16356) );
  OAI21_X1 U18349 ( .B1(n16598), .B2(n22114), .A(n16356), .ZN(P1_U2816) );
  OAI21_X1 U18350 ( .B1(n16439), .B2(n16359), .A(n16358), .ZN(n16607) );
  INV_X1 U18351 ( .A(n16360), .ZN(n16609) );
  NOR3_X1 U18352 ( .A1(n16362), .A2(n22125), .A3(n20422), .ZN(n16361) );
  AOI21_X1 U18353 ( .B1(n20422), .B2(n16362), .A(n16361), .ZN(n16364) );
  NAND2_X1 U18354 ( .A1(n22134), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16363) );
  OAI211_X1 U18355 ( .C1(n22128), .C2(n16609), .A(n16364), .B(n16363), .ZN(
        n16368) );
  NAND2_X1 U18356 ( .A1(n16436), .A2(n16365), .ZN(n16366) );
  NAND2_X1 U18357 ( .A1(n16428), .A2(n16366), .ZN(n22013) );
  NOR2_X1 U18358 ( .A1(n22059), .A2(n22013), .ZN(n16367) );
  AOI211_X1 U18359 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n22118), .A(n16368), .B(
        n16367), .ZN(n16369) );
  OAI21_X1 U18360 ( .B1(n16607), .B2(n22114), .A(n16369), .ZN(P1_U2818) );
  OAI21_X1 U18361 ( .B1(n16370), .B2(n16372), .A(n16371), .ZN(n16625) );
  NAND2_X1 U18362 ( .A1(n22110), .A2(n16628), .ZN(n16375) );
  NAND2_X1 U18363 ( .A1(n22107), .A2(n22096), .ZN(n22122) );
  INV_X1 U18364 ( .A(n22122), .ZN(n16373) );
  OAI21_X1 U18365 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n22106), .A(n16373), 
        .ZN(n16374) );
  OAI211_X1 U18366 ( .C1(n22113), .C2(n16624), .A(n16375), .B(n16374), .ZN(
        n16379) );
  INV_X1 U18367 ( .A(n16434), .ZN(n16376) );
  OAI21_X1 U18368 ( .B1(n16444), .B2(n16377), .A(n16376), .ZN(n16774) );
  NOR2_X1 U18369 ( .A1(n22059), .A2(n16774), .ZN(n16378) );
  AOI211_X1 U18370 ( .C1(P1_EBX_REG_20__SCAN_IN), .C2(n22118), .A(n16379), .B(
        n16378), .ZN(n16380) );
  OAI21_X1 U18371 ( .B1(n16625), .B2(n22114), .A(n16380), .ZN(P1_U2820) );
  OR2_X1 U18372 ( .A1(n16383), .A2(n11250), .ZN(n16384) );
  NAND2_X1 U18373 ( .A1(n16384), .A2(n16445), .ZN(n21980) );
  NOR2_X1 U18374 ( .A1(n22113), .A2(n16630), .ZN(n16385) );
  AOI211_X1 U18375 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n22118), .A(n22100), .B(
        n16385), .ZN(n16386) );
  OAI21_X1 U18376 ( .B1(n22059), .B2(n21980), .A(n16386), .ZN(n16387) );
  AOI21_X1 U18377 ( .B1(n16632), .B2(n22110), .A(n16387), .ZN(n16390) );
  NOR2_X1 U18378 ( .A1(n22125), .A2(n20414), .ZN(n16388) );
  OAI21_X1 U18379 ( .B1(n16388), .B2(n16397), .A(n22094), .ZN(n16389) );
  OAI211_X1 U18380 ( .C1(n16637), .C2(n22114), .A(n16390), .B(n16389), .ZN(
        P1_U2822) );
  NAND2_X1 U18381 ( .A1(n15850), .A2(n16454), .ZN(n16455) );
  NAND2_X1 U18382 ( .A1(n16403), .A2(n16391), .ZN(n16392) );
  AND2_X1 U18383 ( .A1(n16382), .A2(n16392), .ZN(n20506) );
  INV_X1 U18384 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16449) );
  AOI21_X1 U18385 ( .B1(n16393), .B2(n16408), .A(n11250), .ZN(n16790) );
  INV_X1 U18386 ( .A(n16790), .ZN(n16450) );
  AOI21_X1 U18387 ( .B1(n22134), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n22100), .ZN(n16395) );
  NAND2_X1 U18388 ( .A1(n22110), .A2(n20504), .ZN(n16394) );
  OAI211_X1 U18389 ( .C1(n22059), .C2(n16450), .A(n16395), .B(n16394), .ZN(
        n16396) );
  INV_X1 U18390 ( .A(n16396), .ZN(n16400) );
  AOI21_X1 U18391 ( .B1(n20413), .B2(n16412), .A(n16397), .ZN(n16398) );
  NAND2_X1 U18392 ( .A1(n22096), .A2(n16398), .ZN(n16399) );
  OAI211_X1 U18393 ( .C1(n16449), .C2(n22131), .A(n16400), .B(n16399), .ZN(
        n16401) );
  AOI21_X1 U18394 ( .B1(n20506), .B2(n22137), .A(n16401), .ZN(n16402) );
  INV_X1 U18395 ( .A(n16402), .ZN(P1_U2823) );
  INV_X1 U18396 ( .A(n16403), .ZN(n16404) );
  AOI21_X1 U18397 ( .B1(n16405), .B2(n16455), .A(n16404), .ZN(n16648) );
  INV_X1 U18398 ( .A(n16648), .ZN(n16548) );
  AOI21_X1 U18399 ( .B1(n22134), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n22100), .ZN(n16406) );
  OAI21_X1 U18400 ( .B1(n16646), .B2(n22128), .A(n16406), .ZN(n16411) );
  OR2_X1 U18401 ( .A1(n16407), .A2(n16459), .ZN(n16409) );
  NAND2_X1 U18402 ( .A1(n16409), .A2(n16408), .ZN(n21993) );
  NOR2_X1 U18403 ( .A1(n22059), .A2(n21993), .ZN(n16410) );
  AOI211_X1 U18404 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n22118), .A(n16411), .B(
        n16410), .ZN(n16416) );
  NOR2_X1 U18405 ( .A1(n22125), .A2(n20410), .ZN(n16414) );
  OAI21_X1 U18406 ( .B1(n16414), .B2(n16413), .A(n16412), .ZN(n16415) );
  OAI211_X1 U18407 ( .C1(n16548), .C2(n22114), .A(n16416), .B(n16415), .ZN(
        P1_U2824) );
  INV_X1 U18408 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16417) );
  OAI22_X1 U18409 ( .A1(n16418), .A2(n16453), .B1(n16417), .B2(n16451), .ZN(
        P1_U2841) );
  OAI222_X1 U18410 ( .A1(n16419), .A2(n16451), .B1(n16453), .B2(n16700), .C1(
        n16471), .C2(n16425), .ZN(P1_U2843) );
  OAI222_X1 U18411 ( .A1(n16708), .A2(n16453), .B1(n16420), .B2(n16451), .C1(
        n16478), .C2(n16425), .ZN(P1_U2844) );
  INV_X1 U18412 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16421) );
  OAI222_X1 U18413 ( .A1(n16421), .A2(n16451), .B1(n16453), .B2(n16715), .C1(
        n16485), .C2(n16425), .ZN(P1_U2845) );
  OAI222_X1 U18414 ( .A1(n16728), .A2(n16453), .B1(n16422), .B2(n16451), .C1(
        n16578), .C2(n16425), .ZN(P1_U2846) );
  AOI22_X1 U18415 ( .A1(n16423), .A2(n16463), .B1(n16462), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n16424) );
  OAI21_X1 U18416 ( .B1(n16498), .B2(n16425), .A(n16424), .ZN(P1_U2847) );
  OAI222_X1 U18417 ( .A1(n16748), .A2(n16453), .B1(n16426), .B2(n16451), .C1(
        n16598), .C2(n16425), .ZN(P1_U2848) );
  AND2_X1 U18418 ( .A1(n16428), .A2(n16427), .ZN(n16429) );
  NOR2_X1 U18419 ( .A1(n11241), .A2(n16429), .ZN(n22135) );
  INV_X1 U18420 ( .A(n22135), .ZN(n16431) );
  INV_X1 U18421 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n22130) );
  AOI21_X1 U18422 ( .B1(n16430), .B2(n16358), .A(n16346), .ZN(n22138) );
  INV_X1 U18423 ( .A(n22138), .ZN(n16510) );
  OAI222_X1 U18424 ( .A1(n16431), .A2(n16453), .B1(n16451), .B2(n22130), .C1(
        n16425), .C2(n16510), .ZN(P1_U2849) );
  OAI222_X1 U18425 ( .A1(n22013), .A2(n16453), .B1(n16432), .B2(n16451), .C1(
        n16425), .C2(n16607), .ZN(P1_U2850) );
  OR2_X1 U18426 ( .A1(n16434), .A2(n16433), .ZN(n16435) );
  NAND2_X1 U18427 ( .A1(n16436), .A2(n16435), .ZN(n16758) );
  INV_X1 U18428 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n16440) );
  AND2_X1 U18429 ( .A1(n16371), .A2(n16437), .ZN(n16438) );
  OR2_X1 U18430 ( .A1(n16439), .A2(n16438), .ZN(n22115) );
  OAI222_X1 U18431 ( .A1(n16758), .A2(n16453), .B1(n16440), .B2(n16451), .C1(
        n22115), .C2(n16425), .ZN(P1_U2851) );
  OAI222_X1 U18432 ( .A1(n16774), .A2(n16453), .B1(n16441), .B2(n16451), .C1(
        n16625), .C2(n16425), .ZN(P1_U2852) );
  INV_X1 U18433 ( .A(n16442), .ZN(n16443) );
  AOI21_X1 U18434 ( .B1(n16443), .B2(n11190), .A(n16370), .ZN(n22102) );
  INV_X1 U18435 ( .A(n22102), .ZN(n16534) );
  AOI21_X1 U18436 ( .B1(n16446), .B2(n16445), .A(n16444), .ZN(n22101) );
  AOI22_X1 U18437 ( .A1(n16463), .A2(n22101), .B1(n16462), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n16447) );
  OAI21_X1 U18438 ( .B1(n16534), .B2(n16425), .A(n16447), .ZN(P1_U2853) );
  OAI222_X1 U18439 ( .A1(n21980), .A2(n16453), .B1(n16448), .B2(n16451), .C1(
        n16425), .C2(n16637), .ZN(P1_U2854) );
  INV_X1 U18440 ( .A(n20506), .ZN(n16541) );
  OAI222_X1 U18441 ( .A1(n16450), .A2(n16453), .B1(n16451), .B2(n16449), .C1(
        n16425), .C2(n16541), .ZN(P1_U2855) );
  OAI222_X1 U18442 ( .A1(n21993), .A2(n16453), .B1(n16452), .B2(n16451), .C1(
        n16425), .C2(n16548), .ZN(P1_U2856) );
  INV_X1 U18443 ( .A(n16454), .ZN(n16458) );
  INV_X1 U18444 ( .A(n16455), .ZN(n16456) );
  AOI21_X1 U18445 ( .B1(n16458), .B2(n16457), .A(n16456), .ZN(n22090) );
  INV_X1 U18446 ( .A(n22090), .ZN(n16554) );
  AOI21_X1 U18447 ( .B1(n16461), .B2(n16460), .A(n16459), .ZN(n22084) );
  AOI22_X1 U18448 ( .A1(n16463), .A2(n22084), .B1(n16462), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n16464) );
  OAI21_X1 U18449 ( .B1(n16554), .B2(n16425), .A(n16464), .ZN(P1_U2857) );
  NAND3_X1 U18450 ( .A1(n16559), .A2(n22476), .A3(n16523), .ZN(n16466) );
  AOI22_X1 U18451 ( .A1(n16543), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16549), .ZN(n16465) );
  OAI211_X1 U18452 ( .C1(n16526), .C2(n16467), .A(n16466), .B(n16465), .ZN(
        P1_U2873) );
  AOI22_X1 U18453 ( .A1(n16542), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16549), .ZN(n16470) );
  AOI22_X1 U18454 ( .A1(n11159), .A2(n16468), .B1(n16543), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16469) );
  OAI211_X1 U18455 ( .C1(n16471), .C2(n16553), .A(n16470), .B(n16469), .ZN(
        P1_U2875) );
  OAI22_X1 U18456 ( .A1(n16526), .A2(n16473), .B1(n16472), .B2(n16523), .ZN(
        n16474) );
  INV_X1 U18457 ( .A(n16474), .ZN(n16477) );
  AOI22_X1 U18458 ( .A1(n11159), .A2(n16475), .B1(n16543), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16476) );
  OAI211_X1 U18459 ( .C1(n16478), .C2(n16553), .A(n16477), .B(n16476), .ZN(
        P1_U2876) );
  INV_X1 U18460 ( .A(DATAI_27_), .ZN(n16480) );
  OAI22_X1 U18461 ( .A1(n16526), .A2(n16480), .B1(n16479), .B2(n16523), .ZN(
        n16481) );
  INV_X1 U18462 ( .A(n16481), .ZN(n16484) );
  AOI22_X1 U18463 ( .A1(n11159), .A2(n16482), .B1(n16543), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16483) );
  OAI211_X1 U18464 ( .C1(n16485), .C2(n16553), .A(n16484), .B(n16483), .ZN(
        P1_U2877) );
  INV_X1 U18465 ( .A(DATAI_26_), .ZN(n16487) );
  OAI22_X1 U18466 ( .A1(n16526), .A2(n16487), .B1(n16486), .B2(n16523), .ZN(
        n16488) );
  INV_X1 U18467 ( .A(n16488), .ZN(n16491) );
  AOI22_X1 U18468 ( .A1(n11159), .A2(n16489), .B1(n16543), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16490) );
  OAI211_X1 U18469 ( .C1(n16578), .C2(n16553), .A(n16491), .B(n16490), .ZN(
        P1_U2878) );
  INV_X1 U18470 ( .A(DATAI_25_), .ZN(n16493) );
  OAI22_X1 U18471 ( .A1(n16526), .A2(n16493), .B1(n16492), .B2(n16523), .ZN(
        n16494) );
  INV_X1 U18472 ( .A(n16494), .ZN(n16497) );
  AOI22_X1 U18473 ( .A1(n11159), .A2(n16495), .B1(n16543), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16496) );
  OAI211_X1 U18474 ( .C1(n16498), .C2(n16553), .A(n16497), .B(n16496), .ZN(
        P1_U2879) );
  INV_X1 U18475 ( .A(DATAI_24_), .ZN(n16500) );
  OAI22_X1 U18476 ( .A1(n16526), .A2(n16500), .B1(n16499), .B2(n16523), .ZN(
        n16503) );
  NOR2_X1 U18478 ( .A1(n22598), .A2(n16501), .ZN(n16502) );
  AOI211_X1 U18479 ( .C1(n16543), .C2(BUF1_REG_24__SCAN_IN), .A(n16503), .B(
        n16502), .ZN(n16504) );
  OAI21_X1 U18480 ( .B1(n16598), .B2(n16553), .A(n16504), .ZN(P1_U2880) );
  INV_X1 U18481 ( .A(DATAI_23_), .ZN(n16506) );
  OAI22_X1 U18482 ( .A1(n16526), .A2(n16506), .B1(n16505), .B2(n16523), .ZN(
        n16508) );
  NOR2_X1 U18483 ( .A1(n22598), .A2(n22480), .ZN(n16507) );
  AOI211_X1 U18484 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n16543), .A(n16508), .B(
        n16507), .ZN(n16509) );
  OAI21_X1 U18485 ( .B1(n16510), .B2(n16553), .A(n16509), .ZN(P1_U2881) );
  OAI22_X1 U18486 ( .A1(n16526), .A2(n16512), .B1(n16511), .B2(n16523), .ZN(
        n16515) );
  NOR2_X1 U18487 ( .A1(n22598), .A2(n16513), .ZN(n16514) );
  AOI211_X1 U18488 ( .C1(n16543), .C2(BUF1_REG_22__SCAN_IN), .A(n16515), .B(
        n16514), .ZN(n16516) );
  OAI21_X1 U18489 ( .B1(n16607), .B2(n16553), .A(n16516), .ZN(P1_U2882) );
  INV_X1 U18490 ( .A(DATAI_21_), .ZN(n16518) );
  OAI22_X1 U18491 ( .A1(n16526), .A2(n16518), .B1(n16517), .B2(n16523), .ZN(
        n16519) );
  INV_X1 U18492 ( .A(n16519), .ZN(n16522) );
  AOI22_X1 U18493 ( .A1(n11159), .A2(n16520), .B1(n16543), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n16521) );
  OAI211_X1 U18494 ( .C1(n22115), .C2(n16553), .A(n16522), .B(n16521), .ZN(
        P1_U2883) );
  OAI22_X1 U18495 ( .A1(n16526), .A2(n16525), .B1(n16524), .B2(n16523), .ZN(
        n16529) );
  NOR2_X1 U18496 ( .A1(n22598), .A2(n22383), .ZN(n16528) );
  AOI211_X1 U18497 ( .C1(n16543), .C2(BUF1_REG_20__SCAN_IN), .A(n16529), .B(
        n16528), .ZN(n16530) );
  OAI21_X1 U18498 ( .B1(n16625), .B2(n16553), .A(n16530), .ZN(P1_U2884) );
  AOI22_X1 U18499 ( .A1(n16542), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16549), .ZN(n16533) );
  AOI22_X1 U18500 ( .A1(n11159), .A2(n16531), .B1(n16543), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n16532) );
  OAI211_X1 U18501 ( .C1(n16534), .C2(n16553), .A(n16533), .B(n16532), .ZN(
        P1_U2885) );
  AOI22_X1 U18502 ( .A1(n16542), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16549), .ZN(n16537) );
  AOI22_X1 U18503 ( .A1(n11159), .A2(n16535), .B1(n16543), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16536) );
  OAI211_X1 U18504 ( .C1(n16637), .C2(n16553), .A(n16537), .B(n16536), .ZN(
        P1_U2886) );
  AOI22_X1 U18505 ( .A1(n16542), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16549), .ZN(n16540) );
  AOI22_X1 U18506 ( .A1(n11159), .A2(n16538), .B1(n16543), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n16539) );
  OAI211_X1 U18507 ( .C1(n16541), .C2(n16553), .A(n16540), .B(n16539), .ZN(
        P1_U2887) );
  AOI22_X1 U18508 ( .A1(n16542), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16549), .ZN(n16547) );
  AOI22_X1 U18509 ( .A1(n11159), .A2(n16544), .B1(n16543), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n16546) );
  OAI211_X1 U18510 ( .C1(n16548), .C2(n16553), .A(n16547), .B(n16546), .ZN(
        P1_U2888) );
  AOI22_X1 U18511 ( .A1(n16551), .A2(n16550), .B1(P1_EAX_REG_15__SCAN_IN), 
        .B2(n16549), .ZN(n16552) );
  OAI21_X1 U18512 ( .B1(n16554), .B2(n16553), .A(n16552), .ZN(P1_U2889) );
  AOI21_X1 U18513 ( .B1(n20514), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16555), .ZN(n16556) );
  OAI21_X1 U18514 ( .B1(n20522), .B2(n16557), .A(n16556), .ZN(n16558) );
  OAI21_X1 U18515 ( .B1(n22141), .B2(n16561), .A(n16560), .ZN(P1_U2968) );
  XNOR2_X1 U18516 ( .A(n16563), .B(n16562), .ZN(n16704) );
  NOR2_X1 U18517 ( .A1(n22001), .A2(n20433), .ZN(n16696) );
  AOI21_X1 U18518 ( .B1(n20514), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16696), .ZN(n16564) );
  OAI21_X1 U18519 ( .B1(n20522), .B2(n16565), .A(n16564), .ZN(n16566) );
  AOI21_X1 U18520 ( .B1(n16567), .B2(n20519), .A(n16566), .ZN(n16568) );
  OAI21_X1 U18521 ( .B1(n22141), .B2(n16704), .A(n16568), .ZN(P1_U2970) );
  XNOR2_X1 U18522 ( .A(n20516), .B(n16721), .ZN(n16569) );
  XNOR2_X1 U18523 ( .A(n16570), .B(n16569), .ZN(n16724) );
  NAND2_X1 U18524 ( .A1(n22016), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16714) );
  NAND2_X1 U18525 ( .A1(n20514), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16571) );
  OAI211_X1 U18526 ( .C1(n20522), .C2(n16572), .A(n16714), .B(n16571), .ZN(
        n16573) );
  AOI21_X1 U18527 ( .B1(n16574), .B2(n20519), .A(n16573), .ZN(n16575) );
  OAI21_X1 U18528 ( .B1(n16724), .B2(n22141), .A(n16575), .ZN(P1_U2972) );
  NAND2_X1 U18529 ( .A1(n22016), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16727) );
  OAI21_X1 U18530 ( .B1(n16670), .B2(n16577), .A(n16727), .ZN(n16580) );
  NOR2_X1 U18531 ( .A1(n16578), .A2(n20496), .ZN(n16579) );
  AOI211_X1 U18532 ( .C1(n20505), .C2(n16581), .A(n16580), .B(n16579), .ZN(
        n16582) );
  OAI21_X1 U18533 ( .B1(n22141), .B2(n16733), .A(n16582), .ZN(P1_U2973) );
  AOI21_X1 U18534 ( .B1(n16593), .B2(n16583), .A(n16735), .ZN(n16586) );
  MUX2_X1 U18535 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n16584), .S(
        n20516), .Z(n16585) );
  NOR2_X1 U18536 ( .A1(n16586), .A2(n16585), .ZN(n16587) );
  XNOR2_X1 U18537 ( .A(n16587), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16742) );
  NAND2_X1 U18538 ( .A1(n21906), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16736) );
  NAND2_X1 U18539 ( .A1(n20514), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16588) );
  OAI211_X1 U18540 ( .C1(n20522), .C2(n16589), .A(n16736), .B(n16588), .ZN(
        n16590) );
  AOI21_X1 U18541 ( .B1(n16591), .B2(n20519), .A(n16590), .ZN(n16592) );
  OAI21_X1 U18542 ( .B1(n22141), .B2(n16742), .A(n16592), .ZN(P1_U2974) );
  NAND3_X1 U18543 ( .A1(n16593), .A2(n16779), .A3(n20515), .ZN(n16595) );
  NAND3_X1 U18544 ( .A1(n13658), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16778), .ZN(n16594) );
  NAND2_X1 U18545 ( .A1(n16595), .A2(n16594), .ZN(n16596) );
  XNOR2_X1 U18546 ( .A(n16596), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16751) );
  NAND2_X1 U18547 ( .A1(n21906), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16746) );
  OAI21_X1 U18548 ( .B1(n16670), .B2(n16597), .A(n16746), .ZN(n16600) );
  NOR2_X1 U18549 ( .A1(n16598), .A2(n20496), .ZN(n16599) );
  AOI211_X1 U18550 ( .C1(n20505), .C2(n16601), .A(n16600), .B(n16599), .ZN(
        n16602) );
  OAI21_X1 U18551 ( .B1(n16751), .B2(n22141), .A(n16602), .ZN(P1_U2975) );
  NAND2_X1 U18552 ( .A1(n16604), .A2(n16603), .ZN(n16606) );
  XNOR2_X1 U18553 ( .A(n16606), .B(n16605), .ZN(n22005) );
  INV_X1 U18554 ( .A(n16607), .ZN(n16611) );
  AOI22_X1 U18555 ( .A1(n20514), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n22016), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16608) );
  OAI21_X1 U18556 ( .B1(n20522), .B2(n16609), .A(n16608), .ZN(n16610) );
  AOI21_X1 U18557 ( .B1(n16611), .B2(n20519), .A(n16610), .ZN(n16612) );
  OAI21_X1 U18558 ( .B1(n22141), .B2(n22005), .A(n16612), .ZN(P1_U2977) );
  AND2_X1 U18559 ( .A1(n22016), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16759) );
  NOR2_X1 U18560 ( .A1(n20522), .A2(n16613), .ZN(n16614) );
  AOI211_X1 U18561 ( .C1(n20514), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16759), .B(n16614), .ZN(n16620) );
  XNOR2_X1 U18562 ( .A(n20516), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16633) );
  NAND2_X1 U18563 ( .A1(n16634), .A2(n16633), .ZN(n21971) );
  OR2_X1 U18564 ( .A1(n16778), .A2(n16615), .ZN(n16616) );
  MUX2_X1 U18565 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n20511), .S(
        n16779), .Z(n16621) );
  INV_X1 U18566 ( .A(n20511), .ZN(n16622) );
  MUX2_X1 U18567 ( .A(n21995), .B(n16622), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n16617) );
  NAND2_X1 U18568 ( .A1(n16621), .A2(n16617), .ZN(n16618) );
  XNOR2_X1 U18569 ( .A(n16618), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16768) );
  NAND2_X1 U18570 ( .A1(n16768), .A2(n20518), .ZN(n16619) );
  OAI211_X1 U18571 ( .C1(n22115), .C2(n20496), .A(n16620), .B(n16619), .ZN(
        P1_U2978) );
  OAI21_X1 U18572 ( .B1(n21995), .B2(n16622), .A(n16621), .ZN(n16623) );
  XOR2_X1 U18573 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n16623), .Z(
        n16777) );
  NAND2_X1 U18574 ( .A1(n21906), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16772) );
  OAI21_X1 U18575 ( .B1(n16670), .B2(n16624), .A(n16772), .ZN(n16627) );
  NOR2_X1 U18576 ( .A1(n16625), .A2(n20496), .ZN(n16626) );
  AOI211_X1 U18577 ( .C1(n20505), .C2(n16628), .A(n16627), .B(n16626), .ZN(
        n16629) );
  OAI21_X1 U18578 ( .B1(n22141), .B2(n16777), .A(n16629), .ZN(P1_U2979) );
  OAI22_X1 U18579 ( .A1(n16670), .A2(n16630), .B1(n22001), .B2(n20414), .ZN(
        n16631) );
  AOI21_X1 U18580 ( .B1(n16632), .B2(n20505), .A(n16631), .ZN(n16636) );
  OR2_X1 U18581 ( .A1(n16634), .A2(n16633), .ZN(n21972) );
  NAND3_X1 U18582 ( .A1(n21972), .A2(n21971), .A3(n20518), .ZN(n16635) );
  OAI211_X1 U18583 ( .C1(n16637), .C2(n20496), .A(n16636), .B(n16635), .ZN(
        P1_U2981) );
  OAI211_X1 U18584 ( .C1(n16641), .C2(n16640), .A(n16650), .B(n16639), .ZN(
        n16793) );
  NAND2_X1 U18585 ( .A1(n16779), .A2(n16796), .ZN(n16643) );
  NAND3_X1 U18586 ( .A1(n16793), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16778), .ZN(n16642) );
  OAI21_X1 U18587 ( .B1(n16793), .B2(n16643), .A(n16642), .ZN(n16644) );
  XNOR2_X1 U18588 ( .A(n16644), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n21990) );
  NOR2_X1 U18589 ( .A1(n22001), .A2(n20410), .ZN(n21987) );
  AOI21_X1 U18590 ( .B1(n20514), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n21987), .ZN(n16645) );
  OAI21_X1 U18591 ( .B1(n20522), .B2(n16646), .A(n16645), .ZN(n16647) );
  AOI21_X1 U18592 ( .B1(n16648), .B2(n20519), .A(n16647), .ZN(n16649) );
  OAI21_X1 U18593 ( .B1(n21990), .B2(n22141), .A(n16649), .ZN(P1_U2983) );
  INV_X1 U18594 ( .A(n16650), .ZN(n16652) );
  NAND2_X1 U18595 ( .A1(n16654), .A2(n16653), .ZN(n16656) );
  XNOR2_X1 U18596 ( .A(n20516), .B(n21867), .ZN(n16655) );
  XNOR2_X1 U18597 ( .A(n16656), .B(n16655), .ZN(n21872) );
  NAND2_X1 U18598 ( .A1(n21872), .A2(n20518), .ZN(n16660) );
  NOR2_X1 U18599 ( .A1(n22001), .A2(n20407), .ZN(n21871) );
  NOR2_X1 U18600 ( .A1(n20522), .A2(n16657), .ZN(n16658) );
  AOI211_X1 U18601 ( .C1(n20514), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n21871), .B(n16658), .ZN(n16659) );
  OAI211_X1 U18602 ( .C1(n20496), .C2(n16661), .A(n16660), .B(n16659), .ZN(
        P1_U2985) );
  INV_X1 U18603 ( .A(n16662), .ZN(n16663) );
  AND2_X1 U18604 ( .A1(n16665), .A2(n16666), .ZN(n16800) );
  NAND2_X1 U18605 ( .A1(n16801), .A2(n16800), .ZN(n16799) );
  NAND2_X1 U18606 ( .A1(n16799), .A2(n16666), .ZN(n16667) );
  XOR2_X1 U18607 ( .A(n16668), .B(n16667), .Z(n21863) );
  NAND2_X1 U18608 ( .A1(n21863), .A2(n20518), .ZN(n16674) );
  INV_X1 U18609 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16669) );
  OAI22_X1 U18610 ( .A1(n16670), .A2(n16669), .B1(n22001), .B2(n21853), .ZN(
        n16671) );
  AOI21_X1 U18611 ( .B1(n20505), .B2(n16672), .A(n16671), .ZN(n16673) );
  OAI211_X1 U18612 ( .C1(n20496), .C2(n16675), .A(n16674), .B(n16673), .ZN(
        P1_U2986) );
  NOR2_X1 U18613 ( .A1(n16677), .A2(n15658), .ZN(n16813) );
  AOI21_X1 U18614 ( .B1(n15658), .B2(n16677), .A(n16813), .ZN(n21964) );
  NAND2_X1 U18615 ( .A1(n21964), .A2(n20518), .ZN(n16682) );
  NAND2_X1 U18616 ( .A1(n21906), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n21961) );
  INV_X1 U18617 ( .A(n21961), .ZN(n16680) );
  NOR2_X1 U18618 ( .A1(n20522), .A2(n16678), .ZN(n16679) );
  AOI211_X1 U18619 ( .C1(n20514), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16680), .B(n16679), .ZN(n16681) );
  OAI211_X1 U18620 ( .C1(n20496), .C2(n16683), .A(n16682), .B(n16681), .ZN(
        P1_U2989) );
  INV_X1 U18621 ( .A(n16684), .ZN(n16692) );
  OAI21_X1 U18622 ( .B1(n16686), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16685), .ZN(n16691) );
  NAND2_X1 U18623 ( .A1(n16687), .A2(n16716), .ZN(n16695) );
  AOI21_X1 U18624 ( .B1(n16695), .B2(n16689), .A(n16688), .ZN(n16690) );
  AOI211_X1 U18625 ( .C1(n16692), .C2(n22017), .A(n16691), .B(n16690), .ZN(
        n16693) );
  OAI21_X1 U18626 ( .B1(n16694), .B2(n22004), .A(n16693), .ZN(P1_U3001) );
  INV_X1 U18627 ( .A(n16695), .ZN(n16702) );
  INV_X1 U18628 ( .A(n16696), .ZN(n16699) );
  NAND3_X1 U18629 ( .A1(n16722), .A2(n16705), .A3(n16697), .ZN(n16698) );
  OAI211_X1 U18630 ( .C1(n16700), .C2(n22014), .A(n16699), .B(n16698), .ZN(
        n16701) );
  AOI21_X1 U18631 ( .B1(n16702), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16701), .ZN(n16703) );
  OAI21_X1 U18632 ( .B1(n16704), .B2(n22004), .A(n16703), .ZN(P1_U3002) );
  NOR2_X1 U18633 ( .A1(n16706), .A2(n16705), .ZN(n16710) );
  OAI21_X1 U18634 ( .B1(n16708), .B2(n22014), .A(n16707), .ZN(n16709) );
  AOI21_X1 U18635 ( .B1(n16722), .B2(n16710), .A(n16709), .ZN(n16712) );
  INV_X1 U18636 ( .A(n16718), .ZN(n16731) );
  NAND3_X1 U18637 ( .A1(n16731), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16716), .ZN(n16711) );
  OAI211_X1 U18638 ( .C1(n16713), .C2(n22004), .A(n16712), .B(n16711), .ZN(
        P1_U3003) );
  OAI21_X1 U18639 ( .B1(n16715), .B2(n22014), .A(n16714), .ZN(n16720) );
  INV_X1 U18640 ( .A(n16716), .ZN(n16717) );
  NOR3_X1 U18641 ( .A1(n16718), .A2(n16717), .A3(n16721), .ZN(n16719) );
  AOI211_X1 U18642 ( .C1(n16722), .C2(n16721), .A(n16720), .B(n16719), .ZN(
        n16723) );
  OAI21_X1 U18643 ( .B1(n16724), .B2(n22004), .A(n16723), .ZN(P1_U3004) );
  OAI21_X1 U18644 ( .B1(n22022), .B2(n16726), .A(n16725), .ZN(n16730) );
  OAI21_X1 U18645 ( .B1(n16728), .B2(n22014), .A(n16727), .ZN(n16729) );
  AOI21_X1 U18646 ( .B1(n16731), .B2(n16730), .A(n16729), .ZN(n16732) );
  OAI21_X1 U18647 ( .B1(n16733), .B2(n22004), .A(n16732), .ZN(P1_U3005) );
  INV_X1 U18648 ( .A(n16734), .ZN(n16740) );
  INV_X1 U18649 ( .A(n16735), .ZN(n16744) );
  NOR3_X1 U18650 ( .A1(n22022), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n16744), .ZN(n16739) );
  OAI21_X1 U18651 ( .B1(n16737), .B2(n22014), .A(n16736), .ZN(n16738) );
  AOI211_X1 U18652 ( .C1(n16740), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16739), .B(n16738), .ZN(n16741) );
  OAI21_X1 U18653 ( .B1(n16742), .B2(n22004), .A(n16741), .ZN(P1_U3006) );
  INV_X1 U18654 ( .A(n22022), .ZN(n16745) );
  NAND3_X1 U18655 ( .A1(n16745), .A2(n16744), .A3(n16743), .ZN(n16747) );
  OAI211_X1 U18656 ( .C1(n22014), .C2(n16748), .A(n16747), .B(n16746), .ZN(
        n16749) );
  AOI21_X1 U18657 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n22015), .A(
        n16749), .ZN(n16750) );
  OAI21_X1 U18658 ( .B1(n16751), .B2(n22004), .A(n16750), .ZN(P1_U3007) );
  INV_X1 U18659 ( .A(n16770), .ZN(n16754) );
  OR2_X1 U18660 ( .A1(n21932), .A2(n16752), .ZN(n16753) );
  OAI211_X1 U18661 ( .C1(n21884), .C2(n16754), .A(n21880), .B(n16753), .ZN(
        n21997) );
  INV_X1 U18662 ( .A(n16764), .ZN(n16755) );
  OR2_X1 U18663 ( .A1(n21997), .A2(n16755), .ZN(n16757) );
  NAND2_X1 U18664 ( .A1(n16785), .A2(n21880), .ZN(n16756) );
  NAND2_X1 U18665 ( .A1(n16757), .A2(n16756), .ZN(n22008) );
  INV_X1 U18666 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n22003) );
  INV_X1 U18667 ( .A(n16758), .ZN(n22119) );
  AOI21_X1 U18668 ( .B1(n22017), .B2(n22119), .A(n16759), .ZN(n16766) );
  NAND2_X1 U18669 ( .A1(n21952), .A2(n16760), .ZN(n16763) );
  NAND2_X1 U18670 ( .A1(n16761), .A2(n21877), .ZN(n16762) );
  NAND2_X1 U18671 ( .A1(n16763), .A2(n16762), .ZN(n16816) );
  NAND2_X1 U18672 ( .A1(n16816), .A2(n16764), .ZN(n22002) );
  NOR2_X1 U18673 ( .A1(n22002), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n22009) );
  INV_X1 U18674 ( .A(n22009), .ZN(n16765) );
  OAI211_X1 U18675 ( .C1(n22008), .C2(n22003), .A(n16766), .B(n16765), .ZN(
        n16767) );
  AOI21_X1 U18676 ( .B1(n16768), .B2(n22018), .A(n16767), .ZN(n16769) );
  INV_X1 U18677 ( .A(n16769), .ZN(P1_U3010) );
  INV_X1 U18678 ( .A(n16816), .ZN(n16804) );
  NOR2_X1 U18679 ( .A1(n16804), .A2(n16770), .ZN(n21996) );
  XNOR2_X1 U18680 ( .A(n21995), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16771) );
  NAND2_X1 U18681 ( .A1(n21996), .A2(n16771), .ZN(n16773) );
  OAI211_X1 U18682 ( .C1(n22014), .C2(n16774), .A(n16773), .B(n16772), .ZN(
        n16775) );
  AOI21_X1 U18683 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n21997), .A(
        n16775), .ZN(n16776) );
  OAI21_X1 U18684 ( .B1(n16777), .B2(n22004), .A(n16776), .ZN(P1_U3011) );
  NAND2_X1 U18685 ( .A1(n16778), .A2(n21984), .ZN(n16782) );
  AOI21_X1 U18686 ( .B1(n16779), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16793), .ZN(n16780) );
  MUX2_X1 U18687 ( .A(n16782), .B(n16781), .S(n16780), .Z(n16783) );
  XOR2_X1 U18688 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n16783), .Z(
        n20509) );
  NAND3_X1 U18689 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n16816), .ZN(n21973) );
  NOR2_X1 U18690 ( .A1(n21974), .A2(n21973), .ZN(n16794) );
  AOI21_X1 U18691 ( .B1(n21984), .B2(n16794), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16788) );
  INV_X1 U18692 ( .A(n21975), .ZN(n16786) );
  NOR2_X1 U18693 ( .A1(n21873), .A2(n21854), .ZN(n21849) );
  AOI21_X1 U18694 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21849), .A(
        n21932), .ZN(n16784) );
  OAI21_X1 U18695 ( .B1(n21884), .B2(n21856), .A(n21880), .ZN(n21851) );
  AOI211_X1 U18696 ( .C1(n21952), .C2(n21974), .A(n16784), .B(n21851), .ZN(
        n21981) );
  OAI21_X1 U18697 ( .B1(n16786), .B2(n16785), .A(n21981), .ZN(n21970) );
  INV_X1 U18698 ( .A(n21970), .ZN(n16787) );
  OAI22_X1 U18699 ( .A1(n22001), .A2(n20413), .B1(n16788), .B2(n16787), .ZN(
        n16789) );
  AOI21_X1 U18700 ( .B1(n22017), .B2(n16790), .A(n16789), .ZN(n16791) );
  OAI21_X1 U18701 ( .B1(n20509), .B2(n22004), .A(n16791), .ZN(P1_U3014) );
  XNOR2_X1 U18702 ( .A(n12520), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16792) );
  XNOR2_X1 U18703 ( .A(n16793), .B(n16792), .ZN(n20503) );
  INV_X1 U18704 ( .A(n16794), .ZN(n21983) );
  NAND2_X1 U18705 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n21906), .ZN(n16795) );
  OAI221_X1 U18706 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21983), 
        .C1(n16796), .C2(n21981), .A(n16795), .ZN(n16797) );
  AOI21_X1 U18707 ( .B1(n22084), .B2(n22017), .A(n16797), .ZN(n16798) );
  OAI21_X1 U18708 ( .B1(n20503), .B2(n22004), .A(n16798), .ZN(P1_U3016) );
  OAI21_X1 U18709 ( .B1(n16801), .B2(n16800), .A(n16799), .ZN(n16802) );
  INV_X1 U18710 ( .A(n16802), .ZN(n20500) );
  NAND3_X1 U18711 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16803), .A3(
        n16816), .ZN(n16812) );
  NOR2_X1 U18712 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16804), .ZN(
        n16810) );
  INV_X1 U18713 ( .A(n21932), .ZN(n16806) );
  AOI21_X1 U18714 ( .B1(n16805), .B2(n16806), .A(n21934), .ZN(n21949) );
  AOI22_X1 U18715 ( .A1(n21952), .A2(n16807), .B1(n21965), .B2(n16806), .ZN(
        n16808) );
  NAND2_X1 U18716 ( .A1(n21949), .A2(n16808), .ZN(n16817) );
  OAI22_X1 U18717 ( .A1(n20404), .A2(n22001), .B1(n22014), .B2(n22070), .ZN(
        n16809) );
  AOI221_X1 U18718 ( .B1(n16810), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C1(n16817), .C2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16809), .ZN(
        n16811) );
  OAI211_X1 U18719 ( .C1(n20500), .C2(n22004), .A(n16812), .B(n16811), .ZN(
        P1_U3019) );
  MUX2_X1 U18720 ( .A(n11239), .B(n20516), .S(n16813), .Z(n16814) );
  AOI22_X1 U18721 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16817), .B1(
        n16816), .B2(n16815), .ZN(n16819) );
  NOR2_X1 U18722 ( .A1(n22062), .A2(n22001), .ZN(n20494) );
  AOI21_X1 U18723 ( .B1(n22017), .B2(n22057), .A(n20494), .ZN(n16818) );
  OAI211_X1 U18724 ( .C1(n20493), .C2(n22004), .A(n16819), .B(n16818), .ZN(
        P1_U3020) );
  NOR2_X1 U18725 ( .A1(n16820), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16821) );
  OAI22_X1 U18726 ( .A1(n16824), .A2(n16821), .B1(n15410), .B2(n16827), .ZN(
        n16822) );
  MUX2_X1 U18727 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16822), .S(
        n17556), .Z(P1_U3477) );
  MUX2_X1 U18728 ( .A(n16824), .B(n16823), .S(n12463), .Z(n16825) );
  OAI21_X1 U18729 ( .B1(n16827), .B2(n16826), .A(n16825), .ZN(n16828) );
  MUX2_X1 U18730 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n16828), .S(
        n17556), .Z(P1_U3476) );
  OR2_X1 U18731 ( .A1(n15410), .A2(n16829), .ZN(n16835) );
  NOR2_X1 U18732 ( .A1(n11719), .A2(n16830), .ZN(n16838) );
  AOI22_X1 U18733 ( .A1(n16833), .A2(n16832), .B1(n16838), .B2(n16831), .ZN(
        n16834) );
  NAND2_X1 U18734 ( .A1(n16835), .A2(n16834), .ZN(n17516) );
  INV_X1 U18735 ( .A(n17516), .ZN(n16840) );
  NOR2_X1 U18736 ( .A1(n15288), .A2(n21878), .ZN(n16845) );
  AOI22_X1 U18737 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n16836), .B2(n21879), .ZN(
        n16844) );
  INV_X1 U18738 ( .A(n16844), .ZN(n16837) );
  AOI22_X1 U18739 ( .A1(n22156), .A2(n16838), .B1(n16845), .B2(n16837), .ZN(
        n16839) );
  OAI21_X1 U18740 ( .B1(n16840), .B2(n20525), .A(n16839), .ZN(n16841) );
  MUX2_X1 U18741 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16841), .S(
        n22149), .Z(P1_U3473) );
  OAI21_X1 U18742 ( .B1(n16843), .B2(n16842), .A(n22146), .ZN(n16847) );
  NAND2_X1 U18743 ( .A1(n16845), .A2(n16844), .ZN(n16846) );
  OAI211_X1 U18744 ( .C1(n16849), .C2(n16848), .A(n16847), .B(n16846), .ZN(
        n16850) );
  MUX2_X1 U18745 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16850), .S(
        n22149), .Z(P1_U3472) );
  NOR3_X1 U18746 ( .A1(n22411), .A2(n16887), .A3(n22290), .ZN(n16851) );
  NOR2_X1 U18747 ( .A1(n16851), .A2(n22236), .ZN(n16856) );
  INV_X1 U18748 ( .A(n16852), .ZN(n22287) );
  NAND2_X1 U18749 ( .A1(n22287), .A2(n15410), .ZN(n16857) );
  INV_X1 U18750 ( .A(n16853), .ZN(n22241) );
  NOR2_X1 U18751 ( .A1(n22241), .A2(n16854), .ZN(n16860) );
  INV_X1 U18752 ( .A(n16860), .ZN(n22273) );
  OAI22_X1 U18753 ( .A1(n16856), .A2(n16857), .B1(n22289), .B2(n22273), .ZN(
        n22563) );
  OR2_X1 U18754 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16855), .ZN(
        n22561) );
  INV_X1 U18755 ( .A(n16856), .ZN(n16858) );
  AOI22_X1 U18756 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22561), .B1(n16858), 
        .B2(n16857), .ZN(n16859) );
  AOI22_X1 U18757 ( .A1(n16887), .A2(n16861), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n22564), .ZN(n16862) );
  OAI21_X1 U18758 ( .B1(n22266), .B2(n22561), .A(n16862), .ZN(n16863) );
  AOI21_X1 U18759 ( .B1(n22411), .B2(n22299), .A(n16863), .ZN(n16864) );
  OAI21_X1 U18760 ( .B1(n16893), .B2(n16865), .A(n16864), .ZN(P1_U3129) );
  AOI22_X1 U18761 ( .A1(n16887), .A2(n16866), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n22564), .ZN(n16867) );
  OAI21_X1 U18762 ( .B1(n22308), .B2(n22561), .A(n16867), .ZN(n16868) );
  AOI21_X1 U18763 ( .B1(n22411), .B2(n22327), .A(n16868), .ZN(n16869) );
  OAI21_X1 U18764 ( .B1(n16893), .B2(n16870), .A(n16869), .ZN(P1_U3130) );
  INV_X1 U18765 ( .A(n22342), .ZN(n22356) );
  AOI22_X1 U18766 ( .A1(n16887), .A2(n16871), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n22564), .ZN(n16872) );
  OAI21_X1 U18767 ( .B1(n22341), .B2(n22561), .A(n16872), .ZN(n16873) );
  AOI21_X1 U18768 ( .B1(n22411), .B2(n22356), .A(n16873), .ZN(n16874) );
  OAI21_X1 U18769 ( .B1(n16893), .B2(n16875), .A(n16874), .ZN(P1_U3131) );
  AOI22_X1 U18770 ( .A1(n16887), .A2(n16876), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n22564), .ZN(n16877) );
  OAI21_X1 U18771 ( .B1(n22370), .B2(n22561), .A(n16877), .ZN(n16878) );
  AOI21_X1 U18772 ( .B1(n22411), .B2(n22379), .A(n16878), .ZN(n16879) );
  OAI21_X1 U18773 ( .B1(n16893), .B2(n16880), .A(n16879), .ZN(P1_U3132) );
  AOI22_X1 U18774 ( .A1(n16887), .A2(n16881), .B1(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n22564), .ZN(n16882) );
  OAI21_X1 U18775 ( .B1(n22441), .B2(n22561), .A(n16882), .ZN(n16883) );
  AOI21_X1 U18776 ( .B1(n22411), .B2(n22456), .A(n16883), .ZN(n16884) );
  OAI21_X1 U18777 ( .B1(n16893), .B2(n16885), .A(n16884), .ZN(P1_U3134) );
  AOI22_X1 U18778 ( .A1(n16887), .A2(n16886), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n22564), .ZN(n16888) );
  OAI21_X1 U18779 ( .B1(n16889), .B2(n22561), .A(n16888), .ZN(n16890) );
  AOI21_X1 U18780 ( .B1(n22411), .B2(n22470), .A(n16890), .ZN(n16891) );
  OAI21_X1 U18781 ( .B1(n16893), .B2(n16892), .A(n16891), .ZN(P1_U3135) );
  MUX2_X1 U18782 ( .A(n16894), .B(P2_EBX_REG_31__SCAN_IN), .S(n16966), .Z(
        P2_U2856) );
  NAND2_X1 U18783 ( .A1(n16895), .A2(n16896), .ZN(n16898) );
  XNOR2_X1 U18784 ( .A(n16898), .B(n16897), .ZN(n16980) );
  OR2_X1 U18785 ( .A1(n16908), .A2(n16899), .ZN(n16900) );
  NAND2_X1 U18786 ( .A1(n16901), .A2(n16900), .ZN(n17173) );
  NOR2_X1 U18787 ( .A1(n16966), .A2(n17173), .ZN(n16902) );
  AOI21_X1 U18788 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16966), .A(n16902), .ZN(
        n16903) );
  OAI21_X1 U18789 ( .B1(n16980), .B2(n16968), .A(n16903), .ZN(P2_U2859) );
  NAND2_X1 U18790 ( .A1(n16904), .A2(n16895), .ZN(n16906) );
  XNOR2_X1 U18791 ( .A(n16906), .B(n16905), .ZN(n16989) );
  OR2_X1 U18792 ( .A1(n16926), .A2(n16916), .ZN(n16918) );
  AND2_X1 U18793 ( .A1(n16918), .A2(n16907), .ZN(n16909) );
  OR2_X1 U18794 ( .A1(n16909), .A2(n16908), .ZN(n17185) );
  NOR2_X1 U18795 ( .A1(n16966), .A2(n17185), .ZN(n16910) );
  AOI21_X1 U18796 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16966), .A(n16910), .ZN(
        n16911) );
  OAI21_X1 U18797 ( .B1(n16989), .B2(n16968), .A(n16911), .ZN(P2_U2860) );
  OAI21_X1 U18798 ( .B1(n16914), .B2(n16913), .A(n16912), .ZN(n16998) );
  OR2_X1 U18799 ( .A1(n16952), .A2(n16915), .ZN(n16920) );
  NAND2_X1 U18800 ( .A1(n16926), .A2(n16916), .ZN(n16917) );
  NAND2_X1 U18801 ( .A1(n16918), .A2(n16917), .ZN(n18976) );
  NAND2_X1 U18802 ( .A1(n16952), .A2(n17198), .ZN(n16919) );
  OAI211_X1 U18803 ( .C1(n16998), .C2(n16968), .A(n16920), .B(n16919), .ZN(
        P2_U2861) );
  OAI21_X1 U18804 ( .B1(n16921), .B2(n16923), .A(n16922), .ZN(n17007) );
  NAND2_X1 U18805 ( .A1(n16936), .A2(n16924), .ZN(n16925) );
  AND2_X1 U18806 ( .A1(n16926), .A2(n16925), .ZN(n18965) );
  NOR2_X1 U18807 ( .A1(n16952), .A2(n13568), .ZN(n16927) );
  AOI21_X1 U18808 ( .B1(n18965), .B2(n16952), .A(n16927), .ZN(n16928) );
  OAI21_X1 U18809 ( .B1(n17007), .B2(n16968), .A(n16928), .ZN(P2_U2862) );
  OAI21_X1 U18810 ( .B1(n16931), .B2(n16930), .A(n16929), .ZN(n17015) );
  OR2_X1 U18811 ( .A1(n16952), .A2(n16932), .ZN(n16938) );
  OR2_X1 U18812 ( .A1(n16934), .A2(n16933), .ZN(n16935) );
  AND2_X1 U18813 ( .A1(n16936), .A2(n16935), .ZN(n18955) );
  NAND2_X1 U18814 ( .A1(n16952), .A2(n18955), .ZN(n16937) );
  OAI211_X1 U18815 ( .C1(n17015), .C2(n16968), .A(n16938), .B(n16937), .ZN(
        P2_U2863) );
  XNOR2_X1 U18816 ( .A(n16946), .B(n16940), .ZN(n17024) );
  NAND2_X1 U18817 ( .A1(n16941), .A2(n16950), .ZN(n16942) );
  NOR2_X1 U18818 ( .A1(n16966), .A2(n17101), .ZN(n16943) );
  AOI21_X1 U18819 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16966), .A(n16943), .ZN(
        n16944) );
  OAI21_X1 U18820 ( .B1(n17024), .B2(n16968), .A(n16944), .ZN(P2_U2864) );
  OAI21_X1 U18821 ( .B1(n16945), .B2(n16947), .A(n16946), .ZN(n19855) );
  NAND2_X1 U18822 ( .A1(n16966), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16954) );
  OR2_X1 U18823 ( .A1(n16948), .A2(n16949), .ZN(n16951) );
  AND2_X1 U18824 ( .A1(n16951), .A2(n16950), .ZN(n18932) );
  NAND2_X1 U18825 ( .A1(n18932), .A2(n16952), .ZN(n16953) );
  OAI211_X1 U18826 ( .C1(n19855), .C2(n16968), .A(n16954), .B(n16953), .ZN(
        P2_U2865) );
  INV_X1 U18827 ( .A(n16945), .ZN(n16956) );
  OAI21_X1 U18828 ( .B1(n16955), .B2(n16957), .A(n16956), .ZN(n17033) );
  NOR2_X1 U18829 ( .A1(n16959), .A2(n16958), .ZN(n16960) );
  OR2_X1 U18830 ( .A1(n16948), .A2(n16960), .ZN(n17252) );
  NOR2_X1 U18831 ( .A1(n17252), .A2(n16966), .ZN(n16961) );
  AOI21_X1 U18832 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n16966), .A(n16961), .ZN(
        n16962) );
  OAI21_X1 U18833 ( .B1(n17033), .B2(n16968), .A(n16962), .ZN(P2_U2866) );
  AND2_X1 U18834 ( .A1(n16044), .A2(n16963), .ZN(n16964) );
  OR2_X1 U18835 ( .A1(n16964), .A2(n16955), .ZN(n19959) );
  NOR2_X1 U18836 ( .A1(n16966), .A2(n18916), .ZN(n16965) );
  AOI21_X1 U18837 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n16966), .A(n16965), .ZN(
        n16967) );
  OAI21_X1 U18838 ( .B1(n19959), .B2(n16968), .A(n16967), .ZN(P2_U2867) );
  INV_X1 U18839 ( .A(P2_EAX_REG_31__SCAN_IN), .ZN(n16969) );
  OAI22_X1 U18840 ( .A1(n20164), .A2(n19052), .B1(n16969), .B2(n20162), .ZN(
        n16970) );
  AOI21_X1 U18841 ( .B1(n19957), .B2(BUF1_REG_31__SCAN_IN), .A(n16970), .ZN(
        n16971) );
  OAI21_X1 U18842 ( .B1(n16972), .B2(n19200), .A(n16971), .ZN(P2_U2888) );
  OR2_X1 U18843 ( .A1(n16983), .A2(n16973), .ZN(n16974) );
  INV_X1 U18844 ( .A(n19000), .ZN(n16976) );
  OAI22_X1 U18845 ( .A1(n20164), .A2(n16976), .B1(n14112), .B2(n20162), .ZN(
        n16977) );
  AOI21_X1 U18846 ( .B1(n19955), .B2(n19644), .A(n16977), .ZN(n16979) );
  AOI22_X1 U18847 ( .A1(n19956), .A2(BUF2_REG_28__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16978) );
  OAI211_X1 U18848 ( .C1(n16980), .C2(n20115), .A(n16979), .B(n16978), .ZN(
        P2_U2891) );
  NOR2_X1 U18849 ( .A1(n16992), .A2(n16981), .ZN(n16982) );
  OAI22_X1 U18850 ( .A1(n20164), .A2(n18995), .B1(n16984), .B2(n20162), .ZN(
        n16985) );
  AOI21_X1 U18851 ( .B1(n19955), .B2(n16986), .A(n16985), .ZN(n16988) );
  AOI22_X1 U18852 ( .A1(n19956), .A2(BUF2_REG_27__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16987) );
  OAI211_X1 U18853 ( .C1(n16989), .C2(n20115), .A(n16988), .B(n16987), .ZN(
        P2_U2892) );
  NOR2_X1 U18854 ( .A1(n17000), .A2(n16990), .ZN(n16991) );
  OR2_X1 U18855 ( .A1(n16992), .A2(n16991), .ZN(n18975) );
  OAI22_X1 U18856 ( .A1(n20164), .A2(n18975), .B1(n16993), .B2(n20162), .ZN(
        n16994) );
  AOI21_X1 U18857 ( .B1(n19955), .B2(n16995), .A(n16994), .ZN(n16997) );
  AOI22_X1 U18858 ( .A1(n19956), .A2(BUF2_REG_26__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16996) );
  OAI211_X1 U18859 ( .C1(n16998), .C2(n20115), .A(n16997), .B(n16996), .ZN(
        P2_U2893) );
  AND2_X1 U18860 ( .A1(n16999), .A2(n17008), .ZN(n17001) );
  OR2_X1 U18861 ( .A1(n17001), .A2(n17000), .ZN(n18963) );
  OAI22_X1 U18862 ( .A1(n20164), .A2(n18963), .B1(n17002), .B2(n20162), .ZN(
        n17003) );
  AOI21_X1 U18863 ( .B1(n19955), .B2(n17004), .A(n17003), .ZN(n17006) );
  AOI22_X1 U18864 ( .A1(n19956), .A2(BUF2_REG_25__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n17005) );
  OAI211_X1 U18865 ( .C1(n17007), .C2(n20115), .A(n17006), .B(n17005), .ZN(
        P2_U2894) );
  NAND2_X1 U18866 ( .A1(n11298), .A2(n17017), .ZN(n17009) );
  AND2_X1 U18867 ( .A1(n17009), .A2(n17008), .ZN(n18954) );
  INV_X1 U18868 ( .A(n18954), .ZN(n17218) );
  OAI22_X1 U18869 ( .A1(n20164), .A2(n17218), .B1(n17010), .B2(n20162), .ZN(
        n17011) );
  AOI21_X1 U18870 ( .B1(n19955), .B2(n17012), .A(n17011), .ZN(n17014) );
  AOI22_X1 U18871 ( .A1(n19956), .A2(BUF2_REG_24__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n17013) );
  OAI211_X1 U18872 ( .C1(n17015), .C2(n20115), .A(n17014), .B(n17013), .ZN(
        P2_U2895) );
  OAI21_X1 U18873 ( .B1(n17018), .B2(n17016), .A(n17017), .ZN(n18952) );
  OAI22_X1 U18874 ( .A1(n20164), .A2(n18952), .B1(n17019), .B2(n20162), .ZN(
        n17020) );
  AOI21_X1 U18875 ( .B1(n19955), .B2(n17021), .A(n17020), .ZN(n17023) );
  AOI22_X1 U18876 ( .A1(n19956), .A2(BUF2_REG_23__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n17022) );
  OAI211_X1 U18877 ( .C1(n17024), .C2(n20115), .A(n17023), .B(n17022), .ZN(
        P2_U2896) );
  OR2_X1 U18878 ( .A1(n17280), .A2(n17025), .ZN(n17027) );
  NAND2_X1 U18879 ( .A1(n17027), .A2(n17026), .ZN(n18930) );
  OAI22_X1 U18880 ( .A1(n20164), .A2(n18930), .B1(n17028), .B2(n20162), .ZN(
        n17029) );
  AOI21_X1 U18881 ( .B1(n19955), .B2(n17030), .A(n17029), .ZN(n17032) );
  AOI22_X1 U18882 ( .A1(n19956), .A2(BUF2_REG_21__SCAN_IN), .B1(n19957), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n17031) );
  OAI211_X1 U18883 ( .C1(n17033), .C2(n20115), .A(n17032), .B(n17031), .ZN(
        P2_U2898) );
  XNOR2_X1 U18884 ( .A(n17042), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n19047) );
  INV_X1 U18885 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n19025) );
  OAI21_X1 U18886 ( .B1(n17633), .B2(n19025), .A(n17034), .ZN(n17035) );
  AOI21_X1 U18887 ( .B1(n19029), .B2(n17673), .A(n17035), .ZN(n17036) );
  OAI21_X1 U18888 ( .B1(n19047), .B2(n17681), .A(n17036), .ZN(n17037) );
  AOI21_X1 U18889 ( .B1(n17038), .B2(n17671), .A(n17037), .ZN(n17039) );
  OAI21_X1 U18890 ( .B1(n17676), .B2(n17040), .A(n17039), .ZN(P2_U2984) );
  NOR2_X1 U18891 ( .A1(n17056), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17041) );
  OR2_X1 U18892 ( .A1(n17042), .A2(n17041), .ZN(n19018) );
  AOI21_X1 U18893 ( .B1(n17670), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17043), .ZN(n17045) );
  NAND2_X1 U18894 ( .A1(n16252), .A2(n17673), .ZN(n17044) );
  OAI211_X1 U18895 ( .C1(n19018), .C2(n17681), .A(n17045), .B(n17044), .ZN(
        n17046) );
  AOI21_X1 U18896 ( .B1(n17047), .B2(n17671), .A(n17046), .ZN(n17048) );
  OAI21_X1 U18897 ( .B1(n17676), .B2(n11216), .A(n17048), .ZN(P2_U2985) );
  XNOR2_X1 U18898 ( .A(n17072), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17183) );
  NOR2_X1 U18899 ( .A1(n17050), .A2(n17049), .ZN(n17051) );
  NAND2_X1 U18900 ( .A1(n17051), .A2(n11244), .ZN(n17063) );
  NOR2_X1 U18901 ( .A1(n17051), .A2(n11244), .ZN(n17065) );
  AOI21_X1 U18902 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17063), .A(
        n17065), .ZN(n17055) );
  XNOR2_X1 U18903 ( .A(n17053), .B(n17052), .ZN(n17054) );
  XNOR2_X1 U18904 ( .A(n17055), .B(n17054), .ZN(n17181) );
  AND2_X1 U18905 ( .A1(n17067), .A2(n18997), .ZN(n17057) );
  OR2_X1 U18906 ( .A1(n17057), .A2(n17056), .ZN(n19004) );
  NOR2_X1 U18907 ( .A1(n18813), .A2(n17058), .ZN(n17175) );
  NOR2_X1 U18908 ( .A1(n17657), .A2(n17173), .ZN(n17059) );
  AOI211_X1 U18909 ( .C1(n17670), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17175), .B(n17059), .ZN(n17060) );
  OAI21_X1 U18910 ( .B1(n19004), .B2(n17681), .A(n17060), .ZN(n17061) );
  AOI21_X1 U18911 ( .B1(n17181), .B2(n17671), .A(n17061), .ZN(n17062) );
  OAI21_X1 U18912 ( .B1(n17676), .B2(n17183), .A(n17062), .ZN(P2_U2986) );
  INV_X1 U18913 ( .A(n17063), .ZN(n17064) );
  NOR2_X1 U18914 ( .A1(n17065), .A2(n17064), .ZN(n17066) );
  XNOR2_X1 U18915 ( .A(n17066), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17196) );
  INV_X1 U18916 ( .A(n17067), .ZN(n17068) );
  AOI21_X1 U18917 ( .B1(n17069), .B2(n17081), .A(n17068), .ZN(n19002) );
  NOR2_X1 U18918 ( .A1(n18813), .A2(n17742), .ZN(n17187) );
  AOI21_X1 U18919 ( .B1(n17670), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17187), .ZN(n17070) );
  OAI21_X1 U18920 ( .B1(n17657), .B2(n17185), .A(n17070), .ZN(n17071) );
  AOI21_X1 U18921 ( .B1(n19002), .B2(n17640), .A(n17071), .ZN(n17074) );
  AOI21_X1 U18922 ( .B1(n17191), .B2(n17075), .A(n17072), .ZN(n17193) );
  NAND2_X1 U18923 ( .A1(n17193), .A2(n17664), .ZN(n17073) );
  OAI211_X1 U18924 ( .C1(n17196), .C2(n17608), .A(n17074), .B(n17073), .ZN(
        P2_U2987) );
  INV_X1 U18925 ( .A(n17086), .ZN(n17076) );
  OAI21_X1 U18926 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17076), .A(
        n17075), .ZN(n17204) );
  AOI21_X1 U18927 ( .B1(n17077), .B2(n17087), .A(n17088), .ZN(n17079) );
  XNOR2_X1 U18928 ( .A(n17079), .B(n17078), .ZN(n17203) );
  OR2_X1 U18929 ( .A1(n11275), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17080) );
  NAND2_X1 U18930 ( .A1(n17081), .A2(n17080), .ZN(n18980) );
  OR2_X1 U18931 ( .A1(n18813), .A2(n17741), .ZN(n17199) );
  OAI21_X1 U18932 ( .B1(n17633), .B2(n11517), .A(n17199), .ZN(n17082) );
  AOI21_X1 U18933 ( .B1(n17673), .B2(n17198), .A(n17082), .ZN(n17083) );
  OAI21_X1 U18934 ( .B1(n18980), .B2(n17681), .A(n17083), .ZN(n17084) );
  AOI21_X1 U18935 ( .B1(n17203), .B2(n17671), .A(n17084), .ZN(n17085) );
  OAI21_X1 U18936 ( .B1(n17676), .B2(n17204), .A(n17085), .ZN(P2_U2988) );
  OAI21_X1 U18937 ( .B1(n13081), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17086), .ZN(n17214) );
  INV_X1 U18938 ( .A(n17087), .ZN(n17089) );
  NOR2_X1 U18939 ( .A1(n17089), .A2(n17088), .ZN(n17090) );
  XNOR2_X1 U18940 ( .A(n17077), .B(n17090), .ZN(n17212) );
  NAND2_X1 U18941 ( .A1(n17212), .A2(n17671), .ZN(n17095) );
  AOI21_X1 U18942 ( .B1(n17668), .B2(n17092), .A(n11275), .ZN(n18966) );
  NAND2_X1 U18943 ( .A1(n17673), .A2(n18965), .ZN(n17091) );
  OR2_X1 U18944 ( .A1(n18813), .A2(n17740), .ZN(n17205) );
  OAI211_X1 U18945 ( .C1(n17633), .C2(n17092), .A(n17091), .B(n17205), .ZN(
        n17093) );
  AOI21_X1 U18946 ( .B1(n18966), .B2(n17640), .A(n17093), .ZN(n17094) );
  OAI211_X1 U18947 ( .C1(n17214), .C2(n17676), .A(n17095), .B(n17094), .ZN(
        P2_U2989) );
  NAND2_X1 U18948 ( .A1(n11262), .A2(n17096), .ZN(n17097) );
  INV_X1 U18949 ( .A(n17098), .ZN(n17112) );
  NAND2_X1 U18950 ( .A1(n17112), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17100) );
  AOI21_X1 U18951 ( .B1(n17232), .B2(n17100), .A(n17099), .ZN(n17229) );
  NAND2_X1 U18952 ( .A1(n17229), .A2(n17664), .ZN(n17105) );
  AOI21_X1 U18953 ( .B1(n18940), .B2(n17661), .A(n17669), .ZN(n18946) );
  OAI22_X1 U18954 ( .A1(n18940), .A2(n17633), .B1(n13161), .B2(n18813), .ZN(
        n17103) );
  NOR2_X1 U18955 ( .A1(n17657), .A2(n17101), .ZN(n17102) );
  AOI211_X1 U18956 ( .C1(n18946), .C2(n17640), .A(n17103), .B(n17102), .ZN(
        n17104) );
  OAI211_X1 U18957 ( .C1(n17608), .C2(n17238), .A(n17105), .B(n17104), .ZN(
        P2_U2991) );
  INV_X1 U18958 ( .A(n17106), .ZN(n17107) );
  NAND2_X1 U18959 ( .A1(n17109), .A2(n17108), .ZN(n17110) );
  XNOR2_X1 U18960 ( .A(n17111), .B(n17110), .ZN(n17262) );
  AOI21_X1 U18961 ( .B1(n17258), .B2(n17113), .A(n17112), .ZN(n17260) );
  AOI21_X1 U18962 ( .B1(n18918), .B2(n17114), .A(n17662), .ZN(n18924) );
  NAND2_X1 U18963 ( .A1(n19139), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n17253) );
  OAI21_X1 U18964 ( .B1(n17633), .B2(n18918), .A(n17253), .ZN(n17115) );
  AOI21_X1 U18965 ( .B1(n17640), .B2(n18924), .A(n17115), .ZN(n17116) );
  OAI21_X1 U18966 ( .B1(n17657), .B2(n17252), .A(n17116), .ZN(n17117) );
  AOI21_X1 U18967 ( .B1(n17260), .B2(n17664), .A(n17117), .ZN(n17118) );
  OAI21_X1 U18968 ( .B1(n17262), .B2(n17608), .A(n17118), .ZN(P2_U2993) );
  XNOR2_X1 U18969 ( .A(n17300), .B(n17293), .ZN(n17298) );
  AOI21_X1 U18970 ( .B1(n17651), .B2(n17120), .A(n11245), .ZN(n18898) );
  NAND2_X1 U18971 ( .A1(n17673), .A2(n18897), .ZN(n17119) );
  OR2_X1 U18972 ( .A1(n18813), .A2(n18894), .ZN(n17288) );
  OAI211_X1 U18973 ( .C1(n17120), .C2(n17633), .A(n17119), .B(n17288), .ZN(
        n17127) );
  NAND2_X1 U18974 ( .A1(n17121), .A2(n17302), .ZN(n17125) );
  NAND2_X1 U18975 ( .A1(n17123), .A2(n17122), .ZN(n17124) );
  XNOR2_X1 U18976 ( .A(n17125), .B(n17124), .ZN(n17287) );
  NOR2_X1 U18977 ( .A1(n17287), .A2(n17608), .ZN(n17126) );
  AOI211_X1 U18978 ( .C1(n17640), .C2(n18898), .A(n17127), .B(n17126), .ZN(
        n17128) );
  OAI21_X1 U18979 ( .B1(n17676), .B2(n17298), .A(n17128), .ZN(P2_U2995) );
  XNOR2_X1 U18980 ( .A(n19113), .B(n17316), .ZN(n17330) );
  AOI21_X1 U18981 ( .B1(n17615), .B2(n17130), .A(n17632), .ZN(n18840) );
  NAND2_X1 U18982 ( .A1(n17640), .A2(n18840), .ZN(n17129) );
  OR2_X1 U18983 ( .A1(n18813), .A2(n18839), .ZN(n17321) );
  OAI211_X1 U18984 ( .C1(n17130), .C2(n17633), .A(n17129), .B(n17321), .ZN(
        n17141) );
  INV_X1 U18985 ( .A(n17343), .ZN(n17131) );
  AND2_X1 U18986 ( .A1(n17134), .A2(n17133), .ZN(n17332) );
  NAND2_X1 U18987 ( .A1(n17333), .A2(n17332), .ZN(n17331) );
  NAND2_X1 U18988 ( .A1(n17331), .A2(n17134), .ZN(n17618) );
  AND2_X1 U18989 ( .A1(n17136), .A2(n17135), .ZN(n17617) );
  NAND2_X1 U18990 ( .A1(n17618), .A2(n17617), .ZN(n17620) );
  NAND2_X1 U18991 ( .A1(n17620), .A2(n17136), .ZN(n17139) );
  XNOR2_X1 U18992 ( .A(n17137), .B(n17316), .ZN(n17138) );
  XNOR2_X1 U18993 ( .A(n17139), .B(n17138), .ZN(n17325) );
  NOR2_X1 U18994 ( .A1(n17325), .A2(n17608), .ZN(n17140) );
  AOI211_X1 U18995 ( .C1(n17673), .C2(n18844), .A(n17141), .B(n17140), .ZN(
        n17142) );
  OAI21_X1 U18996 ( .B1(n17676), .B2(n17330), .A(n17142), .ZN(P2_U2999) );
  XNOR2_X1 U18997 ( .A(n17579), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17387) );
  NAND2_X1 U18998 ( .A1(n17144), .A2(n17582), .ZN(n17145) );
  XNOR2_X1 U18999 ( .A(n17143), .B(n17145), .ZN(n17385) );
  INV_X1 U19000 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17146) );
  OAI22_X1 U19001 ( .A1(n17146), .A2(n17633), .B1(n17681), .B2(n18780), .ZN(
        n17149) );
  OAI22_X1 U19002 ( .A1(n17657), .A2(n18783), .B1(n18892), .B2(n17147), .ZN(
        n17148) );
  AOI211_X1 U19003 ( .C1(n17385), .C2(n17671), .A(n17149), .B(n17148), .ZN(
        n17150) );
  OAI21_X1 U19004 ( .B1(n17387), .B2(n17676), .A(n17150), .ZN(P2_U3005) );
  NAND2_X1 U19005 ( .A1(n17152), .A2(n17151), .ZN(n17154) );
  XNOR2_X1 U19006 ( .A(n17154), .B(n17153), .ZN(n17399) );
  NOR2_X1 U19007 ( .A1(n17156), .A2(n17155), .ZN(n17158) );
  XOR2_X1 U19008 ( .A(n17158), .B(n17157), .Z(n17397) );
  INV_X1 U19009 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17159) );
  OAI22_X1 U19010 ( .A1(n17159), .A2(n17633), .B1(n17681), .B2(n18757), .ZN(
        n17162) );
  OAI22_X1 U19011 ( .A1(n17657), .A2(n18760), .B1(n18892), .B2(n17160), .ZN(
        n17161) );
  AOI211_X1 U19012 ( .C1(n17397), .C2(n17671), .A(n17162), .B(n17161), .ZN(
        n17163) );
  OAI21_X1 U19013 ( .B1(n17399), .B2(n17676), .A(n17163), .ZN(P2_U3007) );
  XNOR2_X1 U19014 ( .A(n17165), .B(n17164), .ZN(n17408) );
  XNOR2_X1 U19015 ( .A(n17166), .B(n17401), .ZN(n17410) );
  NAND2_X1 U19016 ( .A1(n17410), .A2(n17664), .ZN(n17172) );
  OAI22_X1 U19017 ( .A1(n17167), .A2(n17633), .B1(n13105), .B2(n18813), .ZN(
        n17170) );
  INV_X1 U19018 ( .A(n18751), .ZN(n17168) );
  NOR2_X1 U19019 ( .A1(n17168), .A2(n17657), .ZN(n17169) );
  AOI211_X1 U19020 ( .C1(n17640), .C2(n18750), .A(n17170), .B(n17169), .ZN(
        n17171) );
  OAI211_X1 U19021 ( .C1(n17608), .C2(n17408), .A(n17172), .B(n17171), .ZN(
        P2_U3008) );
  XNOR2_X1 U19022 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17179) );
  NOR2_X1 U19023 ( .A1(n19133), .A2(n17173), .ZN(n17174) );
  NAND2_X1 U19024 ( .A1(n17176), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17177) );
  OAI211_X1 U19025 ( .C1(n17184), .C2(n17179), .A(n17178), .B(n17177), .ZN(
        n17180) );
  AOI21_X1 U19026 ( .B1(n17181), .B2(n19138), .A(n17180), .ZN(n17182) );
  OAI21_X1 U19027 ( .B1(n19134), .B2(n17183), .A(n17182), .ZN(P2_U3018) );
  INV_X1 U19028 ( .A(n17184), .ZN(n17192) );
  INV_X1 U19029 ( .A(n17185), .ZN(n18992) );
  NOR2_X1 U19030 ( .A1(n19119), .A2(n18995), .ZN(n17186) );
  AOI211_X1 U19031 ( .C1(n18992), .C2(n19103), .A(n17187), .B(n17186), .ZN(
        n17188) );
  OAI21_X1 U19032 ( .B1(n17189), .B2(n17191), .A(n17188), .ZN(n17190) );
  AOI21_X1 U19033 ( .B1(n17192), .B2(n17191), .A(n17190), .ZN(n17195) );
  NAND2_X1 U19034 ( .A1(n17193), .A2(n19108), .ZN(n17194) );
  OAI211_X1 U19035 ( .C1(n17196), .C2(n19091), .A(n17195), .B(n17194), .ZN(
        P2_U3019) );
  XNOR2_X1 U19036 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17202) );
  INV_X1 U19037 ( .A(n17197), .ZN(n17208) );
  NAND2_X1 U19038 ( .A1(n19103), .A2(n17198), .ZN(n17200) );
  OAI211_X1 U19039 ( .C1(n19119), .C2(n18975), .A(n17200), .B(n17199), .ZN(
        n17201) );
  NAND2_X1 U19040 ( .A1(n19103), .A2(n18965), .ZN(n17206) );
  OAI211_X1 U19041 ( .C1(n18963), .C2(n19119), .A(n17206), .B(n17205), .ZN(
        n17207) );
  AOI21_X1 U19042 ( .B1(n17208), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17207), .ZN(n17209) );
  OAI21_X1 U19043 ( .B1(n17210), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17209), .ZN(n17211) );
  AOI21_X1 U19044 ( .B1(n17212), .B2(n19138), .A(n17211), .ZN(n17213) );
  OAI21_X1 U19045 ( .B1(n19134), .B2(n17214), .A(n17213), .ZN(P2_U3021) );
  OR2_X1 U19046 ( .A1(n17099), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17215) );
  NAND2_X1 U19047 ( .A1(n17216), .A2(n17215), .ZN(n17677) );
  OAI22_X1 U19048 ( .A1(n19119), .A2(n17218), .B1(n17217), .B2(n18892), .ZN(
        n17223) );
  OAI21_X1 U19049 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17220), .A(
        n17219), .ZN(n17221) );
  INV_X1 U19050 ( .A(n17221), .ZN(n17222) );
  AOI211_X1 U19051 ( .C1(n19103), .C2(n18955), .A(n17223), .B(n17222), .ZN(
        n17228) );
  XNOR2_X1 U19052 ( .A(n17225), .B(n11357), .ZN(n17226) );
  XNOR2_X1 U19053 ( .A(n17224), .B(n17226), .ZN(n17672) );
  NAND2_X1 U19054 ( .A1(n17672), .A2(n19138), .ZN(n17227) );
  OAI211_X1 U19055 ( .C1(n17677), .C2(n19134), .A(n17228), .B(n17227), .ZN(
        P2_U3022) );
  NAND2_X1 U19056 ( .A1(n17229), .A2(n19108), .ZN(n17237) );
  INV_X1 U19057 ( .A(n17257), .ZN(n17235) );
  AOI22_X1 U19058 ( .A1(n19103), .A2(n18945), .B1(n19139), .B2(
        P2_REIP_REG_23__SCAN_IN), .ZN(n17230) );
  OAI21_X1 U19059 ( .B1(n19119), .B2(n18952), .A(n17230), .ZN(n17234) );
  AOI211_X1 U19060 ( .C1(n17244), .C2(n17232), .A(n17231), .B(n17245), .ZN(
        n17233) );
  AOI211_X1 U19061 ( .C1(n17235), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17234), .B(n17233), .ZN(n17236) );
  OAI211_X1 U19062 ( .C1(n17238), .C2(n19091), .A(n17237), .B(n17236), .ZN(
        P2_U3023) );
  XNOR2_X1 U19063 ( .A(n17098), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17663) );
  NAND2_X1 U19064 ( .A1(n17663), .A2(n19108), .ZN(n17250) );
  AOI21_X1 U19065 ( .B1(n17239), .B2(n17026), .A(n17016), .ZN(n19856) );
  AOI22_X1 U19066 ( .A1(n18932), .A2(n19103), .B1(n19129), .B2(n19856), .ZN(
        n17249) );
  XNOR2_X1 U19067 ( .A(n17241), .B(n17244), .ZN(n17242) );
  XNOR2_X1 U19068 ( .A(n13554), .B(n17242), .ZN(n17665) );
  NAND2_X1 U19069 ( .A1(n17665), .A2(n19138), .ZN(n17248) );
  NAND2_X1 U19070 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19139), .ZN(n17243) );
  OAI221_X1 U19071 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17245), 
        .C1(n17244), .C2(n17257), .A(n17243), .ZN(n17246) );
  INV_X1 U19072 ( .A(n17246), .ZN(n17247) );
  NAND4_X1 U19073 ( .A1(n17250), .A2(n17249), .A3(n17248), .A4(n17247), .ZN(
        P2_U3024) );
  NAND2_X1 U19074 ( .A1(n17251), .A2(n17258), .ZN(n17256) );
  INV_X1 U19075 ( .A(n17252), .ZN(n18923) );
  OAI21_X1 U19076 ( .B1(n19119), .B2(n18930), .A(n17253), .ZN(n17254) );
  AOI21_X1 U19077 ( .B1(n19103), .B2(n18923), .A(n17254), .ZN(n17255) );
  OAI211_X1 U19078 ( .C1(n17258), .C2(n17257), .A(n17256), .B(n17255), .ZN(
        n17259) );
  AOI21_X1 U19079 ( .B1(n17260), .B2(n19108), .A(n17259), .ZN(n17261) );
  OAI21_X1 U19080 ( .B1(n17262), .B2(n19091), .A(n17261), .ZN(P2_U3025) );
  NOR3_X1 U19081 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17267), .A3(
        n19112), .ZN(n17306) );
  NAND2_X1 U19082 ( .A1(n17266), .A2(n17265), .ZN(n17317) );
  AOI21_X1 U19083 ( .B1(n17268), .B2(n17317), .A(n17267), .ZN(n17272) );
  INV_X1 U19084 ( .A(n17269), .ZN(n17270) );
  AOI21_X1 U19085 ( .B1(n19106), .B2(n17271), .A(n17270), .ZN(n17318) );
  OAI21_X1 U19086 ( .B1(n19109), .B2(n17272), .A(n17318), .ZN(n17307) );
  NOR2_X1 U19087 ( .A1(n17306), .A2(n17307), .ZN(n17294) );
  INV_X1 U19088 ( .A(n19112), .ZN(n17276) );
  NAND3_X1 U19089 ( .A1(n17276), .A2(n17273), .A3(n17293), .ZN(n17291) );
  AOI21_X1 U19090 ( .B1(n17294), .B2(n17291), .A(n17274), .ZN(n17285) );
  NAND3_X1 U19091 ( .A1(n17276), .A2(n17275), .A3(n17274), .ZN(n17283) );
  NOR2_X1 U19092 ( .A1(n17278), .A2(n17277), .ZN(n17279) );
  OR2_X1 U19093 ( .A1(n17280), .A2(n17279), .ZN(n19958) );
  INV_X1 U19094 ( .A(n19958), .ZN(n18910) );
  AOI21_X1 U19095 ( .B1(n19129), .B2(n18910), .A(n17281), .ZN(n17282) );
  OAI211_X1 U19096 ( .C1(n18916), .C2(n19133), .A(n17283), .B(n17282), .ZN(
        n17284) );
  INV_X1 U19097 ( .A(n17287), .ZN(n17296) );
  INV_X1 U19098 ( .A(n18897), .ZN(n17289) );
  OAI21_X1 U19099 ( .B1(n19133), .B2(n17289), .A(n17288), .ZN(n17290) );
  AOI21_X1 U19100 ( .B1(n19129), .B2(n18896), .A(n17290), .ZN(n17292) );
  OAI211_X1 U19101 ( .C1(n17294), .C2(n17293), .A(n17292), .B(n17291), .ZN(
        n17295) );
  AOI21_X1 U19102 ( .B1(n17296), .B2(n19138), .A(n17295), .ZN(n17297) );
  OAI21_X1 U19103 ( .B1(n19134), .B2(n17298), .A(n17297), .ZN(P2_U3027) );
  OR2_X1 U19104 ( .A1(n17645), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17299) );
  AND2_X1 U19105 ( .A1(n17300), .A2(n17299), .ZN(n17654) );
  INV_X1 U19106 ( .A(n17654), .ZN(n17312) );
  AND2_X1 U19107 ( .A1(n17302), .A2(n17301), .ZN(n17303) );
  XNOR2_X1 U19108 ( .A(n17304), .B(n17303), .ZN(n17653) );
  NOR2_X1 U19109 ( .A1(n13351), .A2(n18813), .ZN(n17305) );
  AOI211_X1 U19110 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n17307), .A(
        n17306), .B(n17305), .ZN(n17308) );
  INV_X1 U19111 ( .A(n17308), .ZN(n17310) );
  OAI22_X1 U19112 ( .A1(n19133), .A2(n18884), .B1(n19119), .B2(n18883), .ZN(
        n17309) );
  AOI211_X1 U19113 ( .C1(n17653), .C2(n19138), .A(n17310), .B(n17309), .ZN(
        n17311) );
  OAI21_X1 U19114 ( .B1(n19134), .B2(n17312), .A(n17311), .ZN(P2_U3028) );
  OR2_X1 U19115 ( .A1(n18829), .A2(n17313), .ZN(n17314) );
  NAND2_X1 U19116 ( .A1(n17315), .A2(n17314), .ZN(n19636) );
  INV_X1 U19117 ( .A(n19636), .ZN(n17328) );
  NOR2_X1 U19118 ( .A1(n17317), .A2(n17316), .ZN(n17320) );
  OAI21_X1 U19119 ( .B1(n17320), .B2(n17319), .A(n17318), .ZN(n19105) );
  INV_X1 U19120 ( .A(n18844), .ZN(n17322) );
  OAI21_X1 U19121 ( .B1(n17322), .B2(n19133), .A(n17321), .ZN(n17323) );
  AOI21_X1 U19122 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n19105), .A(
        n17323), .ZN(n17324) );
  OAI21_X1 U19123 ( .B1(n19112), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17324), .ZN(n17327) );
  NOR2_X1 U19124 ( .A1(n17325), .A2(n19091), .ZN(n17326) );
  AOI211_X1 U19125 ( .C1(n19129), .C2(n17328), .A(n17327), .B(n17326), .ZN(
        n17329) );
  OAI21_X1 U19126 ( .B1(n19134), .B2(n17330), .A(n17329), .ZN(P2_U3031) );
  XNOR2_X1 U19127 ( .A(n17621), .B(n13404), .ZN(n17607) );
  OAI21_X1 U19128 ( .B1(n17333), .B2(n17332), .A(n17331), .ZN(n17606) );
  INV_X1 U19129 ( .A(n17334), .ZN(n17335) );
  AOI21_X1 U19130 ( .B1(n17335), .B2(n17365), .A(n17381), .ZN(n17347) );
  OAI21_X1 U19131 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17349), .A(
        n17347), .ZN(n19096) );
  NOR2_X1 U19132 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17349), .ZN(
        n19097) );
  AOI22_X1 U19133 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19096), .B1(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n19097), .ZN(n17338) );
  INV_X1 U19134 ( .A(n17336), .ZN(n17611) );
  AOI22_X1 U19135 ( .A1(n19103), .A2(n17611), .B1(n19095), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n17337) );
  OAI211_X1 U19136 ( .C1(n19642), .C2(n19119), .A(n17338), .B(n17337), .ZN(
        n17339) );
  AOI21_X1 U19137 ( .B1(n17606), .B2(n19138), .A(n17339), .ZN(n17340) );
  OAI21_X1 U19138 ( .B1(n19134), .B2(n17607), .A(n17340), .ZN(P2_U3033) );
  INV_X1 U19139 ( .A(n17621), .ZN(n17341) );
  AOI21_X1 U19140 ( .B1(n17348), .B2(n17356), .A(n17341), .ZN(n17599) );
  INV_X1 U19141 ( .A(n17599), .ZN(n17354) );
  NAND2_X1 U19142 ( .A1(n17343), .A2(n17342), .ZN(n17344) );
  XNOR2_X1 U19143 ( .A(n17345), .B(n17344), .ZN(n17601) );
  NAND2_X1 U19144 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19139), .ZN(n17346) );
  OAI221_X1 U19145 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17349), 
        .C1(n17348), .C2(n17347), .A(n17346), .ZN(n17352) );
  AOI21_X1 U19146 ( .B1(n17362), .B2(n17350), .A(n15560), .ZN(n18820) );
  INV_X1 U19147 ( .A(n18820), .ZN(n19646) );
  OAI22_X1 U19148 ( .A1(n19646), .A2(n19119), .B1(n19133), .B2(n18823), .ZN(
        n17351) );
  AOI211_X1 U19149 ( .C1(n17601), .C2(n19138), .A(n17352), .B(n17351), .ZN(
        n17353) );
  OAI21_X1 U19150 ( .B1(n17354), .B2(n19134), .A(n17353), .ZN(P2_U3034) );
  INV_X1 U19151 ( .A(n17579), .ZN(n17355) );
  NOR2_X1 U19152 ( .A1(n17355), .A2(n17364), .ZN(n17580) );
  OAI21_X1 U19153 ( .B1(n17580), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17356), .ZN(n17595) );
  NOR2_X1 U19154 ( .A1(n17358), .A2(n17357), .ZN(n17361) );
  NOR2_X1 U19155 ( .A1(n11224), .A2(n17359), .ZN(n17360) );
  XOR2_X1 U19156 ( .A(n17361), .B(n17360), .Z(n17594) );
  NOR2_X1 U19157 ( .A1(n17594), .A2(n19091), .ZN(n17375) );
  OAI21_X1 U19158 ( .B1(n18791), .B2(n17363), .A(n17362), .ZN(n19649) );
  NOR2_X1 U19159 ( .A1(n19649), .A2(n19119), .ZN(n17374) );
  INV_X1 U19160 ( .A(n17367), .ZN(n17383) );
  NOR3_X1 U19161 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17364), .A3(
        n17383), .ZN(n17373) );
  AOI21_X1 U19162 ( .B1(n17366), .B2(n17365), .A(n17381), .ZN(n19080) );
  NAND3_X1 U19163 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17367), .A3(
        n13474), .ZN(n19079) );
  AOI21_X1 U19164 ( .B1(n19080), .B2(n19079), .A(n17368), .ZN(n17369) );
  INV_X1 U19165 ( .A(n17369), .ZN(n17371) );
  AOI22_X1 U19166 ( .A1(n19103), .A2(n18807), .B1(n19139), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n17370) );
  NAND2_X1 U19167 ( .A1(n17371), .A2(n17370), .ZN(n17372) );
  NOR4_X1 U19168 ( .A1(n17375), .A2(n17374), .A3(n17373), .A4(n17372), .ZN(
        n17376) );
  OAI21_X1 U19169 ( .B1(n19134), .B2(n17595), .A(n17376), .ZN(P2_U3035) );
  NOR2_X1 U19170 ( .A1(n19133), .A2(n18783), .ZN(n17380) );
  OR2_X1 U19171 ( .A1(n17377), .A2(n18771), .ZN(n17378) );
  NAND2_X1 U19172 ( .A1(n17378), .A2(n18792), .ZN(n19656) );
  OAI22_X1 U19173 ( .A1(n19119), .A2(n19656), .B1(n17147), .B2(n18813), .ZN(
        n17379) );
  AOI211_X1 U19174 ( .C1(n17381), .C2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17380), .B(n17379), .ZN(n17382) );
  OAI21_X1 U19175 ( .B1(n17383), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17382), .ZN(n17384) );
  AOI21_X1 U19176 ( .B1(n17385), .B2(n19138), .A(n17384), .ZN(n17386) );
  OAI21_X1 U19177 ( .B1(n17387), .B2(n19134), .A(n17386), .ZN(P2_U3037) );
  OAI21_X1 U19178 ( .B1(n19109), .B2(n17389), .A(n17388), .ZN(n19130) );
  NOR2_X1 U19179 ( .A1(n19133), .A2(n18760), .ZN(n17394) );
  OR2_X1 U19180 ( .A1(n17391), .A2(n17390), .ZN(n17392) );
  NAND2_X1 U19181 ( .A1(n17392), .A2(n18772), .ZN(n19663) );
  OAI22_X1 U19182 ( .A1(n19119), .A2(n19663), .B1(n17160), .B2(n18813), .ZN(
        n17393) );
  AOI211_X1 U19183 ( .C1(n19130), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17394), .B(n17393), .ZN(n17395) );
  OAI21_X1 U19184 ( .B1(n19140), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17395), .ZN(n17396) );
  AOI21_X1 U19185 ( .B1(n17397), .B2(n19138), .A(n17396), .ZN(n17398) );
  OAI21_X1 U19186 ( .B1(n17399), .B2(n19134), .A(n17398), .ZN(P2_U3039) );
  NOR2_X1 U19187 ( .A1(n13105), .A2(n18813), .ZN(n17400) );
  AOI221_X1 U19188 ( .B1(n17402), .B2(n17401), .C1(n19130), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n17400), .ZN(n17407) );
  XNOR2_X1 U19189 ( .A(n17403), .B(n17404), .ZN(n19863) );
  NOR2_X1 U19190 ( .A1(n19119), .A2(n19863), .ZN(n17405) );
  AOI21_X1 U19191 ( .B1(n18751), .B2(n19103), .A(n17405), .ZN(n17406) );
  OAI211_X1 U19192 ( .C1(n17408), .C2(n19091), .A(n17407), .B(n17406), .ZN(
        n17409) );
  AOI21_X1 U19193 ( .B1(n17410), .B2(n19108), .A(n17409), .ZN(n17411) );
  INV_X1 U19194 ( .A(n17411), .ZN(P2_U3040) );
  INV_X1 U19195 ( .A(n19148), .ZN(n17416) );
  OAI221_X1 U19196 ( .B1(n17413), .B2(n18778), .C1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17412), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17420) );
  INV_X1 U19197 ( .A(n17420), .ZN(n19056) );
  AOI21_X1 U19198 ( .B1(n18778), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17414), .ZN(n17421) );
  AOI222_X1 U19199 ( .A1(n17416), .A2(n17415), .B1(n19056), .B2(n17421), .C1(
        n19690), .C2(n19162), .ZN(n17418) );
  NAND2_X1 U19200 ( .A1(n19057), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17417) );
  OAI21_X1 U19201 ( .B1(n17418), .B2(n19057), .A(n17417), .ZN(P2_U3600) );
  INV_X1 U19202 ( .A(n19162), .ZN(n19054) );
  OAI222_X1 U19203 ( .A1(n17686), .A2(n19054), .B1(n17421), .B2(n17420), .C1(
        n19148), .C2(n17419), .ZN(n17423) );
  MUX2_X1 U19204 ( .A(n17423), .B(n17422), .S(n19057), .Z(P2_U3599) );
  NOR3_X1 U19205 ( .A1(n20251), .A2(n20259), .A3(n19838), .ZN(n17425) );
  AND2_X1 U19206 ( .A1(n19788), .A2(n22169), .ZN(n19839) );
  NOR2_X1 U19207 ( .A1(n17425), .A2(n19839), .ZN(n17434) );
  INV_X1 U19208 ( .A(n17434), .ZN(n17429) );
  NAND2_X1 U19209 ( .A1(n17426), .A2(n19786), .ZN(n17433) );
  NOR2_X1 U19210 ( .A1(n19757), .A2(n19835), .ZN(n20250) );
  AOI21_X1 U19211 ( .B1(n20250), .B2(n19846), .A(n19841), .ZN(n17428) );
  NAND2_X1 U19212 ( .A1(n12984), .A2(n19842), .ZN(n17427) );
  INV_X1 U19213 ( .A(n20256), .ZN(n17430) );
  NAND2_X1 U19214 ( .A1(n17430), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n17438) );
  AOI22_X1 U19215 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n11151), .ZN(n20153) );
  AOI22_X1 U19216 ( .A1(n20156), .A2(n20259), .B1(n20250), .B2(n20154), .ZN(
        n17437) );
  OAI21_X1 U19217 ( .B1(n12984), .B2(n20250), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17432) );
  NOR2_X2 U19218 ( .A1(n20119), .A2(n20174), .ZN(n20157) );
  NAND2_X1 U19219 ( .A1(n20252), .A2(n20157), .ZN(n17436) );
  AOI22_X1 U19220 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n11151), .ZN(n20160) );
  NAND2_X1 U19221 ( .A1(n20150), .A2(n20251), .ZN(n17435) );
  NAND4_X1 U19222 ( .A1(n17438), .A2(n17437), .A3(n17436), .A4(n17435), .ZN(
        P2_U3081) );
  NAND2_X1 U19223 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19201) );
  AOI221_X1 U19224 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19201), .C1(n17440), 
        .C2(n19201), .A(n17439), .ZN(n18627) );
  INV_X1 U19225 ( .A(n17441), .ZN(n18626) );
  OAI221_X1 U19226 ( .B1(n19241), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19241), .C2(n18626), .A(n17483), .ZN(n17442) );
  AOI22_X1 U19227 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18627), .B1(
        n17442), .B2(n21791), .ZN(P3_U2865) );
  AND2_X1 U19228 ( .A1(n21348), .A2(n18050), .ZN(n17472) );
  NOR2_X1 U19229 ( .A1(n19407), .A2(n21344), .ZN(n17446) );
  NAND2_X1 U19230 ( .A1(n21342), .A2(n21336), .ZN(n17469) );
  INV_X1 U19231 ( .A(n17469), .ZN(n17443) );
  NAND2_X1 U19232 ( .A1(n17443), .A2(n17463), .ZN(n17445) );
  AOI21_X1 U19233 ( .B1(n19535), .B2(n21342), .A(n21283), .ZN(n17470) );
  NOR2_X1 U19234 ( .A1(n17470), .A2(n21293), .ZN(n17444) );
  INV_X1 U19235 ( .A(n17451), .ZN(n17447) );
  INV_X1 U19236 ( .A(n19407), .ZN(n17450) );
  NAND2_X1 U19237 ( .A1(n19535), .A2(n21197), .ZN(n17458) );
  NAND2_X1 U19238 ( .A1(n21160), .A2(n17448), .ZN(n21337) );
  NOR4_X2 U19239 ( .A1(n17450), .A2(n17449), .A3(n17458), .A4(n21337), .ZN(
        n21311) );
  NAND2_X1 U19240 ( .A1(n20665), .A2(n19535), .ZN(n21102) );
  NOR2_X1 U19241 ( .A1(n21102), .A2(n21263), .ZN(n17453) );
  NAND2_X1 U19242 ( .A1(n21311), .A2(n21338), .ZN(n17464) );
  NAND2_X1 U19243 ( .A1(n17464), .A2(n17451), .ZN(n21794) );
  AOI21_X2 U19244 ( .B1(n17487), .B2(n21794), .A(n21808), .ZN(n17484) );
  NOR2_X1 U19245 ( .A1(n19535), .A2(n21341), .ZN(n17488) );
  INV_X1 U19246 ( .A(n21283), .ZN(n17454) );
  NAND2_X1 U19247 ( .A1(n21197), .A2(n17454), .ZN(n21105) );
  NAND2_X1 U19248 ( .A1(n17488), .A2(n21105), .ZN(n17468) );
  OR2_X1 U19249 ( .A1(n21338), .A2(n17487), .ZN(n17466) );
  AOI21_X1 U19250 ( .B1(n21197), .B2(n21337), .A(n21336), .ZN(n17455) );
  AOI21_X1 U19251 ( .B1(n21337), .B2(n17466), .A(n17455), .ZN(n17456) );
  XOR2_X1 U19252 ( .A(n17460), .B(n17459), .Z(n17462) );
  NAND2_X1 U19253 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22224) );
  NAND2_X1 U19254 ( .A1(n21795), .A2(n22224), .ZN(n21343) );
  INV_X2 U19255 ( .A(n22225), .ZN(n22179) );
  INV_X1 U19256 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22214) );
  NOR2_X1 U19257 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n22214), .ZN(n22219) );
  NAND2_X1 U19258 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22179), .ZN(n18711) );
  OAI21_X1 U19259 ( .B1(n22179), .B2(n22219), .A(n18708), .ZN(n21339) );
  NOR3_X1 U19260 ( .A1(n17484), .A2(n21343), .A3(n21339), .ZN(n17471) );
  OAI211_X1 U19261 ( .C1(n21283), .C2(n21336), .A(n17463), .B(n18052), .ZN(
        n17465) );
  OAI21_X1 U19262 ( .B1(n17466), .B2(n17465), .A(n17464), .ZN(n17467) );
  OAI211_X1 U19263 ( .C1(n17470), .C2(n17469), .A(n17468), .B(n17467), .ZN(
        n21345) );
  NAND2_X1 U19264 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21830), .ZN(n19204) );
  OAI211_X1 U19265 ( .C1(n21789), .C2(n21807), .A(n19204), .B(n17473), .ZN(
        n21331) );
  NAND2_X1 U19266 ( .A1(n20664), .A2(n21818), .ZN(n21302) );
  INV_X1 U19267 ( .A(n21302), .ZN(n21329) );
  AND2_X1 U19268 ( .A1(n17475), .A2(n18049), .ZN(n21803) );
  NAND3_X1 U19269 ( .A1(n21331), .A2(n21329), .A3(n21803), .ZN(n17476) );
  OAI21_X1 U19270 ( .B1(n21331), .B2(n21798), .A(n17476), .ZN(P3_U3284) );
  INV_X1 U19271 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17478) );
  OAI21_X1 U19272 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n17477), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18692) );
  INV_X1 U19273 ( .A(BS16), .ZN(n17509) );
  NAND2_X1 U19274 ( .A1(n22214), .A2(n17477), .ZN(n22176) );
  AOI21_X1 U19275 ( .B1(n17509), .B2(n22176), .A(n17479), .ZN(n22174) );
  AOI21_X1 U19276 ( .B1(n17478), .B2(n17479), .A(n22174), .ZN(P3_U3280) );
  AND2_X1 U19277 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17479), .ZN(P3_U3028) );
  AND2_X1 U19278 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17479), .ZN(P3_U3027) );
  AND2_X1 U19279 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17479), .ZN(P3_U3026) );
  AND2_X1 U19280 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17479), .ZN(P3_U3025) );
  AND2_X1 U19281 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17479), .ZN(P3_U3024) );
  AND2_X1 U19282 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17479), .ZN(P3_U3023) );
  AND2_X1 U19283 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17479), .ZN(P3_U3022) );
  AND2_X1 U19284 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17479), .ZN(P3_U3021) );
  AND2_X1 U19285 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17479), .ZN(
        P3_U3020) );
  AND2_X1 U19286 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17479), .ZN(
        P3_U3019) );
  AND2_X1 U19287 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17479), .ZN(
        P3_U3018) );
  AND2_X1 U19288 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17479), .ZN(
        P3_U3017) );
  AND2_X1 U19289 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17479), .ZN(
        P3_U3016) );
  AND2_X1 U19290 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17479), .ZN(
        P3_U3015) );
  AND2_X1 U19291 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17479), .ZN(
        P3_U3014) );
  AND2_X1 U19292 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17479), .ZN(
        P3_U3013) );
  AND2_X1 U19293 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17479), .ZN(
        P3_U3012) );
  AND2_X1 U19294 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17479), .ZN(
        P3_U3011) );
  AND2_X1 U19295 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17479), .ZN(
        P3_U3010) );
  AND2_X1 U19296 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17479), .ZN(
        P3_U3009) );
  AND2_X1 U19297 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17479), .ZN(
        P3_U3008) );
  AND2_X1 U19298 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17479), .ZN(
        P3_U3007) );
  AND2_X1 U19299 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17479), .ZN(
        P3_U3006) );
  AND2_X1 U19300 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17479), .ZN(
        P3_U3005) );
  AND2_X1 U19301 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17479), .ZN(
        P3_U3004) );
  AND2_X1 U19302 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17479), .ZN(
        P3_U3003) );
  AND2_X1 U19303 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17479), .ZN(
        P3_U3002) );
  AND2_X1 U19304 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17479), .ZN(
        P3_U3001) );
  AND2_X1 U19305 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17479), .ZN(
        P3_U3000) );
  AND2_X1 U19306 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17479), .ZN(
        P3_U2999) );
  AOI21_X1 U19307 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17482)
         );
  INV_X1 U19308 ( .A(n22224), .ZN(n22226) );
  NAND4_X1 U19309 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n22226), .A4(n21810), .ZN(n21814) );
  INV_X1 U19310 ( .A(n21814), .ZN(n17480) );
  AOI211_X1 U19311 ( .C1(n18528), .C2(n17482), .A(n17481), .B(n17480), .ZN(
        P3_U2998) );
  NOR2_X1 U19312 ( .A1(n21774), .A2(n17483), .ZN(P3_U2867) );
  NOR2_X1 U19313 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21810), .ZN(n18315) );
  INV_X1 U19314 ( .A(n18315), .ZN(n18620) );
  NOR2_X1 U19315 ( .A1(n20664), .A2(n18620), .ZN(n18681) );
  AND2_X1 U19316 ( .A1(n18685), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U19317 ( .A1(n21818), .A2(n21823), .ZN(n18054) );
  INV_X1 U19318 ( .A(n18054), .ZN(n17486) );
  NOR2_X1 U19319 ( .A1(n17486), .A2(n20670), .ZN(n17491) );
  INV_X1 U19320 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n17490) );
  NOR2_X1 U19321 ( .A1(n17488), .A2(n17487), .ZN(n20604) );
  INV_X1 U19322 ( .A(n20604), .ZN(n17489) );
  AOI22_X1 U19323 ( .A1(n17491), .A2(n17490), .B1(n20670), .B2(n17489), .ZN(
        P3_U3298) );
  INV_X1 U19324 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18652) );
  NAND2_X1 U19325 ( .A1(n19535), .A2(n20670), .ZN(n21100) );
  INV_X1 U19326 ( .A(n21100), .ZN(n20685) );
  AOI21_X1 U19327 ( .B1(n17491), .B2(n18652), .A(n20685), .ZN(P3_U3299) );
  NAND2_X1 U19328 ( .A1(n22205), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22204) );
  OAI21_X1 U19329 ( .B1(n17736), .B2(n22204), .A(n22199), .ZN(n22172) );
  INV_X1 U19330 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17508) );
  NAND2_X1 U19331 ( .A1(n22205), .A2(n17492), .ZN(n22196) );
  AOI21_X1 U19332 ( .B1(n17509), .B2(n22196), .A(n11156), .ZN(n22168) );
  AOI21_X1 U19333 ( .B1(n11157), .B2(n17508), .A(n22168), .ZN(P2_U3591) );
  AND2_X1 U19334 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n11157), .ZN(P2_U3208) );
  AND2_X1 U19335 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n11156), .ZN(P2_U3207) );
  AND2_X1 U19336 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n11157), .ZN(P2_U3206) );
  AND2_X1 U19337 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n11156), .ZN(P2_U3205) );
  AND2_X1 U19338 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n11157), .ZN(P2_U3204) );
  AND2_X1 U19339 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n11156), .ZN(P2_U3203) );
  AND2_X1 U19340 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n11157), .ZN(P2_U3202) );
  AND2_X1 U19341 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n11156), .ZN(P2_U3201) );
  AND2_X1 U19342 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n11156), .ZN(
        P2_U3200) );
  AND2_X1 U19343 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n11157), .ZN(
        P2_U3199) );
  AND2_X1 U19344 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n11156), .ZN(
        P2_U3198) );
  AND2_X1 U19345 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n11157), .ZN(
        P2_U3197) );
  AND2_X1 U19346 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n11156), .ZN(
        P2_U3196) );
  AND2_X1 U19347 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n11157), .ZN(
        P2_U3195) );
  AND2_X1 U19348 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n11156), .ZN(
        P2_U3194) );
  AND2_X1 U19349 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n11157), .ZN(
        P2_U3193) );
  AND2_X1 U19350 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n11156), .ZN(
        P2_U3192) );
  AND2_X1 U19351 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n11157), .ZN(
        P2_U3191) );
  AND2_X1 U19352 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n11157), .ZN(
        P2_U3190) );
  AND2_X1 U19353 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n11156), .ZN(
        P2_U3189) );
  AND2_X1 U19354 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n11157), .ZN(
        P2_U3188) );
  AND2_X1 U19355 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n11156), .ZN(
        P2_U3187) );
  AND2_X1 U19356 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n11156), .ZN(
        P2_U3186) );
  AND2_X1 U19357 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n11157), .ZN(
        P2_U3185) );
  AND2_X1 U19358 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n11156), .ZN(
        P2_U3184) );
  AND2_X1 U19359 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n11157), .ZN(
        P2_U3183) );
  AND2_X1 U19360 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n11156), .ZN(
        P2_U3182) );
  AND2_X1 U19361 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n11157), .ZN(
        P2_U3181) );
  AND2_X1 U19362 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n11156), .ZN(
        P2_U3180) );
  AND2_X1 U19363 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n11157), .ZN(
        P2_U3179) );
  NAND2_X1 U19364 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19164), .ZN(n19149) );
  AOI21_X1 U19365 ( .B1(n17494), .B2(n15635), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17495) );
  AOI221_X1 U19366 ( .B1(n19149), .B2(n17495), .C1(n15237), .C2(n17495), .A(
        n19157), .ZN(P2_U3178) );
  OAI221_X1 U19367 ( .B1(n12689), .B2(n17496), .C1(n19156), .C2(n17496), .A(
        n20174), .ZN(n17695) );
  NOR2_X1 U19368 ( .A1(n17497), .A2(n17695), .ZN(P2_U3047) );
  AND2_X1 U19369 ( .A1(n17722), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19370 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17501) );
  NOR4_X1 U19371 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17500) );
  NOR4_X1 U19372 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17499) );
  NOR4_X1 U19373 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17498) );
  NAND4_X1 U19374 ( .A1(n17501), .A2(n17500), .A3(n17499), .A4(n17498), .ZN(
        n17507) );
  NOR4_X1 U19375 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17505) );
  AOI211_X1 U19376 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17504) );
  NOR4_X1 U19377 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17503) );
  NOR4_X1 U19378 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17502) );
  NAND4_X1 U19379 ( .A1(n17505), .A2(n17504), .A3(n17503), .A4(n17502), .ZN(
        n17506) );
  NOR2_X1 U19380 ( .A1(n17507), .A2(n17506), .ZN(n17704) );
  INV_X1 U19381 ( .A(n17704), .ZN(n17703) );
  NOR2_X1 U19382 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17703), .ZN(n17698) );
  INV_X1 U19383 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22171) );
  NAND3_X1 U19384 ( .A1(n12850), .A2(n22171), .A3(n17508), .ZN(n17702) );
  INV_X1 U19385 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U19386 ( .A1(n17698), .A2(n17702), .B1(n17703), .B2(n17749), .ZN(
        P2_U2821) );
  INV_X1 U19387 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U19388 ( .A1(n17698), .A2(n12850), .B1(n17703), .B2(n17747), .ZN(
        P2_U2820) );
  INV_X1 U19389 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20454) );
  INV_X1 U19390 ( .A(n22180), .ZN(n22188) );
  NAND2_X1 U19391 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20527), .ZN(n22593) );
  OAI21_X1 U19392 ( .B1(n22188), .B2(n20527), .A(n22593), .ZN(n17510) );
  INV_X1 U19393 ( .A(n17510), .ZN(n22167) );
  INV_X1 U19394 ( .A(n22167), .ZN(n17511) );
  AOI221_X1 U19395 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n17509), .C1(
        P1_STATE_REG_2__SCAN_IN), .C2(n17509), .A(n17511), .ZN(n22164) );
  AOI21_X1 U19396 ( .B1(n20454), .B2(n17511), .A(n22164), .ZN(P1_U3464) );
  AND2_X1 U19397 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17511), .ZN(P1_U3193) );
  AND2_X1 U19398 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17511), .ZN(P1_U3192) );
  AND2_X1 U19399 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17511), .ZN(P1_U3191) );
  AND2_X1 U19400 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17511), .ZN(P1_U3190) );
  AND2_X1 U19401 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17511), .ZN(P1_U3189) );
  AND2_X1 U19402 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17511), .ZN(P1_U3188) );
  AND2_X1 U19403 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17511), .ZN(P1_U3187) );
  AND2_X1 U19404 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17511), .ZN(P1_U3186) );
  AND2_X1 U19405 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17511), .ZN(
        P1_U3185) );
  AND2_X1 U19406 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17511), .ZN(
        P1_U3184) );
  AND2_X1 U19407 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17511), .ZN(
        P1_U3183) );
  AND2_X1 U19408 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17511), .ZN(
        P1_U3182) );
  AND2_X1 U19409 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17511), .ZN(
        P1_U3181) );
  AND2_X1 U19410 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17510), .ZN(
        P1_U3180) );
  AND2_X1 U19411 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17510), .ZN(
        P1_U3179) );
  AND2_X1 U19412 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17510), .ZN(
        P1_U3178) );
  AND2_X1 U19413 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17510), .ZN(
        P1_U3177) );
  AND2_X1 U19414 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17510), .ZN(
        P1_U3176) );
  AND2_X1 U19415 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17510), .ZN(
        P1_U3175) );
  AND2_X1 U19416 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17510), .ZN(
        P1_U3174) );
  AND2_X1 U19417 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17510), .ZN(
        P1_U3173) );
  AND2_X1 U19418 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17510), .ZN(
        P1_U3172) );
  AND2_X1 U19419 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17510), .ZN(
        P1_U3171) );
  AND2_X1 U19420 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17510), .ZN(
        P1_U3170) );
  AND2_X1 U19421 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17510), .ZN(
        P1_U3169) );
  AND2_X1 U19422 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17510), .ZN(
        P1_U3168) );
  AND2_X1 U19423 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17510), .ZN(
        P1_U3167) );
  AND2_X1 U19424 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17511), .ZN(
        P1_U3166) );
  AND2_X1 U19425 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17511), .ZN(
        P1_U3165) );
  AND2_X1 U19426 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17511), .ZN(
        P1_U3164) );
  NAND2_X1 U19427 ( .A1(n17524), .A2(n17523), .ZN(n17521) );
  NAND2_X1 U19428 ( .A1(n17512), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17513) );
  OR2_X1 U19429 ( .A1(n17514), .A2(n17513), .ZN(n17518) );
  OAI211_X1 U19430 ( .C1(n17518), .C2(n17517), .A(n17516), .B(n17515), .ZN(
        n17520) );
  NAND2_X1 U19431 ( .A1(n17518), .A2(n17517), .ZN(n17519) );
  NAND3_X1 U19432 ( .A1(n17521), .A2(n17520), .A3(n17519), .ZN(n17522) );
  OAI21_X1 U19433 ( .B1(n17524), .B2(n17523), .A(n17522), .ZN(n17528) );
  INV_X1 U19434 ( .A(n17529), .ZN(n17525) );
  NAND2_X1 U19435 ( .A1(n17528), .A2(n17525), .ZN(n17527) );
  NAND2_X1 U19436 ( .A1(n17527), .A2(n17526), .ZN(n17532) );
  INV_X1 U19437 ( .A(n17528), .ZN(n17530) );
  NAND2_X1 U19438 ( .A1(n17530), .A2(n17529), .ZN(n17531) );
  NAND2_X1 U19439 ( .A1(n17532), .A2(n17531), .ZN(n17543) );
  INV_X1 U19440 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17542) );
  INV_X1 U19441 ( .A(n17533), .ZN(n17540) );
  NAND2_X1 U19442 ( .A1(n17534), .A2(n22142), .ZN(n17535) );
  NAND2_X1 U19443 ( .A1(n17536), .A2(n17535), .ZN(n17537) );
  NAND4_X1 U19444 ( .A1(n17540), .A2(n17539), .A3(n17538), .A4(n17537), .ZN(
        n17541) );
  AOI21_X1 U19445 ( .B1(n17543), .B2(n17542), .A(n17541), .ZN(n22163) );
  INV_X1 U19446 ( .A(n22163), .ZN(n17550) );
  NAND3_X1 U19447 ( .A1(n17546), .A2(n17545), .A3(n17544), .ZN(n17547) );
  OAI221_X1 U19448 ( .B1(n17549), .B2(n22181), .C1(n17549), .C2(n17548), .A(
        n17547), .ZN(n17555) );
  AOI221_X1 U19449 ( .B1(n22153), .B2(n15288), .C1(n17550), .C2(n15288), .A(
        n17555), .ZN(n22155) );
  NOR2_X1 U19450 ( .A1(n22155), .A2(n22153), .ZN(n22154) );
  NAND2_X1 U19451 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22157), .ZN(n17551) );
  OAI211_X1 U19452 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21842), .A(n22154), 
        .B(n17551), .ZN(n22159) );
  NAND4_X1 U19453 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n12293), .A4(n21842), .ZN(n17552) );
  AND2_X1 U19454 ( .A1(n17553), .A2(n17552), .ZN(n22151) );
  NAND2_X1 U19455 ( .A1(n22151), .A2(n22152), .ZN(n17554) );
  AOI22_X1 U19456 ( .A1(n15288), .A2(n22159), .B1(n17555), .B2(n17554), .ZN(
        P1_U3162) );
  NOR2_X1 U19457 ( .A1(n17542), .A2(n17556), .ZN(P1_U3032) );
  AND2_X1 U19458 ( .A1(n20371), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19459 ( .A1(n22188), .A2(n20527), .ZN(n17558) );
  INV_X2 U19460 ( .A(n22593), .ZN(n22596) );
  AOI21_X1 U19461 ( .B1(n17558), .B2(n17557), .A(n22596), .ZN(P1_U2802) );
  INV_X1 U19462 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17560) );
  OAI22_X1 U19463 ( .A1(n18717), .A2(n17560), .B1(n15635), .B2(n17559), .ZN(
        P2_U2816) );
  AOI22_X1 U19464 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17670), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19139), .ZN(n17566) );
  OAI22_X1 U19465 ( .A1(n17562), .A2(n17676), .B1(n17608), .B2(n17561), .ZN(
        n17563) );
  AOI21_X1 U19466 ( .B1(n17673), .B2(n17564), .A(n17563), .ZN(n17565) );
  OAI211_X1 U19467 ( .C1(n17681), .C2(n17567), .A(n17566), .B(n17565), .ZN(
        P2_U3009) );
  AOI22_X1 U19468 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19095), .B1(n17640), 
        .B2(n18770), .ZN(n17577) );
  XOR2_X1 U19469 ( .A(n17569), .B(n17568), .Z(n19131) );
  INV_X1 U19470 ( .A(n19132), .ZN(n17575) );
  INV_X1 U19471 ( .A(n17570), .ZN(n17572) );
  NOR2_X1 U19472 ( .A1(n17572), .A2(n17571), .ZN(n17573) );
  XNOR2_X1 U19473 ( .A(n17574), .B(n17573), .ZN(n19137) );
  AOI222_X1 U19474 ( .A1(n19131), .A2(n17664), .B1(n17673), .B2(n17575), .C1(
        n17671), .C2(n19137), .ZN(n17576) );
  OAI211_X1 U19475 ( .C1(n17578), .C2(n17633), .A(n17577), .B(n17576), .ZN(
        P2_U3006) );
  AOI22_X1 U19476 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17670), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19139), .ZN(n17591) );
  NAND2_X1 U19477 ( .A1(n17579), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17581) );
  AOI21_X1 U19478 ( .B1(n13474), .B2(n17581), .A(n17580), .ZN(n19083) );
  INV_X1 U19479 ( .A(n17582), .ZN(n17583) );
  NOR2_X1 U19480 ( .A1(n17584), .A2(n17583), .ZN(n17588) );
  NAND2_X1 U19481 ( .A1(n17586), .A2(n17585), .ZN(n17587) );
  XNOR2_X1 U19482 ( .A(n17588), .B(n17587), .ZN(n19086) );
  OAI22_X1 U19483 ( .A1(n19086), .A2(n17608), .B1(n17657), .B2(n18800), .ZN(
        n17589) );
  AOI21_X1 U19484 ( .B1(n19083), .B2(n17664), .A(n17589), .ZN(n17590) );
  OAI211_X1 U19485 ( .C1(n17681), .C2(n17592), .A(n17591), .B(n17590), .ZN(
        P2_U3004) );
  AOI22_X1 U19486 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19139), .B1(n17640), 
        .B2(n17593), .ZN(n17598) );
  OAI22_X1 U19487 ( .A1(n17676), .A2(n17595), .B1(n17594), .B2(n17608), .ZN(
        n17596) );
  AOI21_X1 U19488 ( .B1(n17673), .B2(n18807), .A(n17596), .ZN(n17597) );
  OAI211_X1 U19489 ( .C1(n18801), .C2(n17633), .A(n17598), .B(n17597), .ZN(
        P2_U3003) );
  AOI22_X1 U19490 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17670), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19139), .ZN(n17603) );
  INV_X1 U19491 ( .A(n18823), .ZN(n17600) );
  AOI222_X1 U19492 ( .A1(n17601), .A2(n17671), .B1(n17673), .B2(n17600), .C1(
        n17664), .C2(n17599), .ZN(n17602) );
  OAI211_X1 U19493 ( .C1(n17681), .C2(n17604), .A(n17603), .B(n17602), .ZN(
        P2_U3002) );
  AOI22_X1 U19494 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19139), .B1(n17640), 
        .B2(n17605), .ZN(n17613) );
  INV_X1 U19495 ( .A(n17606), .ZN(n17609) );
  OAI22_X1 U19496 ( .A1(n17609), .A2(n17608), .B1(n17676), .B2(n17607), .ZN(
        n17610) );
  AOI21_X1 U19497 ( .B1(n17673), .B2(n17611), .A(n17610), .ZN(n17612) );
  OAI211_X1 U19498 ( .C1(n17614), .C2(n17633), .A(n17613), .B(n17612), .ZN(
        P2_U3001) );
  OAI21_X1 U19499 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17616), .A(
        n17615), .ZN(n18831) );
  AOI22_X1 U19500 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17670), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19139), .ZN(n17627) );
  OR2_X1 U19501 ( .A1(n17618), .A2(n17617), .ZN(n17619) );
  NAND2_X1 U19502 ( .A1(n17620), .A2(n17619), .ZN(n19089) );
  NAND2_X1 U19503 ( .A1(n19089), .A2(n17671), .ZN(n17624) );
  OAI21_X1 U19504 ( .B1(n17621), .B2(n13404), .A(n13497), .ZN(n17622) );
  AND2_X1 U19505 ( .A1(n17622), .A2(n19113), .ZN(n19094) );
  NAND2_X1 U19506 ( .A1(n19094), .A2(n17664), .ZN(n17623) );
  OAI211_X1 U19507 ( .C1(n17657), .C2(n19090), .A(n17624), .B(n17623), .ZN(
        n17625) );
  INV_X1 U19508 ( .A(n17625), .ZN(n17626) );
  OAI211_X1 U19509 ( .C1(n17681), .C2(n18831), .A(n17627), .B(n17626), .ZN(
        P2_U3000) );
  AOI21_X1 U19510 ( .B1(n17630), .B2(n17629), .A(n17628), .ZN(n17631) );
  NOR2_X1 U19511 ( .A1(n11225), .A2(n17631), .ZN(n19125) );
  OAI21_X1 U19512 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17632), .A(
        n17639), .ZN(n18858) );
  NOR2_X1 U19513 ( .A1(n17681), .A2(n18858), .ZN(n17635) );
  INV_X1 U19514 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18852) );
  OR2_X1 U19515 ( .A1(n18813), .A2(n13139), .ZN(n19121) );
  OAI21_X1 U19516 ( .B1(n17633), .B2(n18852), .A(n19121), .ZN(n17634) );
  AOI211_X1 U19517 ( .C1(n19125), .C2(n17671), .A(n17635), .B(n17634), .ZN(
        n17638) );
  OAI211_X1 U19518 ( .C1(n17636), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n17664), .B(n19107), .ZN(n17637) );
  OAI211_X1 U19519 ( .C1(n17657), .C2(n19122), .A(n17638), .B(n17637), .ZN(
        P2_U2998) );
  AOI21_X1 U19520 ( .B1(n18864), .B2(n17639), .A(n17652), .ZN(n18872) );
  AOI22_X1 U19521 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17670), .B1(
        n17640), .B2(n18872), .ZN(n17650) );
  NAND2_X1 U19522 ( .A1(n17642), .A2(n17641), .ZN(n17643) );
  XNOR2_X1 U19523 ( .A(n17644), .B(n17643), .ZN(n19110) );
  AOI22_X1 U19524 ( .A1(n19110), .A2(n17671), .B1(n17673), .B2(n19102), .ZN(
        n17649) );
  INV_X1 U19525 ( .A(n19107), .ZN(n17647) );
  INV_X1 U19526 ( .A(n17645), .ZN(n17646) );
  OAI211_X1 U19527 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17647), .A(
        n17646), .B(n17664), .ZN(n17648) );
  NAND2_X1 U19528 ( .A1(P2_REIP_REG_17__SCAN_IN), .A2(n19095), .ZN(n19116) );
  NAND4_X1 U19529 ( .A1(n17650), .A2(n17649), .A3(n17648), .A4(n19116), .ZN(
        P2_U2997) );
  OAI21_X1 U19530 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17652), .A(
        n17651), .ZN(n18888) );
  AOI22_X1 U19531 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17670), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19139), .ZN(n17660) );
  NAND2_X1 U19532 ( .A1(n17653), .A2(n17671), .ZN(n17656) );
  NAND2_X1 U19533 ( .A1(n17654), .A2(n17664), .ZN(n17655) );
  OAI211_X1 U19534 ( .C1(n17657), .C2(n18884), .A(n17656), .B(n17655), .ZN(
        n17658) );
  INV_X1 U19535 ( .A(n17658), .ZN(n17659) );
  OAI211_X1 U19536 ( .C1(n17681), .C2(n18888), .A(n17660), .B(n17659), .ZN(
        P2_U2996) );
  OAI21_X1 U19537 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17662), .A(
        n17661), .ZN(n18935) );
  AOI22_X1 U19538 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17670), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19139), .ZN(n17667) );
  AOI222_X1 U19539 ( .A1(n17665), .A2(n17671), .B1(n17673), .B2(n18932), .C1(
        n17664), .C2(n17663), .ZN(n17666) );
  OAI211_X1 U19540 ( .C1(n17681), .C2(n18935), .A(n17667), .B(n17666), .ZN(
        P2_U2992) );
  OAI21_X1 U19541 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17669), .A(
        n17668), .ZN(n18957) );
  AOI22_X1 U19542 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17670), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19139), .ZN(n17680) );
  NAND2_X1 U19543 ( .A1(n17672), .A2(n17671), .ZN(n17675) );
  NAND2_X1 U19544 ( .A1(n17673), .A2(n18955), .ZN(n17674) );
  OAI211_X1 U19545 ( .C1(n17677), .C2(n17676), .A(n17675), .B(n17674), .ZN(
        n17678) );
  INV_X1 U19546 ( .A(n17678), .ZN(n17679) );
  OAI211_X1 U19547 ( .C1(n17681), .C2(n18957), .A(n17680), .B(n17679), .ZN(
        P2_U2990) );
  INV_X1 U19548 ( .A(n17695), .ZN(n17697) );
  INV_X1 U19549 ( .A(n17682), .ZN(n18720) );
  OAI22_X1 U19550 ( .A1(n19674), .A2(n18720), .B1(n19734), .B2(n17683), .ZN(
        n17684) );
  AOI21_X1 U19551 ( .B1(n19819), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17684), 
        .ZN(n17685) );
  OAI22_X1 U19552 ( .A1(n19819), .A2(n17695), .B1(n17697), .B2(n17685), .ZN(
        P2_U3605) );
  AND2_X1 U19553 ( .A1(n19690), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19667) );
  NAND2_X1 U19554 ( .A1(n17686), .A2(n19667), .ZN(n19703) );
  INV_X1 U19555 ( .A(n19703), .ZN(n19794) );
  OAI21_X1 U19556 ( .B1(n19667), .B2(n19838), .A(n19148), .ZN(n17692) );
  AOI222_X1 U19557 ( .A1(n20059), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19788), 
        .B2(n19794), .C1(n17692), .C2(n20060), .ZN(n17687) );
  AOI22_X1 U19558 ( .A1(n17697), .A2(n19787), .B1(n17687), .B2(n17695), .ZN(
        P2_U3603) );
  AND2_X1 U19559 ( .A1(n19788), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17693) );
  OR2_X1 U19560 ( .A1(n19690), .A2(n17693), .ZN(n17688) );
  AOI22_X1 U19561 ( .A1(n17692), .A2(n17688), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20111), .ZN(n17689) );
  AOI22_X1 U19562 ( .A1(n17697), .A2(n19807), .B1(n17689), .B2(n17695), .ZN(
        P2_U3604) );
  OAI21_X1 U19563 ( .B1(n19766), .B2(n17690), .A(n19720), .ZN(n17694) );
  AOI222_X1 U19564 ( .A1(n20009), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n17694), 
        .B2(n17693), .C1(n17692), .C2(n17691), .ZN(n17696) );
  AOI22_X1 U19565 ( .A1(n17697), .A2(n19786), .B1(n17696), .B2(n17695), .ZN(
        P2_U3602) );
  NAND2_X1 U19566 ( .A1(n17698), .A2(n22171), .ZN(n17701) );
  OAI21_X1 U19567 ( .B1(n17738), .B2(n12850), .A(n17704), .ZN(n17699) );
  OAI21_X1 U19568 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17704), .A(n17699), 
        .ZN(n17700) );
  OAI221_X1 U19569 ( .B1(n17701), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17701), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17700), .ZN(P2_U2822) );
  INV_X1 U19570 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17752) );
  OAI221_X1 U19571 ( .B1(n17704), .B2(n17752), .C1(n17703), .C2(n17702), .A(
        n17701), .ZN(P2_U2823) );
  INV_X1 U19572 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n17705) );
  AOI22_X1 U19573 ( .A1(n22203), .A2(n17706), .B1(n17705), .B2(n17750), .ZN(
        P2_U3611) );
  INV_X1 U19574 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17707) );
  AOI22_X1 U19575 ( .A1(n22203), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17707), 
        .B2(n17750), .ZN(P2_U3608) );
  INV_X1 U19576 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n17708) );
  OAI21_X1 U19577 ( .B1(n17736), .B2(n17708), .A(n11156), .ZN(P2_U2815) );
  AOI22_X1 U19578 ( .A1(n17733), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17710) );
  OAI21_X1 U19579 ( .B1(n20161), .B2(n17735), .A(n17710), .ZN(P2_U2951) );
  INV_X1 U19580 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17712) );
  AOI22_X1 U19581 ( .A1(n17733), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17711) );
  OAI21_X1 U19582 ( .B1(n17712), .B2(n17735), .A(n17711), .ZN(P2_U2950) );
  INV_X1 U19583 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17714) );
  AOI22_X1 U19584 ( .A1(n17733), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17713) );
  OAI21_X1 U19585 ( .B1(n17714), .B2(n17735), .A(n17713), .ZN(P2_U2949) );
  INV_X1 U19586 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17716) );
  AOI22_X1 U19587 ( .A1(n17725), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17715) );
  OAI21_X1 U19588 ( .B1(n17716), .B2(n17735), .A(n17715), .ZN(P2_U2948) );
  INV_X1 U19589 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U19590 ( .A1(n17733), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17717) );
  OAI21_X1 U19591 ( .B1(n17718), .B2(n17735), .A(n17717), .ZN(P2_U2947) );
  INV_X1 U19592 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U19593 ( .A1(n17725), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17719) );
  OAI21_X1 U19594 ( .B1(n19903), .B2(n17735), .A(n17719), .ZN(P2_U2946) );
  INV_X1 U19595 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U19596 ( .A1(n17725), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17720) );
  OAI21_X1 U19597 ( .B1(n19862), .B2(n17735), .A(n17720), .ZN(P2_U2945) );
  INV_X1 U19598 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19599 ( .A1(n17725), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17721) );
  OAI21_X1 U19600 ( .B1(n19662), .B2(n17735), .A(n17721), .ZN(P2_U2944) );
  INV_X1 U19601 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19659) );
  AOI22_X1 U19602 ( .A1(n17725), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17722), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17723) );
  OAI21_X1 U19603 ( .B1(n19659), .B2(n17735), .A(n17723), .ZN(P2_U2943) );
  INV_X1 U19604 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U19605 ( .A1(n17733), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17724) );
  OAI21_X1 U19606 ( .B1(n19655), .B2(n17735), .A(n17724), .ZN(P2_U2942) );
  INV_X1 U19607 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19652) );
  AOI22_X1 U19608 ( .A1(n17725), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17726) );
  OAI21_X1 U19609 ( .B1(n19652), .B2(n17735), .A(n17726), .ZN(P2_U2941) );
  INV_X1 U19610 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19648) );
  AOI22_X1 U19611 ( .A1(n17733), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17727) );
  OAI21_X1 U19612 ( .B1(n19648), .B2(n17735), .A(n17727), .ZN(P2_U2940) );
  AOI22_X1 U19613 ( .A1(n17733), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17728) );
  OAI21_X1 U19614 ( .B1(n17729), .B2(n17735), .A(n17728), .ZN(P2_U2939) );
  INV_X1 U19615 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U19616 ( .A1(n17733), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17730) );
  OAI21_X1 U19617 ( .B1(n19641), .B2(n17735), .A(n17730), .ZN(P2_U2938) );
  INV_X1 U19618 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U19619 ( .A1(n17733), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17731) );
  OAI21_X1 U19620 ( .B1(n19638), .B2(n17735), .A(n17731), .ZN(P2_U2937) );
  AOI22_X1 U19621 ( .A1(n17733), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17732), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17734) );
  OAI21_X1 U19622 ( .B1(n19635), .B2(n17735), .A(n17734), .ZN(P2_U2936) );
  AOI21_X1 U19623 ( .B1(n22205), .B2(n17736), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17737) );
  AOI22_X1 U19624 ( .A1(n22203), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n17737), 
        .B2(n17750), .ZN(P2_U2817) );
  OAI222_X1 U19625 ( .A1(n17745), .A2(n12868), .B1(n20293), .B2(n22203), .C1(
        n17738), .C2(n17744), .ZN(P2_U3212) );
  INV_X1 U19626 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20295) );
  OAI222_X1 U19627 ( .A1(n17745), .A2(n15481), .B1(n20295), .B2(n22203), .C1(
        n12868), .C2(n17744), .ZN(P2_U3213) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20297) );
  OAI222_X1 U19629 ( .A1(n17745), .A2(n13221), .B1(n20297), .B2(n22203), .C1(
        n15481), .C2(n17744), .ZN(P2_U3214) );
  INV_X1 U19630 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20299) );
  OAI222_X1 U19631 ( .A1(n17745), .A2(n13230), .B1(n20299), .B2(n22203), .C1(
        n13221), .C2(n17744), .ZN(P2_U3215) );
  INV_X1 U19632 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20301) );
  OAI222_X1 U19633 ( .A1(n17745), .A2(n13105), .B1(n20301), .B2(n22203), .C1(
        n13230), .C2(n17744), .ZN(P2_U3216) );
  INV_X1 U19634 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20303) );
  OAI222_X1 U19635 ( .A1(n17745), .A2(n17160), .B1(n20303), .B2(n22203), .C1(
        n13105), .C2(n17744), .ZN(P2_U3217) );
  INV_X1 U19636 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17739) );
  INV_X1 U19637 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20305) );
  OAI222_X1 U19638 ( .A1(n17745), .A2(n17739), .B1(n20305), .B2(n22203), .C1(
        n17160), .C2(n17744), .ZN(P2_U3218) );
  INV_X1 U19639 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20307) );
  OAI222_X1 U19640 ( .A1(n17745), .A2(n17147), .B1(n20307), .B2(n22203), .C1(
        n17739), .C2(n17744), .ZN(P2_U3219) );
  INV_X1 U19641 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20309) );
  OAI222_X1 U19642 ( .A1(n17744), .A2(n17147), .B1(n20309), .B2(n22203), .C1(
        n13264), .C2(n17745), .ZN(P2_U3220) );
  INV_X1 U19643 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20311) );
  OAI222_X1 U19644 ( .A1(n17744), .A2(n13264), .B1(n20311), .B2(n22203), .C1(
        n13123), .C2(n17745), .ZN(P2_U3221) );
  INV_X1 U19645 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20313) );
  OAI222_X1 U19646 ( .A1(n17744), .A2(n13123), .B1(n20313), .B2(n22203), .C1(
        n13301), .C2(n17745), .ZN(P2_U3222) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20315) );
  OAI222_X1 U19648 ( .A1(n17744), .A2(n13301), .B1(n20315), .B2(n22203), .C1(
        n13131), .C2(n17745), .ZN(P2_U3223) );
  INV_X1 U19649 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20317) );
  OAI222_X1 U19650 ( .A1(n17744), .A2(n13131), .B1(n20317), .B2(n22203), .C1(
        n13320), .C2(n17745), .ZN(P2_U3224) );
  INV_X1 U19651 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20319) );
  OAI222_X1 U19652 ( .A1(n17744), .A2(n13320), .B1(n20319), .B2(n22203), .C1(
        n18839), .C2(n17745), .ZN(P2_U3225) );
  INV_X1 U19653 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20321) );
  OAI222_X1 U19654 ( .A1(n17744), .A2(n18839), .B1(n20321), .B2(n22203), .C1(
        n13139), .C2(n17745), .ZN(P2_U3226) );
  INV_X1 U19655 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20323) );
  OAI222_X1 U19656 ( .A1(n17744), .A2(n13139), .B1(n20323), .B2(n22203), .C1(
        n13142), .C2(n17745), .ZN(P2_U3227) );
  INV_X1 U19657 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20325) );
  OAI222_X1 U19658 ( .A1(n17744), .A2(n13142), .B1(n20325), .B2(n22203), .C1(
        n13351), .C2(n17745), .ZN(P2_U3228) );
  INV_X1 U19659 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20327) );
  OAI222_X1 U19660 ( .A1(n17745), .A2(n18894), .B1(n20327), .B2(n22203), .C1(
        n13351), .C2(n17744), .ZN(P2_U3229) );
  INV_X1 U19661 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20329) );
  OAI222_X1 U19662 ( .A1(n17744), .A2(n18894), .B1(n20329), .B2(n22203), .C1(
        n18905), .C2(n17745), .ZN(P2_U3230) );
  INV_X1 U19663 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20331) );
  OAI222_X1 U19664 ( .A1(n17745), .A2(n18917), .B1(n20331), .B2(n22203), .C1(
        n18905), .C2(n17744), .ZN(P2_U3231) );
  INV_X1 U19665 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20333) );
  OAI222_X1 U19666 ( .A1(n17745), .A2(n13360), .B1(n20333), .B2(n22203), .C1(
        n18917), .C2(n17744), .ZN(P2_U3232) );
  INV_X1 U19667 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20335) );
  OAI222_X1 U19668 ( .A1(n17745), .A2(n13161), .B1(n20335), .B2(n22203), .C1(
        n13360), .C2(n17744), .ZN(P2_U3233) );
  INV_X1 U19669 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20337) );
  OAI222_X1 U19670 ( .A1(n17745), .A2(n17217), .B1(n20337), .B2(n22203), .C1(
        n13161), .C2(n17744), .ZN(P2_U3234) );
  INV_X1 U19671 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20339) );
  OAI222_X1 U19672 ( .A1(n17745), .A2(n17740), .B1(n20339), .B2(n22203), .C1(
        n17217), .C2(n17744), .ZN(P2_U3235) );
  INV_X1 U19673 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20342) );
  OAI222_X1 U19674 ( .A1(n17744), .A2(n17740), .B1(n20342), .B2(n22203), .C1(
        n17741), .C2(n17745), .ZN(P2_U3236) );
  INV_X1 U19675 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20344) );
  OAI222_X1 U19676 ( .A1(n17745), .A2(n17742), .B1(n20344), .B2(n22203), .C1(
        n17741), .C2(n17744), .ZN(P2_U3237) );
  INV_X1 U19677 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20346) );
  OAI222_X1 U19678 ( .A1(n17744), .A2(n17742), .B1(n20346), .B2(n22203), .C1(
        n17058), .C2(n17745), .ZN(P2_U3238) );
  INV_X1 U19679 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20348) );
  OAI222_X1 U19680 ( .A1(n17744), .A2(n17058), .B1(n20348), .B2(n22203), .C1(
        n17743), .C2(n17745), .ZN(P2_U3239) );
  INV_X1 U19681 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20350) );
  OAI222_X1 U19682 ( .A1(n17744), .A2(n17743), .B1(n20350), .B2(n22203), .C1(
        n19023), .C2(n17745), .ZN(P2_U3240) );
  INV_X1 U19683 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20353) );
  OAI222_X1 U19684 ( .A1(n17745), .A2(n19042), .B1(n20353), .B2(n22203), .C1(
        n19023), .C2(n17744), .ZN(P2_U3241) );
  INV_X1 U19685 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U19686 ( .A1(n22203), .A2(n17747), .B1(n17746), .B2(n17750), .ZN(
        P2_U3588) );
  INV_X1 U19687 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n17748) );
  AOI22_X1 U19688 ( .A1(n22203), .A2(n17749), .B1(n17748), .B2(n17750), .ZN(
        P2_U3587) );
  MUX2_X1 U19689 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n22203), .Z(P2_U3586) );
  INV_X1 U19690 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U19691 ( .A1(n22203), .A2(n17752), .B1(n17751), .B2(n17750), .ZN(
        P2_U3585) );
  NAND2_X1 U19692 ( .A1(n18039), .A2(n17753), .ZN(n17780) );
  NOR2_X1 U19693 ( .A1(n21197), .A2(n17780), .ZN(n17778) );
  NOR3_X1 U19694 ( .A1(n20705), .A2(n17754), .A3(n18035), .ZN(n17759) );
  AOI21_X1 U19695 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18034), .A(n17759), .ZN(
        n17755) );
  OAI22_X1 U19696 ( .A1(n17778), .A2(n17755), .B1(n18115), .B2(n18034), .ZN(
        P3_U2699) );
  AOI21_X1 U19697 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18034), .A(n17756), .ZN(
        n17758) );
  INV_X1 U19698 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17757) );
  OAI22_X1 U19699 ( .A1(n17759), .A2(n17758), .B1(n17757), .B2(n18034), .ZN(
        P3_U2700) );
  AOI22_X1 U19700 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17770) );
  AOI22_X1 U19701 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U19702 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17760) );
  OAI21_X1 U19703 ( .B1(n11192), .B2(n17761), .A(n17760), .ZN(n17767) );
  AOI22_X1 U19704 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U19705 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17764) );
  AOI22_X1 U19706 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17763) );
  AOI22_X1 U19707 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17762) );
  NAND4_X1 U19708 ( .A1(n17765), .A2(n17764), .A3(n17763), .A4(n17762), .ZN(
        n17766) );
  AOI211_X1 U19709 ( .C1(n11175), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17767), .B(n17766), .ZN(n17768) );
  NAND3_X1 U19710 ( .A1(n17770), .A2(n17769), .A3(n17768), .ZN(n21264) );
  INV_X1 U19711 ( .A(n21264), .ZN(n17773) );
  AND2_X1 U19712 ( .A1(n18039), .A2(n17774), .ZN(n17771) );
  NAND3_X1 U19713 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18039), .A3(n17774), .ZN(
        n17876) );
  OAI21_X1 U19714 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17771), .A(n17876), .ZN(
        n17772) );
  AOI22_X1 U19715 ( .A1(n18037), .A2(n17773), .B1(n17772), .B2(n18034), .ZN(
        P3_U2695) );
  INV_X1 U19716 ( .A(n18039), .ZN(n18027) );
  AOI211_X1 U19717 ( .C1(n20753), .C2(n17775), .A(n17774), .B(n18035), .ZN(
        n17776) );
  AOI21_X1 U19718 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18027), .A(n17776), .ZN(
        n17777) );
  OAI21_X1 U19719 ( .B1(n18060), .B2(n18034), .A(n17777), .ZN(P3_U2696) );
  NAND2_X1 U19720 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17778), .ZN(n17781) );
  INV_X1 U19721 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18131) );
  NAND3_X1 U19722 ( .A1(n17781), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n18034), .ZN(
        n17779) );
  OAI221_X1 U19723 ( .B1(n17781), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n18034), 
        .C2(n18131), .A(n17779), .ZN(P3_U2697) );
  INV_X1 U19724 ( .A(n17780), .ZN(n17782) );
  OAI211_X1 U19725 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17782), .A(n17781), .B(
        n18034), .ZN(n17783) );
  OAI21_X1 U19726 ( .B1(n18034), .B2(n17812), .A(n17783), .ZN(P3_U2698) );
  AOI22_X1 U19727 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U19728 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17786) );
  AOI22_X1 U19729 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17785) );
  AOI22_X1 U19730 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18082), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17784) );
  NAND4_X1 U19731 ( .A1(n17787), .A2(n17786), .A3(n17785), .A4(n17784), .ZN(
        n17793) );
  AOI22_X1 U19732 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17791) );
  AOI22_X1 U19733 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17790) );
  AOI22_X1 U19734 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17789) );
  AOI22_X1 U19735 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17788) );
  NAND4_X1 U19736 ( .A1(n17791), .A2(n17790), .A3(n17789), .A4(n17788), .ZN(
        n17792) );
  NOR2_X1 U19737 ( .A1(n17793), .A2(n17792), .ZN(n21247) );
  INV_X1 U19738 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20872) );
  INV_X1 U19739 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20838) );
  INV_X1 U19740 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20820) );
  NOR2_X1 U19741 ( .A1(n20780), .A2(n17876), .ZN(n17889) );
  NAND2_X1 U19742 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17889), .ZN(n17873) );
  NOR2_X1 U19743 ( .A1(n20820), .A2(n17873), .ZN(n17862) );
  NAND2_X1 U19744 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17862), .ZN(n17848) );
  NOR2_X1 U19745 ( .A1(n20838), .A2(n17848), .ZN(n17824) );
  NAND2_X1 U19746 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17824), .ZN(n17796) );
  NOR2_X1 U19747 ( .A1(n20872), .A2(n17796), .ZN(n17809) );
  NAND2_X1 U19748 ( .A1(n17809), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17794) );
  OAI211_X1 U19749 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17809), .A(n18034), .B(
        n17794), .ZN(n17795) );
  OAI21_X1 U19750 ( .B1(n21247), .B2(n18034), .A(n17795), .ZN(P3_U2687) );
  NAND2_X1 U19751 ( .A1(n20872), .A2(n17796), .ZN(n17797) );
  NAND2_X1 U19752 ( .A1(n17797), .A2(n18034), .ZN(n17808) );
  AOI22_X1 U19753 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14455), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17801) );
  AOI22_X1 U19754 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17800) );
  AOI22_X1 U19755 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U19756 ( .A1(n18105), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17798) );
  NAND4_X1 U19757 ( .A1(n17801), .A2(n17800), .A3(n17799), .A4(n17798), .ZN(
        n17807) );
  AOI22_X1 U19758 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U19759 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17804) );
  AOI22_X1 U19760 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17803) );
  AOI22_X1 U19761 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17802) );
  NAND4_X1 U19762 ( .A1(n17805), .A2(n17804), .A3(n17803), .A4(n17802), .ZN(
        n17806) );
  NOR2_X1 U19763 ( .A1(n17807), .A2(n17806), .ZN(n21261) );
  OAI22_X1 U19764 ( .A1(n17809), .A2(n17808), .B1(n21261), .B2(n18034), .ZN(
        P3_U2688) );
  AOI21_X1 U19765 ( .B1(n20838), .B2(n17848), .A(n18037), .ZN(n17810) );
  INV_X1 U19766 ( .A(n17810), .ZN(n17823) );
  AOI22_X1 U19767 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U19768 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U19769 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17811) );
  OAI21_X1 U19770 ( .B1(n11192), .B2(n17812), .A(n17811), .ZN(n17818) );
  AOI22_X1 U19771 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17816) );
  AOI22_X1 U19772 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17815) );
  AOI22_X1 U19773 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18105), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17814) );
  AOI22_X1 U19774 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17813) );
  NAND4_X1 U19775 ( .A1(n17816), .A2(n17815), .A3(n17814), .A4(n17813), .ZN(
        n17817) );
  AOI211_X1 U19776 ( .C1(n18128), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n17818), .B(n17817), .ZN(n17819) );
  NAND3_X1 U19777 ( .A1(n17821), .A2(n17820), .A3(n17819), .ZN(n21106) );
  INV_X1 U19778 ( .A(n21106), .ZN(n17822) );
  OAI22_X1 U19779 ( .A1(n17824), .A2(n17823), .B1(n17822), .B2(n18034), .ZN(
        P3_U2690) );
  NAND2_X1 U19780 ( .A1(n21263), .A2(n17824), .ZN(n17837) );
  AOI22_X1 U19781 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U19782 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U19783 ( .A1(n18116), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17825) );
  OAI21_X1 U19784 ( .B1(n11192), .B2(n18131), .A(n17825), .ZN(n17831) );
  AOI22_X1 U19785 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17829) );
  AOI22_X1 U19786 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17828) );
  AOI22_X1 U19787 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U19788 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17826) );
  NAND4_X1 U19789 ( .A1(n17829), .A2(n17828), .A3(n17827), .A4(n17826), .ZN(
        n17830) );
  AOI211_X1 U19790 ( .C1(n11175), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17831), .B(n17830), .ZN(n17832) );
  NAND3_X1 U19791 ( .A1(n17834), .A2(n17833), .A3(n17832), .ZN(n21250) );
  INV_X1 U19792 ( .A(n21250), .ZN(n17836) );
  NAND3_X1 U19793 ( .A1(n17837), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n18034), 
        .ZN(n17835) );
  OAI221_X1 U19794 ( .B1(n17837), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n18034), 
        .C2(n17836), .A(n17835), .ZN(P3_U2689) );
  AOI22_X1 U19795 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U19796 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17840) );
  AOI22_X1 U19797 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U19798 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17838) );
  NAND4_X1 U19799 ( .A1(n17841), .A2(n17840), .A3(n17839), .A4(n17838), .ZN(
        n17847) );
  AOI22_X1 U19800 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17845) );
  AOI22_X1 U19801 ( .A1(n18108), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17844) );
  AOI22_X1 U19802 ( .A1(n18095), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17843) );
  AOI22_X1 U19803 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17842) );
  NAND4_X1 U19804 ( .A1(n17845), .A2(n17844), .A3(n17843), .A4(n17842), .ZN(
        n17846) );
  NOR2_X1 U19805 ( .A1(n17847), .A2(n17846), .ZN(n21110) );
  OAI21_X1 U19806 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17862), .A(n17848), .ZN(
        n17849) );
  AOI22_X1 U19807 ( .A1(n18037), .A2(n21110), .B1(n17849), .B2(n18034), .ZN(
        P3_U2691) );
  INV_X1 U19808 ( .A(n17873), .ZN(n17850) );
  OAI21_X1 U19809 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17850), .A(n18034), .ZN(
        n17861) );
  AOI22_X1 U19810 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17854) );
  AOI22_X1 U19811 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U19812 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17852) );
  AOI22_X1 U19813 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17851) );
  NAND4_X1 U19814 ( .A1(n17854), .A2(n17853), .A3(n17852), .A4(n17851), .ZN(
        n17860) );
  AOI22_X1 U19815 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17858) );
  AOI22_X1 U19816 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17857) );
  AOI22_X1 U19817 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17856) );
  AOI22_X1 U19818 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17855) );
  NAND4_X1 U19819 ( .A1(n17858), .A2(n17857), .A3(n17856), .A4(n17855), .ZN(
        n17859) );
  NOR2_X1 U19820 ( .A1(n17860), .A2(n17859), .ZN(n21114) );
  OAI22_X1 U19821 ( .A1(n17862), .A2(n17861), .B1(n21114), .B2(n18034), .ZN(
        P3_U2692) );
  AOI22_X1 U19822 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17872) );
  AOI22_X1 U19823 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14455), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17871) );
  AOI22_X1 U19824 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17863) );
  OAI21_X1 U19825 ( .B1(n11192), .B2(n18094), .A(n17863), .ZN(n17869) );
  AOI22_X1 U19826 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17867) );
  AOI22_X1 U19827 ( .A1(n18071), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17866) );
  AOI22_X1 U19828 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17865) );
  AOI22_X1 U19829 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17864) );
  NAND4_X1 U19830 ( .A1(n17867), .A2(n17866), .A3(n17865), .A4(n17864), .ZN(
        n17868) );
  AOI211_X1 U19831 ( .C1(n18129), .C2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n17869), .B(n17868), .ZN(n17870) );
  NAND3_X1 U19832 ( .A1(n17872), .A2(n17871), .A3(n17870), .ZN(n21118) );
  INV_X1 U19833 ( .A(n21118), .ZN(n17875) );
  OAI21_X1 U19834 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17889), .A(n17873), .ZN(
        n17874) );
  AOI22_X1 U19835 ( .A1(n18037), .A2(n17875), .B1(n17874), .B2(n18034), .ZN(
        P3_U2693) );
  AOI21_X1 U19836 ( .B1(n20780), .B2(n17876), .A(n18037), .ZN(n17877) );
  INV_X1 U19837 ( .A(n17877), .ZN(n17888) );
  AOI22_X1 U19838 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n18116), .ZN(n17881) );
  AOI22_X1 U19839 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18127), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n18108), .ZN(n17880) );
  AOI22_X1 U19840 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n18105), .ZN(n17879) );
  AOI22_X1 U19841 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18148), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18082), .ZN(n17878) );
  NAND4_X1 U19842 ( .A1(n17881), .A2(n17880), .A3(n17879), .A4(n17878), .ZN(
        n17887) );
  AOI22_X1 U19843 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18134), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17885) );
  AOI22_X1 U19844 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11176), .ZN(n17884) );
  AOI22_X1 U19845 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18132), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18155), .ZN(n17883) );
  AOI22_X1 U19846 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18156), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17882) );
  NAND4_X1 U19847 ( .A1(n17885), .A2(n17884), .A3(n17883), .A4(n17882), .ZN(
        n17886) );
  NOR2_X1 U19848 ( .A1(n17887), .A2(n17886), .ZN(n21124) );
  OAI22_X1 U19849 ( .A1(n17889), .A2(n17888), .B1(n21124), .B2(n18034), .ZN(
        P3_U2694) );
  INV_X1 U19850 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21073) );
  INV_X1 U19851 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n21015) );
  INV_X1 U19852 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21006) );
  NOR4_X1 U19853 ( .A1(n21038), .A2(n21030), .A3(n21015), .A4(n21006), .ZN(
        n17943) );
  INV_X1 U19854 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21052) );
  INV_X1 U19855 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20956) );
  NOR4_X1 U19856 ( .A1(n21052), .A2(n20988), .A3(n20956), .A4(n17932), .ZN(
        n17890) );
  NAND4_X1 U19857 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17943), .A4(n17890), .ZN(n17893) );
  NOR2_X1 U19858 ( .A1(n21073), .A2(n17893), .ZN(n17921) );
  NAND2_X1 U19859 ( .A1(n18034), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17892) );
  NAND2_X1 U19860 ( .A1(n17921), .A2(n21263), .ZN(n17891) );
  OAI22_X1 U19861 ( .A1(n17921), .A2(n17892), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17891), .ZN(P3_U2672) );
  NAND2_X1 U19862 ( .A1(n21073), .A2(n17893), .ZN(n17894) );
  NAND2_X1 U19863 ( .A1(n17894), .A2(n18034), .ZN(n17920) );
  AOI22_X1 U19864 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17899) );
  AOI22_X1 U19865 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U19866 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U19867 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17896) );
  NAND4_X1 U19868 ( .A1(n17899), .A2(n17898), .A3(n17897), .A4(n17896), .ZN(
        n17907) );
  AOI22_X1 U19869 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17905) );
  AOI22_X1 U19870 ( .A1(n18071), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17900), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17904) );
  AOI22_X1 U19871 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18105), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17903) );
  AOI22_X1 U19872 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17902) );
  NAND4_X1 U19873 ( .A1(n17905), .A2(n17904), .A3(n17903), .A4(n17902), .ZN(
        n17906) );
  NOR2_X1 U19874 ( .A1(n17907), .A2(n17906), .ZN(n17919) );
  AOI22_X1 U19875 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17918) );
  AOI22_X1 U19876 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17917) );
  AOI22_X1 U19877 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17908) );
  OAI21_X1 U19878 ( .B1(n17909), .B2(n18131), .A(n17908), .ZN(n17915) );
  AOI22_X1 U19879 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U19880 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17912) );
  AOI22_X1 U19881 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17911) );
  AOI22_X1 U19882 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17910) );
  NAND4_X1 U19883 ( .A1(n17913), .A2(n17912), .A3(n17911), .A4(n17910), .ZN(
        n17914) );
  AOI211_X1 U19884 ( .C1(n18129), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17915), .B(n17914), .ZN(n17916) );
  NAND3_X1 U19885 ( .A1(n17918), .A2(n17917), .A3(n17916), .ZN(n17940) );
  NAND2_X1 U19886 ( .A1(n17941), .A2(n17940), .ZN(n17939) );
  XNOR2_X1 U19887 ( .A(n17919), .B(n17939), .ZN(n21214) );
  OAI22_X1 U19888 ( .A1(n17921), .A2(n17920), .B1(n21214), .B2(n18034), .ZN(
        P3_U2673) );
  AOI22_X1 U19889 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17925) );
  AOI22_X1 U19890 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U19891 ( .A1(n18116), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17923) );
  AOI22_X1 U19892 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17922) );
  NAND4_X1 U19893 ( .A1(n17925), .A2(n17924), .A3(n17923), .A4(n17922), .ZN(
        n17931) );
  AOI22_X1 U19894 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17929) );
  AOI22_X1 U19895 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18126), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17928) );
  AOI22_X1 U19896 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17927) );
  AOI22_X1 U19897 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17926) );
  NAND4_X1 U19898 ( .A1(n17929), .A2(n17928), .A3(n17927), .A4(n17926), .ZN(
        n17930) );
  NOR2_X1 U19899 ( .A1(n17931), .A2(n17930), .ZN(n21163) );
  AND2_X1 U19900 ( .A1(n18034), .A2(n17932), .ZN(n17988) );
  AOI22_X1 U19901 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17988), .B1(n17933), 
        .B2(n20956), .ZN(n17934) );
  OAI21_X1 U19902 ( .B1(n21163), .B2(n18034), .A(n17934), .ZN(P3_U2682) );
  OAI21_X1 U19903 ( .B1(n17945), .B2(n17936), .A(n17935), .ZN(n21229) );
  NAND3_X1 U19904 ( .A1(n17938), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18034), 
        .ZN(n17937) );
  OAI221_X1 U19905 ( .B1(n17938), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18034), 
        .C2(n21229), .A(n17937), .ZN(P3_U2676) );
  OAI21_X1 U19906 ( .B1(n17941), .B2(n17940), .A(n17939), .ZN(n21218) );
  OAI222_X1 U19907 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17958), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n17943), .C1(n21052), .C2(n17942), .ZN(
        n17944) );
  OAI21_X1 U19908 ( .B1(n21218), .B2(n18034), .A(n17944), .ZN(P3_U2674) );
  NAND2_X1 U19909 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17958), .ZN(n17951) );
  AOI21_X1 U19910 ( .B1(n17946), .B2(n17949), .A(n17945), .ZN(n21202) );
  NAND2_X1 U19911 ( .A1(n21202), .A2(n18037), .ZN(n17947) );
  OAI221_X1 U19912 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17951), .C1(n21015), 
        .C2(n17948), .A(n17947), .ZN(P3_U2677) );
  OAI21_X1 U19913 ( .B1(n17954), .B2(n17950), .A(n17949), .ZN(n21201) );
  OAI211_X1 U19914 ( .C1(n17958), .C2(P3_EBX_REG_25__SCAN_IN), .A(n18034), .B(
        n17951), .ZN(n17952) );
  OAI21_X1 U19915 ( .B1(n18034), .B2(n21201), .A(n17952), .ZN(P3_U2678) );
  INV_X1 U19916 ( .A(n17953), .ZN(n17964) );
  AOI21_X1 U19917 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18034), .A(n17964), .ZN(
        n17957) );
  AOI21_X1 U19918 ( .B1(n17955), .B2(n17960), .A(n17954), .ZN(n21230) );
  INV_X1 U19919 ( .A(n21230), .ZN(n17956) );
  OAI22_X1 U19920 ( .A1(n17958), .A2(n17957), .B1(n17956), .B2(n18034), .ZN(
        P3_U2679) );
  AOI21_X1 U19921 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18034), .A(n17959), .ZN(
        n17963) );
  OAI21_X1 U19922 ( .B1(n17962), .B2(n17961), .A(n17960), .ZN(n21241) );
  OAI22_X1 U19923 ( .A1(n17964), .A2(n17963), .B1(n21241), .B2(n18034), .ZN(
        P3_U2680) );
  AOI22_X1 U19924 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14388), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U19925 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17973) );
  AOI22_X1 U19926 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17965) );
  OAI21_X1 U19927 ( .B1(n11218), .B2(n18131), .A(n17965), .ZN(n17971) );
  AOI22_X1 U19928 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U19929 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17968) );
  AOI22_X1 U19930 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17967) );
  AOI22_X1 U19931 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17966) );
  NAND4_X1 U19932 ( .A1(n17969), .A2(n17968), .A3(n17967), .A4(n17966), .ZN(
        n17970) );
  AOI211_X1 U19933 ( .C1(n18067), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17971), .B(n17970), .ZN(n17972) );
  NAND3_X1 U19934 ( .A1(n17974), .A2(n17973), .A3(n17972), .ZN(n21173) );
  INV_X1 U19935 ( .A(n21173), .ZN(n17976) );
  NAND3_X1 U19936 ( .A1(n17977), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18034), 
        .ZN(n17975) );
  OAI221_X1 U19937 ( .B1(n17977), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18034), 
        .C2(n17976), .A(n17975), .ZN(P3_U2681) );
  AOI22_X1 U19938 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17981) );
  AOI22_X1 U19939 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18156), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17980) );
  AOI22_X1 U19940 ( .A1(n18071), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17979) );
  AOI22_X1 U19941 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17978) );
  NAND4_X1 U19942 ( .A1(n17981), .A2(n17980), .A3(n17979), .A4(n17978), .ZN(
        n17987) );
  AOI22_X1 U19943 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17985) );
  AOI22_X1 U19944 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U19945 ( .A1(n18134), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17983) );
  AOI22_X1 U19946 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17982) );
  NAND4_X1 U19947 ( .A1(n17985), .A2(n17984), .A3(n17983), .A4(n17982), .ZN(
        n17986) );
  NOR2_X1 U19948 ( .A1(n17987), .A2(n17986), .ZN(n21169) );
  OAI21_X1 U19949 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18016), .A(n17988), .ZN(
        n17989) );
  OAI21_X1 U19950 ( .B1(n21169), .B2(n18034), .A(n17989), .ZN(P3_U2683) );
  AOI22_X1 U19951 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17993) );
  AOI22_X1 U19952 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14388), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U19953 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U19954 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17901), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17990) );
  NAND4_X1 U19955 ( .A1(n17993), .A2(n17992), .A3(n17991), .A4(n17990), .ZN(
        n17999) );
  AOI22_X1 U19956 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17997) );
  AOI22_X1 U19957 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U19958 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17995) );
  AOI22_X1 U19959 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17994) );
  NAND4_X1 U19960 ( .A1(n17997), .A2(n17996), .A3(n17995), .A4(n17994), .ZN(
        n17998) );
  NOR2_X1 U19961 ( .A1(n17999), .A2(n17998), .ZN(n21188) );
  AOI211_X1 U19962 ( .C1(n20912), .C2(n18028), .A(n18000), .B(n18035), .ZN(
        n18001) );
  AOI21_X1 U19963 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n18027), .A(n18001), .ZN(
        n18002) );
  OAI21_X1 U19964 ( .B1(n21188), .B2(n18034), .A(n18002), .ZN(P3_U2685) );
  INV_X1 U19965 ( .A(n18003), .ZN(n18004) );
  OAI21_X1 U19966 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18004), .A(n18034), .ZN(
        n18015) );
  AOI22_X1 U19967 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18128), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18008) );
  AOI22_X1 U19968 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18007) );
  AOI22_X1 U19969 ( .A1(n18116), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18006) );
  AOI22_X1 U19970 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18005) );
  NAND4_X1 U19971 ( .A1(n18008), .A2(n18007), .A3(n18006), .A4(n18005), .ZN(
        n18014) );
  AOI22_X1 U19972 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18012) );
  AOI22_X1 U19973 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18011) );
  AOI22_X1 U19974 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18010) );
  AOI22_X1 U19975 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18009) );
  NAND4_X1 U19976 ( .A1(n18012), .A2(n18011), .A3(n18010), .A4(n18009), .ZN(
        n18013) );
  NOR2_X1 U19977 ( .A1(n18014), .A2(n18013), .ZN(n21184) );
  OAI22_X1 U19978 ( .A1(n18016), .A2(n18015), .B1(n21184), .B2(n18034), .ZN(
        P3_U2684) );
  AOI22_X1 U19979 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18155), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n18116), .ZN(n18020) );
  AOI22_X1 U19980 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U19981 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18105), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n18127), .ZN(n18018) );
  AOI22_X1 U19982 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18082), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n18148), .ZN(n18017) );
  NAND4_X1 U19983 ( .A1(n18020), .A2(n18019), .A3(n18018), .A4(n18017), .ZN(
        n18026) );
  AOI22_X1 U19984 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18158), .ZN(n18024) );
  AOI22_X1 U19985 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11176), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n11174), .ZN(n18023) );
  AOI22_X1 U19986 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14484), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U19987 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18021) );
  NAND4_X1 U19988 ( .A1(n18024), .A2(n18023), .A3(n18022), .A4(n18021), .ZN(
        n18025) );
  NOR2_X1 U19989 ( .A1(n18026), .A2(n18025), .ZN(n21194) );
  NAND2_X1 U19990 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18027), .ZN(n18031) );
  INV_X1 U19991 ( .A(n18035), .ZN(n18036) );
  OAI211_X1 U19992 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n18029), .A(n18036), .B(
        n18028), .ZN(n18030) );
  OAI211_X1 U19993 ( .C1(n21194), .C2(n18034), .A(n18031), .B(n18030), .ZN(
        P3_U2686) );
  INV_X1 U19994 ( .A(n18032), .ZN(n18033) );
  OAI21_X1 U19995 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18033), .ZN(n20677) );
  OAI222_X1 U19996 ( .A1(n20677), .A2(n18035), .B1(n20682), .B2(n18039), .C1(
        n18107), .C2(n18034), .ZN(P3_U2702) );
  AOI22_X1 U19997 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18037), .B1(
        n18036), .B2(n21091), .ZN(n18038) );
  OAI21_X1 U19998 ( .B1(n18039), .B2(n21091), .A(n18038), .ZN(P3_U2703) );
  INV_X1 U19999 ( .A(n21794), .ZN(n18040) );
  OAI21_X1 U20000 ( .B1(n18040), .B2(n20609), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18041) );
  OAI21_X1 U20001 ( .B1(n18054), .B2(n21830), .A(n18041), .ZN(P3_U2634) );
  OAI21_X1 U20002 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18043), .A(n18042), .ZN(
        n21828) );
  OAI21_X1 U20003 ( .B1(n20602), .B2(n18629), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18044) );
  OAI221_X1 U20004 ( .B1(n18629), .B2(n21828), .C1(n18629), .C2(n19202), .A(
        n18044), .ZN(P3_U2863) );
  INV_X1 U20005 ( .A(n21795), .ZN(n18045) );
  AOI21_X1 U20006 ( .B1(n18047), .B2(n18046), .A(n18045), .ZN(n21776) );
  NAND2_X1 U20007 ( .A1(n21352), .A2(n21776), .ZN(n21349) );
  INV_X1 U20008 ( .A(n18051), .ZN(n21292) );
  NOR2_X1 U20009 ( .A1(n20665), .A2(n18052), .ZN(n21290) );
  INV_X1 U20010 ( .A(n21348), .ZN(n21781) );
  AOI21_X4 U20011 ( .B1(n20602), .B2(n21830), .A(n21835), .ZN(n18607) );
  NAND2_X1 U20012 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18466) );
  NOR2_X1 U20013 ( .A1(n18466), .A2(n18470), .ZN(n20863) );
  NAND3_X1 U20014 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18498) );
  NOR2_X1 U20015 ( .A1(n18498), .A2(n20798), .ZN(n20806) );
  NAND2_X1 U20016 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18243) );
  NOR2_X1 U20017 ( .A1(n18451), .A2(n20671), .ZN(n18055) );
  INV_X1 U20018 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20913) );
  INV_X1 U20019 ( .A(n18219), .ZN(n18218) );
  NOR2_X1 U20020 ( .A1(n18218), .A2(n20671), .ZN(n18220) );
  INV_X1 U20021 ( .A(n18220), .ZN(n18053) );
  OAI21_X1 U20022 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18055), .A(
        n18053), .ZN(n20918) );
  NOR2_X1 U20023 ( .A1(n18054), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18279) );
  INV_X2 U20024 ( .A(n11173), .ZN(n21769) );
  AOI21_X1 U20025 ( .B1(n18582), .B2(n18451), .A(n18607), .ZN(n18454) );
  OR3_X1 U20026 ( .A1(n18451), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18406), .ZN(n18056) );
  OAI211_X1 U20027 ( .C1(n18055), .C2(n18620), .A(n18454), .B(n18056), .ZN(
        n18223) );
  NAND2_X1 U20028 ( .A1(n20913), .A2(n18056), .ZN(n18057) );
  AOI22_X1 U20029 ( .A1(n21769), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n18223), 
        .B2(n18057), .ZN(n18217) );
  AOI22_X1 U20030 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18070) );
  AOI22_X1 U20031 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14388), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18069) );
  AOI22_X1 U20032 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18059) );
  OAI21_X1 U20033 ( .B1(n14351), .B2(n18060), .A(n18059), .ZN(n18066) );
  AOI22_X1 U20034 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U20035 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18063) );
  AOI22_X1 U20036 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18062) );
  AOI22_X1 U20037 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18061) );
  NAND4_X1 U20038 ( .A1(n18064), .A2(n18063), .A3(n18062), .A4(n18061), .ZN(
        n18065) );
  AOI211_X1 U20039 ( .C1(n18067), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n18066), .B(n18065), .ZN(n18068) );
  NAND3_X1 U20040 ( .A1(n18070), .A2(n18069), .A3(n18068), .ZN(n21353) );
  AOI22_X1 U20041 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18071), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U20042 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U20043 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18073) );
  AOI22_X1 U20044 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18072) );
  NAND4_X1 U20045 ( .A1(n18075), .A2(n18074), .A3(n18073), .A4(n18072), .ZN(
        n18081) );
  AOI22_X1 U20046 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U20047 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U20048 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18077) );
  AOI22_X1 U20049 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18076) );
  NAND4_X1 U20050 ( .A1(n18079), .A2(n18078), .A3(n18077), .A4(n18076), .ZN(
        n18080) );
  AOI22_X1 U20051 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18086) );
  AOI22_X1 U20052 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18156), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18085) );
  AOI22_X1 U20053 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U20054 ( .A1(n18082), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18083) );
  NAND4_X1 U20055 ( .A1(n18086), .A2(n18085), .A3(n18084), .A4(n18083), .ZN(
        n18092) );
  AOI22_X1 U20056 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18090) );
  AOI22_X1 U20057 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18089) );
  AOI22_X1 U20058 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18088) );
  AOI22_X1 U20059 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18087) );
  NAND4_X1 U20060 ( .A1(n18090), .A2(n18089), .A3(n18088), .A4(n18087), .ZN(
        n18091) );
  INV_X1 U20061 ( .A(n18188), .ZN(n21147) );
  AOI22_X1 U20062 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18116), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18104) );
  AOI22_X1 U20063 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18103) );
  AOI22_X1 U20064 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18093) );
  OAI21_X1 U20065 ( .B1(n14351), .B2(n18094), .A(n18093), .ZN(n18101) );
  AOI22_X1 U20066 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18099) );
  AOI22_X1 U20067 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18095), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18098) );
  AOI22_X1 U20068 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18097) );
  AOI22_X1 U20069 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18096) );
  NAND4_X1 U20070 ( .A1(n18099), .A2(n18098), .A3(n18097), .A4(n18096), .ZN(
        n18100) );
  AOI211_X1 U20071 ( .C1(n18132), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n18101), .B(n18100), .ZN(n18102) );
  NAND3_X1 U20072 ( .A1(n18104), .A2(n18103), .A3(n18102), .ZN(n21151) );
  AOI22_X1 U20073 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18156), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18127), .ZN(n18113) );
  AOI22_X1 U20074 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11168), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18112) );
  AOI22_X1 U20075 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14387), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18111) );
  AOI22_X1 U20076 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18134), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18108), .ZN(n18110) );
  AOI22_X1 U20077 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U20078 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18157), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18124) );
  AOI22_X1 U20079 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18114) );
  OAI21_X1 U20080 ( .B1(n14351), .B2(n18115), .A(n18114), .ZN(n18122) );
  AOI22_X1 U20081 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11176), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U20082 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18155), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U20083 ( .A1(n18126), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18116), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U20084 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18117) );
  NAND4_X1 U20085 ( .A1(n18120), .A2(n18119), .A3(n18118), .A4(n18117), .ZN(
        n18121) );
  AOI211_X1 U20086 ( .C1(n18108), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n18122), .B(n18121), .ZN(n18123) );
  NAND3_X1 U20087 ( .A1(n18125), .A2(n18124), .A3(n18123), .ZN(n21143) );
  AOI22_X1 U20088 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18126), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18143) );
  AOI22_X1 U20089 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18127), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18142) );
  AOI22_X1 U20090 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18148), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18130) );
  OAI21_X1 U20091 ( .B1(n14351), .B2(n18131), .A(n18130), .ZN(n18140) );
  AOI22_X1 U20092 ( .A1(n18133), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18132), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U20093 ( .A1(n11175), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18137) );
  AOI22_X1 U20094 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18136) );
  AOI22_X1 U20095 ( .A1(n11174), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18135) );
  NAND4_X1 U20096 ( .A1(n18138), .A2(n18137), .A3(n18136), .A4(n18135), .ZN(
        n18139) );
  AOI211_X1 U20097 ( .C1(n11176), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n18140), .B(n18139), .ZN(n18141) );
  NAND3_X1 U20098 ( .A1(n18143), .A2(n18142), .A3(n18141), .ZN(n18183) );
  INV_X1 U20099 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18225) );
  NAND2_X1 U20100 ( .A1(n18416), .A2(n18225), .ZN(n18281) );
  INV_X1 U20101 ( .A(n18281), .ZN(n18299) );
  AOI21_X1 U20102 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18492), .A(
        n18299), .ZN(n18182) );
  INV_X1 U20103 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21722) );
  INV_X1 U20104 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21534) );
  INV_X1 U20105 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21733) );
  NAND2_X1 U20106 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21475) );
  INV_X1 U20107 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21484) );
  NOR2_X1 U20108 ( .A1(n21475), .A2(n21484), .ZN(n21492) );
  NAND2_X1 U20109 ( .A1(n21492), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n21502) );
  NOR2_X1 U20110 ( .A1(n21733), .A2(n21502), .ZN(n18234) );
  NAND2_X1 U20111 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18234), .ZN(
        n21535) );
  NOR2_X1 U20112 ( .A1(n21534), .A2(n21535), .ZN(n21696) );
  INV_X1 U20113 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21755) );
  AOI22_X1 U20114 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18416), .B1(
        n18492), .B2(n21755), .ZN(n18527) );
  AOI21_X1 U20115 ( .B1(n21359), .B2(n21637), .A(n18492), .ZN(n18175) );
  INV_X1 U20116 ( .A(n18183), .ZN(n21133) );
  XNOR2_X1 U20117 ( .A(n21133), .B(n18144), .ZN(n18173) );
  NAND2_X1 U20118 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18173), .ZN(
        n18174) );
  XOR2_X1 U20119 ( .A(n21143), .B(n18145), .Z(n18146) );
  NAND2_X1 U20120 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18146), .ZN(
        n18168) );
  INV_X1 U20121 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21419) );
  XNOR2_X1 U20122 ( .A(n21419), .B(n18146), .ZN(n18580) );
  INV_X1 U20123 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21399) );
  XOR2_X1 U20124 ( .A(n21151), .B(n21275), .Z(n18147) );
  XNOR2_X1 U20125 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n18147), .ZN(
        n18600) );
  INV_X1 U20126 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21390) );
  AOI22_X1 U20127 ( .A1(n11176), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11174), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18153) );
  AOI22_X1 U20128 ( .A1(n17895), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18134), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18152) );
  AOI22_X1 U20129 ( .A1(n18148), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18151) );
  AOI22_X1 U20130 ( .A1(n18129), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18149), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18150) );
  NAND4_X1 U20131 ( .A1(n18153), .A2(n18152), .A3(n18151), .A4(n18150), .ZN(
        n18164) );
  AOI22_X1 U20132 ( .A1(n18155), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18154), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U20133 ( .A1(n18128), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11175), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U20134 ( .A1(n18157), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18156), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18160) );
  AOI22_X1 U20135 ( .A1(n18067), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18158), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18159) );
  NAND4_X1 U20136 ( .A1(n18162), .A2(n18161), .A3(n18160), .A4(n18159), .ZN(
        n18163) );
  NOR2_X1 U20137 ( .A1(n18164), .A2(n18163), .ZN(n18194) );
  INV_X1 U20138 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21468) );
  NOR2_X1 U20139 ( .A1(n18194), .A2(n21468), .ZN(n18618) );
  OAI21_X1 U20140 ( .B1(n21390), .B2(n18193), .A(n18609), .ZN(n18599) );
  NAND2_X1 U20141 ( .A1(n18600), .A2(n18599), .ZN(n18598) );
  NAND2_X1 U20142 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18166), .ZN(
        n18167) );
  XNOR2_X1 U20143 ( .A(n18188), .B(n18191), .ZN(n18592) );
  NAND2_X1 U20144 ( .A1(n18580), .A2(n18579), .ZN(n18578) );
  XOR2_X1 U20145 ( .A(n21138), .B(n18169), .Z(n18171) );
  NAND2_X1 U20146 ( .A1(n18171), .A2(n18170), .ZN(n18172) );
  INV_X1 U20147 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21440) );
  XNOR2_X1 U20148 ( .A(n21440), .B(n18173), .ZN(n18554) );
  NAND2_X1 U20149 ( .A1(n18175), .A2(n18232), .ZN(n18176) );
  OAI21_X1 U20150 ( .B1(n18492), .B2(n21755), .A(n18525), .ZN(n18177) );
  NAND2_X1 U20151 ( .A1(n21696), .A2(n18177), .ZN(n18179) );
  NOR2_X1 U20152 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18178) );
  NOR2_X1 U20153 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18504) );
  INV_X1 U20154 ( .A(n18177), .ZN(n18494) );
  INV_X1 U20155 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18268) );
  INV_X1 U20156 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18458) );
  NAND2_X1 U20157 ( .A1(n18457), .A2(n18458), .ZN(n18456) );
  NAND2_X1 U20158 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21575) );
  INV_X1 U20159 ( .A(n18179), .ZN(n18180) );
  NOR2_X1 U20160 ( .A1(n18181), .A2(n18180), .ZN(n18338) );
  OR2_X1 U20161 ( .A1(n21575), .A2(n18338), .ZN(n18224) );
  XNOR2_X1 U20162 ( .A(n18182), .B(n18282), .ZN(n21697) );
  NOR2_X1 U20163 ( .A1(n21275), .A2(n18194), .ZN(n18195) );
  NOR2_X1 U20164 ( .A1(n18188), .A2(n18190), .ZN(n18200) );
  NAND2_X1 U20165 ( .A1(n18200), .A2(n21143), .ZN(n18186) );
  NOR2_X1 U20166 ( .A1(n21138), .A2(n18186), .ZN(n18185) );
  NAND2_X1 U20167 ( .A1(n18185), .A2(n18183), .ZN(n18184) );
  NOR2_X1 U20168 ( .A1(n21359), .A2(n18184), .ZN(n18210) );
  XNOR2_X1 U20169 ( .A(n21353), .B(n18184), .ZN(n18546) );
  XNOR2_X1 U20170 ( .A(n21133), .B(n18185), .ZN(n18203) );
  XOR2_X1 U20171 ( .A(n21138), .B(n18186), .Z(n18187) );
  NAND2_X1 U20172 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18187), .ZN(
        n18202) );
  INV_X1 U20173 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21426) );
  XNOR2_X1 U20174 ( .A(n21426), .B(n18187), .ZN(n18568) );
  XOR2_X1 U20175 ( .A(n18188), .B(n18190), .Z(n18189) );
  NAND2_X1 U20176 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18189), .ZN(
        n18198) );
  INV_X1 U20177 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21420) );
  XNOR2_X1 U20178 ( .A(n21420), .B(n18189), .ZN(n18589) );
  INV_X1 U20179 ( .A(n18194), .ZN(n21276) );
  NAND2_X1 U20180 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18192), .ZN(
        n18197) );
  NOR2_X1 U20181 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18193), .ZN(
        n18196) );
  NAND2_X1 U20182 ( .A1(n18194), .A2(n21468), .ZN(n18616) );
  NOR2_X1 U20183 ( .A1(n18611), .A2(n18616), .ZN(n18610) );
  NOR3_X1 U20184 ( .A1(n18196), .A2(n18195), .A3(n18610), .ZN(n18603) );
  NAND2_X1 U20185 ( .A1(n18604), .A2(n18603), .ZN(n18602) );
  NAND2_X1 U20186 ( .A1(n18197), .A2(n18602), .ZN(n18588) );
  NAND2_X1 U20187 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18199), .ZN(
        n18201) );
  XOR2_X1 U20188 ( .A(n21143), .B(n18200), .Z(n18575) );
  NAND2_X1 U20189 ( .A1(n18201), .A2(n18574), .ZN(n18567) );
  NAND2_X1 U20190 ( .A1(n18568), .A2(n18567), .ZN(n18566) );
  NAND2_X1 U20191 ( .A1(n18202), .A2(n18566), .ZN(n18204) );
  NAND2_X1 U20192 ( .A1(n18203), .A2(n18204), .ZN(n18205) );
  INV_X1 U20193 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21456) );
  NAND2_X1 U20194 ( .A1(n18210), .A2(n18206), .ZN(n18211) );
  INV_X1 U20195 ( .A(n18206), .ZN(n18209) );
  NAND2_X1 U20196 ( .A1(n18546), .A2(n18545), .ZN(n18208) );
  NAND2_X1 U20197 ( .A1(n18210), .A2(n18209), .ZN(n18207) );
  OAI211_X1 U20198 ( .C1(n18210), .C2(n18209), .A(n18208), .B(n18207), .ZN(
        n18524) );
  NAND2_X1 U20199 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18524), .ZN(
        n18523) );
  NOR2_X2 U20200 ( .A1(n21341), .A2(n18212), .ZN(n18549) );
  NOR2_X2 U20201 ( .A1(n18490), .A2(n21755), .ZN(n21701) );
  INV_X1 U20202 ( .A(n21701), .ZN(n21469) );
  INV_X1 U20203 ( .A(n18465), .ZN(n18214) );
  INV_X1 U20204 ( .A(n18234), .ZN(n21506) );
  INV_X1 U20205 ( .A(n21502), .ZN(n18252) );
  NAND2_X1 U20206 ( .A1(n21701), .A2(n18252), .ZN(n21487) );
  OAI22_X1 U20207 ( .A1(n21698), .A2(n18624), .B1(n21517), .B2(n18484), .ZN(
        n18241) );
  AOI21_X1 U20208 ( .B1(n18214), .B2(n21575), .A(n18241), .ZN(n18459) );
  INV_X1 U20209 ( .A(n21575), .ZN(n21699) );
  NAND2_X1 U20210 ( .A1(n21699), .A2(n18225), .ZN(n21711) );
  OAI22_X1 U20211 ( .A1(n18459), .A2(n18225), .B1(n18465), .B2(n21711), .ZN(
        n18215) );
  AOI21_X1 U20212 ( .B1(n18535), .B2(n21697), .A(n18215), .ZN(n18216) );
  OAI211_X1 U20213 ( .C1(n18397), .C2(n20918), .A(n18217), .B(n18216), .ZN(
        P3_U2812) );
  NOR2_X1 U20214 ( .A1(n21575), .A2(n18225), .ZN(n21354) );
  NAND3_X1 U20215 ( .A1(n21354), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21517), .ZN(n21678) );
  NAND3_X1 U20216 ( .A1(n21354), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21698), .ZN(n21677) );
  AOI22_X1 U20217 ( .A1(n18536), .A2(n21678), .B1(n18549), .B2(n21677), .ZN(
        n18311) );
  INV_X1 U20218 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21686) );
  NOR3_X1 U20219 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18406), .A3(
        n18218), .ZN(n18222) );
  INV_X1 U20220 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20934) );
  OAI22_X1 U20221 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18220), .B1(
        n20671), .B2(n18302), .ZN(n20931) );
  OAI22_X1 U20222 ( .A1(n11173), .A2(n20934), .B1(n18397), .B2(n20931), .ZN(
        n18221) );
  AOI211_X1 U20223 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n18223), .A(
        n18222), .B(n18221), .ZN(n18228) );
  NOR2_X1 U20224 ( .A1(n18281), .A2(n18282), .ZN(n18292) );
  NOR3_X1 U20225 ( .A1(n18416), .A2(n18225), .A3(n18224), .ZN(n18298) );
  NOR2_X1 U20226 ( .A1(n18292), .A2(n18298), .ZN(n18226) );
  XNOR2_X1 U20227 ( .A(n18226), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21684) );
  INV_X1 U20228 ( .A(n21354), .ZN(n21355) );
  AOI22_X1 U20229 ( .A1(n18535), .A2(n21684), .B1(n18359), .B2(n21686), .ZN(
        n18227) );
  OAI211_X1 U20230 ( .C1(n18311), .C2(n21686), .A(n18228), .B(n18227), .ZN(
        P3_U2811) );
  INV_X1 U20231 ( .A(n21517), .ZN(n21523) );
  NAND2_X1 U20232 ( .A1(n18536), .A2(n21523), .ZN(n18240) );
  NOR2_X1 U20233 ( .A1(n18229), .A2(n20671), .ZN(n18468) );
  AOI21_X1 U20234 ( .B1(n18582), .B2(n18229), .A(n18607), .ZN(n18479) );
  OAI21_X1 U20235 ( .B1(n18468), .B2(n18620), .A(n18479), .ZN(n18245) );
  INV_X1 U20236 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20878) );
  NOR2_X1 U20237 ( .A1(n11173), .A2(n20878), .ZN(n18231) );
  NAND3_X1 U20238 ( .A1(n18255), .A2(n20863), .A3(n18363), .ZN(n18248) );
  NAND2_X1 U20239 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18468), .ZN(
        n18244) );
  OAI21_X1 U20240 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18468), .A(
        n18244), .ZN(n20869) );
  OAI22_X1 U20241 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18248), .B1(
        n20869), .B2(n18397), .ZN(n18230) );
  AOI211_X1 U20242 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18245), .A(
        n18231), .B(n18230), .ZN(n18239) );
  INV_X1 U20243 ( .A(n18232), .ZN(n18233) );
  NAND2_X1 U20244 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21478) );
  NOR3_X1 U20245 ( .A1(n18233), .A2(n18416), .A3(n21478), .ZN(n18265) );
  NAND2_X1 U20246 ( .A1(n18234), .A2(n18265), .ZN(n18471) );
  NAND2_X1 U20247 ( .A1(n18490), .A2(n18235), .ZN(n18472) );
  INV_X1 U20248 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21516) );
  AOI22_X1 U20249 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18471), .B1(
        n18472), .B2(n21516), .ZN(n18236) );
  XNOR2_X1 U20250 ( .A(n21534), .B(n18236), .ZN(n21527) );
  OAI21_X1 U20251 ( .B1(n21520), .B2(n18624), .A(n21534), .ZN(n18237) );
  AOI22_X1 U20252 ( .A1(n18535), .A2(n21527), .B1(n18241), .B2(n18237), .ZN(
        n18238) );
  OAI211_X1 U20253 ( .C1(n21525), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        P3_U2815) );
  INV_X1 U20254 ( .A(n18241), .ZN(n18251) );
  AOI22_X1 U20255 ( .A1(n18492), .A2(n21722), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18416), .ZN(n18242) );
  XNOR2_X1 U20256 ( .A(n18338), .B(n18242), .ZN(n21725) );
  OAI21_X1 U20257 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18243), .ZN(n18247) );
  INV_X1 U20258 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20885) );
  INV_X1 U20259 ( .A(n18453), .ZN(n20905) );
  NOR2_X1 U20260 ( .A1(n20905), .A2(n20671), .ZN(n18452) );
  AOI21_X1 U20261 ( .B1(n20885), .B2(n18244), .A(n18452), .ZN(n20882) );
  AOI22_X1 U20262 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18245), .B1(
        n18446), .B2(n20882), .ZN(n18246) );
  NAND2_X1 U20263 ( .A1(n18279), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n21726) );
  OAI211_X1 U20264 ( .C1(n18248), .C2(n18247), .A(n18246), .B(n21726), .ZN(
        n18249) );
  AOI21_X1 U20265 ( .B1(n18535), .B2(n21725), .A(n18249), .ZN(n18250) );
  OAI221_X1 U20266 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18465), 
        .C1(n21722), .C2(n18251), .A(n18250), .ZN(P3_U2814) );
  NAND2_X1 U20267 ( .A1(n21492), .A2(n18521), .ZN(n18262) );
  NAND2_X1 U20268 ( .A1(n18252), .A2(n21472), .ZN(n21486) );
  AOI22_X1 U20269 ( .A1(n18549), .A2(n21486), .B1(n18536), .B2(n21487), .ZN(
        n18270) );
  NAND3_X1 U20270 ( .A1(n18490), .A2(n18504), .A3(n21755), .ZN(n18485) );
  INV_X1 U20271 ( .A(n18265), .ZN(n18509) );
  INV_X1 U20272 ( .A(n21492), .ZN(n18253) );
  OAI22_X1 U20273 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18485), .B1(
        n18509), .B2(n18253), .ZN(n18254) );
  XNOR2_X1 U20274 ( .A(n18268), .B(n18254), .ZN(n21493) );
  INV_X1 U20275 ( .A(n18255), .ZN(n18256) );
  NOR2_X1 U20276 ( .A1(n18256), .A2(n20671), .ZN(n18481) );
  NAND2_X1 U20277 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18481), .ZN(
        n18263) );
  OAI21_X1 U20278 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18481), .A(
        n18263), .ZN(n20829) );
  NOR2_X1 U20279 ( .A1(n18397), .A2(n20829), .ZN(n18260) );
  INV_X1 U20280 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20833) );
  NOR2_X1 U20281 ( .A1(n18256), .A2(n18406), .ZN(n18272) );
  AOI21_X1 U20282 ( .B1(n18256), .B2(n18582), .A(n18315), .ZN(n18257) );
  OAI21_X1 U20283 ( .B1(n18481), .B2(n18257), .A(n18619), .ZN(n18264) );
  INV_X1 U20284 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20848) );
  NOR2_X1 U20285 ( .A1(n11173), .A2(n20848), .ZN(n21494) );
  AOI221_X1 U20286 ( .B1(n20833), .B2(n18272), .C1(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18264), .A(n21494), .ZN(
        n18258) );
  INV_X1 U20287 ( .A(n18258), .ZN(n18259) );
  AOI211_X1 U20288 ( .C1(n18535), .C2(n21493), .A(n18260), .B(n18259), .ZN(
        n18261) );
  OAI221_X1 U20289 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18262), 
        .C1(n18268), .C2(n18270), .A(n18261), .ZN(P3_U2818) );
  INV_X1 U20290 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20839) );
  NOR2_X1 U20291 ( .A1(n20839), .A2(n18263), .ZN(n20835) );
  AOI21_X1 U20292 ( .B1(n20839), .B2(n18263), .A(n20835), .ZN(n20843) );
  AOI22_X1 U20293 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18264), .B1(
        n18446), .B2(n20843), .ZN(n18275) );
  NOR2_X1 U20294 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21502), .ZN(
        n21736) );
  NAND2_X1 U20295 ( .A1(n21492), .A2(n18265), .ZN(n18266) );
  AOI22_X1 U20296 ( .A1(n18492), .A2(n18268), .B1(n18267), .B2(n18266), .ZN(
        n18269) );
  XNOR2_X1 U20297 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18269), .ZN(
        n21739) );
  OAI22_X1 U20298 ( .A1(n18270), .A2(n21733), .B1(n18508), .B2(n21739), .ZN(
        n18271) );
  AOI21_X1 U20299 ( .B1(n21736), .B2(n18521), .A(n18271), .ZN(n18274) );
  NAND2_X1 U20300 ( .A1(n21769), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n21737) );
  OAI211_X1 U20301 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18272), .B(n18466), .ZN(n18273) );
  NAND4_X1 U20302 ( .A1(n18275), .A2(n18274), .A3(n21737), .A4(n18273), .ZN(
        P3_U2817) );
  INV_X1 U20303 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18278) );
  INV_X1 U20304 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n20941) );
  NAND2_X1 U20305 ( .A1(n11274), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18303) );
  NOR2_X1 U20306 ( .A1(n18278), .A2(n18303), .ZN(n18276) );
  OAI22_X1 U20307 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18276), .B1(
        n20671), .B2(n18313), .ZN(n20970) );
  NOR2_X1 U20308 ( .A1(n18302), .A2(n20671), .ZN(n18304) );
  OAI22_X1 U20309 ( .A1(n11274), .A2(n18528), .B1(n18304), .B2(n18620), .ZN(
        n18277) );
  NOR2_X1 U20310 ( .A1(n18607), .A2(n18277), .ZN(n18301) );
  OAI21_X1 U20311 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18407), .A(
        n18301), .ZN(n18291) );
  INV_X1 U20312 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20964) );
  NAND2_X1 U20313 ( .A1(n11274), .A2(n18363), .ZN(n18289) );
  AOI221_X1 U20314 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n20964), .C2(n18278), .A(
        n18289), .ZN(n18280) );
  INV_X1 U20315 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18704) );
  NOR2_X1 U20316 ( .A1(n11173), .A2(n18704), .ZN(n21543) );
  AOI211_X1 U20317 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n18291), .A(
        n18280), .B(n21543), .ZN(n18288) );
  NOR4_X1 U20318 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n18281), .ZN(n18323) );
  NAND2_X1 U20319 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21366) );
  INV_X1 U20320 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21533) );
  NOR2_X1 U20321 ( .A1(n21366), .A2(n21533), .ZN(n21538) );
  OAI21_X1 U20322 ( .B1(n18323), .B2(n18341), .A(n18340), .ZN(n18324) );
  XNOR2_X1 U20323 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18324), .ZN(
        n21544) );
  NAND2_X1 U20324 ( .A1(n21354), .A2(n21538), .ZN(n18283) );
  NOR2_X1 U20325 ( .A1(n18465), .A2(n18283), .ZN(n18285) );
  NAND3_X1 U20326 ( .A1(n21354), .A2(n21538), .A3(n21517), .ZN(n21363) );
  NAND3_X1 U20327 ( .A1(n21354), .A2(n21538), .A3(n21698), .ZN(n21362) );
  AOI22_X1 U20328 ( .A1(n18536), .A2(n21363), .B1(n18549), .B2(n21362), .ZN(
        n18297) );
  INV_X1 U20329 ( .A(n18297), .ZN(n18284) );
  MUX2_X1 U20330 ( .A(n18285), .B(n18284), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n18286) );
  AOI21_X1 U20331 ( .B1(n18535), .B2(n21544), .A(n18286), .ZN(n18287) );
  OAI211_X1 U20332 ( .C1(n18397), .C2(n20970), .A(n18288), .B(n18287), .ZN(
        P3_U2808) );
  INV_X1 U20333 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20952) );
  NOR2_X1 U20334 ( .A1(n11173), .A2(n20952), .ZN(n21369) );
  XOR2_X1 U20335 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n18303), .Z(
        n20955) );
  OAI22_X1 U20336 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18289), .B1(
        n20955), .B2(n18397), .ZN(n18290) );
  AOI211_X1 U20337 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n18291), .A(
        n21369), .B(n18290), .ZN(n18296) );
  INV_X1 U20338 ( .A(n21366), .ZN(n21365) );
  NOR2_X1 U20339 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18293) );
  AOI22_X1 U20340 ( .A1(n21365), .A2(n18298), .B1(n18293), .B2(n18292), .ZN(
        n18294) );
  XNOR2_X1 U20341 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18294), .ZN(
        n21370) );
  NOR2_X1 U20342 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21366), .ZN(
        n21335) );
  AOI22_X1 U20343 ( .A1(n18535), .A2(n21370), .B1(n18359), .B2(n21335), .ZN(
        n18295) );
  OAI211_X1 U20344 ( .C1(n18297), .C2(n21533), .A(n18296), .B(n18295), .ZN(
        P3_U2809) );
  INV_X1 U20345 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18310) );
  OAI221_X1 U20346 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18299), 
        .C1(n21686), .C2(n18298), .A(n18340), .ZN(n18300) );
  XNOR2_X1 U20347 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18300), .ZN(
        n21690) );
  AOI221_X1 U20348 ( .B1(n18302), .B2(n20941), .C1(n19324), .C2(n20941), .A(
        n18301), .ZN(n18306) );
  OAI21_X1 U20349 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18304), .A(
        n18303), .ZN(n20946) );
  NAND2_X1 U20350 ( .A1(n21769), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21692) );
  OAI221_X1 U20351 ( .B1(n20946), .B2(n18397), .C1(n20946), .C2(n18407), .A(
        n21692), .ZN(n18305) );
  AOI211_X1 U20352 ( .C1(n21690), .C2(n18535), .A(n18306), .B(n18305), .ZN(
        n18309) );
  NAND2_X1 U20353 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18310), .ZN(
        n21694) );
  INV_X1 U20354 ( .A(n21694), .ZN(n18307) );
  NAND2_X1 U20355 ( .A1(n18359), .A2(n18307), .ZN(n18308) );
  OAI211_X1 U20356 ( .C1(n18311), .C2(n18310), .A(n18309), .B(n18308), .ZN(
        P3_U2810) );
  NAND2_X1 U20357 ( .A1(n21538), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18400) );
  INV_X1 U20358 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21665) );
  NOR2_X1 U20359 ( .A1(n18400), .A2(n21665), .ZN(n18358) );
  NAND2_X1 U20360 ( .A1(n21354), .A2(n18358), .ZN(n18337) );
  INV_X1 U20361 ( .A(n18337), .ZN(n18312) );
  NAND2_X1 U20362 ( .A1(n18312), .A2(n21698), .ZN(n21657) );
  NAND2_X1 U20363 ( .A1(n18312), .A2(n21517), .ZN(n21658) );
  AOI22_X1 U20364 ( .A1(n18549), .A2(n21657), .B1(n18536), .B2(n21658), .ZN(
        n18357) );
  INV_X1 U20365 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18317) );
  NOR2_X1 U20366 ( .A1(n18331), .A2(n19324), .ZN(n18320) );
  INV_X1 U20367 ( .A(n18313), .ZN(n18319) );
  INV_X1 U20368 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18705) );
  NOR2_X1 U20369 ( .A1(n11173), .A2(n18705), .ZN(n21667) );
  NOR2_X1 U20370 ( .A1(n18313), .A2(n20671), .ZN(n18316) );
  INV_X1 U20371 ( .A(n18316), .ZN(n18314) );
  AOI211_X1 U20372 ( .C1(n18315), .C2(n18314), .A(n18607), .B(n18320), .ZN(
        n18329) );
  NAND2_X1 U20373 ( .A1(n18331), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18346) );
  OAI21_X1 U20374 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18316), .A(
        n18346), .ZN(n20979) );
  OAI22_X1 U20375 ( .A1(n18329), .A2(n18317), .B1(n18605), .B2(n20979), .ZN(
        n18318) );
  AOI211_X1 U20376 ( .C1(n18320), .C2(n18319), .A(n21667), .B(n18318), .ZN(
        n18328) );
  NAND2_X1 U20377 ( .A1(n18549), .A2(n21657), .ZN(n18322) );
  NAND2_X1 U20378 ( .A1(n18536), .A2(n21658), .ZN(n18321) );
  OAI22_X1 U20379 ( .A1(n21362), .A2(n18322), .B1(n21363), .B2(n18321), .ZN(
        n18326) );
  INV_X1 U20380 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21546) );
  NAND2_X1 U20381 ( .A1(n18323), .A2(n21546), .ZN(n18336) );
  AOI221_X1 U20382 ( .B1(n18416), .B2(n18336), .C1(n21546), .C2(n18336), .A(
        n18324), .ZN(n18325) );
  XNOR2_X1 U20383 ( .A(n18325), .B(n21665), .ZN(n21668) );
  AOI22_X1 U20384 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18326), .B1(
        n18535), .B2(n21668), .ZN(n18327) );
  OAI211_X1 U20385 ( .C1(n18357), .C2(n21665), .A(n18328), .B(n18327), .ZN(
        P3_U2807) );
  INV_X1 U20386 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18356) );
  XOR2_X1 U20387 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18361), .Z(
        n21553) );
  INV_X1 U20388 ( .A(n21553), .ZN(n18345) );
  OAI21_X1 U20389 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18407), .A(
        n18329), .ZN(n18350) );
  INV_X1 U20390 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18330) );
  INV_X1 U20391 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20989) );
  NAND2_X1 U20392 ( .A1(n18331), .A2(n18363), .ZN(n18347) );
  AOI221_X1 U20393 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n18330), .C2(n20989), .A(
        n18347), .ZN(n18335) );
  INV_X1 U20394 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21001) );
  NOR2_X1 U20395 ( .A1(n20989), .A2(n18346), .ZN(n18333) );
  NAND3_X1 U20396 ( .A1(n18331), .A2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18394) );
  NOR2_X1 U20397 ( .A1(n18394), .A2(n20671), .ZN(n18396) );
  INV_X1 U20398 ( .A(n18396), .ZN(n18332) );
  OAI21_X1 U20399 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18333), .A(
        n18332), .ZN(n21005) );
  OAI22_X1 U20400 ( .A1(n11173), .A2(n21001), .B1(n18397), .B2(n21005), .ZN(
        n18334) );
  AOI211_X1 U20401 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18350), .A(
        n18335), .B(n18334), .ZN(n18344) );
  NOR2_X1 U20402 ( .A1(n18356), .A2(n21657), .ZN(n18360) );
  INV_X1 U20403 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21565) );
  XNOR2_X1 U20404 ( .A(n18360), .B(n21565), .ZN(n21554) );
  OAI22_X1 U20405 ( .A1(n18338), .A2(n18337), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18336), .ZN(n18339) );
  NAND2_X1 U20406 ( .A1(n18416), .A2(n18351), .ZN(n18390) );
  OAI21_X1 U20407 ( .B1(n18416), .B2(n18391), .A(n18390), .ZN(n18342) );
  XNOR2_X1 U20408 ( .A(n18342), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21555) );
  AOI22_X1 U20409 ( .A1(n18549), .A2(n21554), .B1(n18535), .B2(n21555), .ZN(
        n18343) );
  OAI211_X1 U20410 ( .C1(n18484), .C2(n18345), .A(n18344), .B(n18343), .ZN(
        P3_U2805) );
  INV_X1 U20411 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21000) );
  NOR2_X1 U20412 ( .A1(n11173), .A2(n21000), .ZN(n18349) );
  XOR2_X1 U20413 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n18346), .Z(
        n20995) );
  OAI22_X1 U20414 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18347), .B1(
        n20995), .B2(n18397), .ZN(n18348) );
  AOI211_X1 U20415 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n18350), .A(
        n18349), .B(n18348), .ZN(n18355) );
  OAI21_X1 U20416 ( .B1(n18352), .B2(n18356), .A(n18351), .ZN(n21670) );
  NAND2_X1 U20417 ( .A1(n18358), .A2(n18356), .ZN(n21676) );
  INV_X1 U20418 ( .A(n21676), .ZN(n18353) );
  AOI22_X1 U20419 ( .A1(n18535), .A2(n21670), .B1(n18359), .B2(n18353), .ZN(
        n18354) );
  OAI211_X1 U20420 ( .C1(n18357), .C2(n18356), .A(n18355), .B(n18354), .ZN(
        P3_U2806) );
  NAND2_X1 U20421 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21573) );
  NAND2_X1 U20422 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18358), .ZN(
        n21550) );
  NOR2_X1 U20423 ( .A1(n21573), .A2(n21550), .ZN(n21589) );
  INV_X1 U20424 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21606) );
  NAND2_X1 U20425 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21606), .ZN(
        n21639) );
  INV_X1 U20426 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21039) );
  INV_X1 U20427 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21016) );
  OR2_X1 U20428 ( .A1(n18368), .A2(n20671), .ZN(n18379) );
  AND2_X1 U20429 ( .A1(n18442), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18444) );
  AOI21_X1 U20430 ( .B1(n21039), .B2(n18379), .A(n18444), .ZN(n21058) );
  INV_X1 U20431 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21596) );
  INV_X1 U20432 ( .A(n21573), .ZN(n18362) );
  NAND2_X1 U20433 ( .A1(n18362), .A2(n18360), .ZN(n21580) );
  INV_X1 U20434 ( .A(n21580), .ZN(n21559) );
  NAND2_X1 U20435 ( .A1(n18362), .A2(n18361), .ZN(n21603) );
  INV_X1 U20436 ( .A(n21603), .ZN(n18430) );
  OAI22_X1 U20437 ( .A1(n21559), .A2(n18624), .B1(n18430), .B2(n18484), .ZN(
        n18402) );
  NOR2_X1 U20438 ( .A1(n21596), .A2(n18402), .ZN(n18389) );
  AOI211_X1 U20439 ( .C1(n18484), .C2(n18624), .A(n18389), .B(n21606), .ZN(
        n18370) );
  NAND2_X1 U20440 ( .A1(n21039), .A2(n18363), .ZN(n18367) );
  NAND2_X1 U20441 ( .A1(n21769), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21652) );
  INV_X1 U20442 ( .A(n18364), .ZN(n18395) );
  NOR3_X1 U20443 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18406), .A3(
        n18395), .ZN(n18381) );
  OAI22_X1 U20444 ( .A1(n18364), .A2(n18528), .B1(n18396), .B2(n18620), .ZN(
        n18365) );
  NOR2_X1 U20445 ( .A1(n18607), .A2(n18365), .ZN(n18393) );
  OAI21_X1 U20446 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18407), .A(
        n18393), .ZN(n18385) );
  OAI21_X1 U20447 ( .B1(n18381), .B2(n18385), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18366) );
  OAI211_X1 U20448 ( .C1(n18368), .C2(n18367), .A(n21652), .B(n18366), .ZN(
        n18369) );
  AOI211_X1 U20449 ( .C1(n18446), .C2(n21058), .A(n18370), .B(n18369), .ZN(
        n18378) );
  NOR2_X1 U20450 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18492), .ZN(
        n18413) );
  AOI21_X1 U20451 ( .B1(n18492), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18413), .ZN(n21650) );
  INV_X1 U20452 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21562) );
  AOI21_X1 U20453 ( .B1(n21562), .B2(n21565), .A(n18492), .ZN(n18371) );
  INV_X1 U20454 ( .A(n18371), .ZN(n18372) );
  INV_X1 U20455 ( .A(n18374), .ZN(n18375) );
  NAND2_X1 U20456 ( .A1(n18375), .A2(n21596), .ZN(n21651) );
  INV_X1 U20457 ( .A(n21651), .ZN(n18414) );
  NOR2_X1 U20458 ( .A1(n18375), .A2(n21596), .ZN(n18418) );
  NOR2_X1 U20459 ( .A1(n18414), .A2(n18418), .ZN(n18384) );
  NAND2_X1 U20460 ( .A1(n18384), .A2(n18492), .ZN(n18383) );
  NAND2_X1 U20461 ( .A1(n18383), .A2(n21651), .ZN(n18376) );
  NAND2_X1 U20462 ( .A1(n21650), .A2(n18376), .ZN(n21635) );
  OAI211_X1 U20463 ( .C1(n21650), .C2(n18376), .A(n18535), .B(n21635), .ZN(
        n18377) );
  OAI211_X1 U20464 ( .C1(n18429), .C2(n21639), .A(n18378), .B(n18377), .ZN(
        P3_U2802) );
  AND2_X1 U20465 ( .A1(n21596), .A2(n18429), .ZN(n18388) );
  NOR2_X1 U20466 ( .A1(n18395), .A2(n20671), .ZN(n18380) );
  OAI21_X1 U20467 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18380), .A(
        n18379), .ZN(n21029) );
  INV_X1 U20468 ( .A(n21029), .ZN(n18382) );
  INV_X1 U20469 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21026) );
  NOR2_X1 U20470 ( .A1(n11173), .A2(n21026), .ZN(n21586) );
  AOI211_X1 U20471 ( .C1(n18446), .C2(n18382), .A(n18381), .B(n21586), .ZN(
        n18387) );
  OAI21_X1 U20472 ( .B1(n18492), .B2(n18384), .A(n18383), .ZN(n21587) );
  AOI22_X1 U20473 ( .A1(n18535), .A2(n21587), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18385), .ZN(n18386) );
  OAI211_X1 U20474 ( .C1(n18389), .C2(n18388), .A(n18387), .B(n18386), .ZN(
        P3_U2803) );
  OAI221_X1 U20475 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18416), 
        .C1(n21565), .C2(n18391), .A(n18390), .ZN(n18392) );
  XNOR2_X1 U20476 ( .A(n21562), .B(n18392), .ZN(n21571) );
  AOI221_X1 U20477 ( .B1(n18394), .B2(n21016), .C1(n19324), .C2(n21016), .A(
        n18393), .ZN(n18399) );
  OAI22_X1 U20478 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18396), .B1(
        n20671), .B2(n18395), .ZN(n21021) );
  AOI21_X1 U20479 ( .B1(n18397), .B2(n18407), .A(n21021), .ZN(n18398) );
  AOI211_X1 U20480 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n18279), .A(n18399), 
        .B(n18398), .ZN(n18404) );
  INV_X1 U20481 ( .A(n18400), .ZN(n21564) );
  NAND2_X1 U20482 ( .A1(n21354), .A2(n21564), .ZN(n21576) );
  NAND2_X1 U20483 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21572) );
  NOR4_X1 U20484 ( .A1(n21565), .A2(n21576), .A3(n21572), .A4(n18465), .ZN(
        n18401) );
  AOI22_X1 U20485 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18402), .B1(
        n18401), .B2(n21562), .ZN(n18403) );
  OAI211_X1 U20486 ( .C1(n18508), .C2(n21571), .A(n18404), .B(n18403), .ZN(
        P3_U2804) );
  INV_X1 U20487 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21615) );
  NOR2_X1 U20488 ( .A1(n18415), .A2(n21615), .ZN(n21625) );
  NAND2_X1 U20489 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21590) );
  NAND2_X1 U20490 ( .A1(n21625), .A2(n21646), .ZN(n18405) );
  XOR2_X1 U20491 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n18405), .Z(
        n21628) );
  INV_X1 U20492 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21081) );
  NOR2_X1 U20493 ( .A1(n11173), .A2(n21081), .ZN(n21622) );
  OR2_X1 U20494 ( .A1(n18408), .A2(n18406), .ZN(n18428) );
  XOR2_X1 U20495 ( .A(n11549), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n18410) );
  NOR2_X1 U20496 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18407), .ZN(
        n18447) );
  INV_X2 U20497 ( .A(n19324), .ZN(n19531) );
  AOI21_X1 U20498 ( .B1(n19531), .B2(n18408), .A(n18607), .ZN(n18409) );
  OAI21_X1 U20499 ( .B1(n18444), .B2(n18620), .A(n18409), .ZN(n18441) );
  NOR2_X1 U20500 ( .A1(n18447), .A2(n18441), .ZN(n18427) );
  OAI22_X1 U20501 ( .A1(n18428), .A2(n18410), .B1(n18427), .B2(n11549), .ZN(
        n18411) );
  AOI211_X1 U20502 ( .C1(n21065), .C2(n18446), .A(n21622), .B(n18411), .ZN(
        n18425) );
  NOR2_X1 U20503 ( .A1(n21590), .A2(n21580), .ZN(n21645) );
  NAND2_X1 U20504 ( .A1(n21625), .A2(n21645), .ZN(n18412) );
  XOR2_X1 U20505 ( .A(n18412), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n21634) );
  INV_X1 U20506 ( .A(n21634), .ZN(n18423) );
  NAND2_X1 U20507 ( .A1(n18414), .A2(n18413), .ZN(n18435) );
  NAND2_X1 U20508 ( .A1(n21615), .A2(n18415), .ZN(n18420) );
  NOR2_X1 U20509 ( .A1(n21606), .A2(n18416), .ZN(n18417) );
  NAND2_X1 U20510 ( .A1(n18418), .A2(n18417), .ZN(n21641) );
  INV_X1 U20511 ( .A(n21625), .ZN(n18419) );
  OAI22_X1 U20512 ( .A1(n18435), .A2(n18420), .B1(n21641), .B2(n18419), .ZN(
        n18422) );
  AOI22_X1 U20513 ( .A1(n18423), .A2(n18549), .B1(n21629), .B2(n18535), .ZN(
        n18424) );
  OAI211_X1 U20514 ( .C1(n21628), .C2(n18484), .A(n18425), .B(n18424), .ZN(
        P3_U2799) );
  OAI22_X1 U20515 ( .A1(n18415), .A2(n21641), .B1(n18435), .B2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18426) );
  XNOR2_X1 U20516 ( .A(n18426), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n21621) );
  XOR2_X1 U20517 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n18443), .Z(
        n21077) );
  NAND2_X1 U20518 ( .A1(n21769), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21620) );
  OAI221_X1 U20519 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18428), .C1(
        n11550), .C2(n18427), .A(n21620), .ZN(n18433) );
  NOR2_X1 U20520 ( .A1(n21590), .A2(n18415), .ZN(n21612) );
  INV_X1 U20521 ( .A(n21612), .ZN(n21602) );
  NAND2_X1 U20522 ( .A1(n21559), .A2(n21612), .ZN(n21604) );
  AOI21_X1 U20523 ( .B1(n18430), .B2(n21612), .A(n18484), .ZN(n18440) );
  AOI21_X1 U20524 ( .B1(n18549), .B2(n21604), .A(n18440), .ZN(n18438) );
  INV_X1 U20525 ( .A(n18438), .ZN(n18431) );
  AOI211_X1 U20526 ( .C1(n18446), .C2(n21077), .A(n18433), .B(n18432), .ZN(
        n18434) );
  OAI21_X1 U20527 ( .B1(n21621), .B2(n18508), .A(n18434), .ZN(P3_U2800) );
  AOI21_X1 U20528 ( .B1(n21645), .B2(n18549), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18437) );
  NAND2_X1 U20529 ( .A1(n18435), .A2(n21641), .ZN(n18436) );
  XNOR2_X1 U20530 ( .A(n18436), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21610) );
  OAI22_X1 U20531 ( .A1(n18438), .A2(n18437), .B1(n21610), .B2(n18508), .ZN(
        n18439) );
  AOI21_X1 U20532 ( .B1(n21646), .B2(n18440), .A(n18439), .ZN(n18450) );
  NAND2_X1 U20533 ( .A1(n21769), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n21608) );
  OAI221_X1 U20534 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18442), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19531), .A(n18441), .ZN(
        n18449) );
  OAI21_X1 U20535 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18444), .A(
        n11551), .ZN(n21060) );
  INV_X1 U20536 ( .A(n21060), .ZN(n18445) );
  OAI21_X1 U20537 ( .B1(n18447), .B2(n18446), .A(n18445), .ZN(n18448) );
  NAND4_X1 U20538 ( .A1(n18450), .A2(n21608), .A3(n18449), .A4(n18448), .ZN(
        P3_U2801) );
  NAND2_X1 U20539 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18458), .ZN(
        n21718) );
  OAI22_X1 U20540 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18452), .B1(
        n20671), .B2(n18451), .ZN(n20907) );
  INV_X1 U20541 ( .A(n20907), .ZN(n18463) );
  AOI21_X1 U20542 ( .B1(n18453), .B2(n19531), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18455) );
  NAND2_X1 U20543 ( .A1(n18279), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21716) );
  OAI21_X1 U20544 ( .B1(n18455), .B2(n18454), .A(n21716), .ZN(n18462) );
  OAI21_X1 U20545 ( .B1(n18457), .B2(n18458), .A(n18456), .ZN(n21714) );
  INV_X1 U20546 ( .A(n21714), .ZN(n18460) );
  OAI22_X1 U20547 ( .A1(n18460), .A2(n18508), .B1(n18459), .B2(n18458), .ZN(
        n18461) );
  AOI211_X1 U20548 ( .C1(n18463), .C2(n18613), .A(n18462), .B(n18461), .ZN(
        n18464) );
  OAI21_X1 U20549 ( .B1(n18465), .B2(n21718), .A(n18464), .ZN(P3_U2813) );
  NAND3_X1 U20550 ( .A1(n11539), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n19531), .ZN(n18483) );
  OAI21_X1 U20551 ( .B1(n18466), .B2(n18483), .A(n18470), .ZN(n18467) );
  INV_X1 U20552 ( .A(n18467), .ZN(n18480) );
  INV_X1 U20553 ( .A(n20835), .ZN(n18469) );
  AOI21_X1 U20554 ( .B1(n18470), .B2(n18469), .A(n18468), .ZN(n20854) );
  AOI22_X1 U20555 ( .A1(n21769), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n20854), 
        .B2(n18613), .ZN(n18478) );
  NAND2_X1 U20556 ( .A1(n18472), .A2(n18471), .ZN(n18473) );
  XNOR2_X1 U20557 ( .A(n18473), .B(n21516), .ZN(n21499) );
  OAI21_X1 U20558 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18474), .A(
        n21525), .ZN(n21511) );
  OAI21_X1 U20559 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18475), .A(
        n21520), .ZN(n21510) );
  OAI22_X1 U20560 ( .A1(n18484), .A2(n21511), .B1(n18624), .B2(n21510), .ZN(
        n18476) );
  AOI21_X1 U20561 ( .B1(n18535), .B2(n21499), .A(n18476), .ZN(n18477) );
  OAI211_X1 U20562 ( .C1(n18480), .C2(n18479), .A(n18478), .B(n18477), .ZN(
        P3_U2816) );
  NAND2_X1 U20563 ( .A1(n11539), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18499) );
  AOI21_X1 U20564 ( .B1(n20826), .B2(n18499), .A(n18481), .ZN(n20808) );
  NOR2_X1 U20565 ( .A1(n18607), .A2(n18582), .ZN(n18556) );
  OAI22_X1 U20566 ( .A1(n18556), .A2(n20826), .B1(n18497), .B2(n19324), .ZN(
        n18482) );
  AOI22_X1 U20567 ( .A1(n20808), .A2(n18613), .B1(n18483), .B2(n18482), .ZN(
        n18489) );
  OAI22_X1 U20568 ( .A1(n21701), .A2(n18484), .B1(n18624), .B2(n21472), .ZN(
        n18520) );
  OAI21_X1 U20569 ( .B1(n18509), .B2(n21475), .A(n18485), .ZN(n18486) );
  XNOR2_X1 U20570 ( .A(n18486), .B(n21484), .ZN(n21481) );
  AOI22_X1 U20571 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18520), .B1(
        n18535), .B2(n21481), .ZN(n18488) );
  NAND2_X1 U20572 ( .A1(n21769), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n21482) );
  NOR2_X1 U20573 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21475), .ZN(
        n21480) );
  OAI221_X1 U20574 ( .B1(n21480), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), 
        .C1(n21480), .C2(n21475), .A(n18521), .ZN(n18487) );
  NAND4_X1 U20575 ( .A1(n18489), .A2(n18488), .A3(n21482), .A4(n18487), .ZN(
        P3_U2819) );
  NAND2_X1 U20576 ( .A1(n18490), .A2(n21755), .ZN(n18510) );
  INV_X1 U20577 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21762) );
  INV_X1 U20578 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18491) );
  OAI221_X1 U20579 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18510), .C1(
        n21762), .C2(n18509), .A(n18491), .ZN(n18496) );
  OAI21_X1 U20580 ( .B1(n18492), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18509), .ZN(n18493) );
  OAI211_X1 U20581 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18494), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18493), .ZN(n18495) );
  NAND2_X1 U20582 ( .A1(n18496), .A2(n18495), .ZN(n21751) );
  INV_X1 U20583 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20795) );
  NOR2_X1 U20584 ( .A1(n11173), .A2(n20795), .ZN(n18503) );
  NOR2_X1 U20585 ( .A1(n18497), .A2(n19324), .ZN(n18501) );
  INV_X1 U20586 ( .A(n18556), .ZN(n18614) );
  NOR2_X1 U20587 ( .A1(n18557), .A2(n19324), .ZN(n18555) );
  NAND2_X1 U20588 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18555), .ZN(
        n18542) );
  NOR2_X1 U20589 ( .A1(n18498), .A2(n18542), .ZN(n18515) );
  AOI21_X1 U20590 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18614), .A(
        n18515), .ZN(n18500) );
  INV_X1 U20591 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20778) );
  NAND2_X1 U20592 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18540), .ZN(
        n20767) );
  NOR2_X1 U20593 ( .A1(n20671), .A2(n20767), .ZN(n18541) );
  NAND2_X1 U20594 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18541), .ZN(
        n20776) );
  NOR2_X1 U20595 ( .A1(n20778), .A2(n20776), .ZN(n20791) );
  OAI21_X1 U20596 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20791), .A(
        n18499), .ZN(n20792) );
  OAI22_X1 U20597 ( .A1(n18501), .A2(n18500), .B1(n18605), .B2(n20792), .ZN(
        n18502) );
  AOI211_X1 U20598 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n18520), .A(
        n18503), .B(n18502), .ZN(n18507) );
  INV_X1 U20599 ( .A(n18504), .ZN(n18505) );
  NAND3_X1 U20600 ( .A1(n21475), .A2(n18505), .A3(n18521), .ZN(n18506) );
  OAI211_X1 U20601 ( .C1(n21751), .C2(n18508), .A(n18507), .B(n18506), .ZN(
        P3_U2820) );
  NAND2_X1 U20602 ( .A1(n18510), .A2(n18509), .ZN(n18511) );
  XNOR2_X1 U20603 ( .A(n18511), .B(n21762), .ZN(n21764) );
  INV_X1 U20604 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21767) );
  NOR2_X1 U20605 ( .A1(n11173), .A2(n21767), .ZN(n18517) );
  INV_X1 U20606 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18530) );
  INV_X1 U20607 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20756) );
  NOR2_X1 U20608 ( .A1(n18530), .A2(n20756), .ZN(n18529) );
  INV_X1 U20609 ( .A(n18542), .ZN(n18512) );
  AOI22_X1 U20610 ( .A1(n18529), .A2(n18512), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18614), .ZN(n18514) );
  AOI21_X1 U20611 ( .B1(n20778), .B2(n20776), .A(n20791), .ZN(n18513) );
  INV_X1 U20612 ( .A(n18513), .ZN(n20779) );
  OAI22_X1 U20613 ( .A1(n18515), .A2(n18514), .B1(n18605), .B2(n20779), .ZN(
        n18516) );
  AOI211_X1 U20614 ( .C1(n18535), .C2(n21764), .A(n18517), .B(n18516), .ZN(
        n18518) );
  INV_X1 U20615 ( .A(n18518), .ZN(n18519) );
  AOI221_X1 U20616 ( .B1(n21762), .B2(n18521), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18520), .A(n18519), .ZN(
        n18522) );
  INV_X1 U20617 ( .A(n18522), .ZN(P3_U2821) );
  OAI21_X1 U20618 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18524), .A(
        n18523), .ZN(n21467) );
  OAI21_X1 U20619 ( .B1(n18527), .B2(n18526), .A(n18525), .ZN(n21462) );
  INV_X1 U20620 ( .A(n21462), .ZN(n18534) );
  OAI21_X1 U20621 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18541), .A(
        n20776), .ZN(n20769) );
  OAI21_X1 U20622 ( .B1(n18540), .B2(n18528), .A(n18619), .ZN(n18548) );
  AOI211_X1 U20623 ( .C1(n18530), .C2(n20767), .A(n18529), .B(n19324), .ZN(
        n18531) );
  AOI21_X1 U20624 ( .B1(n18548), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n18531), .ZN(n18532) );
  NAND2_X1 U20625 ( .A1(n21769), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n21465) );
  OAI211_X1 U20626 ( .C1(n18605), .C2(n20769), .A(n18532), .B(n21465), .ZN(
        n18533) );
  AOI221_X1 U20627 ( .B1(n18536), .B2(n21462), .C1(n18535), .C2(n18534), .A(
        n18533), .ZN(n18537) );
  OAI21_X1 U20628 ( .B1(n18624), .B2(n21467), .A(n18537), .ZN(P3_U2822) );
  OAI21_X1 U20629 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18539), .A(
        n18538), .ZN(n21455) );
  NAND2_X1 U20630 ( .A1(n18540), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20739) );
  AOI21_X1 U20631 ( .B1(n20756), .B2(n20739), .A(n18541), .ZN(n20751) );
  INV_X1 U20632 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n21442) );
  OAI22_X1 U20633 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18542), .B1(
        n11173), .B2(n21442), .ZN(n18543) );
  AOI21_X1 U20634 ( .B1(n20751), .B2(n18613), .A(n18543), .ZN(n18551) );
  AOI21_X1 U20635 ( .B1(n18546), .B2(n18545), .A(n18544), .ZN(n18547) );
  XNOR2_X1 U20636 ( .A(n18547), .B(n21456), .ZN(n21452) );
  AOI22_X1 U20637 ( .A1(n18549), .A2(n21452), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18548), .ZN(n18550) );
  OAI211_X1 U20638 ( .C1(n18623), .C2(n21455), .A(n18551), .B(n18550), .ZN(
        P3_U2823) );
  OAI21_X1 U20639 ( .B1(n18554), .B2(n18553), .A(n18552), .ZN(n21434) );
  AOI22_X1 U20640 ( .A1(n21769), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18555), 
        .B2(n20742), .ZN(n18562) );
  NOR2_X1 U20641 ( .A1(n18556), .A2(n18555), .ZN(n18570) );
  NOR2_X1 U20642 ( .A1(n18557), .A2(n20671), .ZN(n18565) );
  OAI21_X1 U20643 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18565), .A(
        n20739), .ZN(n20744) );
  OAI21_X1 U20644 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18559), .A(
        n18558), .ZN(n21435) );
  OAI22_X1 U20645 ( .A1(n18605), .A2(n20744), .B1(n18624), .B2(n21435), .ZN(
        n18560) );
  AOI21_X1 U20646 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18570), .A(
        n18560), .ZN(n18561) );
  OAI211_X1 U20647 ( .C1(n18623), .C2(n21434), .A(n18562), .B(n18561), .ZN(
        P3_U2824) );
  OAI21_X1 U20648 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18564), .A(
        n18563), .ZN(n21431) );
  INV_X1 U20649 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20737) );
  NAND2_X1 U20650 ( .A1(n20717), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18573) );
  AOI21_X1 U20651 ( .B1(n20737), .B2(n18573), .A(n18565), .ZN(n20728) );
  INV_X1 U20652 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20724) );
  OAI21_X1 U20653 ( .B1(n18568), .B2(n18567), .A(n18566), .ZN(n21425) );
  OAI22_X1 U20654 ( .A1(n11173), .A2(n20724), .B1(n18624), .B2(n21425), .ZN(
        n18569) );
  AOI21_X1 U20655 ( .B1(n20728), .B2(n18613), .A(n18569), .ZN(n18572) );
  OAI221_X1 U20656 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20717), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18619), .A(n18570), .ZN(n18571) );
  OAI211_X1 U20657 ( .C1(n18623), .C2(n21431), .A(n18572), .B(n18571), .ZN(
        P3_U2825) );
  NOR2_X1 U20658 ( .A1(n18581), .A2(n20671), .ZN(n18590) );
  OAI21_X1 U20659 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18590), .A(
        n18573), .ZN(n20718) );
  OAI21_X1 U20660 ( .B1(n18576), .B2(n18575), .A(n18574), .ZN(n21413) );
  NAND2_X1 U20661 ( .A1(n19531), .A2(n18583), .ZN(n18577) );
  OAI22_X1 U20662 ( .A1(n18624), .A2(n21413), .B1(n18581), .B2(n18577), .ZN(
        n18585) );
  OAI21_X1 U20663 ( .B1(n18580), .B2(n18579), .A(n18578), .ZN(n21412) );
  AOI21_X1 U20664 ( .B1(n18582), .B2(n18581), .A(n18607), .ZN(n18594) );
  OAI22_X1 U20665 ( .A1(n18623), .A2(n21412), .B1(n18583), .B2(n18594), .ZN(
        n18584) );
  AOI211_X1 U20666 ( .C1(n18279), .C2(P3_REIP_REG_4__SCAN_IN), .A(n18585), .B(
        n18584), .ZN(n18586) );
  OAI21_X1 U20667 ( .B1(n18605), .B2(n20718), .A(n18586), .ZN(P3_U2826) );
  OAI21_X1 U20668 ( .B1(n18589), .B2(n18588), .A(n18587), .ZN(n21407) );
  INV_X1 U20669 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20709) );
  NAND2_X1 U20670 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18601) );
  AOI21_X1 U20671 ( .B1(n20709), .B2(n18601), .A(n18590), .ZN(n20699) );
  AOI21_X1 U20672 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18619), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18595) );
  OAI21_X1 U20673 ( .B1(n18593), .B2(n18592), .A(n18591), .ZN(n21406) );
  OAI22_X1 U20674 ( .A1(n18595), .A2(n18594), .B1(n18623), .B2(n21406), .ZN(
        n18596) );
  AOI21_X1 U20675 ( .B1(n20699), .B2(n18613), .A(n18596), .ZN(n18597) );
  NAND2_X1 U20676 ( .A1(n21769), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21409) );
  OAI211_X1 U20677 ( .C1(n18624), .C2(n21407), .A(n18597), .B(n21409), .ZN(
        P3_U2827) );
  OAI21_X1 U20678 ( .B1(n18600), .B2(n18599), .A(n18598), .ZN(n21393) );
  INV_X1 U20679 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20691) );
  OAI21_X1 U20680 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n18601), .ZN(n20694) );
  OAI21_X1 U20681 ( .B1(n18604), .B2(n18603), .A(n18602), .ZN(n21394) );
  OAI22_X1 U20682 ( .A1(n18605), .A2(n20694), .B1(n18624), .B2(n21394), .ZN(
        n18606) );
  AOI221_X1 U20683 ( .B1(n18607), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19531), .C2(n20691), .A(n18606), .ZN(n18608) );
  NAND2_X1 U20684 ( .A1(n21769), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21397) );
  OAI211_X1 U20685 ( .C1(n18623), .C2(n21393), .A(n18608), .B(n21397), .ZN(
        P3_U2828) );
  OAI21_X1 U20686 ( .B1(n18618), .B2(n18611), .A(n18609), .ZN(n21382) );
  AOI21_X1 U20687 ( .B1(n18611), .B2(n18616), .A(n18610), .ZN(n21383) );
  INV_X1 U20688 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20668) );
  OAI22_X1 U20689 ( .A1(n21383), .A2(n18624), .B1(n11173), .B2(n20668), .ZN(
        n18612) );
  AOI221_X1 U20690 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18614), .C1(
        n20671), .C2(n18613), .A(n18612), .ZN(n18615) );
  OAI21_X1 U20691 ( .B1(n18623), .B2(n21382), .A(n18615), .ZN(P3_U2829) );
  INV_X1 U20692 ( .A(n18616), .ZN(n18617) );
  NOR2_X1 U20693 ( .A1(n18618), .A2(n18617), .ZN(n21378) );
  INV_X1 U20694 ( .A(n21378), .ZN(n21377) );
  NAND3_X1 U20695 ( .A1(n20664), .A2(n18620), .A3(n18619), .ZN(n18621) );
  AOI22_X1 U20696 ( .A1(n18279), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18621), .ZN(n18622) );
  OAI221_X1 U20697 ( .B1(n21378), .B2(n18624), .C1(n21377), .C2(n18623), .A(
        n18622), .ZN(P3_U2830) );
  NOR2_X1 U20698 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19201), .ZN(
        n19240) );
  INV_X1 U20699 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21773) );
  NAND2_X1 U20700 ( .A1(n21791), .A2(n21773), .ZN(n19267) );
  INV_X1 U20701 ( .A(n19267), .ZN(n19269) );
  INV_X1 U20702 ( .A(n19241), .ZN(n19246) );
  NOR2_X1 U20703 ( .A1(n19269), .A2(n19246), .ZN(n18625) );
  NAND2_X1 U20704 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19203) );
  AOI22_X1 U20705 ( .A1(n19240), .A2(n18626), .B1(n18625), .B2(n19203), .ZN(
        n18628) );
  OAI22_X1 U20706 ( .A1(n18629), .A2(n18628), .B1(n18627), .B2(n21773), .ZN(
        P3_U2866) );
  NOR4_X1 U20707 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18633) );
  NOR4_X1 U20708 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18632) );
  NOR4_X1 U20709 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18631) );
  NOR4_X1 U20710 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18630) );
  NAND4_X1 U20711 ( .A1(n18633), .A2(n18632), .A3(n18631), .A4(n18630), .ZN(
        n18639) );
  NOR4_X1 U20712 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18637) );
  AOI211_X1 U20713 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18636) );
  NOR4_X1 U20714 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18635) );
  NOR4_X1 U20715 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18634) );
  NAND4_X1 U20716 ( .A1(n18637), .A2(n18636), .A3(n18635), .A4(n18634), .ZN(
        n18638) );
  NOR2_X1 U20717 ( .A1(n18639), .A2(n18638), .ZN(n18645) );
  NAND2_X1 U20718 ( .A1(n18645), .A2(n20668), .ZN(n18651) );
  INV_X1 U20719 ( .A(n18651), .ZN(n18647) );
  INV_X1 U20720 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n21373) );
  INV_X1 U20721 ( .A(n18645), .ZN(n18648) );
  INV_X1 U20722 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18640) );
  AOI22_X1 U20723 ( .A1(n18647), .A2(n21373), .B1(n18648), .B2(n18640), .ZN(
        P3_U3293) );
  NOR2_X1 U20724 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18644) );
  AOI211_X1 U20725 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(n21373), .A(n18644), 
        .B(n18651), .ZN(n18643) );
  NAND3_X1 U20726 ( .A1(n18645), .A2(P3_REIP_REG_1__SCAN_IN), .A3(n21373), 
        .ZN(n18641) );
  OAI21_X1 U20727 ( .B1(n18645), .B2(P3_BYTEENABLE_REG_2__SCAN_IN), .A(n18641), 
        .ZN(n18642) );
  NOR2_X1 U20728 ( .A1(n18643), .A2(n18642), .ZN(P3_U3292) );
  NOR2_X1 U20729 ( .A1(n18645), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18646)
         );
  NAND3_X1 U20730 ( .A1(n18645), .A2(n18644), .A3(n21373), .ZN(n18650) );
  OAI21_X1 U20731 ( .B1(n18647), .B2(n18646), .A(n18650), .ZN(P3_U2638) );
  NAND2_X1 U20732 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18648), .ZN(n18649) );
  OAI211_X1 U20733 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(n18651), .A(n18650), 
        .B(n18649), .ZN(P3_U2639) );
  INV_X1 U20734 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18714) );
  AOI22_X1 U20735 ( .A1(n22179), .A2(n18652), .B1(n18714), .B2(n22225), .ZN(
        P3_U3297) );
  INV_X1 U20736 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18653) );
  AOI22_X1 U20737 ( .A1(n22179), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18653), 
        .B2(n22225), .ZN(P3_U3294) );
  INV_X1 U20738 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22216) );
  AOI21_X1 U20739 ( .B1(n22214), .B2(n22216), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18654) );
  AOI22_X1 U20740 ( .A1(n22179), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18654), 
        .B2(n22225), .ZN(P3_U2635) );
  INV_X1 U20741 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21281) );
  AOI22_X1 U20742 ( .A1(n21770), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18655) );
  OAI21_X1 U20743 ( .B1(n21281), .B2(n18671), .A(n18655), .ZN(P3_U2767) );
  INV_X1 U20744 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20637) );
  AOI22_X1 U20745 ( .A1(n21770), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18656) );
  OAI21_X1 U20746 ( .B1(n20637), .B2(n18671), .A(n18656), .ZN(P3_U2766) );
  INV_X1 U20747 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20639) );
  AOI22_X1 U20748 ( .A1(n21770), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18657) );
  OAI21_X1 U20749 ( .B1(n20639), .B2(n18671), .A(n18657), .ZN(P3_U2765) );
  INV_X1 U20750 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n21149) );
  AOI22_X1 U20751 ( .A1(n21770), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18658) );
  OAI21_X1 U20752 ( .B1(n21149), .B2(n18671), .A(n18658), .ZN(P3_U2764) );
  INV_X1 U20753 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21145) );
  AOI22_X1 U20754 ( .A1(n21770), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18659) );
  OAI21_X1 U20755 ( .B1(n21145), .B2(n18671), .A(n18659), .ZN(P3_U2763) );
  INV_X1 U20756 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20643) );
  AOI22_X1 U20757 ( .A1(n21770), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18660) );
  OAI21_X1 U20758 ( .B1(n20643), .B2(n18671), .A(n18660), .ZN(P3_U2762) );
  INV_X1 U20759 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20645) );
  AOI22_X1 U20760 ( .A1(n21770), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18661) );
  OAI21_X1 U20761 ( .B1(n20645), .B2(n18671), .A(n18661), .ZN(P3_U2761) );
  INV_X1 U20762 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n21129) );
  AOI22_X1 U20763 ( .A1(n21770), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18662) );
  OAI21_X1 U20764 ( .B1(n21129), .B2(n18671), .A(n18662), .ZN(P3_U2760) );
  INV_X1 U20765 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21267) );
  AOI22_X1 U20766 ( .A1(n21770), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18663) );
  OAI21_X1 U20767 ( .B1(n21267), .B2(n18671), .A(n18663), .ZN(P3_U2759) );
  INV_X1 U20768 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21156) );
  AOI22_X1 U20769 ( .A1(n18681), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18664) );
  OAI21_X1 U20770 ( .B1(n21156), .B2(n18671), .A(n18664), .ZN(P3_U2758) );
  INV_X1 U20771 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U20772 ( .A1(n18681), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18665) );
  OAI21_X1 U20773 ( .B1(n20650), .B2(n18671), .A(n18665), .ZN(P3_U2757) );
  INV_X1 U20774 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21112) );
  AOI22_X1 U20775 ( .A1(n18681), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18666) );
  OAI21_X1 U20776 ( .B1(n21112), .B2(n18671), .A(n18666), .ZN(P3_U2756) );
  INV_X1 U20777 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20654) );
  AOI22_X1 U20778 ( .A1(n18681), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18667) );
  OAI21_X1 U20779 ( .B1(n20654), .B2(n18671), .A(n18667), .ZN(P3_U2755) );
  INV_X1 U20780 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20656) );
  AOI22_X1 U20781 ( .A1(n18681), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18668) );
  OAI21_X1 U20782 ( .B1(n20656), .B2(n18671), .A(n18668), .ZN(P3_U2754) );
  INV_X1 U20783 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21253) );
  AOI22_X1 U20784 ( .A1(n18681), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18669) );
  OAI21_X1 U20785 ( .B1(n21253), .B2(n18671), .A(n18669), .ZN(P3_U2753) );
  INV_X1 U20786 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21257) );
  AOI22_X1 U20787 ( .A1(n18681), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18670) );
  OAI21_X1 U20788 ( .B1(n21257), .B2(n18671), .A(n18670), .ZN(P3_U2752) );
  INV_X1 U20789 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20613) );
  NAND2_X1 U20790 ( .A1(n18672), .A2(n20666), .ZN(n18691) );
  AOI22_X1 U20791 ( .A1(n18681), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18673) );
  OAI21_X1 U20792 ( .B1(n20613), .B2(n18691), .A(n18673), .ZN(P3_U2751) );
  INV_X1 U20793 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21159) );
  AOI22_X1 U20794 ( .A1(n18681), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18674) );
  OAI21_X1 U20795 ( .B1(n21159), .B2(n18691), .A(n18674), .ZN(P3_U2750) );
  INV_X1 U20796 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20616) );
  AOI22_X1 U20797 ( .A1(n18681), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18675) );
  OAI21_X1 U20798 ( .B1(n20616), .B2(n18691), .A(n18675), .ZN(P3_U2749) );
  INV_X1 U20799 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21180) );
  AOI22_X1 U20800 ( .A1(n21770), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18676) );
  OAI21_X1 U20801 ( .B1(n21180), .B2(n18691), .A(n18676), .ZN(P3_U2748) );
  INV_X1 U20802 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21170) );
  AOI22_X1 U20803 ( .A1(n21770), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18677) );
  OAI21_X1 U20804 ( .B1(n21170), .B2(n18691), .A(n18677), .ZN(P3_U2747) );
  INV_X1 U20805 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21171) );
  AOI22_X1 U20806 ( .A1(n21770), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18678) );
  OAI21_X1 U20807 ( .B1(n21171), .B2(n18691), .A(n18678), .ZN(P3_U2746) );
  INV_X1 U20808 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n21195) );
  AOI22_X1 U20809 ( .A1(n21770), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18679) );
  OAI21_X1 U20810 ( .B1(n21195), .B2(n18691), .A(n18679), .ZN(P3_U2745) );
  INV_X1 U20811 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20623) );
  AOI22_X1 U20812 ( .A1(n21770), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18680) );
  OAI21_X1 U20813 ( .B1(n20623), .B2(n18691), .A(n18680), .ZN(P3_U2744) );
  AOI22_X1 U20814 ( .A1(n18681), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18682) );
  OAI21_X1 U20815 ( .B1(n11384), .B2(n18691), .A(n18682), .ZN(P3_U2743) );
  INV_X1 U20816 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20626) );
  AOI22_X1 U20817 ( .A1(n21770), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18683) );
  OAI21_X1 U20818 ( .B1(n20626), .B2(n18691), .A(n18683), .ZN(P3_U2742) );
  INV_X1 U20819 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21204) );
  AOI22_X1 U20820 ( .A1(n21770), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18684) );
  OAI21_X1 U20821 ( .B1(n21204), .B2(n18691), .A(n18684), .ZN(P3_U2741) );
  INV_X1 U20822 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20629) );
  AOI22_X1 U20823 ( .A1(n21770), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18685), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18686) );
  OAI21_X1 U20824 ( .B1(n20629), .B2(n18691), .A(n18686), .ZN(P3_U2740) );
  INV_X1 U20825 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n21220) );
  AOI22_X1 U20826 ( .A1(n21770), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18687) );
  OAI21_X1 U20827 ( .B1(n21220), .B2(n18691), .A(n18687), .ZN(P3_U2739) );
  INV_X1 U20828 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20632) );
  AOI22_X1 U20829 ( .A1(n21770), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18688) );
  OAI21_X1 U20830 ( .B1(n20632), .B2(n18691), .A(n18688), .ZN(P3_U2738) );
  INV_X1 U20831 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20634) );
  AOI22_X1 U20832 ( .A1(n21770), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18689), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18690) );
  OAI21_X1 U20833 ( .B1(n20634), .B2(n18691), .A(n18690), .ZN(P3_U2737) );
  NOR2_X1 U20834 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18692), .ZN(n18693) );
  NOR2_X1 U20835 ( .A1(n22179), .A2(n18693), .ZN(P3_U2633) );
  NOR2_X1 U20836 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22225), .ZN(n18706) );
  AOI22_X1 U20837 ( .A1(n18706), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n22225), .ZN(n18694) );
  OAI21_X1 U20838 ( .B1(n18708), .B2(n20668), .A(n18694), .ZN(P3_U3032) );
  INV_X1 U20839 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20695) );
  AOI22_X1 U20840 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18709), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n22225), .ZN(n18695) );
  OAI21_X1 U20841 ( .B1(n20695), .B2(n18712), .A(n18695), .ZN(P3_U3033) );
  INV_X1 U20842 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n21418) );
  INV_X1 U20843 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20298) );
  OAI222_X1 U20844 ( .A1(n18712), .A2(n21418), .B1(n20298), .B2(n22179), .C1(
        n20695), .C2(n18708), .ZN(P3_U3034) );
  INV_X1 U20845 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20300) );
  OAI222_X1 U20846 ( .A1(n18712), .A2(n20724), .B1(n20300), .B2(n22179), .C1(
        n21418), .C2(n18711), .ZN(P3_U3035) );
  AOI22_X1 U20847 ( .A1(n18706), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n22225), .ZN(n18696) );
  OAI21_X1 U20848 ( .B1(n18708), .B2(n20724), .A(n18696), .ZN(P3_U3036) );
  AOI22_X1 U20849 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18709), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n22225), .ZN(n18697) );
  OAI21_X1 U20850 ( .B1(n21442), .B2(n18712), .A(n18697), .ZN(P3_U3037) );
  AOI22_X1 U20851 ( .A1(n18706), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n22225), .ZN(n18698) );
  OAI21_X1 U20852 ( .B1(n18708), .B2(n21442), .A(n18698), .ZN(P3_U3038) );
  AOI22_X1 U20853 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18709), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n22225), .ZN(n18699) );
  OAI21_X1 U20854 ( .B1(n21767), .B2(n18712), .A(n18699), .ZN(P3_U3039) );
  INV_X1 U20855 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20310) );
  OAI222_X1 U20856 ( .A1(n18712), .A2(n20795), .B1(n20310), .B2(n22179), .C1(
        n21767), .C2(n18708), .ZN(P3_U3040) );
  INV_X1 U20857 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20824) );
  INV_X1 U20858 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20312) );
  OAI222_X1 U20859 ( .A1(n18712), .A2(n20824), .B1(n20312), .B2(n22179), .C1(
        n20795), .C2(n18711), .ZN(P3_U3041) );
  INV_X1 U20860 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20314) );
  OAI222_X1 U20861 ( .A1(n18712), .A2(n20848), .B1(n20314), .B2(n22179), .C1(
        n20824), .C2(n18711), .ZN(P3_U3042) );
  INV_X1 U20862 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20849) );
  INV_X1 U20863 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20316) );
  OAI222_X1 U20864 ( .A1(n18712), .A2(n20849), .B1(n20316), .B2(n22179), .C1(
        n20848), .C2(n18711), .ZN(P3_U3043) );
  AOI22_X1 U20865 ( .A1(n18706), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n22225), .ZN(n18700) );
  OAI21_X1 U20866 ( .B1(n18708), .B2(n20849), .A(n18700), .ZN(P3_U3044) );
  AOI22_X1 U20867 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18709), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n22225), .ZN(n18701) );
  OAI21_X1 U20868 ( .B1(n20878), .B2(n18712), .A(n18701), .ZN(P3_U3045) );
  AOI22_X1 U20869 ( .A1(n18706), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n22225), .ZN(n18702) );
  OAI21_X1 U20870 ( .B1(n18708), .B2(n20878), .A(n18702), .ZN(P3_U3046) );
  INV_X1 U20871 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20910) );
  AOI22_X1 U20872 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18709), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n22225), .ZN(n18703) );
  OAI21_X1 U20873 ( .B1(n20910), .B2(n18712), .A(n18703), .ZN(P3_U3047) );
  INV_X1 U20874 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20326) );
  INV_X1 U20875 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20923) );
  OAI222_X1 U20876 ( .A1(n20910), .A2(n18708), .B1(n20326), .B2(n22179), .C1(
        n20923), .C2(n18712), .ZN(P3_U3048) );
  INV_X1 U20877 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20328) );
  OAI222_X1 U20878 ( .A1(n20923), .A2(n18708), .B1(n20328), .B2(n22179), .C1(
        n20934), .C2(n18712), .ZN(P3_U3049) );
  INV_X1 U20879 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20936) );
  INV_X1 U20880 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20330) );
  OAI222_X1 U20881 ( .A1(n18712), .A2(n20936), .B1(n20330), .B2(n22179), .C1(
        n20934), .C2(n18711), .ZN(P3_U3050) );
  INV_X1 U20882 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20332) );
  OAI222_X1 U20883 ( .A1(n18712), .A2(n20952), .B1(n20332), .B2(n22179), .C1(
        n20936), .C2(n18711), .ZN(P3_U3051) );
  INV_X1 U20884 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20334) );
  OAI222_X1 U20885 ( .A1(n18712), .A2(n18704), .B1(n20334), .B2(n22179), .C1(
        n20952), .C2(n18711), .ZN(P3_U3052) );
  INV_X1 U20886 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20336) );
  OAI222_X1 U20887 ( .A1(n18712), .A2(n18705), .B1(n20336), .B2(n22179), .C1(
        n18704), .C2(n18711), .ZN(P3_U3053) );
  INV_X1 U20888 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20338) );
  OAI222_X1 U20889 ( .A1(n18712), .A2(n21000), .B1(n20338), .B2(n22179), .C1(
        n18705), .C2(n18711), .ZN(P3_U3054) );
  INV_X1 U20890 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20340) );
  OAI222_X1 U20891 ( .A1(n18712), .A2(n21001), .B1(n20340), .B2(n22179), .C1(
        n21000), .C2(n18711), .ZN(P3_U3055) );
  INV_X1 U20892 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21025) );
  INV_X1 U20893 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20343) );
  OAI222_X1 U20894 ( .A1(n18712), .A2(n21025), .B1(n20343), .B2(n22179), .C1(
        n21001), .C2(n18708), .ZN(P3_U3056) );
  INV_X1 U20895 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20345) );
  OAI222_X1 U20896 ( .A1(n21025), .A2(n18708), .B1(n20345), .B2(n22179), .C1(
        n21026), .C2(n18712), .ZN(P3_U3057) );
  AOI22_X1 U20897 ( .A1(n18706), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n22225), .ZN(n18707) );
  OAI21_X1 U20898 ( .B1(n18708), .B2(n21026), .A(n18707), .ZN(P3_U3058) );
  INV_X1 U20899 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21063) );
  AOI22_X1 U20900 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18709), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n22225), .ZN(n18710) );
  OAI21_X1 U20901 ( .B1(n21063), .B2(n18712), .A(n18710), .ZN(P3_U3059) );
  INV_X1 U20902 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21079) );
  INV_X1 U20903 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20351) );
  OAI222_X1 U20904 ( .A1(n18712), .A2(n21079), .B1(n20351), .B2(n22179), .C1(
        n21063), .C2(n18711), .ZN(P3_U3060) );
  INV_X1 U20905 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20354) );
  OAI222_X1 U20906 ( .A1(n18712), .A2(n21081), .B1(n20354), .B2(n22179), .C1(
        n21079), .C2(n18711), .ZN(P3_U3061) );
  OAI22_X1 U20907 ( .A1(n22225), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n22179), .ZN(n18713) );
  INV_X1 U20908 ( .A(n18713), .ZN(P3_U3277) );
  MUX2_X1 U20909 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n22179), .Z(P3_U3276) );
  MUX2_X1 U20910 ( .A(P3_BE_N_REG_2__SCAN_IN), .B(P3_BYTEENABLE_REG_2__SCAN_IN), .S(n22179), .Z(P3_U3275) );
  MUX2_X1 U20911 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n22179), .Z(P3_U3274) );
  NOR4_X1 U20912 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18716)
         );
  NOR4_X1 U20913 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18714), .ZN(n18715) );
  INV_X2 U20914 ( .A(n19487), .ZN(U215) );
  NAND3_X1 U20915 ( .A1(n18716), .A2(n18715), .A3(U215), .ZN(U213) );
  INV_X1 U20916 ( .A(n18717), .ZN(n18719) );
  NAND4_X1 U20917 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n15635), .A4(n19164), .ZN(n18718) );
  OAI211_X1 U20918 ( .C1(n19160), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        n18728) );
  INV_X1 U20919 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22200) );
  AOI211_X1 U20920 ( .C1(n18722), .C2(P2_STATEBS16_REG_SCAN_IN), .A(n15635), 
        .B(n18721), .ZN(n18726) );
  NOR2_X1 U20921 ( .A1(n22197), .A2(n19734), .ZN(n18724) );
  INV_X1 U20922 ( .A(n18722), .ZN(n22207) );
  NAND4_X1 U20923 ( .A1(n20177), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n22207), 
        .A4(n19060), .ZN(n18723) );
  OAI21_X1 U20924 ( .B1(n18724), .B2(n19165), .A(n18723), .ZN(n18725) );
  OAI21_X1 U20925 ( .B1(n18726), .B2(n18725), .A(n18728), .ZN(n18727) );
  OAI21_X1 U20926 ( .B1(n18728), .B2(n22200), .A(n18727), .ZN(P2_U3610) );
  INV_X1 U20927 ( .A(n18729), .ZN(n19905) );
  OAI21_X1 U20928 ( .B1(n19036), .B2(n15510), .A(n18813), .ZN(n18732) );
  OAI22_X1 U20929 ( .A1(n19051), .A2(n18730), .B1(n13221), .B2(n19041), .ZN(
        n18731) );
  AOI211_X1 U20930 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n19013), .A(n18732), .B(
        n18731), .ZN(n18733) );
  OAI21_X1 U20931 ( .B1(n18734), .B2(n19037), .A(n18733), .ZN(n18735) );
  AOI21_X1 U20932 ( .B1(n19905), .B2(n18736), .A(n18735), .ZN(n18742) );
  AND2_X1 U20933 ( .A1(n11188), .A2(n18737), .ZN(n18739) );
  AOI21_X1 U20934 ( .B1(n18740), .B2(n18739), .A(n19154), .ZN(n18738) );
  OAI21_X1 U20935 ( .B1(n18740), .B2(n18739), .A(n18738), .ZN(n18741) );
  OAI211_X1 U20936 ( .C1(n18743), .C2(n19008), .A(n18742), .B(n18741), .ZN(
        P2_U2851) );
  OAI21_X1 U20937 ( .B1(n13105), .B2(n19041), .A(n18813), .ZN(n18747) );
  OAI22_X1 U20938 ( .A1(n19037), .A2(n18745), .B1(n18744), .B2(n19040), .ZN(
        n18746) );
  AOI211_X1 U20939 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19012), .A(
        n18747), .B(n18746), .ZN(n18754) );
  NAND2_X1 U20940 ( .A1(n11188), .A2(n18748), .ZN(n18749) );
  XNOR2_X1 U20941 ( .A(n18750), .B(n18749), .ZN(n18752) );
  AOI22_X1 U20942 ( .A1(n19003), .A2(n18752), .B1(n19045), .B2(n18751), .ZN(
        n18753) );
  OAI211_X1 U20943 ( .C1(n19051), .C2(n19863), .A(n18754), .B(n18753), .ZN(
        P2_U2849) );
  NOR2_X1 U20944 ( .A1(n18778), .A2(n18755), .ZN(n18756) );
  XOR2_X1 U20945 ( .A(n18757), .B(n18756), .Z(n18764) );
  AOI22_X1 U20946 ( .A1(n19009), .A2(n18758), .B1(n19013), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n18759) );
  OAI211_X1 U20947 ( .C1(n17160), .C2(n19041), .A(n18759), .B(n18813), .ZN(
        n18762) );
  OAI22_X1 U20948 ( .A1(n19051), .A2(n19663), .B1(n19008), .B2(n18760), .ZN(
        n18761) );
  AOI211_X1 U20949 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19012), .A(
        n18762), .B(n18761), .ZN(n18763) );
  OAI21_X1 U20950 ( .B1(n19154), .B2(n18764), .A(n18763), .ZN(P2_U2848) );
  AOI22_X1 U20951 ( .A1(n19013), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19012), .ZN(n18765) );
  OAI21_X1 U20952 ( .B1(n18766), .B2(n19037), .A(n18765), .ZN(n18767) );
  AOI211_X1 U20953 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19011), .A(n19139), .B(
        n18767), .ZN(n18776) );
  NAND2_X1 U20954 ( .A1(n17412), .A2(n18768), .ZN(n18769) );
  XNOR2_X1 U20955 ( .A(n18770), .B(n18769), .ZN(n18774) );
  AOI21_X1 U20956 ( .B1(n18773), .B2(n18772), .A(n18771), .ZN(n19657) );
  AOI22_X1 U20957 ( .A1(n19003), .A2(n18774), .B1(n19014), .B2(n19657), .ZN(
        n18775) );
  OAI211_X1 U20958 ( .C1(n19008), .C2(n19132), .A(n18776), .B(n18775), .ZN(
        P2_U2847) );
  NOR2_X1 U20959 ( .A1(n18778), .A2(n18777), .ZN(n18779) );
  XOR2_X1 U20960 ( .A(n18780), .B(n18779), .Z(n18787) );
  AOI22_X1 U20961 ( .A1(n18781), .A2(n19009), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19013), .ZN(n18782) );
  OAI211_X1 U20962 ( .C1(n17147), .C2(n19041), .A(n18782), .B(n18892), .ZN(
        n18785) );
  OAI22_X1 U20963 ( .A1(n19051), .A2(n19656), .B1(n19008), .B2(n18783), .ZN(
        n18784) );
  AOI211_X1 U20964 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19012), .A(
        n18785), .B(n18784), .ZN(n18786) );
  OAI21_X1 U20965 ( .B1(n19154), .B2(n18787), .A(n18786), .ZN(P2_U2846) );
  AOI22_X1 U20966 ( .A1(n19013), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19012), .ZN(n18788) );
  OAI21_X1 U20967 ( .B1(n18789), .B2(n19037), .A(n18788), .ZN(n18790) );
  AOI211_X1 U20968 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19011), .A(n19139), 
        .B(n18790), .ZN(n18799) );
  AOI21_X1 U20969 ( .B1(n18793), .B2(n18792), .A(n18791), .ZN(n19650) );
  NAND2_X1 U20970 ( .A1(n17412), .A2(n18794), .ZN(n18795) );
  XNOR2_X1 U20971 ( .A(n18796), .B(n18795), .ZN(n18797) );
  AOI22_X1 U20972 ( .A1(n19650), .A2(n19014), .B1(n19003), .B2(n18797), .ZN(
        n18798) );
  OAI211_X1 U20973 ( .C1(n18800), .C2(n19008), .A(n18799), .B(n18798), .ZN(
        P2_U2845) );
  OAI22_X1 U20974 ( .A1(n19040), .A2(n13475), .B1(n19036), .B2(n18801), .ZN(
        n18806) );
  INV_X1 U20975 ( .A(n19649), .ZN(n18802) );
  AOI22_X1 U20976 ( .A1(n18803), .A2(n19009), .B1(n18802), .B2(n19014), .ZN(
        n18804) );
  OAI211_X1 U20977 ( .C1(n13123), .C2(n19041), .A(n18804), .B(n18813), .ZN(
        n18805) );
  AOI211_X1 U20978 ( .C1(n18807), .C2(n19045), .A(n18806), .B(n18805), .ZN(
        n18810) );
  OAI211_X1 U20979 ( .C1(n18808), .C2(n18811), .A(n19048), .B(n18816), .ZN(
        n18809) );
  OAI211_X1 U20980 ( .C1(n18875), .C2(n18811), .A(n18810), .B(n18809), .ZN(
        P2_U2844) );
  AOI22_X1 U20981 ( .A1(n18812), .A2(n19009), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19013), .ZN(n18814) );
  OAI211_X1 U20982 ( .C1(n13301), .C2(n19041), .A(n18814), .B(n18813), .ZN(
        n18815) );
  AOI21_X1 U20983 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19012), .A(
        n18815), .ZN(n18822) );
  NAND2_X1 U20984 ( .A1(n17412), .A2(n18816), .ZN(n18817) );
  XNOR2_X1 U20985 ( .A(n18818), .B(n18817), .ZN(n18819) );
  AOI22_X1 U20986 ( .A1(n18820), .A2(n19014), .B1(n19003), .B2(n18819), .ZN(
        n18821) );
  OAI211_X1 U20987 ( .C1(n18823), .C2(n19008), .A(n18822), .B(n18821), .ZN(
        P2_U2843) );
  AOI22_X1 U20988 ( .A1(n19013), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19012), .ZN(n18824) );
  OAI21_X1 U20989 ( .B1(n18825), .B2(n19037), .A(n18824), .ZN(n18826) );
  AOI211_X1 U20990 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19011), .A(n19139), 
        .B(n18826), .ZN(n18837) );
  AND2_X1 U20991 ( .A1(n18828), .A2(n18827), .ZN(n18830) );
  OR2_X1 U20992 ( .A1(n18830), .A2(n18829), .ZN(n19639) );
  INV_X1 U20993 ( .A(n19639), .ZN(n19088) );
  INV_X1 U20994 ( .A(n18831), .ZN(n18846) );
  NAND2_X1 U20995 ( .A1(n18833), .A2(n18832), .ZN(n18845) );
  NAND2_X1 U20996 ( .A1(n11188), .A2(n18845), .ZN(n18834) );
  XNOR2_X1 U20997 ( .A(n18846), .B(n18834), .ZN(n18835) );
  AOI22_X1 U20998 ( .A1(n19088), .A2(n19014), .B1(n19003), .B2(n18835), .ZN(
        n18836) );
  OAI211_X1 U20999 ( .C1(n19090), .C2(n19008), .A(n18837), .B(n18836), .ZN(
        P2_U2841) );
  AOI22_X1 U21000 ( .A1(n19013), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19012), .ZN(n18838) );
  OAI211_X1 U21001 ( .C1(n18839), .C2(n19041), .A(n18838), .B(n18892), .ZN(
        n18843) );
  INV_X1 U21002 ( .A(n18840), .ZN(n18848) );
  OAI22_X1 U21003 ( .A1(n18841), .A2(n19037), .B1(n18848), .B2(n18875), .ZN(
        n18842) );
  AOI211_X1 U21004 ( .C1(n18844), .C2(n19045), .A(n18843), .B(n18842), .ZN(
        n18851) );
  NOR2_X1 U21005 ( .A1(n18846), .A2(n18845), .ZN(n18849) );
  NAND2_X1 U21006 ( .A1(n18849), .A2(n18848), .ZN(n18870) );
  NAND2_X1 U21007 ( .A1(n17412), .A2(n18870), .ZN(n18859) );
  INV_X1 U21008 ( .A(n18859), .ZN(n18847) );
  OAI211_X1 U21009 ( .C1(n18849), .C2(n18848), .A(n19003), .B(n18847), .ZN(
        n18850) );
  OAI211_X1 U21010 ( .C1(n19051), .C2(n19636), .A(n18851), .B(n18850), .ZN(
        P2_U2840) );
  OAI21_X1 U21011 ( .B1(n18852), .B2(n19036), .A(n18892), .ZN(n18853) );
  AOI21_X1 U21012 ( .B1(n19013), .B2(P2_EBX_REG_16__SCAN_IN), .A(n18853), .ZN(
        n18855) );
  NAND2_X1 U21013 ( .A1(n19011), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n18854) );
  OAI211_X1 U21014 ( .C1(n18856), .C2(n19037), .A(n18855), .B(n18854), .ZN(
        n18857) );
  INV_X1 U21015 ( .A(n18857), .ZN(n18863) );
  INV_X1 U21016 ( .A(n19122), .ZN(n18861) );
  INV_X1 U21017 ( .A(n18858), .ZN(n18871) );
  XNOR2_X1 U21018 ( .A(n18871), .B(n18859), .ZN(n18860) );
  AOI22_X1 U21019 ( .A1(n18861), .A2(n19045), .B1(n19003), .B2(n18860), .ZN(
        n18862) );
  OAI211_X1 U21020 ( .C1(n19120), .C2(n19051), .A(n18863), .B(n18862), .ZN(
        P2_U2839) );
  INV_X1 U21021 ( .A(n19102), .ZN(n18880) );
  OAI21_X1 U21022 ( .B1(n19036), .B2(n18864), .A(n18813), .ZN(n18865) );
  AOI21_X1 U21023 ( .B1(n19013), .B2(P2_EBX_REG_17__SCAN_IN), .A(n18865), .ZN(
        n18867) );
  NAND2_X1 U21024 ( .A1(n19011), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n18866) );
  OAI211_X1 U21025 ( .C1(n18868), .C2(n19037), .A(n18867), .B(n18866), .ZN(
        n18869) );
  INV_X1 U21026 ( .A(n18869), .ZN(n18879) );
  NOR2_X1 U21027 ( .A1(n18871), .A2(n18870), .ZN(n18873) );
  INV_X1 U21028 ( .A(n18872), .ZN(n18876) );
  NAND2_X1 U21029 ( .A1(n18873), .A2(n18876), .ZN(n18887) );
  OAI21_X1 U21030 ( .B1(n18876), .B2(n18873), .A(n19048), .ZN(n18874) );
  OAI21_X1 U21031 ( .B1(n18876), .B2(n18875), .A(n18874), .ZN(n18877) );
  AOI22_X1 U21032 ( .A1(n19104), .A2(n19014), .B1(n18887), .B2(n18877), .ZN(
        n18878) );
  OAI211_X1 U21033 ( .C1(n18880), .C2(n19008), .A(n18879), .B(n18878), .ZN(
        P2_U2838) );
  AOI22_X1 U21034 ( .A1(n18881), .A2(n19009), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19013), .ZN(n18882) );
  OAI211_X1 U21035 ( .C1(n13351), .C2(n19041), .A(n18882), .B(n18892), .ZN(
        n18886) );
  OAI22_X1 U21036 ( .A1(n18884), .A2(n19008), .B1(n18883), .B2(n19051), .ZN(
        n18885) );
  AOI211_X1 U21037 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19012), .A(
        n18886), .B(n18885), .ZN(n18890) );
  NAND2_X1 U21038 ( .A1(n18890), .A2(n18889), .ZN(P2_U2837) );
  AOI22_X1 U21039 ( .A1(n18891), .A2(n19009), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n19013), .ZN(n18893) );
  OAI211_X1 U21040 ( .C1(n18894), .C2(n19041), .A(n18893), .B(n18892), .ZN(
        n18895) );
  AOI21_X1 U21041 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19012), .A(
        n18895), .ZN(n18904) );
  AOI22_X1 U21042 ( .A1(n18897), .A2(n19045), .B1(n18896), .B2(n19014), .ZN(
        n18903) );
  INV_X1 U21043 ( .A(n18898), .ZN(n18901) );
  NAND2_X1 U21044 ( .A1(n18899), .A2(n11188), .ZN(n18900) );
  NAND2_X1 U21045 ( .A1(n18900), .A2(n18901), .ZN(n18911) );
  OAI211_X1 U21046 ( .C1(n18901), .C2(n18900), .A(n19003), .B(n18911), .ZN(
        n18902) );
  NAND3_X1 U21047 ( .A1(n18904), .A2(n18903), .A3(n18902), .ZN(P2_U2836) );
  OAI22_X1 U21048 ( .A1(n11513), .A2(n19036), .B1(n18905), .B2(n19041), .ZN(
        n18909) );
  INV_X1 U21049 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n18906) );
  OAI22_X1 U21050 ( .A1(n18907), .A2(n19037), .B1(n18906), .B2(n19040), .ZN(
        n18908) );
  AOI211_X1 U21051 ( .C1(n18910), .C2(n19014), .A(n18909), .B(n18908), .ZN(
        n18915) );
  NAND2_X1 U21052 ( .A1(n18912), .A2(n18913), .ZN(n18925) );
  OAI211_X1 U21053 ( .C1(n18913), .C2(n18912), .A(n19003), .B(n18925), .ZN(
        n18914) );
  OAI211_X1 U21054 ( .C1(n19008), .C2(n18916), .A(n18915), .B(n18914), .ZN(
        P2_U2835) );
  OAI22_X1 U21055 ( .A1(n18918), .A2(n19036), .B1(n18917), .B2(n19041), .ZN(
        n18922) );
  INV_X1 U21056 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n18919) );
  OAI22_X1 U21057 ( .A1(n18920), .A2(n19037), .B1(n18919), .B2(n19040), .ZN(
        n18921) );
  AOI211_X1 U21058 ( .C1(n18923), .C2(n19045), .A(n18922), .B(n18921), .ZN(
        n18929) );
  INV_X1 U21059 ( .A(n18924), .ZN(n18927) );
  NAND2_X1 U21060 ( .A1(n17412), .A2(n18925), .ZN(n18926) );
  NAND2_X1 U21061 ( .A1(n18926), .A2(n18927), .ZN(n18933) );
  OAI211_X1 U21062 ( .C1(n18927), .C2(n18926), .A(n19003), .B(n18933), .ZN(
        n18928) );
  OAI211_X1 U21063 ( .C1(n19051), .C2(n18930), .A(n18929), .B(n18928), .ZN(
        P2_U2834) );
  AOI22_X1 U21064 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19012), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19011), .ZN(n18939) );
  AOI22_X1 U21065 ( .A1(n18931), .A2(n19009), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n19013), .ZN(n18938) );
  AOI22_X1 U21066 ( .A1(n18932), .A2(n19045), .B1(n19856), .B2(n19014), .ZN(
        n18937) );
  NAND2_X1 U21067 ( .A1(n17412), .A2(n18933), .ZN(n18934) );
  NAND2_X1 U21068 ( .A1(n18934), .A2(n18935), .ZN(n18947) );
  OAI211_X1 U21069 ( .C1(n18935), .C2(n18934), .A(n19003), .B(n18947), .ZN(
        n18936) );
  NAND4_X1 U21070 ( .A1(n18939), .A2(n18938), .A3(n18937), .A4(n18936), .ZN(
        P2_U2833) );
  OAI22_X1 U21071 ( .A1(n18940), .A2(n19036), .B1(n13161), .B2(n19041), .ZN(
        n18944) );
  INV_X1 U21072 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n18941) );
  OAI22_X1 U21073 ( .A1(n18942), .A2(n19037), .B1(n18941), .B2(n19040), .ZN(
        n18943) );
  AOI211_X1 U21074 ( .C1(n18945), .C2(n19045), .A(n18944), .B(n18943), .ZN(
        n18951) );
  INV_X1 U21075 ( .A(n18946), .ZN(n18949) );
  NAND2_X1 U21076 ( .A1(n17412), .A2(n18947), .ZN(n18948) );
  OAI211_X1 U21077 ( .C1(n19051), .C2(n18952), .A(n18951), .B(n18950), .ZN(
        P2_U2832) );
  AOI22_X1 U21078 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19011), .B1(n18953), 
        .B2(n19009), .ZN(n18961) );
  AOI22_X1 U21079 ( .A1(n19013), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19012), .ZN(n18960) );
  AOI22_X1 U21080 ( .A1(n18955), .A2(n19045), .B1(n18954), .B2(n19014), .ZN(
        n18959) );
  NAND2_X1 U21081 ( .A1(n18956), .A2(n18957), .ZN(n18967) );
  OAI211_X1 U21082 ( .C1(n18957), .C2(n18956), .A(n19003), .B(n18967), .ZN(
        n18958) );
  NAND4_X1 U21083 ( .A1(n18961), .A2(n18960), .A3(n18959), .A4(n18958), .ZN(
        P2_U2831) );
  AOI22_X1 U21084 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19012), .B1(
        n18962), .B2(n19009), .ZN(n18973) );
  AOI22_X1 U21085 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19011), .B1(n19013), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n18972) );
  INV_X1 U21086 ( .A(n18963), .ZN(n18964) );
  AOI22_X1 U21087 ( .A1(n18965), .A2(n19045), .B1(n18964), .B2(n19014), .ZN(
        n18971) );
  INV_X1 U21088 ( .A(n18966), .ZN(n18969) );
  NAND2_X1 U21089 ( .A1(n17412), .A2(n18967), .ZN(n18968) );
  NAND2_X1 U21090 ( .A1(n18968), .A2(n18969), .ZN(n18978) );
  OAI211_X1 U21091 ( .C1(n18969), .C2(n18968), .A(n19003), .B(n18978), .ZN(
        n18970) );
  NAND4_X1 U21092 ( .A1(n18973), .A2(n18972), .A3(n18971), .A4(n18970), .ZN(
        P2_U2830) );
  AOI22_X1 U21093 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19011), .B1(n18974), 
        .B2(n19009), .ZN(n18984) );
  AOI22_X1 U21094 ( .A1(n19013), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19012), .ZN(n18983) );
  OAI22_X1 U21095 ( .A1(n18976), .A2(n19008), .B1(n18975), .B2(n19051), .ZN(
        n18977) );
  INV_X1 U21096 ( .A(n18977), .ZN(n18982) );
  NAND2_X1 U21097 ( .A1(n17412), .A2(n18978), .ZN(n18979) );
  OAI211_X1 U21098 ( .C1(n18980), .C2(n18979), .A(n19003), .B(n19001), .ZN(
        n18981) );
  NAND4_X1 U21099 ( .A1(n18984), .A2(n18983), .A3(n18982), .A4(n18981), .ZN(
        P2_U2829) );
  INV_X1 U21100 ( .A(n18985), .ZN(n18989) );
  INV_X1 U21101 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n18987) );
  AOI22_X1 U21102 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19012), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19011), .ZN(n18986) );
  OAI21_X1 U21103 ( .B1(n19040), .B2(n18987), .A(n18986), .ZN(n18988) );
  AOI21_X1 U21104 ( .B1(n18989), .B2(n19009), .A(n18988), .ZN(n18994) );
  NAND2_X1 U21105 ( .A1(n19001), .A2(n11188), .ZN(n18990) );
  XNOR2_X1 U21106 ( .A(n18990), .B(n19002), .ZN(n18991) );
  AOI22_X1 U21107 ( .A1(n18992), .A2(n19045), .B1(n19003), .B2(n18991), .ZN(
        n18993) );
  OAI211_X1 U21108 ( .C1(n18995), .C2(n19051), .A(n18994), .B(n18993), .ZN(
        P2_U2828) );
  INV_X1 U21109 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18997) );
  OAI22_X1 U21110 ( .A1(n18997), .A2(n19036), .B1(n18996), .B2(n19037), .ZN(
        n18999) );
  OAI22_X1 U21111 ( .A1(n17058), .A2(n19041), .B1(n19040), .B2(n13584), .ZN(
        n18998) );
  AOI211_X1 U21112 ( .C1(n19000), .C2(n19014), .A(n18999), .B(n18998), .ZN(
        n19007) );
  NAND2_X1 U21113 ( .A1(n19005), .A2(n19004), .ZN(n19016) );
  OAI211_X1 U21114 ( .C1(n19005), .C2(n19004), .A(n19003), .B(n19016), .ZN(
        n19006) );
  OAI211_X1 U21115 ( .C1(n19008), .C2(n17173), .A(n19007), .B(n19006), .ZN(
        P2_U2827) );
  AOI22_X1 U21116 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19011), .B1(n19010), 
        .B2(n19009), .ZN(n19022) );
  AOI22_X1 U21117 ( .A1(n19013), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19012), .ZN(n19021) );
  AOI22_X1 U21118 ( .A1(n16252), .A2(n19045), .B1(n19015), .B2(n19014), .ZN(
        n19020) );
  NAND2_X1 U21119 ( .A1(n19016), .A2(n17412), .ZN(n19017) );
  NAND2_X1 U21120 ( .A1(n19017), .A2(n19018), .ZN(n19030) );
  OAI211_X1 U21121 ( .C1(n19018), .C2(n19017), .A(n19003), .B(n19030), .ZN(
        n19019) );
  NAND4_X1 U21122 ( .A1(n19022), .A2(n19021), .A3(n19020), .A4(n19019), .ZN(
        P2_U2826) );
  OAI22_X1 U21123 ( .A1(n19024), .A2(n19037), .B1(n19023), .B2(n19041), .ZN(
        n19028) );
  OAI22_X1 U21124 ( .A1(n19040), .A2(n19026), .B1(n19036), .B2(n19025), .ZN(
        n19027) );
  AOI211_X1 U21125 ( .C1(n19029), .C2(n19045), .A(n19028), .B(n19027), .ZN(
        n19033) );
  NAND2_X1 U21126 ( .A1(n17412), .A2(n19030), .ZN(n19046) );
  AOI21_X1 U21127 ( .B1(n19047), .B2(n19046), .A(n19154), .ZN(n19031) );
  OAI21_X1 U21128 ( .B1(n19047), .B2(n19046), .A(n19031), .ZN(n19032) );
  OAI211_X1 U21129 ( .C1(n19034), .C2(n19051), .A(n19033), .B(n19032), .ZN(
        P2_U2825) );
  INV_X1 U21130 ( .A(n19035), .ZN(n19038) );
  OAI22_X1 U21131 ( .A1(n19038), .A2(n19037), .B1(n15224), .B2(n19036), .ZN(
        n19044) );
  OAI22_X1 U21132 ( .A1(n19042), .A2(n19041), .B1(n19040), .B2(n19039), .ZN(
        n19043) );
  AOI211_X1 U21133 ( .C1(n19045), .C2(n16894), .A(n19044), .B(n19043), .ZN(
        n19050) );
  NAND3_X1 U21134 ( .A1(n19048), .A2(n19047), .A3(n19046), .ZN(n19049) );
  OAI211_X1 U21135 ( .C1(n19052), .C2(n19051), .A(n19050), .B(n19049), .ZN(
        P2_U2824) );
  AOI21_X1 U21136 ( .B1(n19053), .B2(n19733), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19055) );
  OAI22_X1 U21137 ( .A1(n19056), .A2(n19055), .B1(n19054), .B2(n19674), .ZN(
        n19058) );
  MUX2_X1 U21138 ( .A(n19058), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n19057), .Z(P2_U3601) );
  INV_X1 U21139 ( .A(n19059), .ZN(n19061) );
  NOR4_X1 U21140 ( .A1(n19062), .A2(n19061), .A3(n19060), .A4(n19148), .ZN(
        n19063) );
  NAND2_X1 U21141 ( .A1(n19066), .A2(n19063), .ZN(n19064) );
  OAI21_X1 U21142 ( .B1(n19066), .B2(n19065), .A(n19064), .ZN(P2_U3595) );
  INV_X1 U21143 ( .A(n20163), .ZN(n20169) );
  AOI22_X1 U21144 ( .A1(n19129), .A2(n20169), .B1(n19138), .B2(n19067), .ZN(
        n19077) );
  AOI21_X1 U21145 ( .B1(n19103), .B2(n19069), .A(n19068), .ZN(n19072) );
  NAND2_X1 U21146 ( .A1(n19108), .A2(n19070), .ZN(n19071) );
  OAI211_X1 U21147 ( .C1(n19074), .C2(n19073), .A(n19072), .B(n19071), .ZN(
        n19075) );
  INV_X1 U21148 ( .A(n19075), .ZN(n19076) );
  OAI211_X1 U21149 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19109), .A(
        n19077), .B(n19076), .ZN(P2_U3046) );
  NAND2_X1 U21150 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19139), .ZN(n19078) );
  OAI211_X1 U21151 ( .C1(n19080), .C2(n13474), .A(n19079), .B(n19078), .ZN(
        n19081) );
  AOI21_X1 U21152 ( .B1(n19129), .B2(n19650), .A(n19081), .ZN(n19085) );
  AOI22_X1 U21153 ( .A1(n19083), .A2(n19108), .B1(n19103), .B2(n19082), .ZN(
        n19084) );
  OAI211_X1 U21154 ( .C1(n19086), .C2(n19091), .A(n19085), .B(n19084), .ZN(
        P2_U3036) );
  AOI22_X1 U21155 ( .A1(n19088), .A2(n19129), .B1(n19087), .B2(n13497), .ZN(
        n19101) );
  INV_X1 U21156 ( .A(n19089), .ZN(n19092) );
  OAI22_X1 U21157 ( .A1(n19092), .A2(n19091), .B1(n19133), .B2(n19090), .ZN(
        n19093) );
  AOI21_X1 U21158 ( .B1(n19108), .B2(n19094), .A(n19093), .ZN(n19100) );
  NAND2_X1 U21159 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19095), .ZN(n19099) );
  OAI21_X1 U21160 ( .B1(n19097), .B2(n19096), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19098) );
  NAND4_X1 U21161 ( .A1(n19101), .A2(n19100), .A3(n19099), .A4(n19098), .ZN(
        P2_U3032) );
  AOI22_X1 U21162 ( .A1(n19129), .A2(n19104), .B1(n19103), .B2(n19102), .ZN(
        n19118) );
  OAI21_X1 U21163 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19109), .A(
        n19127), .ZN(n19111) );
  AOI22_X1 U21164 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n19111), .B1(
        n19138), .B2(n19110), .ZN(n19117) );
  OAI21_X1 U21165 ( .B1(n19113), .B2(n19134), .A(n19112), .ZN(n19114) );
  NAND2_X1 U21166 ( .A1(n19114), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19128) );
  NAND4_X1 U21167 ( .A1(n19118), .A2(n19117), .A3(n19116), .A4(n19115), .ZN(
        P2_U3029) );
  NOR2_X1 U21168 ( .A1(n19120), .A2(n19119), .ZN(n19124) );
  OAI21_X1 U21169 ( .B1(n19122), .B2(n19133), .A(n19121), .ZN(n19123) );
  AOI211_X1 U21170 ( .C1(n19125), .C2(n19138), .A(n19124), .B(n19123), .ZN(
        n19126) );
  OAI221_X1 U21171 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19128), 
        .C1(n13487), .C2(n19127), .A(n19126), .ZN(P2_U3030) );
  AOI22_X1 U21172 ( .A1(n19130), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19129), .B2(n19657), .ZN(n19146) );
  INV_X1 U21173 ( .A(n19131), .ZN(n19135) );
  OAI22_X1 U21174 ( .A1(n19135), .A2(n19134), .B1(n19133), .B2(n19132), .ZN(
        n19136) );
  AOI21_X1 U21175 ( .B1(n19138), .B2(n19137), .A(n19136), .ZN(n19145) );
  NAND2_X1 U21176 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19139), .ZN(n19144) );
  INV_X1 U21177 ( .A(n19140), .ZN(n19142) );
  OAI211_X1 U21178 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n19142), .B(n19141), .ZN(n19143) );
  NAND4_X1 U21179 ( .A1(n19146), .A2(n19145), .A3(n19144), .A4(n19143), .ZN(
        P2_U3038) );
  NAND2_X1 U21180 ( .A1(n19161), .A2(n19147), .ZN(n19163) );
  OAI21_X1 U21181 ( .B1(n19149), .B2(n19148), .A(n19171), .ZN(n19153) );
  INV_X1 U21182 ( .A(n19158), .ZN(n19151) );
  NAND2_X1 U21183 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n22197), .ZN(n19150) );
  AOI21_X1 U21184 ( .B1(n19151), .B2(n19163), .A(n19150), .ZN(n19152) );
  AOI21_X1 U21185 ( .B1(n19163), .B2(n19153), .A(n19152), .ZN(n19155) );
  NAND2_X1 U21186 ( .A1(n19155), .A2(n19154), .ZN(P2_U3177) );
  AOI22_X1 U21187 ( .A1(n19158), .A2(n22197), .B1(n19157), .B2(n19156), .ZN(
        n19170) );
  AOI22_X1 U21188 ( .A1(n19161), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19160), 
        .B2(n19159), .ZN(n19169) );
  NOR2_X1 U21189 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19162), .ZN(n19166) );
  OAI22_X1 U21190 ( .A1(n19166), .A2(n19165), .B1(n19164), .B2(n19163), .ZN(
        n19167) );
  NAND4_X1 U21191 ( .A1(n19170), .A2(n19169), .A3(n19168), .A4(n19167), .ZN(
        P2_U3176) );
  NOR2_X1 U21192 ( .A1(n19172), .A2(n19171), .ZN(n19175) );
  MUX2_X1 U21193 ( .A(P2_MORE_REG_SCAN_IN), .B(n19173), .S(n19175), .Z(
        P2_U3609) );
  OAI21_X1 U21194 ( .B1(n19175), .B2(n12689), .A(n19174), .ZN(P2_U2819) );
  INV_X1 U21195 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20598) );
  AOI22_X1 U21196 ( .A1(n19487), .A2(n20598), .B1(n19200), .B2(U215), .ZN(U282) );
  OAI22_X1 U21197 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19487), .ZN(n19176) );
  INV_X1 U21198 ( .A(n19176), .ZN(U281) );
  INV_X1 U21199 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n19177) );
  INV_X1 U21200 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19913) );
  AOI22_X1 U21201 ( .A1(n19487), .A2(n19177), .B1(n19913), .B2(U215), .ZN(U280) );
  OAI22_X1 U21202 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19487), .ZN(n19178) );
  INV_X1 U21203 ( .A(n19178), .ZN(U279) );
  OAI22_X1 U21204 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19487), .ZN(n19179) );
  INV_X1 U21205 ( .A(n19179), .ZN(U278) );
  OAI22_X1 U21206 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19487), .ZN(n19180) );
  INV_X1 U21207 ( .A(n19180), .ZN(U277) );
  OAI22_X1 U21208 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19529), .ZN(n19181) );
  INV_X1 U21209 ( .A(n19181), .ZN(U276) );
  OAI22_X1 U21210 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19529), .ZN(n19182) );
  INV_X1 U21211 ( .A(n19182), .ZN(U275) );
  OAI22_X1 U21212 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19529), .ZN(n19183) );
  INV_X1 U21213 ( .A(n19183), .ZN(U274) );
  OAI22_X1 U21214 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19529), .ZN(n19184) );
  INV_X1 U21215 ( .A(n19184), .ZN(U273) );
  INV_X1 U21216 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n19185) );
  INV_X1 U21217 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21162) );
  AOI22_X1 U21218 ( .A1(n19529), .A2(n19185), .B1(n21162), .B2(U215), .ZN(U272) );
  INV_X1 U21219 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n19186) );
  INV_X1 U21220 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19964) );
  AOI22_X1 U21221 ( .A1(n19487), .A2(n19186), .B1(n19964), .B2(U215), .ZN(U271) );
  OAI22_X1 U21222 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19487), .ZN(n19187) );
  INV_X1 U21223 ( .A(n19187), .ZN(U270) );
  INV_X1 U21224 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n19188) );
  INV_X1 U21225 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n20066) );
  AOI22_X1 U21226 ( .A1(n19487), .A2(n19188), .B1(n20066), .B2(U215), .ZN(U269) );
  OAI22_X1 U21227 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19529), .ZN(n19189) );
  INV_X1 U21228 ( .A(n19189), .ZN(U268) );
  OAI22_X1 U21229 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19487), .ZN(n19190) );
  INV_X1 U21230 ( .A(n19190), .ZN(U267) );
  OAI22_X1 U21231 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19487), .ZN(n19191) );
  INV_X1 U21232 ( .A(n19191), .ZN(U266) );
  OAI22_X1 U21233 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19487), .ZN(n19192) );
  INV_X1 U21234 ( .A(n19192), .ZN(U265) );
  OAI22_X1 U21235 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19487), .ZN(n19193) );
  INV_X1 U21236 ( .A(n19193), .ZN(U264) );
  INV_X1 U21237 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n19194) );
  INV_X1 U21238 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21224) );
  AOI22_X1 U21239 ( .A1(n19487), .A2(n19194), .B1(n21224), .B2(U215), .ZN(U263) );
  INV_X1 U21240 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n19195) );
  INV_X1 U21241 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21117) );
  AOI22_X1 U21242 ( .A1(n19487), .A2(n19195), .B1(n21117), .B2(U215), .ZN(U262) );
  OAI22_X1 U21243 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19487), .ZN(n19196) );
  INV_X1 U21244 ( .A(n19196), .ZN(U261) );
  INV_X1 U21245 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n19197) );
  INV_X1 U21246 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21127) );
  AOI22_X1 U21247 ( .A1(n19529), .A2(n19197), .B1(n21127), .B2(U215), .ZN(U260) );
  INV_X1 U21248 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n19198) );
  INV_X1 U21249 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n21235) );
  AOI22_X1 U21250 ( .A1(n19529), .A2(n19198), .B1(n21235), .B2(U215), .ZN(U259) );
  OAI22_X1 U21251 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19487), .ZN(n19199) );
  INV_X1 U21252 ( .A(n19199), .ZN(U258) );
  NOR2_X1 U21253 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19203), .ZN(
        n19213) );
  NAND2_X1 U21254 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19213), .ZN(
        n19491) );
  NAND2_X1 U21255 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19531), .ZN(n19226) );
  INV_X1 U21256 ( .A(n19213), .ZN(n19212) );
  NOR2_X2 U21257 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19212), .ZN(
        n19552) );
  NOR2_X2 U21258 ( .A1(n19200), .A2(n19324), .ZN(n19280) );
  NAND2_X1 U21259 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21810), .ZN(n21811) );
  NOR2_X1 U21260 ( .A1(n21773), .A2(n19201), .ZN(n19271) );
  AND2_X1 U21261 ( .A1(n21811), .A2(n19271), .ZN(n19533) );
  AND2_X1 U21262 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n19532), .ZN(n19274) );
  AOI22_X1 U21263 ( .A1(n19552), .A2(n19280), .B1(n19533), .B2(n19274), .ZN(
        n19208) );
  NAND2_X1 U21264 ( .A1(n19202), .A2(n19532), .ZN(n19232) );
  INV_X1 U21265 ( .A(n19232), .ZN(n19222) );
  AOI22_X1 U21266 ( .A1(n19531), .A2(n19213), .B1(n19271), .B2(n19222), .ZN(
        n19536) );
  NAND2_X1 U21267 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21783) );
  NOR2_X2 U21268 ( .A1(n21783), .A2(n19203), .ZN(n19617) );
  INV_X1 U21269 ( .A(n19204), .ZN(n19205) );
  NAND2_X1 U21270 ( .A1(n19206), .A2(n19205), .ZN(n19534) );
  NOR2_X1 U21271 ( .A1(n21263), .A2(n19534), .ZN(n19223) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n19223), .ZN(n19207) );
  OAI211_X1 U21273 ( .C1(n19491), .C2(n19226), .A(n19208), .B(n19207), .ZN(
        P3_U2995) );
  INV_X1 U21274 ( .A(n19223), .ZN(n19283) );
  NAND2_X1 U21275 ( .A1(n19271), .A2(n19234), .ZN(n19633) );
  INV_X1 U21276 ( .A(n19226), .ZN(n19275) );
  INV_X1 U21277 ( .A(n21811), .ZN(n20669) );
  INV_X1 U21278 ( .A(n19491), .ZN(n19626) );
  INV_X1 U21279 ( .A(n19633), .ZN(n19540) );
  NOR2_X1 U21280 ( .A1(n19626), .A2(n19540), .ZN(n19276) );
  NOR2_X1 U21281 ( .A1(n20669), .A2(n19276), .ZN(n19539) );
  AOI22_X1 U21282 ( .A1(n19275), .A2(n19552), .B1(n19274), .B2(n19539), .ZN(
        n19211) );
  NAND2_X1 U21283 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21791), .ZN(
        n19231) );
  NOR2_X1 U21284 ( .A1(n21783), .A2(n19231), .ZN(n19558) );
  CLKBUF_X1 U21285 ( .A(n19558), .Z(n19546) );
  NOR2_X1 U21286 ( .A1(n19552), .A2(n19546), .ZN(n19216) );
  OAI21_X1 U21287 ( .B1(n19216), .B2(n19246), .A(n19276), .ZN(n19209) );
  OAI211_X1 U21288 ( .C1(n19540), .C2(n21818), .A(n19532), .B(n19209), .ZN(
        n19541) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19541), .B1(
        n19280), .B2(n19546), .ZN(n19210) );
  OAI211_X1 U21290 ( .C1(n19283), .C2(n19633), .A(n19211), .B(n19210), .ZN(
        P3_U2987) );
  NOR2_X1 U21291 ( .A1(n20669), .A2(n19212), .ZN(n19545) );
  AOI22_X1 U21292 ( .A1(n19275), .A2(n19546), .B1(n19274), .B2(n19545), .ZN(
        n19215) );
  NOR2_X1 U21293 ( .A1(n21784), .A2(n19231), .ZN(n19221) );
  AOI22_X1 U21294 ( .A1(n19531), .A2(n19221), .B1(n19213), .B2(n19222), .ZN(
        n19547) );
  INV_X1 U21295 ( .A(n19221), .ZN(n19220) );
  NOR2_X2 U21296 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19220), .ZN(
        n19565) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19547), .B1(
        n19280), .B2(n19565), .ZN(n19214) );
  OAI211_X1 U21298 ( .C1(n19491), .C2(n19283), .A(n19215), .B(n19214), .ZN(
        P3_U2979) );
  INV_X1 U21299 ( .A(n19552), .ZN(n19544) );
  NOR2_X1 U21300 ( .A1(n20669), .A2(n19216), .ZN(n19551) );
  AOI22_X1 U21301 ( .A1(n19275), .A2(n19565), .B1(n19274), .B2(n19551), .ZN(
        n19219) );
  INV_X1 U21302 ( .A(n19565), .ZN(n19550) );
  INV_X1 U21303 ( .A(n19231), .ZN(n19233) );
  NOR2_X1 U21304 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19234), .ZN(
        n19255) );
  NAND2_X1 U21305 ( .A1(n19233), .A2(n19255), .ZN(n19556) );
  NAND2_X1 U21306 ( .A1(n19550), .A2(n19556), .ZN(n19228) );
  AOI21_X1 U21307 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19366), .ZN(n19278) );
  INV_X1 U21308 ( .A(n19216), .ZN(n19217) );
  AOI22_X1 U21309 ( .A1(n19531), .A2(n19228), .B1(n19278), .B2(n19217), .ZN(
        n19553) );
  INV_X1 U21310 ( .A(n19556), .ZN(n19570) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19553), .B1(
        n19280), .B2(n19570), .ZN(n19218) );
  OAI211_X1 U21312 ( .C1(n19283), .C2(n19544), .A(n19219), .B(n19218), .ZN(
        P3_U2971) );
  NAND2_X1 U21313 ( .A1(n21784), .A2(n19234), .ZN(n21787) );
  NOR2_X2 U21314 ( .A1(n21787), .A2(n19231), .ZN(n19575) );
  NOR2_X1 U21315 ( .A1(n20669), .A2(n19220), .ZN(n19557) );
  AOI22_X1 U21316 ( .A1(n19280), .A2(n19575), .B1(n19274), .B2(n19557), .ZN(
        n19225) );
  AOI22_X1 U21317 ( .A1(n19531), .A2(n19233), .B1(n19222), .B2(n19221), .ZN(
        n19559) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19559), .B1(
        n19223), .B2(n19558), .ZN(n19224) );
  OAI211_X1 U21319 ( .C1(n19226), .C2(n19556), .A(n19225), .B(n19224), .ZN(
        P3_U2963) );
  INV_X1 U21320 ( .A(n19575), .ZN(n19562) );
  INV_X1 U21321 ( .A(n21783), .ZN(n19227) );
  NOR2_X1 U21322 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21791), .ZN(
        n19252) );
  NAND2_X1 U21323 ( .A1(n19227), .A2(n19252), .ZN(n19568) );
  NAND2_X1 U21324 ( .A1(n19562), .A2(n19568), .ZN(n19237) );
  OAI221_X1 U21325 ( .B1(n19228), .B2(n19241), .C1(n19228), .C2(n19237), .A(
        n19278), .ZN(n19564) );
  AND2_X1 U21326 ( .A1(n21811), .A2(n19228), .ZN(n19563) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19564), .B1(
        n19274), .B2(n19563), .ZN(n19230) );
  INV_X1 U21328 ( .A(n19568), .ZN(n19582) );
  AOI22_X1 U21329 ( .A1(n19275), .A2(n19575), .B1(n19280), .B2(n19582), .ZN(
        n19229) );
  OAI211_X1 U21330 ( .C1(n19283), .C2(n19550), .A(n19230), .B(n19229), .ZN(
        P3_U2955) );
  NAND2_X1 U21331 ( .A1(n21784), .A2(n21811), .ZN(n19268) );
  NOR2_X1 U21332 ( .A1(n19231), .A2(n19268), .ZN(n19569) );
  AOI22_X1 U21333 ( .A1(n19275), .A2(n19582), .B1(n19274), .B2(n19569), .ZN(
        n19236) );
  NOR2_X1 U21334 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19232), .ZN(
        n19270) );
  AOI22_X1 U21335 ( .A1(n19531), .A2(n19240), .B1(n19233), .B2(n19270), .ZN(
        n19571) );
  NAND2_X1 U21336 ( .A1(n19234), .A2(n19240), .ZN(n19579) );
  INV_X1 U21337 ( .A(n19579), .ZN(n19587) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19571), .B1(
        n19280), .B2(n19587), .ZN(n19235) );
  OAI211_X1 U21339 ( .C1(n19283), .C2(n19556), .A(n19236), .B(n19235), .ZN(
        P3_U2947) );
  NAND2_X1 U21340 ( .A1(n19255), .A2(n19252), .ZN(n19508) );
  INV_X1 U21341 ( .A(n19508), .ZN(n19593) );
  AND2_X1 U21342 ( .A1(n21811), .A2(n19237), .ZN(n19574) );
  AOI22_X1 U21343 ( .A1(n19280), .A2(n19593), .B1(n19274), .B2(n19574), .ZN(
        n19239) );
  NAND2_X1 U21344 ( .A1(n19579), .A2(n19508), .ZN(n19245) );
  AOI22_X1 U21345 ( .A1(n19531), .A2(n19245), .B1(n19278), .B2(n19237), .ZN(
        n19576) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19576), .B1(
        n19275), .B2(n19587), .ZN(n19238) );
  OAI211_X1 U21347 ( .C1(n19283), .C2(n19562), .A(n19239), .B(n19238), .ZN(
        P3_U2939) );
  AND2_X1 U21348 ( .A1(n21811), .A2(n19240), .ZN(n19580) );
  AOI22_X1 U21349 ( .A1(n19275), .A2(n19593), .B1(n19274), .B2(n19580), .ZN(
        n19244) );
  OAI21_X1 U21350 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19241), .A(
        n19532), .ZN(n19242) );
  AOI21_X1 U21351 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n21783), .A(n19242), 
        .ZN(n19261) );
  NAND2_X1 U21352 ( .A1(n19252), .A2(n19261), .ZN(n19581) );
  INV_X1 U21353 ( .A(n19252), .ZN(n19251) );
  NOR2_X2 U21354 ( .A1(n21787), .A2(n19251), .ZN(n19599) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19581), .B1(
        n19280), .B2(n19599), .ZN(n19243) );
  OAI211_X1 U21356 ( .C1(n19283), .C2(n19568), .A(n19244), .B(n19243), .ZN(
        P3_U2931) );
  NOR2_X2 U21357 ( .A1(n21783), .A2(n19267), .ZN(n19605) );
  NOR2_X1 U21358 ( .A1(n19599), .A2(n19605), .ZN(n19256) );
  INV_X1 U21359 ( .A(n19245), .ZN(n19248) );
  OAI21_X1 U21360 ( .B1(n19256), .B2(n19246), .A(n19248), .ZN(n19247) );
  OAI211_X1 U21361 ( .C1(n19587), .C2(n21818), .A(n19532), .B(n19247), .ZN(
        n19588) );
  NOR2_X1 U21362 ( .A1(n20669), .A2(n19248), .ZN(n19586) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19588), .B1(
        n19274), .B2(n19586), .ZN(n19250) );
  AOI22_X1 U21364 ( .A1(n19275), .A2(n19599), .B1(n19280), .B2(n19605), .ZN(
        n19249) );
  OAI211_X1 U21365 ( .C1(n19283), .C2(n19579), .A(n19250), .B(n19249), .ZN(
        P3_U2923) );
  NOR2_X1 U21366 ( .A1(n19251), .A2(n19268), .ZN(n19592) );
  AOI22_X1 U21367 ( .A1(n19275), .A2(n19605), .B1(n19274), .B2(n19592), .ZN(
        n19254) );
  NOR2_X1 U21368 ( .A1(n21784), .A2(n19267), .ZN(n19260) );
  AOI22_X1 U21369 ( .A1(n19531), .A2(n19260), .B1(n19252), .B2(n19270), .ZN(
        n19594) );
  NOR3_X4 U21370 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21784), .A3(
        n19267), .ZN(n19610) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19594), .B1(
        n19280), .B2(n19610), .ZN(n19253) );
  OAI211_X1 U21372 ( .C1(n19283), .C2(n19508), .A(n19254), .B(n19253), .ZN(
        P3_U2915) );
  INV_X1 U21373 ( .A(n19599), .ZN(n19585) );
  NOR2_X1 U21374 ( .A1(n20669), .A2(n19256), .ZN(n19598) );
  AOI22_X1 U21375 ( .A1(n19275), .A2(n19610), .B1(n19274), .B2(n19598), .ZN(
        n19259) );
  INV_X1 U21376 ( .A(n19610), .ZN(n19597) );
  NAND2_X1 U21377 ( .A1(n19255), .A2(n19269), .ZN(n19603) );
  NAND2_X1 U21378 ( .A1(n19597), .A2(n19603), .ZN(n19264) );
  INV_X1 U21379 ( .A(n19256), .ZN(n19257) );
  AOI22_X1 U21380 ( .A1(n19531), .A2(n19264), .B1(n19278), .B2(n19257), .ZN(
        n19600) );
  INV_X1 U21381 ( .A(n19603), .ZN(n19618) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19600), .B1(
        n19280), .B2(n19618), .ZN(n19258) );
  OAI211_X1 U21383 ( .C1(n19283), .C2(n19585), .A(n19259), .B(n19258), .ZN(
        P3_U2907) );
  INV_X1 U21384 ( .A(n19605), .ZN(n19591) );
  AND2_X1 U21385 ( .A1(n21811), .A2(n19260), .ZN(n19604) );
  AOI22_X1 U21386 ( .A1(n19275), .A2(n19618), .B1(n19274), .B2(n19604), .ZN(
        n19263) );
  NAND2_X1 U21387 ( .A1(n19261), .A2(n19269), .ZN(n19606) );
  NOR2_X2 U21388 ( .A1(n21787), .A2(n19267), .ZN(n19628) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19606), .B1(
        n19280), .B2(n19628), .ZN(n19262) );
  OAI211_X1 U21390 ( .C1(n19283), .C2(n19591), .A(n19263), .B(n19262), .ZN(
        P3_U2899) );
  AND2_X1 U21391 ( .A1(n21811), .A2(n19264), .ZN(n19609) );
  AOI22_X1 U21392 ( .A1(n19275), .A2(n19628), .B1(n19274), .B2(n19609), .ZN(
        n19266) );
  INV_X1 U21393 ( .A(n19617), .ZN(n19480) );
  INV_X1 U21394 ( .A(n19628), .ZN(n19614) );
  NAND2_X1 U21395 ( .A1(n19480), .A2(n19614), .ZN(n19277) );
  AOI22_X1 U21396 ( .A1(n19531), .A2(n19277), .B1(n19278), .B2(n19264), .ZN(
        n19611) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19611), .B1(
        n19617), .B2(n19280), .ZN(n19265) );
  OAI211_X1 U21398 ( .C1(n19283), .C2(n19597), .A(n19266), .B(n19265), .ZN(
        P3_U2891) );
  NOR2_X1 U21399 ( .A1(n19268), .A2(n19267), .ZN(n19615) );
  AOI22_X1 U21400 ( .A1(n19275), .A2(n19617), .B1(n19274), .B2(n19615), .ZN(
        n19273) );
  AOI22_X1 U21401 ( .A1(n19531), .A2(n19271), .B1(n19270), .B2(n19269), .ZN(
        n19619) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19619), .B1(
        n19280), .B2(n19540), .ZN(n19272) );
  OAI211_X1 U21403 ( .C1(n19283), .C2(n19603), .A(n19273), .B(n19272), .ZN(
        P3_U2883) );
  AND2_X1 U21404 ( .A1(n21811), .A2(n19277), .ZN(n19624) );
  AOI22_X1 U21405 ( .A1(n19275), .A2(n19540), .B1(n19274), .B2(n19624), .ZN(
        n19282) );
  INV_X1 U21406 ( .A(n19276), .ZN(n19279) );
  AOI22_X1 U21407 ( .A1(n19531), .A2(n19279), .B1(n19278), .B2(n19277), .ZN(
        n19629) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19629), .B1(
        n19626), .B2(n19280), .ZN(n19281) );
  OAI211_X1 U21409 ( .C1(n19283), .C2(n19614), .A(n19282), .B(n19281), .ZN(
        P3_U2875) );
  INV_X1 U21410 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n19284) );
  AOI22_X1 U21411 ( .A1(n19487), .A2(n19284), .B1(n21136), .B2(U215), .ZN(U257) );
  NAND2_X1 U21412 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19531), .ZN(n19322) );
  NAND2_X1 U21413 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19531), .ZN(n19316) );
  INV_X1 U21414 ( .A(n19316), .ZN(n19318) );
  NOR2_X2 U21415 ( .A1(n21136), .A2(n19366), .ZN(n19317) );
  AOI22_X1 U21416 ( .A1(n19552), .A2(n19318), .B1(n19533), .B2(n19317), .ZN(
        n19286) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n11161), .ZN(n19285) );
  OAI211_X1 U21418 ( .C1(n19491), .C2(n19322), .A(n19286), .B(n19285), .ZN(
        P3_U2994) );
  AOI22_X1 U21419 ( .A1(n19546), .A2(n19318), .B1(n19539), .B2(n19317), .ZN(
        n19288) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n11161), .ZN(n19287) );
  OAI211_X1 U21421 ( .C1(n19544), .C2(n19322), .A(n19288), .B(n19287), .ZN(
        P3_U2986) );
  INV_X1 U21422 ( .A(n19322), .ZN(n19313) );
  AOI22_X1 U21423 ( .A1(n19546), .A2(n19313), .B1(n19545), .B2(n19317), .ZN(
        n19290) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19547), .B1(
        n19626), .B2(n11161), .ZN(n19289) );
  OAI211_X1 U21425 ( .C1(n19550), .C2(n19316), .A(n19290), .B(n19289), .ZN(
        P3_U2978) );
  AOI22_X1 U21426 ( .A1(n19570), .A2(n19318), .B1(n19551), .B2(n19317), .ZN(
        n19292) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n11161), .ZN(n19291) );
  OAI211_X1 U21428 ( .C1(n19550), .C2(n19322), .A(n19292), .B(n19291), .ZN(
        P3_U2970) );
  AOI22_X1 U21429 ( .A1(n19575), .A2(n19318), .B1(n19557), .B2(n19317), .ZN(
        n19294) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19559), .B1(
        n19558), .B2(n11161), .ZN(n19293) );
  OAI211_X1 U21431 ( .C1(n19556), .C2(n19322), .A(n19294), .B(n19293), .ZN(
        P3_U2962) );
  AOI22_X1 U21432 ( .A1(n19582), .A2(n19318), .B1(n19563), .B2(n19317), .ZN(
        n19296) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19564), .B1(
        n19565), .B2(n11161), .ZN(n19295) );
  OAI211_X1 U21434 ( .C1(n19562), .C2(n19322), .A(n19296), .B(n19295), .ZN(
        P3_U2954) );
  AOI22_X1 U21435 ( .A1(n19582), .A2(n19313), .B1(n19569), .B2(n19317), .ZN(
        n19298) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19571), .B1(
        n19570), .B2(n11161), .ZN(n19297) );
  OAI211_X1 U21437 ( .C1(n19579), .C2(n19316), .A(n19298), .B(n19297), .ZN(
        P3_U2946) );
  AOI22_X1 U21438 ( .A1(n19587), .A2(n19313), .B1(n19574), .B2(n19317), .ZN(
        n19300) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19576), .B1(
        n19575), .B2(n11161), .ZN(n19299) );
  OAI211_X1 U21440 ( .C1(n19508), .C2(n19316), .A(n19300), .B(n19299), .ZN(
        P3_U2938) );
  AOI22_X1 U21441 ( .A1(n19599), .A2(n19318), .B1(n19580), .B2(n19317), .ZN(
        n19302) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19581), .B1(
        n19582), .B2(n11161), .ZN(n19301) );
  OAI211_X1 U21443 ( .C1(n19508), .C2(n19322), .A(n19302), .B(n19301), .ZN(
        P3_U2930) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19588), .B1(
        n19586), .B2(n19317), .ZN(n19304) );
  AOI22_X1 U21445 ( .A1(n19587), .A2(n11161), .B1(n19605), .B2(n19318), .ZN(
        n19303) );
  OAI211_X1 U21446 ( .C1(n19585), .C2(n19322), .A(n19304), .B(n19303), .ZN(
        P3_U2922) );
  AOI22_X1 U21447 ( .A1(n19605), .A2(n19313), .B1(n19592), .B2(n19317), .ZN(
        n19306) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n11161), .ZN(n19305) );
  OAI211_X1 U21449 ( .C1(n19597), .C2(n19316), .A(n19306), .B(n19305), .ZN(
        P3_U2914) );
  AOI22_X1 U21450 ( .A1(n19610), .A2(n19313), .B1(n19598), .B2(n19317), .ZN(
        n19308) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n11161), .ZN(n19307) );
  OAI211_X1 U21452 ( .C1(n19603), .C2(n19316), .A(n19308), .B(n19307), .ZN(
        P3_U2906) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19606), .B1(
        n19604), .B2(n19317), .ZN(n19310) );
  AOI22_X1 U21454 ( .A1(n19605), .A2(n11161), .B1(n19618), .B2(n19313), .ZN(
        n19309) );
  OAI211_X1 U21455 ( .C1(n19614), .C2(n19316), .A(n19310), .B(n19309), .ZN(
        P3_U2898) );
  AOI22_X1 U21456 ( .A1(n19628), .A2(n19313), .B1(n19609), .B2(n19317), .ZN(
        n19312) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n11161), .ZN(n19311) );
  OAI211_X1 U21458 ( .C1(n19480), .C2(n19316), .A(n19312), .B(n19311), .ZN(
        P3_U2890) );
  AOI22_X1 U21459 ( .A1(n19617), .A2(n19313), .B1(n19615), .B2(n19317), .ZN(
        n19315) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n11161), .ZN(n19314) );
  OAI211_X1 U21461 ( .C1(n19633), .C2(n19316), .A(n19315), .B(n19314), .ZN(
        P3_U2882) );
  AOI22_X1 U21462 ( .A1(n19626), .A2(n19318), .B1(n19624), .B2(n19317), .ZN(
        n19321) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n11161), .ZN(n19320) );
  OAI211_X1 U21464 ( .C1(n19633), .C2(n19322), .A(n19321), .B(n19320), .ZN(
        P3_U2874) );
  INV_X1 U21465 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n19323) );
  INV_X1 U21466 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21142) );
  AOI22_X1 U21467 ( .A1(n19487), .A2(n19323), .B1(n21142), .B2(U215), .ZN(U256) );
  NAND2_X1 U21468 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19531), .ZN(n19343) );
  NOR2_X2 U21469 ( .A1(n19913), .A2(n19324), .ZN(n19360) );
  NOR2_X2 U21470 ( .A1(n21142), .A2(n19366), .ZN(n19358) );
  AOI22_X1 U21471 ( .A1(n19552), .A2(n19360), .B1(n19533), .B2(n19358), .ZN(
        n19327) );
  NOR2_X1 U21472 ( .A1(n19325), .A2(n19534), .ZN(n19340) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n19340), .ZN(n19326) );
  OAI211_X1 U21474 ( .C1(n19491), .C2(n19343), .A(n19327), .B(n19326), .ZN(
        P3_U2993) );
  INV_X1 U21475 ( .A(n19343), .ZN(n19359) );
  AOI22_X1 U21476 ( .A1(n19552), .A2(n19359), .B1(n19539), .B2(n19358), .ZN(
        n19329) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19541), .B1(
        n19558), .B2(n19360), .ZN(n19328) );
  OAI211_X1 U21478 ( .C1(n19633), .C2(n19363), .A(n19329), .B(n19328), .ZN(
        P3_U2985) );
  AOI22_X1 U21479 ( .A1(n19565), .A2(n19360), .B1(n19545), .B2(n19358), .ZN(
        n19331) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19547), .B1(
        n19558), .B2(n19359), .ZN(n19330) );
  OAI211_X1 U21481 ( .C1(n19491), .C2(n19363), .A(n19331), .B(n19330), .ZN(
        P3_U2977) );
  AOI22_X1 U21482 ( .A1(n19565), .A2(n19359), .B1(n19551), .B2(n19358), .ZN(
        n19333) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19553), .B1(
        n19570), .B2(n19360), .ZN(n19332) );
  OAI211_X1 U21484 ( .C1(n19544), .C2(n19363), .A(n19333), .B(n19332), .ZN(
        P3_U2969) );
  AOI22_X1 U21485 ( .A1(n19575), .A2(n19360), .B1(n19557), .B2(n19358), .ZN(
        n19335) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19559), .B1(
        n19558), .B2(n19340), .ZN(n19334) );
  OAI211_X1 U21487 ( .C1(n19556), .C2(n19343), .A(n19335), .B(n19334), .ZN(
        P3_U2961) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19564), .B1(
        n19563), .B2(n19358), .ZN(n19337) );
  AOI22_X1 U21489 ( .A1(n19565), .A2(n19340), .B1(n19582), .B2(n19360), .ZN(
        n19336) );
  OAI211_X1 U21490 ( .C1(n19562), .C2(n19343), .A(n19337), .B(n19336), .ZN(
        P3_U2953) );
  AOI22_X1 U21491 ( .A1(n19582), .A2(n19359), .B1(n19569), .B2(n19358), .ZN(
        n19339) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19571), .B1(
        n19587), .B2(n19360), .ZN(n19338) );
  OAI211_X1 U21493 ( .C1(n19556), .C2(n19363), .A(n19339), .B(n19338), .ZN(
        P3_U2945) );
  AOI22_X1 U21494 ( .A1(n19593), .A2(n19360), .B1(n19574), .B2(n19358), .ZN(
        n19342) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19576), .B1(
        n19575), .B2(n19340), .ZN(n19341) );
  OAI211_X1 U21496 ( .C1(n19579), .C2(n19343), .A(n19342), .B(n19341), .ZN(
        P3_U2937) );
  AOI22_X1 U21497 ( .A1(n19593), .A2(n19359), .B1(n19580), .B2(n19358), .ZN(
        n19345) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19581), .B1(
        n19599), .B2(n19360), .ZN(n19344) );
  OAI211_X1 U21499 ( .C1(n19568), .C2(n19363), .A(n19345), .B(n19344), .ZN(
        P3_U2929) );
  AOI22_X1 U21500 ( .A1(n19599), .A2(n19359), .B1(n19586), .B2(n19358), .ZN(
        n19347) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19588), .B1(
        n19605), .B2(n19360), .ZN(n19346) );
  OAI211_X1 U21502 ( .C1(n19579), .C2(n19363), .A(n19347), .B(n19346), .ZN(
        P3_U2921) );
  AOI22_X1 U21503 ( .A1(n19605), .A2(n19359), .B1(n19592), .B2(n19358), .ZN(
        n19349) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19594), .B1(
        n19610), .B2(n19360), .ZN(n19348) );
  OAI211_X1 U21505 ( .C1(n19508), .C2(n19363), .A(n19349), .B(n19348), .ZN(
        P3_U2913) );
  AOI22_X1 U21506 ( .A1(n19610), .A2(n19359), .B1(n19598), .B2(n19358), .ZN(
        n19351) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19600), .B1(
        n19618), .B2(n19360), .ZN(n19350) );
  OAI211_X1 U21508 ( .C1(n19585), .C2(n19363), .A(n19351), .B(n19350), .ZN(
        P3_U2905) );
  AOI22_X1 U21509 ( .A1(n19618), .A2(n19359), .B1(n19604), .B2(n19358), .ZN(
        n19353) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19606), .B1(
        n19628), .B2(n19360), .ZN(n19352) );
  OAI211_X1 U21511 ( .C1(n19591), .C2(n19363), .A(n19353), .B(n19352), .ZN(
        P3_U2897) );
  AOI22_X1 U21512 ( .A1(n19628), .A2(n19359), .B1(n19609), .B2(n19358), .ZN(
        n19355) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19611), .B1(
        n19617), .B2(n19360), .ZN(n19354) );
  OAI211_X1 U21514 ( .C1(n19597), .C2(n19363), .A(n19355), .B(n19354), .ZN(
        P3_U2889) );
  AOI22_X1 U21515 ( .A1(n19617), .A2(n19359), .B1(n19615), .B2(n19358), .ZN(
        n19357) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19619), .B1(
        n19540), .B2(n19360), .ZN(n19356) );
  OAI211_X1 U21517 ( .C1(n19603), .C2(n19363), .A(n19357), .B(n19356), .ZN(
        P3_U2881) );
  AOI22_X1 U21518 ( .A1(n19540), .A2(n19359), .B1(n19624), .B2(n19358), .ZN(
        n19362) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19629), .B1(
        n19626), .B2(n19360), .ZN(n19361) );
  OAI211_X1 U21520 ( .C1(n19614), .C2(n19363), .A(n19362), .B(n19361), .ZN(
        P3_U2873) );
  INV_X1 U21521 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n19365) );
  AOI22_X1 U21522 ( .A1(n19529), .A2(n19365), .B1(n19367), .B2(U215), .ZN(U255) );
  NAND2_X1 U21523 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19531), .ZN(n19399) );
  AND2_X1 U21524 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19531), .ZN(n19402) );
  NOR2_X2 U21525 ( .A1(n19367), .A2(n19366), .ZN(n19400) );
  AOI22_X1 U21526 ( .A1(n19552), .A2(n19402), .B1(n19533), .B2(n19400), .ZN(
        n19369) );
  NOR2_X1 U21527 ( .A1(n21336), .A2(n19534), .ZN(n19396) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n19396), .ZN(n19368) );
  OAI211_X1 U21529 ( .C1(n19491), .C2(n19399), .A(n19369), .B(n19368), .ZN(
        P3_U2992) );
  INV_X1 U21530 ( .A(n19396), .ZN(n19405) );
  INV_X1 U21531 ( .A(n19399), .ZN(n19401) );
  AOI22_X1 U21532 ( .A1(n19552), .A2(n19401), .B1(n19539), .B2(n19400), .ZN(
        n19371) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19541), .B1(
        n19558), .B2(n19402), .ZN(n19370) );
  OAI211_X1 U21534 ( .C1(n19633), .C2(n19405), .A(n19371), .B(n19370), .ZN(
        P3_U2984) );
  AOI22_X1 U21535 ( .A1(n19565), .A2(n19402), .B1(n19545), .B2(n19400), .ZN(
        n19373) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19547), .B1(
        n19558), .B2(n19401), .ZN(n19372) );
  OAI211_X1 U21537 ( .C1(n19491), .C2(n19405), .A(n19373), .B(n19372), .ZN(
        P3_U2976) );
  AOI22_X1 U21538 ( .A1(n19570), .A2(n19402), .B1(n19551), .B2(n19400), .ZN(
        n19375) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19396), .ZN(n19374) );
  OAI211_X1 U21540 ( .C1(n19550), .C2(n19399), .A(n19375), .B(n19374), .ZN(
        P3_U2968) );
  AOI22_X1 U21541 ( .A1(n19575), .A2(n19402), .B1(n19557), .B2(n19400), .ZN(
        n19377) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19559), .B1(
        n19558), .B2(n19396), .ZN(n19376) );
  OAI211_X1 U21543 ( .C1(n19556), .C2(n19399), .A(n19377), .B(n19376), .ZN(
        P3_U2960) );
  AOI22_X1 U21544 ( .A1(n19582), .A2(n19402), .B1(n19563), .B2(n19400), .ZN(
        n19379) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19564), .B1(
        n19565), .B2(n19396), .ZN(n19378) );
  OAI211_X1 U21546 ( .C1(n19562), .C2(n19399), .A(n19379), .B(n19378), .ZN(
        P3_U2952) );
  AOI22_X1 U21547 ( .A1(n19582), .A2(n19401), .B1(n19569), .B2(n19400), .ZN(
        n19381) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19571), .B1(
        n19587), .B2(n19402), .ZN(n19380) );
  OAI211_X1 U21549 ( .C1(n19556), .C2(n19405), .A(n19381), .B(n19380), .ZN(
        P3_U2944) );
  AOI22_X1 U21550 ( .A1(n19587), .A2(n19401), .B1(n19574), .B2(n19400), .ZN(
        n19383) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19576), .B1(
        n19593), .B2(n19402), .ZN(n19382) );
  OAI211_X1 U21552 ( .C1(n19562), .C2(n19405), .A(n19383), .B(n19382), .ZN(
        P3_U2936) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19581), .B1(
        n19580), .B2(n19400), .ZN(n19385) );
  AOI22_X1 U21554 ( .A1(n19582), .A2(n19396), .B1(n19599), .B2(n19402), .ZN(
        n19384) );
  OAI211_X1 U21555 ( .C1(n19508), .C2(n19399), .A(n19385), .B(n19384), .ZN(
        P3_U2928) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19588), .B1(
        n19586), .B2(n19400), .ZN(n19387) );
  AOI22_X1 U21557 ( .A1(n19587), .A2(n19396), .B1(n19605), .B2(n19402), .ZN(
        n19386) );
  OAI211_X1 U21558 ( .C1(n19585), .C2(n19399), .A(n19387), .B(n19386), .ZN(
        P3_U2920) );
  AOI22_X1 U21559 ( .A1(n19610), .A2(n19402), .B1(n19592), .B2(n19400), .ZN(
        n19389) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19396), .ZN(n19388) );
  OAI211_X1 U21561 ( .C1(n19591), .C2(n19399), .A(n19389), .B(n19388), .ZN(
        P3_U2912) );
  AOI22_X1 U21562 ( .A1(n19610), .A2(n19401), .B1(n19598), .B2(n19400), .ZN(
        n19391) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19600), .B1(
        n19618), .B2(n19402), .ZN(n19390) );
  OAI211_X1 U21564 ( .C1(n19585), .C2(n19405), .A(n19391), .B(n19390), .ZN(
        P3_U2904) );
  AOI22_X1 U21565 ( .A1(n19628), .A2(n19402), .B1(n19604), .B2(n19400), .ZN(
        n19393) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19396), .ZN(n19392) );
  OAI211_X1 U21567 ( .C1(n19603), .C2(n19399), .A(n19393), .B(n19392), .ZN(
        P3_U2896) );
  AOI22_X1 U21568 ( .A1(n19617), .A2(n19402), .B1(n19609), .B2(n19400), .ZN(
        n19395) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19396), .ZN(n19394) );
  OAI211_X1 U21570 ( .C1(n19614), .C2(n19399), .A(n19395), .B(n19394), .ZN(
        P3_U2888) );
  AOI22_X1 U21571 ( .A1(n19540), .A2(n19402), .B1(n19615), .B2(n19400), .ZN(
        n19398) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19396), .ZN(n19397) );
  OAI211_X1 U21573 ( .C1(n19480), .C2(n19399), .A(n19398), .B(n19397), .ZN(
        P3_U2880) );
  AOI22_X1 U21574 ( .A1(n19540), .A2(n19401), .B1(n19624), .B2(n19400), .ZN(
        n19404) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19629), .B1(
        n19626), .B2(n19402), .ZN(n19403) );
  OAI211_X1 U21576 ( .C1(n19614), .C2(n19405), .A(n19404), .B(n19403), .ZN(
        P3_U2872) );
  OAI22_X1 U21577 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19487), .ZN(n19406) );
  INV_X1 U21578 ( .A(n19406), .ZN(U254) );
  NAND2_X1 U21579 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19531), .ZN(n19439) );
  NAND2_X1 U21580 ( .A1(n19531), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19445) );
  INV_X1 U21581 ( .A(n19445), .ZN(n19436) );
  AND2_X1 U21582 ( .A1(n19532), .A2(BUF2_REG_3__SCAN_IN), .ZN(n19440) );
  AOI22_X1 U21583 ( .A1(n19626), .A2(n19436), .B1(n19533), .B2(n19440), .ZN(
        n19409) );
  NOR2_X2 U21584 ( .A1(n19407), .A2(n19534), .ZN(n19442) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n19442), .ZN(n19408) );
  OAI211_X1 U21586 ( .C1(n19544), .C2(n19439), .A(n19409), .B(n19408), .ZN(
        P3_U2991) );
  INV_X1 U21587 ( .A(n19439), .ZN(n19441) );
  AOI22_X1 U21588 ( .A1(n19546), .A2(n19441), .B1(n19539), .B2(n19440), .ZN(
        n19411) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19442), .ZN(n19410) );
  OAI211_X1 U21590 ( .C1(n19544), .C2(n19445), .A(n19411), .B(n19410), .ZN(
        P3_U2983) );
  INV_X1 U21591 ( .A(n19558), .ZN(n19453) );
  AOI22_X1 U21592 ( .A1(n19565), .A2(n19441), .B1(n19545), .B2(n19440), .ZN(
        n19413) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19547), .B1(
        n19626), .B2(n19442), .ZN(n19412) );
  OAI211_X1 U21594 ( .C1(n19453), .C2(n19445), .A(n19413), .B(n19412), .ZN(
        P3_U2975) );
  AOI22_X1 U21595 ( .A1(n19570), .A2(n19441), .B1(n19551), .B2(n19440), .ZN(
        n19415) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19442), .ZN(n19414) );
  OAI211_X1 U21597 ( .C1(n19550), .C2(n19445), .A(n19415), .B(n19414), .ZN(
        P3_U2967) );
  AOI22_X1 U21598 ( .A1(n19570), .A2(n19436), .B1(n19557), .B2(n19440), .ZN(
        n19417) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19559), .B1(
        n19546), .B2(n19442), .ZN(n19416) );
  OAI211_X1 U21600 ( .C1(n19562), .C2(n19439), .A(n19417), .B(n19416), .ZN(
        P3_U2959) );
  AOI22_X1 U21601 ( .A1(n19582), .A2(n19441), .B1(n19563), .B2(n19440), .ZN(
        n19419) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19564), .B1(
        n19565), .B2(n19442), .ZN(n19418) );
  OAI211_X1 U21603 ( .C1(n19562), .C2(n19445), .A(n19419), .B(n19418), .ZN(
        P3_U2951) );
  AOI22_X1 U21604 ( .A1(n19582), .A2(n19436), .B1(n19569), .B2(n19440), .ZN(
        n19421) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19571), .B1(
        n19570), .B2(n19442), .ZN(n19420) );
  OAI211_X1 U21606 ( .C1(n19579), .C2(n19439), .A(n19421), .B(n19420), .ZN(
        P3_U2943) );
  AOI22_X1 U21607 ( .A1(n19587), .A2(n19436), .B1(n19574), .B2(n19440), .ZN(
        n19423) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19576), .B1(
        n19575), .B2(n19442), .ZN(n19422) );
  OAI211_X1 U21609 ( .C1(n19508), .C2(n19439), .A(n19423), .B(n19422), .ZN(
        P3_U2935) );
  AOI22_X1 U21610 ( .A1(n19599), .A2(n19441), .B1(n19580), .B2(n19440), .ZN(
        n19425) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19581), .B1(
        n19582), .B2(n19442), .ZN(n19424) );
  OAI211_X1 U21612 ( .C1(n19508), .C2(n19445), .A(n19425), .B(n19424), .ZN(
        P3_U2927) );
  AOI22_X1 U21613 ( .A1(n19599), .A2(n19436), .B1(n19586), .B2(n19440), .ZN(
        n19427) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19442), .ZN(n19426) );
  OAI211_X1 U21615 ( .C1(n19591), .C2(n19439), .A(n19427), .B(n19426), .ZN(
        P3_U2919) );
  AOI22_X1 U21616 ( .A1(n19605), .A2(n19436), .B1(n19592), .B2(n19440), .ZN(
        n19429) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19442), .ZN(n19428) );
  OAI211_X1 U21618 ( .C1(n19597), .C2(n19439), .A(n19429), .B(n19428), .ZN(
        P3_U2911) );
  AOI22_X1 U21619 ( .A1(n19610), .A2(n19436), .B1(n19598), .B2(n19440), .ZN(
        n19431) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19442), .ZN(n19430) );
  OAI211_X1 U21621 ( .C1(n19603), .C2(n19439), .A(n19431), .B(n19430), .ZN(
        P3_U2903) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19606), .B1(
        n19604), .B2(n19440), .ZN(n19433) );
  AOI22_X1 U21623 ( .A1(n19605), .A2(n19442), .B1(n19628), .B2(n19441), .ZN(
        n19432) );
  OAI211_X1 U21624 ( .C1(n19603), .C2(n19445), .A(n19433), .B(n19432), .ZN(
        P3_U2895) );
  AOI22_X1 U21625 ( .A1(n19617), .A2(n19441), .B1(n19609), .B2(n19440), .ZN(
        n19435) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19442), .ZN(n19434) );
  OAI211_X1 U21627 ( .C1(n19614), .C2(n19445), .A(n19435), .B(n19434), .ZN(
        P3_U2887) );
  AOI22_X1 U21628 ( .A1(n19617), .A2(n19436), .B1(n19615), .B2(n19440), .ZN(
        n19438) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19442), .ZN(n19437) );
  OAI211_X1 U21630 ( .C1(n19633), .C2(n19439), .A(n19438), .B(n19437), .ZN(
        P3_U2879) );
  AOI22_X1 U21631 ( .A1(n19626), .A2(n19441), .B1(n19624), .B2(n19440), .ZN(
        n19444) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19442), .ZN(n19443) );
  OAI211_X1 U21633 ( .C1(n19633), .C2(n19445), .A(n19444), .B(n19443), .ZN(
        P3_U2871) );
  OAI22_X1 U21634 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19487), .ZN(n19446) );
  INV_X1 U21635 ( .A(n19446), .ZN(U253) );
  NAND2_X1 U21636 ( .A1(n19531), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19486) );
  NAND2_X1 U21637 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19531), .ZN(n19477) );
  INV_X1 U21638 ( .A(n19477), .ZN(n19482) );
  AND2_X1 U21639 ( .A1(n19532), .A2(BUF2_REG_2__SCAN_IN), .ZN(n19481) );
  AOI22_X1 U21640 ( .A1(n19552), .A2(n19482), .B1(n19533), .B2(n19481), .ZN(
        n19448) );
  NOR2_X2 U21641 ( .A1(n21342), .A2(n19534), .ZN(n19483) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n19483), .ZN(n19447) );
  OAI211_X1 U21643 ( .C1(n19491), .C2(n19486), .A(n19448), .B(n19447), .ZN(
        P3_U2990) );
  INV_X1 U21644 ( .A(n19486), .ZN(n19474) );
  AOI22_X1 U21645 ( .A1(n19552), .A2(n19474), .B1(n19539), .B2(n19481), .ZN(
        n19450) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19483), .ZN(n19449) );
  OAI211_X1 U21647 ( .C1(n19453), .C2(n19477), .A(n19450), .B(n19449), .ZN(
        P3_U2982) );
  AOI22_X1 U21648 ( .A1(n19565), .A2(n19482), .B1(n19545), .B2(n19481), .ZN(
        n19452) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19547), .B1(
        n19626), .B2(n19483), .ZN(n19451) );
  OAI211_X1 U21650 ( .C1(n19453), .C2(n19486), .A(n19452), .B(n19451), .ZN(
        P3_U2974) );
  AOI22_X1 U21651 ( .A1(n19565), .A2(n19474), .B1(n19551), .B2(n19481), .ZN(
        n19455) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19483), .ZN(n19454) );
  OAI211_X1 U21653 ( .C1(n19556), .C2(n19477), .A(n19455), .B(n19454), .ZN(
        P3_U2966) );
  AOI22_X1 U21654 ( .A1(n19575), .A2(n19482), .B1(n19557), .B2(n19481), .ZN(
        n19457) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19559), .B1(
        n19558), .B2(n19483), .ZN(n19456) );
  OAI211_X1 U21656 ( .C1(n19556), .C2(n19486), .A(n19457), .B(n19456), .ZN(
        P3_U2958) );
  AOI22_X1 U21657 ( .A1(n19575), .A2(n19474), .B1(n19563), .B2(n19481), .ZN(
        n19459) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19564), .B1(
        n19565), .B2(n19483), .ZN(n19458) );
  OAI211_X1 U21659 ( .C1(n19568), .C2(n19477), .A(n19459), .B(n19458), .ZN(
        P3_U2950) );
  AOI22_X1 U21660 ( .A1(n19587), .A2(n19482), .B1(n19569), .B2(n19481), .ZN(
        n19461) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19571), .B1(
        n19570), .B2(n19483), .ZN(n19460) );
  OAI211_X1 U21662 ( .C1(n19568), .C2(n19486), .A(n19461), .B(n19460), .ZN(
        P3_U2942) );
  AOI22_X1 U21663 ( .A1(n19587), .A2(n19474), .B1(n19574), .B2(n19481), .ZN(
        n19463) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19576), .B1(
        n19575), .B2(n19483), .ZN(n19462) );
  OAI211_X1 U21665 ( .C1(n19508), .C2(n19477), .A(n19463), .B(n19462), .ZN(
        P3_U2934) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19581), .B1(
        n19580), .B2(n19481), .ZN(n19465) );
  AOI22_X1 U21667 ( .A1(n19582), .A2(n19483), .B1(n19593), .B2(n19474), .ZN(
        n19464) );
  OAI211_X1 U21668 ( .C1(n19585), .C2(n19477), .A(n19465), .B(n19464), .ZN(
        P3_U2926) );
  AOI22_X1 U21669 ( .A1(n19605), .A2(n19482), .B1(n19586), .B2(n19481), .ZN(
        n19467) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19483), .ZN(n19466) );
  OAI211_X1 U21671 ( .C1(n19585), .C2(n19486), .A(n19467), .B(n19466), .ZN(
        P3_U2918) );
  AOI22_X1 U21672 ( .A1(n19610), .A2(n19482), .B1(n19592), .B2(n19481), .ZN(
        n19469) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19483), .ZN(n19468) );
  OAI211_X1 U21674 ( .C1(n19591), .C2(n19486), .A(n19469), .B(n19468), .ZN(
        P3_U2910) );
  AOI22_X1 U21675 ( .A1(n19610), .A2(n19474), .B1(n19598), .B2(n19481), .ZN(
        n19471) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19483), .ZN(n19470) );
  OAI211_X1 U21677 ( .C1(n19603), .C2(n19477), .A(n19471), .B(n19470), .ZN(
        P3_U2902) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19606), .B1(
        n19604), .B2(n19481), .ZN(n19473) );
  AOI22_X1 U21679 ( .A1(n19605), .A2(n19483), .B1(n19628), .B2(n19482), .ZN(
        n19472) );
  OAI211_X1 U21680 ( .C1(n19603), .C2(n19486), .A(n19473), .B(n19472), .ZN(
        P3_U2894) );
  AOI22_X1 U21681 ( .A1(n19628), .A2(n19474), .B1(n19609), .B2(n19481), .ZN(
        n19476) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19483), .ZN(n19475) );
  OAI211_X1 U21683 ( .C1(n19480), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        P3_U2886) );
  AOI22_X1 U21684 ( .A1(n19540), .A2(n19482), .B1(n19615), .B2(n19481), .ZN(
        n19479) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19483), .ZN(n19478) );
  OAI211_X1 U21686 ( .C1(n19480), .C2(n19486), .A(n19479), .B(n19478), .ZN(
        P3_U2878) );
  AOI22_X1 U21687 ( .A1(n19626), .A2(n19482), .B1(n19624), .B2(n19481), .ZN(
        n19485) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19483), .ZN(n19484) );
  OAI211_X1 U21689 ( .C1(n19633), .C2(n19486), .A(n19485), .B(n19484), .ZN(
        P3_U2870) );
  OAI22_X1 U21690 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19487), .ZN(n19488) );
  INV_X1 U21691 ( .A(n19488), .ZN(U252) );
  NAND2_X1 U21692 ( .A1(n19531), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19528) );
  NAND2_X1 U21693 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19531), .ZN(n19522) );
  INV_X1 U21694 ( .A(n19522), .ZN(n19524) );
  AND2_X1 U21695 ( .A1(n19532), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19523) );
  AOI22_X1 U21696 ( .A1(n19552), .A2(n19524), .B1(n19533), .B2(n19523), .ZN(
        n19490) );
  NOR2_X2 U21697 ( .A1(n20665), .A2(n19534), .ZN(n19525) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n19525), .ZN(n19489) );
  OAI211_X1 U21699 ( .C1(n19491), .C2(n19528), .A(n19490), .B(n19489), .ZN(
        P3_U2989) );
  AOI22_X1 U21700 ( .A1(n19546), .A2(n19524), .B1(n19539), .B2(n19523), .ZN(
        n19493) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19525), .ZN(n19492) );
  OAI211_X1 U21702 ( .C1(n19544), .C2(n19528), .A(n19493), .B(n19492), .ZN(
        P3_U2981) );
  INV_X1 U21703 ( .A(n19528), .ZN(n19519) );
  AOI22_X1 U21704 ( .A1(n19546), .A2(n19519), .B1(n19545), .B2(n19523), .ZN(
        n19495) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19547), .B1(
        n19626), .B2(n19525), .ZN(n19494) );
  OAI211_X1 U21706 ( .C1(n19550), .C2(n19522), .A(n19495), .B(n19494), .ZN(
        P3_U2973) );
  AOI22_X1 U21707 ( .A1(n19570), .A2(n19524), .B1(n19551), .B2(n19523), .ZN(
        n19497) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19525), .ZN(n19496) );
  OAI211_X1 U21709 ( .C1(n19550), .C2(n19528), .A(n19497), .B(n19496), .ZN(
        P3_U2965) );
  AOI22_X1 U21710 ( .A1(n19575), .A2(n19524), .B1(n19557), .B2(n19523), .ZN(
        n19499) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19559), .B1(
        n19546), .B2(n19525), .ZN(n19498) );
  OAI211_X1 U21712 ( .C1(n19556), .C2(n19528), .A(n19499), .B(n19498), .ZN(
        P3_U2957) );
  AOI22_X1 U21713 ( .A1(n19575), .A2(n19519), .B1(n19563), .B2(n19523), .ZN(
        n19501) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19564), .B1(
        n19565), .B2(n19525), .ZN(n19500) );
  OAI211_X1 U21715 ( .C1(n19568), .C2(n19522), .A(n19501), .B(n19500), .ZN(
        P3_U2949) );
  AOI22_X1 U21716 ( .A1(n19582), .A2(n19519), .B1(n19569), .B2(n19523), .ZN(
        n19503) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19571), .B1(
        n19570), .B2(n19525), .ZN(n19502) );
  OAI211_X1 U21718 ( .C1(n19579), .C2(n19522), .A(n19503), .B(n19502), .ZN(
        P3_U2941) );
  AOI22_X1 U21719 ( .A1(n19587), .A2(n19519), .B1(n19574), .B2(n19523), .ZN(
        n19505) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19576), .B1(
        n19575), .B2(n19525), .ZN(n19504) );
  OAI211_X1 U21721 ( .C1(n19508), .C2(n19522), .A(n19505), .B(n19504), .ZN(
        P3_U2933) );
  AOI22_X1 U21722 ( .A1(n19599), .A2(n19524), .B1(n19580), .B2(n19523), .ZN(
        n19507) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19581), .B1(
        n19582), .B2(n19525), .ZN(n19506) );
  OAI211_X1 U21724 ( .C1(n19508), .C2(n19528), .A(n19507), .B(n19506), .ZN(
        P3_U2925) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19588), .B1(
        n19586), .B2(n19523), .ZN(n19510) );
  AOI22_X1 U21726 ( .A1(n19587), .A2(n19525), .B1(n19605), .B2(n19524), .ZN(
        n19509) );
  OAI211_X1 U21727 ( .C1(n19585), .C2(n19528), .A(n19510), .B(n19509), .ZN(
        P3_U2917) );
  AOI22_X1 U21728 ( .A1(n19610), .A2(n19524), .B1(n19592), .B2(n19523), .ZN(
        n19512) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19525), .ZN(n19511) );
  OAI211_X1 U21730 ( .C1(n19591), .C2(n19528), .A(n19512), .B(n19511), .ZN(
        P3_U2909) );
  AOI22_X1 U21731 ( .A1(n19610), .A2(n19519), .B1(n19598), .B2(n19523), .ZN(
        n19514) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19525), .ZN(n19513) );
  OAI211_X1 U21733 ( .C1(n19603), .C2(n19522), .A(n19514), .B(n19513), .ZN(
        P3_U2901) );
  AOI22_X1 U21734 ( .A1(n19618), .A2(n19519), .B1(n19604), .B2(n19523), .ZN(
        n19516) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19525), .ZN(n19515) );
  OAI211_X1 U21736 ( .C1(n19614), .C2(n19522), .A(n19516), .B(n19515), .ZN(
        P3_U2893) );
  AOI22_X1 U21737 ( .A1(n19617), .A2(n19524), .B1(n19609), .B2(n19523), .ZN(
        n19518) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19525), .ZN(n19517) );
  OAI211_X1 U21739 ( .C1(n19614), .C2(n19528), .A(n19518), .B(n19517), .ZN(
        P3_U2885) );
  AOI22_X1 U21740 ( .A1(n19617), .A2(n19519), .B1(n19615), .B2(n19523), .ZN(
        n19521) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19525), .ZN(n19520) );
  OAI211_X1 U21742 ( .C1(n19633), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P3_U2877) );
  AOI22_X1 U21743 ( .A1(n19626), .A2(n19524), .B1(n19624), .B2(n19523), .ZN(
        n19527) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19525), .ZN(n19526) );
  OAI211_X1 U21745 ( .C1(n19633), .C2(n19528), .A(n19527), .B(n19526), .ZN(
        P3_U2869) );
  OAI22_X1 U21746 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19529), .ZN(n19530) );
  INV_X1 U21747 ( .A(n19530), .ZN(U251) );
  NAND2_X1 U21748 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19531), .ZN(n19622) );
  NAND2_X1 U21749 ( .A1(n19531), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19632) );
  INV_X1 U21750 ( .A(n19632), .ZN(n19616) );
  AND2_X1 U21751 ( .A1(n19532), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19623) );
  AOI22_X1 U21752 ( .A1(n19626), .A2(n19616), .B1(n19533), .B2(n19623), .ZN(
        n19538) );
  NOR2_X2 U21753 ( .A1(n19535), .A2(n19534), .ZN(n19627) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19536), .B1(
        n19617), .B2(n19627), .ZN(n19537) );
  OAI211_X1 U21755 ( .C1(n19544), .C2(n19622), .A(n19538), .B(n19537), .ZN(
        P3_U2988) );
  INV_X1 U21756 ( .A(n19622), .ZN(n19625) );
  AOI22_X1 U21757 ( .A1(n19546), .A2(n19625), .B1(n19539), .B2(n19623), .ZN(
        n19543) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19627), .ZN(n19542) );
  OAI211_X1 U21759 ( .C1(n19544), .C2(n19632), .A(n19543), .B(n19542), .ZN(
        P3_U2980) );
  AOI22_X1 U21760 ( .A1(n19546), .A2(n19616), .B1(n19545), .B2(n19623), .ZN(
        n19549) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19547), .B1(
        n19626), .B2(n19627), .ZN(n19548) );
  OAI211_X1 U21762 ( .C1(n19550), .C2(n19622), .A(n19549), .B(n19548), .ZN(
        P3_U2972) );
  AOI22_X1 U21763 ( .A1(n19565), .A2(n19616), .B1(n19551), .B2(n19623), .ZN(
        n19555) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19627), .ZN(n19554) );
  OAI211_X1 U21765 ( .C1(n19556), .C2(n19622), .A(n19555), .B(n19554), .ZN(
        P3_U2964) );
  AOI22_X1 U21766 ( .A1(n19570), .A2(n19616), .B1(n19557), .B2(n19623), .ZN(
        n19561) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19559), .B1(
        n19558), .B2(n19627), .ZN(n19560) );
  OAI211_X1 U21768 ( .C1(n19562), .C2(n19622), .A(n19561), .B(n19560), .ZN(
        P3_U2956) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19564), .B1(
        n19563), .B2(n19623), .ZN(n19567) );
  AOI22_X1 U21770 ( .A1(n19565), .A2(n19627), .B1(n19575), .B2(n19616), .ZN(
        n19566) );
  OAI211_X1 U21771 ( .C1(n19568), .C2(n19622), .A(n19567), .B(n19566), .ZN(
        P3_U2948) );
  AOI22_X1 U21772 ( .A1(n19582), .A2(n19616), .B1(n19569), .B2(n19623), .ZN(
        n19573) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19571), .B1(
        n19570), .B2(n19627), .ZN(n19572) );
  OAI211_X1 U21774 ( .C1(n19579), .C2(n19622), .A(n19573), .B(n19572), .ZN(
        P3_U2940) );
  AOI22_X1 U21775 ( .A1(n19593), .A2(n19625), .B1(n19574), .B2(n19623), .ZN(
        n19578) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19576), .B1(
        n19575), .B2(n19627), .ZN(n19577) );
  OAI211_X1 U21777 ( .C1(n19579), .C2(n19632), .A(n19578), .B(n19577), .ZN(
        P3_U2932) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19581), .B1(
        n19580), .B2(n19623), .ZN(n19584) );
  AOI22_X1 U21779 ( .A1(n19582), .A2(n19627), .B1(n19593), .B2(n19616), .ZN(
        n19583) );
  OAI211_X1 U21780 ( .C1(n19585), .C2(n19622), .A(n19584), .B(n19583), .ZN(
        P3_U2924) );
  AOI22_X1 U21781 ( .A1(n19599), .A2(n19616), .B1(n19586), .B2(n19623), .ZN(
        n19590) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19588), .B1(
        n19587), .B2(n19627), .ZN(n19589) );
  OAI211_X1 U21783 ( .C1(n19591), .C2(n19622), .A(n19590), .B(n19589), .ZN(
        P3_U2916) );
  AOI22_X1 U21784 ( .A1(n19605), .A2(n19616), .B1(n19592), .B2(n19623), .ZN(
        n19596) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19594), .B1(
        n19593), .B2(n19627), .ZN(n19595) );
  OAI211_X1 U21786 ( .C1(n19597), .C2(n19622), .A(n19596), .B(n19595), .ZN(
        P3_U2908) );
  AOI22_X1 U21787 ( .A1(n19610), .A2(n19616), .B1(n19598), .B2(n19623), .ZN(
        n19602) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19600), .B1(
        n19599), .B2(n19627), .ZN(n19601) );
  OAI211_X1 U21789 ( .C1(n19603), .C2(n19622), .A(n19602), .B(n19601), .ZN(
        P3_U2900) );
  AOI22_X1 U21790 ( .A1(n19618), .A2(n19616), .B1(n19604), .B2(n19623), .ZN(
        n19608) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19606), .B1(
        n19605), .B2(n19627), .ZN(n19607) );
  OAI211_X1 U21792 ( .C1(n19614), .C2(n19622), .A(n19608), .B(n19607), .ZN(
        P3_U2892) );
  AOI22_X1 U21793 ( .A1(n19617), .A2(n19625), .B1(n19609), .B2(n19623), .ZN(
        n19613) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19627), .ZN(n19612) );
  OAI211_X1 U21795 ( .C1(n19614), .C2(n19632), .A(n19613), .B(n19612), .ZN(
        P3_U2884) );
  AOI22_X1 U21796 ( .A1(n19617), .A2(n19616), .B1(n19615), .B2(n19623), .ZN(
        n19621) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19619), .B1(
        n19618), .B2(n19627), .ZN(n19620) );
  OAI211_X1 U21798 ( .C1(n19633), .C2(n19622), .A(n19621), .B(n19620), .ZN(
        P3_U2876) );
  AOI22_X1 U21799 ( .A1(n19626), .A2(n19625), .B1(n19624), .B2(n19623), .ZN(
        n19631) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19629), .B1(
        n19628), .B2(n19627), .ZN(n19630) );
  OAI211_X1 U21801 ( .C1(n19633), .C2(n19632), .A(n19631), .B(n19630), .ZN(
        P3_U2868) );
  OAI222_X1 U21802 ( .A1(n19636), .A2(n19910), .B1(n19635), .B2(n20162), .C1(
        n19634), .C2(n20173), .ZN(P2_U2904) );
  OAI222_X1 U21803 ( .A1(n19639), .A2(n19910), .B1(n19638), .B2(n20162), .C1(
        n20173), .C2(n19637), .ZN(P2_U2905) );
  OAI222_X1 U21804 ( .A1(n19642), .A2(n19910), .B1(n19641), .B2(n20162), .C1(
        n20173), .C2(n19640), .ZN(P2_U2906) );
  AOI22_X1 U21805 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n20110), .B1(n19644), 
        .B2(n19643), .ZN(n19645) );
  OAI21_X1 U21806 ( .B1(n19910), .B2(n19646), .A(n19645), .ZN(P2_U2907) );
  OAI222_X1 U21807 ( .A1(n19649), .A2(n19910), .B1(n19648), .B2(n20162), .C1(
        n20173), .C2(n19647), .ZN(P2_U2908) );
  INV_X1 U21808 ( .A(n19650), .ZN(n19653) );
  OAI222_X1 U21809 ( .A1(n19653), .A2(n19910), .B1(n19652), .B2(n20162), .C1(
        n20173), .C2(n19651), .ZN(P2_U2909) );
  OAI222_X1 U21810 ( .A1(n19656), .A2(n19910), .B1(n19655), .B2(n20162), .C1(
        n20173), .C2(n19654), .ZN(P2_U2910) );
  INV_X1 U21811 ( .A(n19657), .ZN(n19660) );
  OAI222_X1 U21812 ( .A1(n19660), .A2(n19910), .B1(n19659), .B2(n20162), .C1(
        n20173), .C2(n19658), .ZN(P2_U2911) );
  OAI222_X1 U21813 ( .A1(n19663), .A2(n19910), .B1(n19662), .B2(n20162), .C1(
        n20173), .C2(n19661), .ZN(P2_U2912) );
  NAND3_X1 U21814 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19677) );
  NOR2_X1 U21815 ( .A1(n19664), .A2(n19786), .ZN(n20178) );
  OAI21_X1 U21816 ( .B1(n19668), .B2(n20178), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19665) );
  OAI21_X1 U21817 ( .B1(n19677), .B2(n19838), .A(n19665), .ZN(n20179) );
  AOI22_X1 U21818 ( .A1(n20179), .A2(n15675), .B1(n19836), .B2(n20178), .ZN(
        n19673) );
  INV_X1 U21819 ( .A(n19667), .ZN(n19744) );
  OAI21_X1 U21820 ( .B1(n19691), .B2(n19744), .A(n19677), .ZN(n19671) );
  INV_X1 U21821 ( .A(n20178), .ZN(n19844) );
  NAND2_X1 U21822 ( .A1(n19668), .A2(n19842), .ZN(n19669) );
  OAI211_X1 U21823 ( .C1(n20174), .C2(n19844), .A(n19669), .B(n19799), .ZN(
        n19670) );
  NAND2_X1 U21824 ( .A1(n19671), .A2(n19670), .ZN(n20182) );
  AOI22_X1 U21825 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n19837), .ZN(n19672) );
  OAI211_X1 U21826 ( .C1(n19853), .C2(n20289), .A(n19673), .B(n19672), .ZN(
        P2_U3175) );
  INV_X1 U21827 ( .A(n15675), .ZN(n19806) );
  INV_X1 U21828 ( .A(n20186), .ZN(n19675) );
  NAND3_X1 U21829 ( .A1(n19920), .A2(n19675), .A3(n19788), .ZN(n19676) );
  INV_X1 U21830 ( .A(n19839), .ZN(n19731) );
  NAND2_X1 U21831 ( .A1(n19676), .A2(n19731), .ZN(n19685) );
  INV_X1 U21832 ( .A(n19682), .ZN(n19678) );
  NOR2_X1 U21833 ( .A1(n19677), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20185) );
  INV_X1 U21834 ( .A(n20185), .ZN(n19679) );
  AOI21_X1 U21835 ( .B1(n19678), .B2(n19679), .A(n19734), .ZN(n19681) );
  NOR2_X1 U21836 ( .A1(n19819), .A2(n19692), .ZN(n20191) );
  INV_X1 U21837 ( .A(n20191), .ZN(n19684) );
  NAND2_X1 U21838 ( .A1(n19679), .A2(n19684), .ZN(n19680) );
  AOI22_X1 U21839 ( .A1(n19803), .A2(n20186), .B1(n19836), .B2(n20185), .ZN(
        n19688) );
  AOI21_X1 U21840 ( .B1(n19682), .B2(n19842), .A(n19841), .ZN(n19683) );
  AOI21_X1 U21841 ( .B1(n19685), .B2(n19684), .A(n19683), .ZN(n19686) );
  AOI22_X1 U21842 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20187), .B1(
        n20193), .B2(n19837), .ZN(n19687) );
  OAI211_X1 U21843 ( .C1(n19806), .C2(n20190), .A(n19688), .B(n19687), .ZN(
        P2_U3167) );
  OAI21_X1 U21844 ( .B1(n12994), .B2(n20191), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19689) );
  OAI21_X1 U21845 ( .B1(n19692), .B2(n19838), .A(n19689), .ZN(n20192) );
  AOI22_X1 U21846 ( .A1(n20192), .A2(n15675), .B1(n19836), .B2(n20191), .ZN(
        n19699) );
  OR2_X1 U21847 ( .A1(n19690), .A2(n22169), .ZN(n19827) );
  NOR2_X1 U21848 ( .A1(n19691), .A2(n19827), .ZN(n19697) );
  INV_X1 U21849 ( .A(n19692), .ZN(n19696) );
  INV_X1 U21850 ( .A(n12994), .ZN(n19694) );
  OAI21_X1 U21851 ( .B1(n19788), .B2(n20191), .A(n19846), .ZN(n19693) );
  OAI21_X1 U21852 ( .B1(n19694), .B2(n19823), .A(n19693), .ZN(n19695) );
  OAI21_X1 U21853 ( .B1(n19697), .B2(n19696), .A(n19695), .ZN(n20194) );
  AOI22_X1 U21854 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20194), .B1(
        n20200), .B2(n19837), .ZN(n19698) );
  OAI211_X1 U21855 ( .C1(n19853), .C2(n19920), .A(n19699), .B(n19698), .ZN(
        P2_U3159) );
  NAND3_X1 U21856 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19787), .ZN(n19709) );
  NOR2_X1 U21857 ( .A1(n19819), .A2(n19709), .ZN(n20205) );
  OAI21_X1 U21858 ( .B1(n13027), .B2(n20205), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19700) );
  OAI21_X1 U21859 ( .B1(n19709), .B2(n19838), .A(n19700), .ZN(n20206) );
  AOI22_X1 U21860 ( .A1(n20206), .A2(n15675), .B1(n19836), .B2(n20205), .ZN(
        n19708) );
  INV_X1 U21861 ( .A(n20205), .ZN(n19701) );
  AOI21_X1 U21862 ( .B1(n19701), .B2(n19838), .A(n20174), .ZN(n19706) );
  NOR2_X1 U21863 ( .A1(n19702), .A2(n19823), .ZN(n19705) );
  OAI21_X1 U21864 ( .B1(n19795), .B2(n19703), .A(n19709), .ZN(n19704) );
  OAI21_X1 U21865 ( .B1(n19706), .B2(n19705), .A(n19704), .ZN(n20207) );
  AOI22_X1 U21866 ( .A1(n19837), .A2(n20130), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n20207), .ZN(n19707) );
  OAI211_X1 U21867 ( .C1(n19853), .C2(n20204), .A(n19708), .B(n19707), .ZN(
        P2_U3143) );
  NOR2_X1 U21868 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19709), .ZN(
        n20211) );
  AOI22_X1 U21869 ( .A1(n19837), .A2(n20212), .B1(n19836), .B2(n20211), .ZN(
        n19717) );
  NOR3_X1 U21870 ( .A1(n12995), .A2(n20211), .A3(n19734), .ZN(n19712) );
  OAI21_X1 U21871 ( .B1(n20212), .B2(n20130), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19710) );
  NAND2_X1 U21872 ( .A1(n19710), .A2(n19788), .ZN(n19715) );
  NAND3_X1 U21873 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19807), .A3(
        n19787), .ZN(n19730) );
  NOR2_X1 U21874 ( .A1(n19819), .A2(n19730), .ZN(n20218) );
  NOR2_X1 U21875 ( .A1(n20218), .A2(n20211), .ZN(n19714) );
  OAI21_X1 U21876 ( .B1(n12995), .B2(n20211), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19713) );
  AOI22_X1 U21877 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20214), .B1(
        n15675), .B2(n20213), .ZN(n19716) );
  OAI211_X1 U21878 ( .C1(n19853), .C2(n20217), .A(n19717), .B(n19716), .ZN(
        P2_U3135) );
  AOI22_X1 U21879 ( .A1(n19837), .A2(n20225), .B1(n19836), .B2(n20218), .ZN(
        n19728) );
  OAI21_X1 U21880 ( .B1(n19720), .B2(n19827), .A(n19788), .ZN(n19726) );
  INV_X1 U21881 ( .A(n19730), .ZN(n19724) );
  INV_X1 U21882 ( .A(n20218), .ZN(n19722) );
  NAND2_X1 U21883 ( .A1(n12985), .A2(n19842), .ZN(n19721) );
  OAI211_X1 U21884 ( .C1(n20174), .C2(n19722), .A(n19721), .B(n19799), .ZN(
        n19723) );
  OAI21_X1 U21885 ( .B1(n19726), .B2(n19724), .A(n19723), .ZN(n20220) );
  OAI21_X1 U21886 ( .B1(n12985), .B2(n20218), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19725) );
  OAI21_X1 U21887 ( .B1(n19726), .B2(n19730), .A(n19725), .ZN(n20219) );
  AOI22_X1 U21888 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20220), .B1(
        n15675), .B2(n20219), .ZN(n19727) );
  OAI211_X1 U21889 ( .C1(n19853), .C2(n20223), .A(n19728), .B(n19727), .ZN(
        P2_U3127) );
  NOR2_X1 U21890 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19730), .ZN(
        n20224) );
  AOI22_X1 U21891 ( .A1(n19837), .A2(n20233), .B1(n19836), .B2(n20224), .ZN(
        n19741) );
  NAND2_X1 U21892 ( .A1(n20137), .A2(n19788), .ZN(n19732) );
  OAI21_X1 U21893 ( .B1(n19732), .B2(n20233), .A(n19731), .ZN(n19737) );
  OAI21_X1 U21894 ( .B1(n12983), .B2(n19734), .A(n19733), .ZN(n19735) );
  AOI21_X1 U21895 ( .B1(n19737), .B2(n19746), .A(n19735), .ZN(n19736) );
  INV_X1 U21896 ( .A(n19746), .ZN(n20231) );
  OAI21_X1 U21897 ( .B1(n20231), .B2(n20224), .A(n19737), .ZN(n19739) );
  OAI21_X1 U21898 ( .B1(n12983), .B2(n20224), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19738) );
  NAND2_X1 U21899 ( .A1(n19739), .A2(n19738), .ZN(n20226) );
  AOI22_X1 U21900 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n15675), .ZN(n19740) );
  OAI211_X1 U21901 ( .C1(n19853), .C2(n20137), .A(n19741), .B(n19740), .ZN(
        P2_U3119) );
  NAND2_X1 U21902 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19769), .ZN(
        n19743) );
  OAI21_X1 U21903 ( .B1(n19745), .B2(n20231), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19742) );
  OAI21_X1 U21904 ( .B1(n19743), .B2(n19838), .A(n19742), .ZN(n20232) );
  AOI22_X1 U21905 ( .A1(n20232), .A2(n15675), .B1(n20231), .B2(n19836), .ZN(
        n19752) );
  OAI22_X1 U21906 ( .A1(n19766), .A2(n19744), .B1(n19807), .B2(n19757), .ZN(
        n19749) );
  INV_X1 U21907 ( .A(n19745), .ZN(n19747) );
  OAI211_X1 U21908 ( .C1(n19747), .C2(n19823), .A(n19746), .B(n19838), .ZN(
        n19748) );
  NAND3_X1 U21909 ( .A1(n19749), .A2(n19846), .A3(n19748), .ZN(n20234) );
  AOI22_X1 U21910 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20234), .B1(
        n20138), .B2(n19837), .ZN(n19751) );
  OAI211_X1 U21911 ( .C1(n19853), .C2(n20230), .A(n19752), .B(n19751), .ZN(
        P2_U3111) );
  NOR3_X2 U21912 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19807), .A3(
        n19757), .ZN(n20237) );
  OAI21_X1 U21913 ( .B1(n19759), .B2(n20237), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19753) );
  OAI21_X1 U21914 ( .B1(n19757), .B2(n19810), .A(n19753), .ZN(n20238) );
  AOI22_X1 U21915 ( .A1(n20238), .A2(n15675), .B1(n19836), .B2(n20237), .ZN(
        n19765) );
  INV_X1 U21916 ( .A(n19754), .ZN(n19758) );
  NOR2_X2 U21917 ( .A1(n19766), .A2(n19755), .ZN(n20239) );
  OAI21_X1 U21918 ( .B1(n20239), .B2(n20138), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19756) );
  OAI21_X1 U21919 ( .B1(n19758), .B2(n19757), .A(n19756), .ZN(n19763) );
  INV_X1 U21920 ( .A(n20237), .ZN(n19761) );
  NAND2_X1 U21921 ( .A1(n19759), .A2(n19842), .ZN(n19760) );
  OAI211_X1 U21922 ( .C1(n20174), .C2(n19761), .A(n19760), .B(n19799), .ZN(
        n19762) );
  NAND2_X1 U21923 ( .A1(n19763), .A2(n19762), .ZN(n20240) );
  AOI22_X1 U21924 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n19837), .ZN(n19764) );
  OAI211_X1 U21925 ( .C1(n19853), .C2(n20243), .A(n19765), .B(n19764), .ZN(
        P2_U3103) );
  INV_X1 U21926 ( .A(n19766), .ZN(n19768) );
  INV_X1 U21927 ( .A(n19827), .ZN(n19767) );
  NAND2_X1 U21928 ( .A1(n19768), .A2(n19767), .ZN(n19770) );
  NAND2_X1 U21929 ( .A1(n19769), .A2(n19807), .ZN(n19775) );
  NAND2_X1 U21930 ( .A1(n19770), .A2(n19775), .ZN(n19774) );
  NAND2_X1 U21931 ( .A1(n19777), .A2(n19842), .ZN(n19772) );
  NOR2_X1 U21932 ( .A1(n19819), .A2(n19775), .ZN(n20244) );
  OAI21_X1 U21933 ( .B1(n19788), .B2(n20244), .A(n19846), .ZN(n19771) );
  NAND2_X1 U21934 ( .A1(n19772), .A2(n19771), .ZN(n19773) );
  INV_X1 U21935 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U21936 ( .A1(n19803), .A2(n20239), .B1(n19836), .B2(n20244), .ZN(
        n19781) );
  INV_X1 U21937 ( .A(n19775), .ZN(n19776) );
  NAND2_X1 U21938 ( .A1(n19776), .A2(n19788), .ZN(n19779) );
  OAI21_X1 U21939 ( .B1(n19777), .B2(n20244), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19778) );
  NAND2_X1 U21940 ( .A1(n19779), .A2(n19778), .ZN(n20245) );
  AOI22_X1 U21941 ( .A1(n15675), .A2(n20245), .B1(n20251), .B2(n19837), .ZN(
        n19780) );
  OAI211_X1 U21942 ( .C1(n20039), .C2(n19782), .A(n19781), .B(n19780), .ZN(
        P2_U3095) );
  INV_X1 U21943 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U21944 ( .A1(n19803), .A2(n20251), .B1(n19836), .B2(n20250), .ZN(
        n19784) );
  AOI22_X1 U21945 ( .A1(n15675), .A2(n20252), .B1(n20259), .B2(n19837), .ZN(
        n19783) );
  OAI211_X1 U21946 ( .C1(n20256), .C2(n19785), .A(n19784), .B(n19783), .ZN(
        P2_U3087) );
  NAND2_X1 U21947 ( .A1(n19787), .A2(n19786), .ZN(n19834) );
  NOR2_X1 U21948 ( .A1(n19807), .A2(n19834), .ZN(n19793) );
  NAND2_X1 U21949 ( .A1(n19793), .A2(n19788), .ZN(n19791) );
  NOR2_X1 U21950 ( .A1(n19789), .A2(n19834), .ZN(n20257) );
  OAI21_X1 U21951 ( .B1(n19798), .B2(n20257), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19790) );
  AOI22_X1 U21952 ( .A1(n19837), .A2(n20258), .B1(n19836), .B2(n20257), .ZN(
        n19805) );
  INV_X1 U21953 ( .A(n19793), .ZN(n19797) );
  NAND2_X1 U21954 ( .A1(n19795), .A2(n19794), .ZN(n19796) );
  NAND2_X1 U21955 ( .A1(n19797), .A2(n19796), .ZN(n19802) );
  AOI21_X1 U21956 ( .B1(n19798), .B2(n19842), .A(n20257), .ZN(n19800) );
  OAI21_X1 U21957 ( .B1(n19800), .B2(n20174), .A(n19799), .ZN(n19801) );
  NAND2_X1 U21958 ( .A1(n19802), .A2(n19801), .ZN(n20260) );
  AOI22_X1 U21959 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20260), .B1(
        n20259), .B2(n19803), .ZN(n19804) );
  OAI211_X1 U21960 ( .C1(n20264), .C2(n19806), .A(n19805), .B(n19804), .ZN(
        P2_U3079) );
  NOR3_X2 U21961 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19807), .A3(
        n19834), .ZN(n20265) );
  OAI21_X1 U21962 ( .B1(n12993), .B2(n20265), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19808) );
  OAI21_X1 U21963 ( .B1(n19834), .B2(n19810), .A(n19808), .ZN(n20266) );
  AOI22_X1 U21964 ( .A1(n20266), .A2(n15675), .B1(n19836), .B2(n20265), .ZN(
        n19818) );
  OR2_X1 U21965 ( .A1(n19810), .A2(n19834), .ZN(n19811) );
  OAI221_X1 U21966 ( .B1(n22169), .B2(n20053), .C1(n22169), .C2(n20271), .A(
        n19811), .ZN(n19815) );
  INV_X1 U21967 ( .A(n12993), .ZN(n19813) );
  INV_X1 U21968 ( .A(n20265), .ZN(n19812) );
  OAI21_X1 U21969 ( .B1(n19813), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19812), 
        .ZN(n19814) );
  MUX2_X1 U21970 ( .A(n19815), .B(n19814), .S(n19838), .Z(n19816) );
  NAND2_X1 U21971 ( .A1(n19816), .A2(n19846), .ZN(n20268) );
  AOI22_X1 U21972 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n19837), .ZN(n19817) );
  OAI211_X1 U21973 ( .C1(n19853), .C2(n20271), .A(n19818), .B(n19817), .ZN(
        P2_U3071) );
  OR2_X1 U21974 ( .A1(n19834), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19826) );
  NOR2_X1 U21975 ( .A1(n19819), .A2(n19826), .ZN(n20273) );
  OAI21_X1 U21976 ( .B1(n12982), .B2(n20273), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19820) );
  OAI21_X1 U21977 ( .B1(n19826), .B2(n19838), .A(n19820), .ZN(n20274) );
  AOI22_X1 U21978 ( .A1(n20274), .A2(n15675), .B1(n19836), .B2(n20273), .ZN(
        n19833) );
  INV_X1 U21979 ( .A(n20273), .ZN(n19822) );
  AOI21_X1 U21980 ( .B1(n19822), .B2(n19838), .A(n20174), .ZN(n19831) );
  NOR2_X1 U21981 ( .A1(n19824), .A2(n19823), .ZN(n19830) );
  INV_X1 U21982 ( .A(n19825), .ZN(n19828) );
  OAI21_X1 U21983 ( .B1(n19828), .B2(n19827), .A(n19826), .ZN(n19829) );
  OAI21_X1 U21984 ( .B1(n19831), .B2(n19830), .A(n19829), .ZN(n20275) );
  AOI22_X1 U21985 ( .A1(n19837), .A2(n20282), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n20275), .ZN(n19832) );
  OAI211_X1 U21986 ( .C1(n19853), .C2(n20053), .A(n19833), .B(n19832), .ZN(
        P2_U3063) );
  NOR2_X1 U21987 ( .A1(n19835), .A2(n19834), .ZN(n20280) );
  AOI22_X1 U21988 ( .A1(n19837), .A2(n20155), .B1(n19836), .B2(n20280), .ZN(
        n19852) );
  NOR3_X1 U21989 ( .A1(n20282), .A2(n20155), .A3(n19838), .ZN(n19840) );
  NOR2_X1 U21990 ( .A1(n19840), .A2(n19839), .ZN(n19850) );
  INV_X1 U21991 ( .A(n19850), .ZN(n19845) );
  AOI21_X1 U21992 ( .B1(n12992), .B2(n19842), .A(n19841), .ZN(n19843) );
  AOI21_X1 U21993 ( .B1(n19845), .B2(n19844), .A(n19843), .ZN(n19847) );
  NOR2_X1 U21994 ( .A1(n20178), .A2(n20280), .ZN(n19849) );
  OAI21_X1 U21995 ( .B1(n12992), .B2(n20280), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19848) );
  AOI22_X1 U21996 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20286), .B1(
        n15675), .B2(n20285), .ZN(n19851) );
  OAI211_X1 U21997 ( .C1(n19853), .C2(n20279), .A(n19852), .B(n19851), .ZN(
        P2_U3055) );
  AOI22_X1 U21998 ( .A1(n19955), .A2(n19854), .B1(n20110), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n19860) );
  AOI22_X1 U21999 ( .A1(n19957), .A2(BUF1_REG_22__SCAN_IN), .B1(n19956), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n19859) );
  INV_X1 U22000 ( .A(n19855), .ZN(n19857) );
  AOI22_X1 U22001 ( .A1(n19857), .A2(n20167), .B1(n20112), .B2(n19856), .ZN(
        n19858) );
  NAND3_X1 U22002 ( .A1(n19860), .A2(n19859), .A3(n19858), .ZN(P2_U2897) );
  OAI222_X1 U22003 ( .A1(n19863), .A2(n19910), .B1(n19862), .B2(n20162), .C1(
        n20173), .C2(n19861), .ZN(P2_U2913) );
  AOI22_X1 U22004 ( .A1(n20179), .A2(n15648), .B1(n19898), .B2(n20178), .ZN(
        n19866) );
  AOI22_X1 U22005 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n19892), .ZN(n19865) );
  OAI211_X1 U22006 ( .C1(n19895), .C2(n20289), .A(n19866), .B(n19865), .ZN(
        P2_U3174) );
  INV_X1 U22007 ( .A(n15648), .ZN(n19891) );
  AOI22_X1 U22008 ( .A1(n19892), .A2(n20193), .B1(n19898), .B2(n20185), .ZN(
        n19868) );
  AOI22_X1 U22009 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n19899), .ZN(n19867) );
  OAI211_X1 U22010 ( .C1(n19891), .C2(n20190), .A(n19868), .B(n19867), .ZN(
        P2_U3166) );
  AOI22_X1 U22011 ( .A1(n20192), .A2(n15648), .B1(n19898), .B2(n20191), .ZN(
        n19870) );
  AOI22_X1 U22012 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20194), .B1(
        n20200), .B2(n19892), .ZN(n19869) );
  OAI211_X1 U22013 ( .C1(n19895), .C2(n19920), .A(n19870), .B(n19869), .ZN(
        P2_U3158) );
  AOI22_X1 U22014 ( .A1(n20206), .A2(n15648), .B1(n19898), .B2(n20205), .ZN(
        n19872) );
  AOI22_X1 U22015 ( .A1(n19899), .A2(n20208), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n20207), .ZN(n19871) );
  OAI211_X1 U22016 ( .C1(n19902), .C2(n20217), .A(n19872), .B(n19871), .ZN(
        P2_U3142) );
  AOI22_X1 U22017 ( .A1(n19892), .A2(n20212), .B1(n19898), .B2(n20211), .ZN(
        n19874) );
  AOI22_X1 U22018 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20214), .B1(
        n15648), .B2(n20213), .ZN(n19873) );
  OAI211_X1 U22019 ( .C1(n19895), .C2(n20217), .A(n19874), .B(n19873), .ZN(
        P2_U3134) );
  AOI22_X1 U22020 ( .A1(n19892), .A2(n20225), .B1(n19898), .B2(n20218), .ZN(
        n19876) );
  AOI22_X1 U22021 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20220), .B1(
        n15648), .B2(n20219), .ZN(n19875) );
  OAI211_X1 U22022 ( .C1(n19895), .C2(n20223), .A(n19876), .B(n19875), .ZN(
        P2_U3126) );
  AOI22_X1 U22023 ( .A1(n19892), .A2(n20233), .B1(n19898), .B2(n20224), .ZN(
        n19878) );
  AOI22_X1 U22024 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n15648), .ZN(n19877) );
  OAI211_X1 U22025 ( .C1(n19895), .C2(n20137), .A(n19878), .B(n19877), .ZN(
        P2_U3118) );
  AOI22_X1 U22026 ( .A1(n20232), .A2(n15648), .B1(n20231), .B2(n19898), .ZN(
        n19880) );
  AOI22_X1 U22027 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20234), .B1(
        n20233), .B2(n19899), .ZN(n19879) );
  OAI211_X1 U22028 ( .C1(n19902), .C2(n20243), .A(n19880), .B(n19879), .ZN(
        P2_U3110) );
  AOI22_X1 U22029 ( .A1(n20238), .A2(n15648), .B1(n19898), .B2(n20237), .ZN(
        n19882) );
  AOI22_X1 U22030 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n19892), .ZN(n19881) );
  OAI211_X1 U22031 ( .C1(n19895), .C2(n20243), .A(n19882), .B(n19881), .ZN(
        P2_U3102) );
  INV_X1 U22032 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U22033 ( .A1(n19899), .A2(n20239), .B1(n19898), .B2(n20244), .ZN(
        n19884) );
  AOI22_X1 U22034 ( .A1(n15648), .A2(n20245), .B1(n20251), .B2(n19892), .ZN(
        n19883) );
  OAI211_X1 U22035 ( .C1(n20039), .C2(n19885), .A(n19884), .B(n19883), .ZN(
        P2_U3094) );
  INV_X1 U22036 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U22037 ( .A1(n19899), .A2(n20251), .B1(n19898), .B2(n20250), .ZN(
        n19887) );
  AOI22_X1 U22038 ( .A1(n15648), .A2(n20252), .B1(n20259), .B2(n19892), .ZN(
        n19886) );
  OAI211_X1 U22039 ( .C1(n20256), .C2(n19888), .A(n19887), .B(n19886), .ZN(
        P2_U3086) );
  AOI22_X1 U22040 ( .A1(n19892), .A2(n20258), .B1(n19898), .B2(n20257), .ZN(
        n19890) );
  AOI22_X1 U22041 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20260), .B1(
        n20259), .B2(n19899), .ZN(n19889) );
  OAI211_X1 U22042 ( .C1(n20264), .C2(n19891), .A(n19890), .B(n19889), .ZN(
        P2_U3078) );
  AOI22_X1 U22043 ( .A1(n20266), .A2(n15648), .B1(n19898), .B2(n20265), .ZN(
        n19894) );
  AOI22_X1 U22044 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n19892), .ZN(n19893) );
  OAI211_X1 U22045 ( .C1(n19895), .C2(n20271), .A(n19894), .B(n19893), .ZN(
        P2_U3070) );
  AOI22_X1 U22046 ( .A1(n20274), .A2(n15648), .B1(n19898), .B2(n20273), .ZN(
        n19897) );
  AOI22_X1 U22047 ( .A1(n19899), .A2(n20276), .B1(n20275), .B2(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n19896) );
  OAI211_X1 U22048 ( .C1(n19902), .C2(n20279), .A(n19897), .B(n19896), .ZN(
        P2_U3062) );
  AOI22_X1 U22049 ( .A1(n19899), .A2(n20282), .B1(n19898), .B2(n20280), .ZN(
        n19901) );
  AOI22_X1 U22050 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n15648), .ZN(n19900) );
  OAI211_X1 U22051 ( .C1(n19902), .C2(n20289), .A(n19901), .B(n19900), .ZN(
        P2_U3054) );
  OAI22_X1 U22052 ( .A1(n19903), .A2(n20162), .B1(n19911), .B2(n20173), .ZN(
        n19904) );
  INV_X1 U22053 ( .A(n19904), .ZN(n19908) );
  NAND3_X1 U22054 ( .A1(n19906), .A2(n19905), .A3(n20167), .ZN(n19907) );
  OAI211_X1 U22055 ( .C1(n19910), .C2(n19909), .A(n19908), .B(n19907), .ZN(
        P2_U2914) );
  AOI22_X1 U22056 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n11151), .ZN(n19954) );
  NOR2_X2 U22057 ( .A1(n13479), .A2(n20176), .ZN(n19950) );
  AOI22_X1 U22058 ( .A1(n20179), .A2(n19912), .B1(n20178), .B2(n19950), .ZN(
        n19915) );
  INV_X1 U22059 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20592) );
  OAI22_X2 U22060 ( .A1(n20592), .A2(n22599), .B1(n19913), .B2(n20065), .ZN(
        n19951) );
  AOI22_X1 U22061 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n19951), .ZN(n19914) );
  OAI211_X1 U22062 ( .C1(n19954), .C2(n20289), .A(n19915), .B(n19914), .ZN(
        P2_U3173) );
  INV_X1 U22063 ( .A(n19912), .ZN(n19945) );
  AOI22_X1 U22064 ( .A1(n19951), .A2(n20193), .B1(n19950), .B2(n20185), .ZN(
        n19917) );
  INV_X1 U22065 ( .A(n19954), .ZN(n19942) );
  AOI22_X1 U22066 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n19942), .ZN(n19916) );
  OAI211_X1 U22067 ( .C1(n19945), .C2(n20190), .A(n19917), .B(n19916), .ZN(
        P2_U3165) );
  AOI22_X1 U22068 ( .A1(n20192), .A2(n19912), .B1(n19950), .B2(n20191), .ZN(
        n19919) );
  AOI22_X1 U22069 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20194), .B1(
        n20200), .B2(n19951), .ZN(n19918) );
  OAI211_X1 U22070 ( .C1(n19954), .C2(n19920), .A(n19919), .B(n19918), .ZN(
        P2_U3157) );
  INV_X1 U22071 ( .A(n19951), .ZN(n19933) );
  AOI22_X1 U22072 ( .A1(n20199), .A2(n19912), .B1(n20198), .B2(n19950), .ZN(
        n19922) );
  AOI22_X1 U22073 ( .A1(n20201), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20200), .B2(n19942), .ZN(n19921) );
  OAI211_X1 U22074 ( .C1(n19933), .C2(n20204), .A(n19922), .B(n19921), .ZN(
        P2_U3149) );
  AOI22_X1 U22075 ( .A1(n20206), .A2(n19912), .B1(n19950), .B2(n20205), .ZN(
        n19924) );
  AOI22_X1 U22076 ( .A1(n19951), .A2(n20130), .B1(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .B2(n20207), .ZN(n19923) );
  OAI211_X1 U22077 ( .C1(n19954), .C2(n20204), .A(n19924), .B(n19923), .ZN(
        P2_U3141) );
  AOI22_X1 U22078 ( .A1(n19942), .A2(n20130), .B1(n19950), .B2(n20211), .ZN(
        n19926) );
  AOI22_X1 U22079 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20214), .B1(
        n19912), .B2(n20213), .ZN(n19925) );
  OAI211_X1 U22080 ( .C1(n19933), .C2(n20223), .A(n19926), .B(n19925), .ZN(
        P2_U3133) );
  AOI22_X1 U22081 ( .A1(n19942), .A2(n20212), .B1(n20218), .B2(n19950), .ZN(
        n19928) );
  AOI22_X1 U22082 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20220), .B1(
        n19912), .B2(n20219), .ZN(n19927) );
  OAI211_X1 U22083 ( .C1(n19933), .C2(n20137), .A(n19928), .B(n19927), .ZN(
        P2_U3125) );
  AOI22_X1 U22084 ( .A1(n19951), .A2(n20233), .B1(n20224), .B2(n19950), .ZN(
        n19930) );
  AOI22_X1 U22085 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n19912), .ZN(n19929) );
  OAI211_X1 U22086 ( .C1(n19954), .C2(n20137), .A(n19930), .B(n19929), .ZN(
        P2_U3117) );
  AOI22_X1 U22087 ( .A1(n20232), .A2(n19912), .B1(n20231), .B2(n19950), .ZN(
        n19932) );
  AOI22_X1 U22088 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20234), .B1(
        n20233), .B2(n19942), .ZN(n19931) );
  OAI211_X1 U22089 ( .C1(n19933), .C2(n20243), .A(n19932), .B(n19931), .ZN(
        P2_U3109) );
  AOI22_X1 U22090 ( .A1(n20238), .A2(n19912), .B1(n20237), .B2(n19950), .ZN(
        n19935) );
  AOI22_X1 U22091 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n19951), .ZN(n19934) );
  OAI211_X1 U22092 ( .C1(n19954), .C2(n20243), .A(n19935), .B(n19934), .ZN(
        P2_U3101) );
  INV_X1 U22093 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n19938) );
  AOI22_X1 U22094 ( .A1(n19942), .A2(n20239), .B1(n19950), .B2(n20244), .ZN(
        n19937) );
  AOI22_X1 U22095 ( .A1(n19912), .A2(n20245), .B1(n20251), .B2(n19951), .ZN(
        n19936) );
  OAI211_X1 U22096 ( .C1(n20039), .C2(n19938), .A(n19937), .B(n19936), .ZN(
        P2_U3093) );
  INV_X1 U22097 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n19941) );
  AOI22_X1 U22098 ( .A1(n19942), .A2(n20251), .B1(n20250), .B2(n19950), .ZN(
        n19940) );
  AOI22_X1 U22099 ( .A1(n19912), .A2(n20252), .B1(n20259), .B2(n19951), .ZN(
        n19939) );
  OAI211_X1 U22100 ( .C1(n20256), .C2(n19941), .A(n19940), .B(n19939), .ZN(
        P2_U3085) );
  AOI22_X1 U22101 ( .A1(n19942), .A2(n20259), .B1(n19950), .B2(n20257), .ZN(
        n19944) );
  AOI22_X1 U22102 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20260), .B1(
        n20258), .B2(n19951), .ZN(n19943) );
  OAI211_X1 U22103 ( .C1(n20264), .C2(n19945), .A(n19944), .B(n19943), .ZN(
        P2_U3077) );
  AOI22_X1 U22104 ( .A1(n20266), .A2(n19912), .B1(n19950), .B2(n20265), .ZN(
        n19947) );
  AOI22_X1 U22105 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n19951), .ZN(n19946) );
  OAI211_X1 U22106 ( .C1(n19954), .C2(n20271), .A(n19947), .B(n19946), .ZN(
        P2_U3069) );
  AOI22_X1 U22107 ( .A1(n20274), .A2(n19912), .B1(n19950), .B2(n20273), .ZN(
        n19949) );
  AOI22_X1 U22108 ( .A1(n19951), .A2(n20282), .B1(
        P2_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n20275), .ZN(n19948) );
  OAI211_X1 U22109 ( .C1(n19954), .C2(n20053), .A(n19949), .B(n19948), .ZN(
        P2_U3061) );
  AOI22_X1 U22110 ( .A1(n19951), .A2(n20155), .B1(n19950), .B2(n20280), .ZN(
        n19953) );
  AOI22_X1 U22111 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n19912), .ZN(n19952) );
  OAI211_X1 U22112 ( .C1(n19954), .C2(n20279), .A(n19953), .B(n19952), .ZN(
        P2_U3053) );
  AOI22_X1 U22113 ( .A1(n19955), .A2(n19965), .B1(n20110), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U22114 ( .A1(n19957), .A2(BUF1_REG_20__SCAN_IN), .B1(n19956), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n19962) );
  OAI22_X1 U22115 ( .A1(n19959), .A2(n20115), .B1(n20164), .B2(n19958), .ZN(
        n19960) );
  INV_X1 U22116 ( .A(n19960), .ZN(n19961) );
  NAND3_X1 U22117 ( .A1(n19963), .A2(n19962), .A3(n19961), .ZN(P2_U2899) );
  INV_X1 U22118 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20573) );
  INV_X1 U22119 ( .A(n19965), .ZN(n19966) );
  NOR2_X2 U22120 ( .A1(n19966), .A2(n20174), .ZN(n20005) );
  NOR2_X2 U22121 ( .A1(n19967), .A2(n20176), .ZN(n20003) );
  AOI22_X1 U22122 ( .A1(n20179), .A2(n20005), .B1(n20178), .B2(n20003), .ZN(
        n19969) );
  AOI22_X1 U22123 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n11151), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n11154), .ZN(n20002) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n20004), .ZN(n19968) );
  OAI211_X1 U22125 ( .C1(n20008), .C2(n20289), .A(n19969), .B(n19968), .ZN(
        P2_U3172) );
  INV_X1 U22126 ( .A(n20005), .ZN(n19996) );
  AOI22_X1 U22127 ( .A1(n19999), .A2(n20186), .B1(n20003), .B2(n20185), .ZN(
        n19971) );
  AOI22_X1 U22128 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20187), .B1(
        n20193), .B2(n20004), .ZN(n19970) );
  OAI211_X1 U22129 ( .C1(n19996), .C2(n20190), .A(n19971), .B(n19970), .ZN(
        P2_U3164) );
  AOI22_X1 U22130 ( .A1(n20192), .A2(n20005), .B1(n20003), .B2(n20191), .ZN(
        n19973) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n19999), .ZN(n19972) );
  OAI211_X1 U22132 ( .C1(n20002), .C2(n20197), .A(n19973), .B(n19972), .ZN(
        P2_U3156) );
  AOI22_X1 U22133 ( .A1(n20199), .A2(n20005), .B1(n20198), .B2(n20003), .ZN(
        n19975) );
  AOI22_X1 U22134 ( .A1(n20201), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20200), .B2(n19999), .ZN(n19974) );
  OAI211_X1 U22135 ( .C1(n20002), .C2(n20204), .A(n19975), .B(n19974), .ZN(
        P2_U3148) );
  AOI22_X1 U22136 ( .A1(n20206), .A2(n20005), .B1(n20003), .B2(n20205), .ZN(
        n19977) );
  AOI22_X1 U22137 ( .A1(n20004), .A2(n20130), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n20207), .ZN(n19976) );
  OAI211_X1 U22138 ( .C1(n20008), .C2(n20204), .A(n19977), .B(n19976), .ZN(
        P2_U3140) );
  AOI22_X1 U22139 ( .A1(n20004), .A2(n20212), .B1(n20003), .B2(n20211), .ZN(
        n19979) );
  AOI22_X1 U22140 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20214), .B1(
        n20005), .B2(n20213), .ZN(n19978) );
  OAI211_X1 U22141 ( .C1(n20008), .C2(n20217), .A(n19979), .B(n19978), .ZN(
        P2_U3132) );
  AOI22_X1 U22142 ( .A1(n20004), .A2(n20225), .B1(n20218), .B2(n20003), .ZN(
        n19981) );
  AOI22_X1 U22143 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20220), .B1(
        n20005), .B2(n20219), .ZN(n19980) );
  OAI211_X1 U22144 ( .C1(n20008), .C2(n20223), .A(n19981), .B(n19980), .ZN(
        P2_U3124) );
  AOI22_X1 U22145 ( .A1(n19999), .A2(n20225), .B1(n20224), .B2(n20003), .ZN(
        n19983) );
  AOI22_X1 U22146 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n20005), .ZN(n19982) );
  OAI211_X1 U22147 ( .C1(n20002), .C2(n20230), .A(n19983), .B(n19982), .ZN(
        P2_U3116) );
  AOI22_X1 U22148 ( .A1(n20232), .A2(n20005), .B1(n20231), .B2(n20003), .ZN(
        n19985) );
  AOI22_X1 U22149 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20234), .B1(
        n20138), .B2(n20004), .ZN(n19984) );
  OAI211_X1 U22150 ( .C1(n20008), .C2(n20230), .A(n19985), .B(n19984), .ZN(
        P2_U3108) );
  AOI22_X1 U22151 ( .A1(n20238), .A2(n20005), .B1(n20237), .B2(n20003), .ZN(
        n19987) );
  AOI22_X1 U22152 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n20004), .ZN(n19986) );
  OAI211_X1 U22153 ( .C1(n20008), .C2(n20243), .A(n19987), .B(n19986), .ZN(
        P2_U3100) );
  INV_X1 U22154 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19990) );
  AOI22_X1 U22155 ( .A1(n19999), .A2(n20239), .B1(n20003), .B2(n20244), .ZN(
        n19989) );
  AOI22_X1 U22156 ( .A1(n20005), .A2(n20245), .B1(n20251), .B2(n20004), .ZN(
        n19988) );
  OAI211_X1 U22157 ( .C1(n20039), .C2(n19990), .A(n19989), .B(n19988), .ZN(
        P2_U3092) );
  INV_X1 U22158 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U22159 ( .A1(n19999), .A2(n20251), .B1(n20250), .B2(n20003), .ZN(
        n19992) );
  AOI22_X1 U22160 ( .A1(n20005), .A2(n20252), .B1(n20259), .B2(n20004), .ZN(
        n19991) );
  OAI211_X1 U22161 ( .C1(n20256), .C2(n19993), .A(n19992), .B(n19991), .ZN(
        P2_U3084) );
  AOI22_X1 U22162 ( .A1(n20004), .A2(n20258), .B1(n20003), .B2(n20257), .ZN(
        n19995) );
  AOI22_X1 U22163 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20260), .B1(
        n20259), .B2(n19999), .ZN(n19994) );
  OAI211_X1 U22164 ( .C1(n20264), .C2(n19996), .A(n19995), .B(n19994), .ZN(
        P2_U3076) );
  AOI22_X1 U22165 ( .A1(n20266), .A2(n20005), .B1(n20003), .B2(n20265), .ZN(
        n19998) );
  AOI22_X1 U22166 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n20004), .ZN(n19997) );
  OAI211_X1 U22167 ( .C1(n20008), .C2(n20271), .A(n19998), .B(n19997), .ZN(
        P2_U3068) );
  AOI22_X1 U22168 ( .A1(n20274), .A2(n20005), .B1(n20003), .B2(n20273), .ZN(
        n20001) );
  AOI22_X1 U22169 ( .A1(n19999), .A2(n20276), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n20275), .ZN(n20000) );
  OAI211_X1 U22170 ( .C1(n20002), .C2(n20279), .A(n20001), .B(n20000), .ZN(
        P2_U3060) );
  AOI22_X1 U22171 ( .A1(n20004), .A2(n20155), .B1(n20003), .B2(n20280), .ZN(
        n20007) );
  AOI22_X1 U22172 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20005), .ZN(n20006) );
  OAI211_X1 U22173 ( .C1(n20008), .C2(n20279), .A(n20007), .B(n20006), .ZN(
        P2_U3052) );
  AOI22_X1 U22174 ( .A1(n20009), .A2(n20112), .B1(n20110), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n20015) );
  AOI21_X1 U22175 ( .B1(n20012), .B2(n20011), .A(n20010), .ZN(n20013) );
  OR2_X1 U22176 ( .A1(n20013), .A2(n20115), .ZN(n20014) );
  OAI211_X1 U22177 ( .C1(n20016), .C2(n20173), .A(n20015), .B(n20014), .ZN(
        P2_U2916) );
  AOI22_X1 U22178 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n11151), .ZN(n20058) );
  NOR2_X2 U22179 ( .A1(n12745), .A2(n20176), .ZN(n20054) );
  AOI22_X1 U22180 ( .A1(n20179), .A2(n20017), .B1(n20178), .B2(n20054), .ZN(
        n20019) );
  AOI22_X1 U22181 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n11151), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n11154), .ZN(n20036) );
  AOI22_X1 U22182 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n20055), .ZN(n20018) );
  OAI211_X1 U22183 ( .C1(n20058), .C2(n20289), .A(n20019), .B(n20018), .ZN(
        P2_U3171) );
  INV_X1 U22184 ( .A(n20017), .ZN(n20048) );
  AOI22_X1 U22185 ( .A1(n20045), .A2(n20186), .B1(n20054), .B2(n20185), .ZN(
        n20021) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20187), .B1(
        n20193), .B2(n20055), .ZN(n20020) );
  OAI211_X1 U22187 ( .C1(n20048), .C2(n20190), .A(n20021), .B(n20020), .ZN(
        P2_U3163) );
  AOI22_X1 U22188 ( .A1(n20192), .A2(n20017), .B1(n20054), .B2(n20191), .ZN(
        n20023) );
  AOI22_X1 U22189 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20045), .ZN(n20022) );
  OAI211_X1 U22190 ( .C1(n20036), .C2(n20197), .A(n20023), .B(n20022), .ZN(
        P2_U3155) );
  AOI22_X1 U22191 ( .A1(n20199), .A2(n20017), .B1(n20198), .B2(n20054), .ZN(
        n20025) );
  AOI22_X1 U22192 ( .A1(n20201), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20200), .B2(n20045), .ZN(n20024) );
  OAI211_X1 U22193 ( .C1(n20036), .C2(n20204), .A(n20025), .B(n20024), .ZN(
        P2_U3147) );
  AOI22_X1 U22194 ( .A1(n20206), .A2(n20017), .B1(n20054), .B2(n20205), .ZN(
        n20027) );
  AOI22_X1 U22195 ( .A1(n20045), .A2(n20208), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n20207), .ZN(n20026) );
  OAI211_X1 U22196 ( .C1(n20036), .C2(n20217), .A(n20027), .B(n20026), .ZN(
        P2_U3139) );
  AOI22_X1 U22197 ( .A1(n20045), .A2(n20130), .B1(n20054), .B2(n20211), .ZN(
        n20029) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20214), .B1(
        n20017), .B2(n20213), .ZN(n20028) );
  OAI211_X1 U22199 ( .C1(n20036), .C2(n20223), .A(n20029), .B(n20028), .ZN(
        P2_U3131) );
  AOI22_X1 U22200 ( .A1(n20055), .A2(n20225), .B1(n20218), .B2(n20054), .ZN(
        n20031) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20220), .B1(
        n20017), .B2(n20219), .ZN(n20030) );
  OAI211_X1 U22202 ( .C1(n20058), .C2(n20223), .A(n20031), .B(n20030), .ZN(
        P2_U3123) );
  AOI22_X1 U22203 ( .A1(n20045), .A2(n20225), .B1(n20224), .B2(n20054), .ZN(
        n20033) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n20017), .ZN(n20032) );
  OAI211_X1 U22205 ( .C1(n20036), .C2(n20230), .A(n20033), .B(n20032), .ZN(
        P2_U3115) );
  AOI22_X1 U22206 ( .A1(n20232), .A2(n20017), .B1(n20231), .B2(n20054), .ZN(
        n20035) );
  AOI22_X1 U22207 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20234), .B1(
        n20233), .B2(n20045), .ZN(n20034) );
  OAI211_X1 U22208 ( .C1(n20036), .C2(n20243), .A(n20035), .B(n20034), .ZN(
        P2_U3107) );
  AOI22_X1 U22209 ( .A1(n20238), .A2(n20017), .B1(n20237), .B2(n20054), .ZN(
        n20038) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n20055), .ZN(n20037) );
  OAI211_X1 U22211 ( .C1(n20058), .C2(n20243), .A(n20038), .B(n20037), .ZN(
        P2_U3099) );
  INV_X1 U22212 ( .A(n20239), .ZN(n20249) );
  AOI22_X1 U22213 ( .A1(n20055), .A2(n20251), .B1(n20054), .B2(n20244), .ZN(
        n20041) );
  INV_X1 U22214 ( .A(n20039), .ZN(n20246) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20246), .B1(
        n20017), .B2(n20245), .ZN(n20040) );
  OAI211_X1 U22216 ( .C1(n20058), .C2(n20249), .A(n20041), .B(n20040), .ZN(
        P2_U3091) );
  INV_X1 U22217 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n20044) );
  AOI22_X1 U22218 ( .A1(n20045), .A2(n20251), .B1(n20250), .B2(n20054), .ZN(
        n20043) );
  AOI22_X1 U22219 ( .A1(n20017), .A2(n20252), .B1(n20259), .B2(n20055), .ZN(
        n20042) );
  OAI211_X1 U22220 ( .C1(n20256), .C2(n20044), .A(n20043), .B(n20042), .ZN(
        P2_U3083) );
  AOI22_X1 U22221 ( .A1(n20055), .A2(n20258), .B1(n20054), .B2(n20257), .ZN(
        n20047) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20260), .B1(
        n20259), .B2(n20045), .ZN(n20046) );
  OAI211_X1 U22223 ( .C1(n20264), .C2(n20048), .A(n20047), .B(n20046), .ZN(
        P2_U3075) );
  AOI22_X1 U22224 ( .A1(n20266), .A2(n20017), .B1(n20054), .B2(n20265), .ZN(
        n20050) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n20055), .ZN(n20049) );
  OAI211_X1 U22226 ( .C1(n20058), .C2(n20271), .A(n20050), .B(n20049), .ZN(
        P2_U3067) );
  AOI22_X1 U22227 ( .A1(n20274), .A2(n20017), .B1(n20054), .B2(n20273), .ZN(
        n20052) );
  AOI22_X1 U22228 ( .A1(n20282), .A2(n20055), .B1(n20275), .B2(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20051) );
  OAI211_X1 U22229 ( .C1(n20058), .C2(n20053), .A(n20052), .B(n20051), .ZN(
        P2_U3059) );
  AOI22_X1 U22230 ( .A1(n20055), .A2(n20155), .B1(n20054), .B2(n20280), .ZN(
        n20057) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20017), .ZN(n20056) );
  OAI211_X1 U22232 ( .C1(n20058), .C2(n20279), .A(n20057), .B(n20056), .ZN(
        P2_U3051) );
  AOI22_X1 U22233 ( .A1(n20112), .A2(n20059), .B1(n20110), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n20064) );
  XNOR2_X1 U22234 ( .A(n20061), .B(n20060), .ZN(n20062) );
  NAND2_X1 U22235 ( .A1(n20062), .A2(n20167), .ZN(n20063) );
  OAI211_X1 U22236 ( .C1(n20068), .C2(n20173), .A(n20064), .B(n20063), .ZN(
        P2_U2917) );
  INV_X1 U22237 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20569) );
  INV_X1 U22238 ( .A(n20100), .ZN(n20109) );
  NOR2_X2 U22239 ( .A1(n20068), .A2(n20174), .ZN(n20106) );
  NOR2_X2 U22240 ( .A1(n20069), .A2(n20176), .ZN(n20104) );
  AOI22_X1 U22241 ( .A1(n20179), .A2(n20106), .B1(n20178), .B2(n20104), .ZN(
        n20071) );
  AOI22_X1 U22242 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n11151), .ZN(n20103) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n20105), .ZN(n20070) );
  OAI211_X1 U22244 ( .C1(n20109), .C2(n20289), .A(n20071), .B(n20070), .ZN(
        P2_U3170) );
  INV_X1 U22245 ( .A(n20106), .ZN(n20097) );
  AOI22_X1 U22246 ( .A1(n20105), .A2(n20193), .B1(n20104), .B2(n20185), .ZN(
        n20073) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n20100), .ZN(n20072) );
  OAI211_X1 U22248 ( .C1(n20097), .C2(n20190), .A(n20073), .B(n20072), .ZN(
        P2_U3162) );
  AOI22_X1 U22249 ( .A1(n20192), .A2(n20106), .B1(n20104), .B2(n20191), .ZN(
        n20075) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20100), .ZN(n20074) );
  OAI211_X1 U22251 ( .C1(n20103), .C2(n20197), .A(n20075), .B(n20074), .ZN(
        P2_U3154) );
  AOI22_X1 U22252 ( .A1(n20199), .A2(n20106), .B1(n20198), .B2(n20104), .ZN(
        n20077) );
  AOI22_X1 U22253 ( .A1(n20201), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20200), .B2(n20100), .ZN(n20076) );
  OAI211_X1 U22254 ( .C1(n20103), .C2(n20204), .A(n20077), .B(n20076), .ZN(
        P2_U3146) );
  AOI22_X1 U22255 ( .A1(n20206), .A2(n20106), .B1(n20104), .B2(n20205), .ZN(
        n20079) );
  AOI22_X1 U22256 ( .A1(n20105), .A2(n20130), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n20207), .ZN(n20078) );
  OAI211_X1 U22257 ( .C1(n20109), .C2(n20204), .A(n20079), .B(n20078), .ZN(
        P2_U3138) );
  AOI22_X1 U22258 ( .A1(n20100), .A2(n20130), .B1(n20104), .B2(n20211), .ZN(
        n20081) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20214), .B1(
        n20106), .B2(n20213), .ZN(n20080) );
  OAI211_X1 U22260 ( .C1(n20103), .C2(n20223), .A(n20081), .B(n20080), .ZN(
        P2_U3130) );
  AOI22_X1 U22261 ( .A1(n20100), .A2(n20212), .B1(n20218), .B2(n20104), .ZN(
        n20083) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20220), .B1(
        n20106), .B2(n20219), .ZN(n20082) );
  OAI211_X1 U22263 ( .C1(n20103), .C2(n20137), .A(n20083), .B(n20082), .ZN(
        P2_U3122) );
  AOI22_X1 U22264 ( .A1(n20100), .A2(n20225), .B1(n20224), .B2(n20104), .ZN(
        n20085) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n20106), .ZN(n20084) );
  OAI211_X1 U22266 ( .C1(n20103), .C2(n20230), .A(n20085), .B(n20084), .ZN(
        P2_U3114) );
  AOI22_X1 U22267 ( .A1(n20232), .A2(n20106), .B1(n20231), .B2(n20104), .ZN(
        n20087) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20234), .B1(
        n20138), .B2(n20105), .ZN(n20086) );
  OAI211_X1 U22269 ( .C1(n20109), .C2(n20230), .A(n20087), .B(n20086), .ZN(
        P2_U3106) );
  AOI22_X1 U22270 ( .A1(n20238), .A2(n20106), .B1(n20237), .B2(n20104), .ZN(
        n20089) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n20105), .ZN(n20088) );
  OAI211_X1 U22272 ( .C1(n20109), .C2(n20243), .A(n20089), .B(n20088), .ZN(
        P2_U3098) );
  AOI22_X1 U22273 ( .A1(n20105), .A2(n20251), .B1(n20244), .B2(n20104), .ZN(
        n20091) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20246), .B1(
        n20106), .B2(n20245), .ZN(n20090) );
  OAI211_X1 U22275 ( .C1(n20109), .C2(n20249), .A(n20091), .B(n20090), .ZN(
        P2_U3090) );
  INV_X1 U22276 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20094) );
  AOI22_X1 U22277 ( .A1(n20100), .A2(n20251), .B1(n20250), .B2(n20104), .ZN(
        n20093) );
  AOI22_X1 U22278 ( .A1(n20106), .A2(n20252), .B1(n20259), .B2(n20105), .ZN(
        n20092) );
  OAI211_X1 U22279 ( .C1(n20256), .C2(n20094), .A(n20093), .B(n20092), .ZN(
        P2_U3082) );
  AOI22_X1 U22280 ( .A1(n20105), .A2(n20258), .B1(n20104), .B2(n20257), .ZN(
        n20096) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20260), .B1(
        n20259), .B2(n20100), .ZN(n20095) );
  OAI211_X1 U22282 ( .C1(n20264), .C2(n20097), .A(n20096), .B(n20095), .ZN(
        P2_U3074) );
  AOI22_X1 U22283 ( .A1(n20266), .A2(n20106), .B1(n20104), .B2(n20265), .ZN(
        n20099) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n20105), .ZN(n20098) );
  OAI211_X1 U22285 ( .C1(n20109), .C2(n20271), .A(n20099), .B(n20098), .ZN(
        P2_U3066) );
  AOI22_X1 U22286 ( .A1(n20274), .A2(n20106), .B1(n20104), .B2(n20273), .ZN(
        n20102) );
  AOI22_X1 U22287 ( .A1(n20100), .A2(n20276), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n20275), .ZN(n20101) );
  OAI211_X1 U22288 ( .C1(n20103), .C2(n20279), .A(n20102), .B(n20101), .ZN(
        P2_U3058) );
  AOI22_X1 U22289 ( .A1(n20105), .A2(n20155), .B1(n20104), .B2(n20280), .ZN(
        n20108) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20106), .ZN(n20107) );
  OAI211_X1 U22291 ( .C1(n20109), .C2(n20279), .A(n20108), .B(n20107), .ZN(
        P2_U3050) );
  AOI22_X1 U22292 ( .A1(n20112), .A2(n20111), .B1(n20110), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n20118) );
  AOI21_X1 U22293 ( .B1(n20166), .B2(n20114), .A(n20113), .ZN(n20116) );
  OR2_X1 U22294 ( .A1(n20116), .A2(n20115), .ZN(n20117) );
  OAI211_X1 U22295 ( .C1(n20119), .C2(n20173), .A(n20118), .B(n20117), .ZN(
        P2_U2918) );
  AOI22_X1 U22296 ( .A1(n20179), .A2(n20157), .B1(n20154), .B2(n20178), .ZN(
        n20121) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n20156), .ZN(n20120) );
  OAI211_X1 U22298 ( .C1(n20160), .C2(n20289), .A(n20121), .B(n20120), .ZN(
        P2_U3169) );
  INV_X1 U22299 ( .A(n20157), .ZN(n20147) );
  AOI22_X1 U22300 ( .A1(n20156), .A2(n20193), .B1(n20154), .B2(n20185), .ZN(
        n20123) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20187), .B1(
        n20186), .B2(n20150), .ZN(n20122) );
  OAI211_X1 U22302 ( .C1(n20147), .C2(n20190), .A(n20123), .B(n20122), .ZN(
        P2_U3161) );
  AOI22_X1 U22303 ( .A1(n20192), .A2(n20157), .B1(n20154), .B2(n20191), .ZN(
        n20125) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20150), .ZN(n20124) );
  OAI211_X1 U22305 ( .C1(n20153), .C2(n20197), .A(n20125), .B(n20124), .ZN(
        P2_U3153) );
  AOI22_X1 U22306 ( .A1(n20199), .A2(n20157), .B1(n20198), .B2(n20154), .ZN(
        n20127) );
  AOI22_X1 U22307 ( .A1(n20201), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20200), .B2(n20150), .ZN(n20126) );
  OAI211_X1 U22308 ( .C1(n20153), .C2(n20204), .A(n20127), .B(n20126), .ZN(
        P2_U3145) );
  AOI22_X1 U22309 ( .A1(n20206), .A2(n20157), .B1(n20154), .B2(n20205), .ZN(
        n20129) );
  AOI22_X1 U22310 ( .A1(n20150), .A2(n20208), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n20207), .ZN(n20128) );
  OAI211_X1 U22311 ( .C1(n20153), .C2(n20217), .A(n20129), .B(n20128), .ZN(
        P2_U3137) );
  AOI22_X1 U22312 ( .A1(n20150), .A2(n20130), .B1(n20154), .B2(n20211), .ZN(
        n20132) );
  AOI22_X1 U22313 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20214), .B1(
        n20157), .B2(n20213), .ZN(n20131) );
  OAI211_X1 U22314 ( .C1(n20153), .C2(n20223), .A(n20132), .B(n20131), .ZN(
        P2_U3129) );
  AOI22_X1 U22315 ( .A1(n20150), .A2(n20212), .B1(n20154), .B2(n20218), .ZN(
        n20134) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20220), .B1(
        n20157), .B2(n20219), .ZN(n20133) );
  OAI211_X1 U22317 ( .C1(n20153), .C2(n20137), .A(n20134), .B(n20133), .ZN(
        P2_U3121) );
  AOI22_X1 U22318 ( .A1(n20156), .A2(n20233), .B1(n20154), .B2(n20224), .ZN(
        n20136) );
  AOI22_X1 U22319 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n20157), .ZN(n20135) );
  OAI211_X1 U22320 ( .C1(n20160), .C2(n20137), .A(n20136), .B(n20135), .ZN(
        P2_U3113) );
  AOI22_X1 U22321 ( .A1(n20232), .A2(n20157), .B1(n20231), .B2(n20154), .ZN(
        n20140) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20234), .B1(
        n20138), .B2(n20156), .ZN(n20139) );
  OAI211_X1 U22323 ( .C1(n20160), .C2(n20230), .A(n20140), .B(n20139), .ZN(
        P2_U3105) );
  AOI22_X1 U22324 ( .A1(n20238), .A2(n20157), .B1(n20237), .B2(n20154), .ZN(
        n20142) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n20156), .ZN(n20141) );
  OAI211_X1 U22326 ( .C1(n20160), .C2(n20243), .A(n20142), .B(n20141), .ZN(
        P2_U3097) );
  AOI22_X1 U22327 ( .A1(n20156), .A2(n20251), .B1(n20154), .B2(n20244), .ZN(
        n20144) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20246), .B1(
        n20157), .B2(n20245), .ZN(n20143) );
  OAI211_X1 U22329 ( .C1(n20160), .C2(n20249), .A(n20144), .B(n20143), .ZN(
        P2_U3089) );
  AOI22_X1 U22330 ( .A1(n20156), .A2(n20258), .B1(n20154), .B2(n20257), .ZN(
        n20146) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20260), .B1(
        n20259), .B2(n20150), .ZN(n20145) );
  OAI211_X1 U22332 ( .C1(n20264), .C2(n20147), .A(n20146), .B(n20145), .ZN(
        P2_U3073) );
  AOI22_X1 U22333 ( .A1(n20266), .A2(n20157), .B1(n20154), .B2(n20265), .ZN(
        n20149) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n20156), .ZN(n20148) );
  OAI211_X1 U22335 ( .C1(n20160), .C2(n20271), .A(n20149), .B(n20148), .ZN(
        P2_U3065) );
  AOI22_X1 U22336 ( .A1(n20274), .A2(n20157), .B1(n20154), .B2(n20273), .ZN(
        n20152) );
  AOI22_X1 U22337 ( .A1(n20150), .A2(n20276), .B1(n20275), .B2(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n20151) );
  OAI211_X1 U22338 ( .C1(n20153), .C2(n20279), .A(n20152), .B(n20151), .ZN(
        P2_U3057) );
  AOI22_X1 U22339 ( .A1(n20156), .A2(n20155), .B1(n20154), .B2(n20280), .ZN(
        n20159) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20157), .ZN(n20158) );
  OAI211_X1 U22341 ( .C1(n20160), .C2(n20279), .A(n20159), .B(n20158), .ZN(
        P2_U3049) );
  OAI22_X1 U22342 ( .A1(n20164), .A2(n20163), .B1(n20162), .B2(n20161), .ZN(
        n20165) );
  INV_X1 U22343 ( .A(n20165), .ZN(n20172) );
  INV_X1 U22344 ( .A(n20166), .ZN(n20168) );
  OAI211_X1 U22345 ( .C1(n20170), .C2(n20169), .A(n20168), .B(n20167), .ZN(
        n20171) );
  OAI211_X1 U22346 ( .C1(n20175), .C2(n20173), .A(n20172), .B(n20171), .ZN(
        P2_U2919) );
  AOI22_X1 U22347 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n11151), .ZN(n20272) );
  NOR2_X2 U22348 ( .A1(n20175), .A2(n20174), .ZN(n20284) );
  NOR2_X2 U22349 ( .A1(n20177), .A2(n20176), .ZN(n20281) );
  AOI22_X1 U22350 ( .A1(n20179), .A2(n20284), .B1(n20178), .B2(n20281), .ZN(
        n20184) );
  AOI22_X1 U22351 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n11154), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n11151), .ZN(n20290) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20182), .B1(
        n20186), .B2(n20267), .ZN(n20183) );
  OAI211_X1 U22353 ( .C1(n20272), .C2(n20289), .A(n20184), .B(n20183), .ZN(
        P2_U3168) );
  INV_X1 U22354 ( .A(n20284), .ZN(n20263) );
  AOI22_X1 U22355 ( .A1(n20283), .A2(n20186), .B1(n20281), .B2(n20185), .ZN(
        n20189) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20187), .B1(
        n20193), .B2(n20267), .ZN(n20188) );
  OAI211_X1 U22357 ( .C1(n20263), .C2(n20190), .A(n20189), .B(n20188), .ZN(
        P2_U3160) );
  AOI22_X1 U22358 ( .A1(n20192), .A2(n20284), .B1(n20281), .B2(n20191), .ZN(
        n20196) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20194), .B1(
        n20193), .B2(n20283), .ZN(n20195) );
  OAI211_X1 U22360 ( .C1(n20290), .C2(n20197), .A(n20196), .B(n20195), .ZN(
        P2_U3152) );
  AOI22_X1 U22361 ( .A1(n20199), .A2(n20284), .B1(n20198), .B2(n20281), .ZN(
        n20203) );
  AOI22_X1 U22362 ( .A1(n20201), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20200), .B2(n20283), .ZN(n20202) );
  OAI211_X1 U22363 ( .C1(n20290), .C2(n20204), .A(n20203), .B(n20202), .ZN(
        P2_U3144) );
  AOI22_X1 U22364 ( .A1(n20206), .A2(n20284), .B1(n20281), .B2(n20205), .ZN(
        n20210) );
  AOI22_X1 U22365 ( .A1(n20283), .A2(n20208), .B1(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n20207), .ZN(n20209) );
  OAI211_X1 U22366 ( .C1(n20290), .C2(n20217), .A(n20210), .B(n20209), .ZN(
        P2_U3136) );
  AOI22_X1 U22367 ( .A1(n20267), .A2(n20212), .B1(n20281), .B2(n20211), .ZN(
        n20216) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20214), .B1(
        n20284), .B2(n20213), .ZN(n20215) );
  OAI211_X1 U22369 ( .C1(n20272), .C2(n20217), .A(n20216), .B(n20215), .ZN(
        P2_U3128) );
  AOI22_X1 U22370 ( .A1(n20267), .A2(n20225), .B1(n20218), .B2(n20281), .ZN(
        n20222) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20220), .B1(
        n20284), .B2(n20219), .ZN(n20221) );
  OAI211_X1 U22372 ( .C1(n20272), .C2(n20223), .A(n20222), .B(n20221), .ZN(
        P2_U3120) );
  AOI22_X1 U22373 ( .A1(n20283), .A2(n20225), .B1(n20224), .B2(n20281), .ZN(
        n20229) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20227), .B1(
        n20226), .B2(n20284), .ZN(n20228) );
  OAI211_X1 U22375 ( .C1(n20290), .C2(n20230), .A(n20229), .B(n20228), .ZN(
        P2_U3112) );
  AOI22_X1 U22376 ( .A1(n20232), .A2(n20284), .B1(n20231), .B2(n20281), .ZN(
        n20236) );
  AOI22_X1 U22377 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20234), .B1(
        n20233), .B2(n20283), .ZN(n20235) );
  OAI211_X1 U22378 ( .C1(n20290), .C2(n20243), .A(n20236), .B(n20235), .ZN(
        P2_U3104) );
  AOI22_X1 U22379 ( .A1(n20238), .A2(n20284), .B1(n20237), .B2(n20281), .ZN(
        n20242) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20240), .B1(
        n20239), .B2(n20267), .ZN(n20241) );
  OAI211_X1 U22381 ( .C1(n20272), .C2(n20243), .A(n20242), .B(n20241), .ZN(
        P2_U3096) );
  AOI22_X1 U22382 ( .A1(n20267), .A2(n20251), .B1(n20244), .B2(n20281), .ZN(
        n20248) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20246), .B1(
        n20284), .B2(n20245), .ZN(n20247) );
  OAI211_X1 U22384 ( .C1(n20272), .C2(n20249), .A(n20248), .B(n20247), .ZN(
        P2_U3088) );
  INV_X1 U22385 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n20255) );
  AOI22_X1 U22386 ( .A1(n20283), .A2(n20251), .B1(n20250), .B2(n20281), .ZN(
        n20254) );
  AOI22_X1 U22387 ( .A1(n20284), .A2(n20252), .B1(n20259), .B2(n20267), .ZN(
        n20253) );
  OAI211_X1 U22388 ( .C1(n20256), .C2(n20255), .A(n20254), .B(n20253), .ZN(
        P2_U3080) );
  AOI22_X1 U22389 ( .A1(n20267), .A2(n20258), .B1(n20281), .B2(n20257), .ZN(
        n20262) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20260), .B1(
        n20259), .B2(n20283), .ZN(n20261) );
  OAI211_X1 U22391 ( .C1(n20264), .C2(n20263), .A(n20262), .B(n20261), .ZN(
        P2_U3072) );
  AOI22_X1 U22392 ( .A1(n20266), .A2(n20284), .B1(n20281), .B2(n20265), .ZN(
        n20270) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20268), .B1(
        n20276), .B2(n20267), .ZN(n20269) );
  OAI211_X1 U22394 ( .C1(n20272), .C2(n20271), .A(n20270), .B(n20269), .ZN(
        P2_U3064) );
  AOI22_X1 U22395 ( .A1(n20274), .A2(n20284), .B1(n20281), .B2(n20273), .ZN(
        n20278) );
  AOI22_X1 U22396 ( .A1(n20283), .A2(n20276), .B1(n20275), .B2(
        P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20277) );
  OAI211_X1 U22397 ( .C1(n20290), .C2(n20279), .A(n20278), .B(n20277), .ZN(
        P2_U3056) );
  AOI22_X1 U22398 ( .A1(n20283), .A2(n20282), .B1(n20281), .B2(n20280), .ZN(
        n20288) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20286), .B1(
        n20285), .B2(n20284), .ZN(n20287) );
  OAI211_X1 U22400 ( .C1(n20290), .C2(n20289), .A(n20288), .B(n20287), .ZN(
        P2_U3048) );
  INV_X1 U22401 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20595) );
  INV_X1 U22402 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20291) );
  AOI222_X1 U22403 ( .A1(n20595), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20598), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20291), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20292) );
  INV_X2 U22404 ( .A(n20292), .ZN(n20352) );
  INV_X1 U22405 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20294) );
  AOI22_X1 U22406 ( .A1(n20341), .A2(n20294), .B1(n20293), .B2(n20352), .ZN(
        U376) );
  INV_X1 U22407 ( .A(n20352), .ZN(n20355) );
  INV_X1 U22408 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20296) );
  AOI22_X1 U22409 ( .A1(n20355), .A2(n20296), .B1(n20295), .B2(n20352), .ZN(
        U365) );
  AOI22_X1 U22410 ( .A1(n20341), .A2(n20298), .B1(n20297), .B2(n20352), .ZN(
        U354) );
  AOI22_X1 U22411 ( .A1(n20341), .A2(n20300), .B1(n20299), .B2(n20352), .ZN(
        U353) );
  INV_X1 U22412 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20302) );
  AOI22_X1 U22413 ( .A1(n20341), .A2(n20302), .B1(n20301), .B2(n20352), .ZN(
        U352) );
  INV_X1 U22414 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20304) );
  AOI22_X1 U22415 ( .A1(n20341), .A2(n20304), .B1(n20303), .B2(n20352), .ZN(
        U351) );
  INV_X1 U22416 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20306) );
  AOI22_X1 U22417 ( .A1(n20355), .A2(n20306), .B1(n20305), .B2(n20352), .ZN(
        U350) );
  INV_X1 U22418 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20308) );
  AOI22_X1 U22419 ( .A1(n20341), .A2(n20308), .B1(n20307), .B2(n20352), .ZN(
        U349) );
  AOI22_X1 U22420 ( .A1(n20341), .A2(n20310), .B1(n20309), .B2(n20352), .ZN(
        U348) );
  AOI22_X1 U22421 ( .A1(n20341), .A2(n20312), .B1(n20311), .B2(n20352), .ZN(
        U347) );
  AOI22_X1 U22422 ( .A1(n20341), .A2(n20314), .B1(n20313), .B2(n20352), .ZN(
        U375) );
  AOI22_X1 U22423 ( .A1(n20341), .A2(n20316), .B1(n20315), .B2(n20352), .ZN(
        U374) );
  INV_X1 U22424 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20318) );
  AOI22_X1 U22425 ( .A1(n20341), .A2(n20318), .B1(n20317), .B2(n20352), .ZN(
        U373) );
  INV_X1 U22426 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20320) );
  AOI22_X1 U22427 ( .A1(n20341), .A2(n20320), .B1(n20319), .B2(n20352), .ZN(
        U372) );
  INV_X1 U22428 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20322) );
  AOI22_X1 U22429 ( .A1(n20341), .A2(n20322), .B1(n20321), .B2(n20352), .ZN(
        U371) );
  INV_X1 U22430 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20324) );
  AOI22_X1 U22431 ( .A1(n20341), .A2(n20324), .B1(n20323), .B2(n20352), .ZN(
        U370) );
  AOI22_X1 U22432 ( .A1(n20341), .A2(n20326), .B1(n20325), .B2(n20352), .ZN(
        U369) );
  AOI22_X1 U22433 ( .A1(n20341), .A2(n20328), .B1(n20327), .B2(n20352), .ZN(
        U368) );
  AOI22_X1 U22434 ( .A1(n20341), .A2(n20330), .B1(n20329), .B2(n20352), .ZN(
        U367) );
  AOI22_X1 U22435 ( .A1(n20341), .A2(n20332), .B1(n20331), .B2(n20352), .ZN(
        U366) );
  AOI22_X1 U22436 ( .A1(n20341), .A2(n20334), .B1(n20333), .B2(n20352), .ZN(
        U364) );
  AOI22_X1 U22437 ( .A1(n20341), .A2(n20336), .B1(n20335), .B2(n20352), .ZN(
        U363) );
  AOI22_X1 U22438 ( .A1(n20341), .A2(n20338), .B1(n20337), .B2(n20352), .ZN(
        U362) );
  AOI22_X1 U22439 ( .A1(n20341), .A2(n20340), .B1(n20339), .B2(n20352), .ZN(
        U361) );
  AOI22_X1 U22440 ( .A1(n20355), .A2(n20343), .B1(n20342), .B2(n20352), .ZN(
        U360) );
  AOI22_X1 U22441 ( .A1(n20355), .A2(n20345), .B1(n20344), .B2(n20352), .ZN(
        U359) );
  INV_X1 U22442 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20347) );
  AOI22_X1 U22443 ( .A1(n20355), .A2(n20347), .B1(n20346), .B2(n20352), .ZN(
        U358) );
  INV_X1 U22444 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20349) );
  AOI22_X1 U22445 ( .A1(n20355), .A2(n20349), .B1(n20348), .B2(n20352), .ZN(
        U357) );
  AOI22_X1 U22446 ( .A1(n20355), .A2(n20351), .B1(n20350), .B2(n20352), .ZN(
        U356) );
  AOI22_X1 U22447 ( .A1(n20355), .A2(n20354), .B1(n20353), .B2(n20352), .ZN(
        U355) );
  AOI22_X1 U22448 ( .A1(n21841), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20357) );
  OAI21_X1 U22449 ( .B1(n20358), .B2(n20384), .A(n20357), .ZN(P1_U2936) );
  AOI22_X1 U22450 ( .A1(n21841), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20359) );
  OAI21_X1 U22451 ( .B1(n11920), .B2(n20384), .A(n20359), .ZN(P1_U2935) );
  AOI22_X1 U22452 ( .A1(n21841), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20360) );
  OAI21_X1 U22453 ( .B1(n11966), .B2(n20384), .A(n20360), .ZN(P1_U2934) );
  AOI22_X1 U22454 ( .A1(n20376), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20361) );
  OAI21_X1 U22455 ( .B1(n11997), .B2(n20384), .A(n20361), .ZN(P1_U2933) );
  AOI22_X1 U22456 ( .A1(n20376), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20362) );
  OAI21_X1 U22457 ( .B1(n20363), .B2(n20384), .A(n20362), .ZN(P1_U2932) );
  AOI22_X1 U22458 ( .A1(n20376), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20364) );
  OAI21_X1 U22459 ( .B1(n20365), .B2(n20384), .A(n20364), .ZN(P1_U2931) );
  AOI22_X1 U22460 ( .A1(n20376), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20366) );
  OAI21_X1 U22461 ( .B1(n15270), .B2(n20384), .A(n20366), .ZN(P1_U2930) );
  AOI22_X1 U22462 ( .A1(n20376), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20367) );
  OAI21_X1 U22463 ( .B1(n12073), .B2(n20384), .A(n20367), .ZN(P1_U2929) );
  AOI22_X1 U22464 ( .A1(n20376), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20368) );
  OAI21_X1 U22465 ( .B1(n15479), .B2(n20384), .A(n20368), .ZN(P1_U2928) );
  AOI22_X1 U22466 ( .A1(n20376), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20369) );
  OAI21_X1 U22467 ( .B1(n20370), .B2(n20384), .A(n20369), .ZN(P1_U2927) );
  AOI22_X1 U22468 ( .A1(n20376), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20372) );
  OAI21_X1 U22469 ( .B1(n20373), .B2(n20384), .A(n20372), .ZN(P1_U2926) );
  AOI22_X1 U22470 ( .A1(n20376), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20374) );
  OAI21_X1 U22471 ( .B1(n20375), .B2(n20384), .A(n20374), .ZN(P1_U2925) );
  AOI22_X1 U22472 ( .A1(n20376), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20377) );
  OAI21_X1 U22473 ( .B1(n20378), .B2(n20384), .A(n20377), .ZN(P1_U2924) );
  AOI22_X1 U22474 ( .A1(n21841), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20379) );
  OAI21_X1 U22475 ( .B1(n20380), .B2(n20384), .A(n20379), .ZN(P1_U2923) );
  AOI22_X1 U22476 ( .A1(n21841), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20381) );
  OAI21_X1 U22477 ( .B1(n20382), .B2(n20384), .A(n20381), .ZN(P1_U2922) );
  INV_X1 U22478 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20385) );
  AOI22_X1 U22479 ( .A1(n21841), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20371), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20383) );
  OAI21_X1 U22480 ( .B1(n20385), .B2(n20384), .A(n20383), .ZN(P1_U2921) );
  AND2_X1 U22481 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22596), .ZN(n20418) );
  INV_X2 U22482 ( .A(n20418), .ZN(n20438) );
  INV_X1 U22483 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21885) );
  AND2_X1 U22484 ( .A1(n22596), .A2(n20528), .ZN(n20416) );
  OAI222_X1 U22485 ( .A1(n20438), .A2(n20387), .B1(n20386), .B2(n22596), .C1(
        n21885), .C2(n11172), .ZN(P1_U3197) );
  INV_X1 U22486 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20388) );
  OAI222_X1 U22487 ( .A1(n11172), .A2(n20390), .B1(n20388), .B2(n22596), .C1(
        n21885), .C2(n20438), .ZN(P1_U3198) );
  INV_X1 U22488 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20389) );
  OAI222_X1 U22489 ( .A1(n20438), .A2(n20390), .B1(n20389), .B2(n22596), .C1(
        n20392), .C2(n11172), .ZN(P1_U3199) );
  INV_X1 U22490 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20391) );
  INV_X1 U22491 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20394) );
  OAI222_X1 U22492 ( .A1(n20438), .A2(n20392), .B1(n20391), .B2(n22596), .C1(
        n20394), .C2(n11172), .ZN(P1_U3200) );
  INV_X1 U22493 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20393) );
  OAI222_X1 U22494 ( .A1(n20438), .A2(n20394), .B1(n20393), .B2(n22596), .C1(
        n22039), .C2(n11172), .ZN(P1_U3201) );
  INV_X1 U22495 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20395) );
  OAI222_X1 U22496 ( .A1(n20438), .A2(n22039), .B1(n20395), .B2(n22596), .C1(
        n22050), .C2(n11172), .ZN(P1_U3202) );
  INV_X1 U22497 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20396) );
  OAI222_X1 U22498 ( .A1(n20438), .A2(n22050), .B1(n20396), .B2(n22596), .C1(
        n20398), .C2(n11172), .ZN(P1_U3203) );
  INV_X1 U22499 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20397) );
  OAI222_X1 U22500 ( .A1(n20438), .A2(n20398), .B1(n20397), .B2(n22596), .C1(
        n20400), .C2(n11172), .ZN(P1_U3204) );
  INV_X1 U22501 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20399) );
  OAI222_X1 U22502 ( .A1(n20438), .A2(n20400), .B1(n20399), .B2(n22596), .C1(
        n22064), .C2(n11172), .ZN(P1_U3205) );
  INV_X1 U22503 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20401) );
  OAI222_X1 U22504 ( .A1(n20438), .A2(n22064), .B1(n20401), .B2(n22596), .C1(
        n22062), .C2(n11172), .ZN(P1_U3206) );
  INV_X1 U22505 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20402) );
  OAI222_X1 U22506 ( .A1(n20438), .A2(n22062), .B1(n20402), .B2(n22596), .C1(
        n20404), .C2(n11172), .ZN(P1_U3207) );
  INV_X1 U22507 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20403) );
  OAI222_X1 U22508 ( .A1(n20438), .A2(n20404), .B1(n20403), .B2(n22596), .C1(
        n21853), .C2(n11172), .ZN(P1_U3208) );
  INV_X1 U22509 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20405) );
  OAI222_X1 U22510 ( .A1(n11172), .A2(n20407), .B1(n20405), .B2(n22596), .C1(
        n21853), .C2(n20438), .ZN(P1_U3209) );
  INV_X1 U22511 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20406) );
  OAI222_X1 U22512 ( .A1(n20438), .A2(n20407), .B1(n20406), .B2(n22596), .C1(
        n20408), .C2(n11172), .ZN(P1_U3210) );
  INV_X1 U22513 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20409) );
  OAI222_X1 U22514 ( .A1(n11172), .A2(n20410), .B1(n20409), .B2(n22596), .C1(
        n20408), .C2(n20438), .ZN(P1_U3211) );
  INV_X1 U22515 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20411) );
  OAI222_X1 U22516 ( .A1(n11172), .A2(n20413), .B1(n20411), .B2(n22596), .C1(
        n20410), .C2(n20438), .ZN(P1_U3212) );
  INV_X1 U22517 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20412) );
  OAI222_X1 U22518 ( .A1(n20438), .A2(n20413), .B1(n20412), .B2(n22596), .C1(
        n20414), .C2(n11172), .ZN(P1_U3213) );
  INV_X1 U22519 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20415) );
  OAI222_X1 U22520 ( .A1(n11172), .A2(n22000), .B1(n20415), .B2(n22596), .C1(
        n20414), .C2(n20438), .ZN(P1_U3214) );
  AOI22_X1 U22521 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n20416), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n22593), .ZN(n20417) );
  OAI21_X1 U22522 ( .B1(n22000), .B2(n20438), .A(n20417), .ZN(P1_U3215) );
  AOI22_X1 U22523 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n20418), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n22593), .ZN(n20419) );
  OAI21_X1 U22524 ( .B1(n22123), .B2(n11172), .A(n20419), .ZN(P1_U3216) );
  INV_X1 U22525 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20420) );
  OAI222_X1 U22526 ( .A1(n20438), .A2(n22123), .B1(n20420), .B2(n22596), .C1(
        n20422), .C2(n11172), .ZN(P1_U3217) );
  INV_X1 U22527 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20421) );
  INV_X1 U22528 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n22127) );
  OAI222_X1 U22529 ( .A1(n20438), .A2(n20422), .B1(n20421), .B2(n22596), .C1(
        n22127), .C2(n11172), .ZN(P1_U3218) );
  INV_X1 U22530 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20423) );
  OAI222_X1 U22531 ( .A1(n11172), .A2(n11382), .B1(n20423), .B2(n22596), .C1(
        n22127), .C2(n20438), .ZN(P1_U3219) );
  INV_X1 U22532 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20424) );
  OAI222_X1 U22533 ( .A1(n20438), .A2(n11382), .B1(n20424), .B2(n22596), .C1(
        n20425), .C2(n11172), .ZN(P1_U3220) );
  INV_X1 U22534 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20426) );
  OAI222_X1 U22535 ( .A1(n11172), .A2(n20428), .B1(n20426), .B2(n22596), .C1(
        n20425), .C2(n20438), .ZN(P1_U3221) );
  INV_X1 U22536 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20427) );
  OAI222_X1 U22537 ( .A1(n20438), .A2(n20428), .B1(n20427), .B2(n22596), .C1(
        n20430), .C2(n11172), .ZN(P1_U3222) );
  INV_X1 U22538 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20429) );
  OAI222_X1 U22539 ( .A1(n20438), .A2(n20430), .B1(n20429), .B2(n22596), .C1(
        n20431), .C2(n11172), .ZN(P1_U3223) );
  INV_X1 U22540 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20432) );
  OAI222_X1 U22541 ( .A1(n11172), .A2(n20433), .B1(n20432), .B2(n22596), .C1(
        n20431), .C2(n20438), .ZN(P1_U3224) );
  INV_X1 U22542 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20434) );
  OAI222_X1 U22543 ( .A1(n11172), .A2(n20437), .B1(n20434), .B2(n22596), .C1(
        n20433), .C2(n20438), .ZN(P1_U3225) );
  INV_X1 U22544 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20436) );
  OAI222_X1 U22545 ( .A1(n20438), .A2(n20437), .B1(n20436), .B2(n22596), .C1(
        n20435), .C2(n11172), .ZN(P1_U3226) );
  INV_X1 U22546 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20451) );
  INV_X1 U22547 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20439) );
  AOI22_X1 U22548 ( .A1(n22596), .A2(n20451), .B1(n20439), .B2(n22593), .ZN(
        P1_U3458) );
  NOR4_X1 U22549 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20443) );
  NOR4_X1 U22550 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20442) );
  NOR4_X1 U22551 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20441) );
  NOR4_X1 U22552 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20440) );
  NAND4_X1 U22553 ( .A1(n20443), .A2(n20442), .A3(n20441), .A4(n20440), .ZN(
        n20449) );
  NOR4_X1 U22554 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20447) );
  AOI211_X1 U22555 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20446) );
  NOR4_X1 U22556 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20445) );
  NOR4_X1 U22557 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20444) );
  NAND4_X1 U22558 ( .A1(n20447), .A2(n20446), .A3(n20445), .A4(n20444), .ZN(
        n20448) );
  NOR2_X1 U22559 ( .A1(n20449), .A2(n20448), .ZN(n20466) );
  NOR3_X1 U22560 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20459) );
  NOR2_X1 U22561 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20455) );
  OAI21_X1 U22562 ( .B1(n20459), .B2(n20455), .A(n20466), .ZN(n20450) );
  OAI21_X1 U22563 ( .B1(n20466), .B2(n20451), .A(n20450), .ZN(P1_U2808) );
  INV_X1 U22564 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20456) );
  INV_X1 U22565 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20452) );
  AOI22_X1 U22566 ( .A1(n22596), .A2(n20456), .B1(n20452), .B2(n22593), .ZN(
        P1_U3459) );
  NOR3_X1 U22567 ( .A1(n20454), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20453) );
  AOI221_X1 U22568 ( .B1(n20455), .B2(n20454), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20453), .ZN(n20457) );
  INV_X1 U22569 ( .A(n20466), .ZN(n20463) );
  AOI22_X1 U22570 ( .A1(n20466), .A2(n20457), .B1(n20456), .B2(n20463), .ZN(
        P1_U3481) );
  INV_X1 U22571 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20461) );
  INV_X1 U22572 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20458) );
  AOI22_X1 U22573 ( .A1(n22596), .A2(n20461), .B1(n20458), .B2(n22593), .ZN(
        P1_U3460) );
  OAI21_X1 U22574 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20459), .A(n20466), .ZN(
        n20460) );
  OAI21_X1 U22575 ( .B1(n20466), .B2(n20461), .A(n20460), .ZN(P1_U2807) );
  INV_X1 U22576 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20464) );
  INV_X1 U22577 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20462) );
  AOI22_X1 U22578 ( .A1(n22596), .A2(n20464), .B1(n20462), .B2(n22593), .ZN(
        P1_U3461) );
  NOR2_X1 U22579 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20465) );
  AOI22_X1 U22580 ( .A1(n20466), .A2(n20465), .B1(n20464), .B2(n20463), .ZN(
        P1_U3482) );
  AOI22_X1 U22581 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20514), .ZN(n20473) );
  OAI21_X1 U22582 ( .B1(n20469), .B2(n20468), .A(n20467), .ZN(n20470) );
  INV_X1 U22583 ( .A(n20470), .ZN(n21899) );
  AOI22_X1 U22584 ( .A1(n21899), .A2(n20518), .B1(n20471), .B2(n20519), .ZN(
        n20472) );
  OAI211_X1 U22585 ( .C1(n20522), .C2(n20474), .A(n20473), .B(n20472), .ZN(
        P1_U2995) );
  AOI22_X1 U22586 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20514), .ZN(n20480) );
  OAI21_X1 U22587 ( .B1(n20477), .B2(n20476), .A(n20475), .ZN(n20478) );
  INV_X1 U22588 ( .A(n20478), .ZN(n21925) );
  AOI22_X1 U22589 ( .A1(n21925), .A2(n20518), .B1(n20519), .B2(n22031), .ZN(
        n20479) );
  OAI211_X1 U22590 ( .C1(n20522), .C2(n22034), .A(n20480), .B(n20479), .ZN(
        P1_U2994) );
  AOI22_X1 U22591 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20514), .ZN(n20486) );
  OAI21_X1 U22592 ( .B1(n20483), .B2(n20482), .A(n20481), .ZN(n20484) );
  INV_X1 U22593 ( .A(n20484), .ZN(n21919) );
  AOI22_X1 U22594 ( .A1(n21919), .A2(n20518), .B1(n20519), .B2(n22042), .ZN(
        n20485) );
  OAI211_X1 U22595 ( .C1(n20522), .C2(n22045), .A(n20486), .B(n20485), .ZN(
        P1_U2993) );
  AOI22_X1 U22596 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20514), .ZN(n20492) );
  OAI21_X1 U22597 ( .B1(n20489), .B2(n20488), .A(n20487), .ZN(n20490) );
  INV_X1 U22598 ( .A(n20490), .ZN(n21937) );
  AOI22_X1 U22599 ( .A1(n21937), .A2(n20518), .B1(n20519), .B2(n22053), .ZN(
        n20491) );
  OAI211_X1 U22600 ( .C1(n20522), .C2(n22056), .A(n20492), .B(n20491), .ZN(
        P1_U2992) );
  AOI22_X1 U22601 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20514), .ZN(n20499) );
  INV_X1 U22602 ( .A(n22083), .ZN(n20497) );
  AOI22_X1 U22603 ( .A1(n20505), .A2(n22080), .B1(n20519), .B2(n20497), .ZN(
        n20498) );
  OAI211_X1 U22604 ( .C1(n20500), .C2(n22141), .A(n20499), .B(n20498), .ZN(
        P1_U2987) );
  AOI22_X1 U22605 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20514), .ZN(n20502) );
  AOI22_X1 U22606 ( .A1(n22090), .A2(n20519), .B1(n20505), .B2(n22089), .ZN(
        n20501) );
  OAI211_X1 U22607 ( .C1(n22141), .C2(n20503), .A(n20502), .B(n20501), .ZN(
        P1_U2984) );
  AOI22_X1 U22608 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20514), .ZN(n20508) );
  AOI22_X1 U22609 ( .A1(n20506), .A2(n20519), .B1(n20505), .B2(n20504), .ZN(
        n20507) );
  OAI211_X1 U22610 ( .C1(n20509), .C2(n22141), .A(n20508), .B(n20507), .ZN(
        P1_U2982) );
  AOI22_X1 U22611 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20514), .ZN(n20513) );
  XNOR2_X1 U22612 ( .A(n20516), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n20510) );
  XNOR2_X1 U22613 ( .A(n20511), .B(n20510), .ZN(n21994) );
  AOI22_X1 U22614 ( .A1(n22102), .A2(n20519), .B1(n20518), .B2(n21994), .ZN(
        n20512) );
  OAI211_X1 U22615 ( .C1(n20522), .C2(n22097), .A(n20513), .B(n20512), .ZN(
        P1_U2980) );
  AOI22_X1 U22616 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n22016), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20514), .ZN(n20521) );
  XNOR2_X1 U22617 ( .A(n20516), .B(n20515), .ZN(n20517) );
  XNOR2_X1 U22618 ( .A(n13658), .B(n20517), .ZN(n22019) );
  AOI22_X1 U22619 ( .A1(n22138), .A2(n20519), .B1(n20518), .B2(n22019), .ZN(
        n20520) );
  OAI211_X1 U22620 ( .C1(n20522), .C2(n22129), .A(n20521), .B(n20520), .ZN(
        P1_U2976) );
  NAND2_X1 U22621 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12293), .ZN(n20526) );
  OAI21_X1 U22622 ( .B1(n20523), .B2(n22162), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20524) );
  OAI21_X1 U22623 ( .B1(n20526), .B2(n20525), .A(n20524), .ZN(P1_U2803) );
  OAI21_X1 U22624 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20528), .A(n20527), 
        .ZN(n20529) );
  AOI22_X1 U22625 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22596), .B1(n20530), 
        .B2(n20529), .ZN(P1_U2804) );
  AOI22_X1 U22626 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n11170), .ZN(n20532) );
  OAI21_X1 U22627 ( .B1(n20533), .B2(n20597), .A(n20532), .ZN(U247) );
  AOI22_X1 U22628 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n11170), .ZN(n20534) );
  OAI21_X1 U22629 ( .B1(n20535), .B2(n20597), .A(n20534), .ZN(U246) );
  AOI22_X1 U22630 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n11170), .ZN(n20536) );
  OAI21_X1 U22631 ( .B1(n20537), .B2(n20597), .A(n20536), .ZN(U245) );
  AOI22_X1 U22632 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n11170), .ZN(n20538) );
  OAI21_X1 U22633 ( .B1(n20539), .B2(n20597), .A(n20538), .ZN(U244) );
  AOI22_X1 U22634 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n11170), .ZN(n20540) );
  OAI21_X1 U22635 ( .B1(n20541), .B2(n20597), .A(n20540), .ZN(U243) );
  AOI22_X1 U22636 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n11170), .ZN(n20542) );
  OAI21_X1 U22637 ( .B1(n20543), .B2(n20597), .A(n20542), .ZN(U242) );
  AOI22_X1 U22638 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n11170), .ZN(n20544) );
  OAI21_X1 U22639 ( .B1(n20545), .B2(n20597), .A(n20544), .ZN(U241) );
  AOI22_X1 U22640 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n11170), .ZN(n20546) );
  OAI21_X1 U22641 ( .B1(n20547), .B2(n20597), .A(n20546), .ZN(U240) );
  AOI22_X1 U22642 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n11170), .ZN(n20548) );
  OAI21_X1 U22643 ( .B1(n20549), .B2(n20597), .A(n20548), .ZN(U239) );
  INV_X1 U22644 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20551) );
  AOI22_X1 U22645 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n11170), .ZN(n20550) );
  OAI21_X1 U22646 ( .B1(n20551), .B2(n20597), .A(n20550), .ZN(U238) );
  AOI22_X1 U22647 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n11170), .ZN(n20552) );
  OAI21_X1 U22648 ( .B1(n20553), .B2(n20597), .A(n20552), .ZN(U237) );
  INV_X1 U22649 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U22650 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n11170), .ZN(n20554) );
  OAI21_X1 U22651 ( .B1(n20555), .B2(n20597), .A(n20554), .ZN(U236) );
  AOI22_X1 U22652 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11170), .ZN(n20556) );
  OAI21_X1 U22653 ( .B1(n20557), .B2(n20597), .A(n20556), .ZN(U235) );
  INV_X1 U22654 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20559) );
  AOI22_X1 U22655 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n11170), .ZN(n20558) );
  OAI21_X1 U22656 ( .B1(n20559), .B2(n20597), .A(n20558), .ZN(U234) );
  AOI22_X1 U22657 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n11170), .ZN(n20560) );
  OAI21_X1 U22658 ( .B1(n20561), .B2(n20597), .A(n20560), .ZN(U233) );
  INV_X1 U22659 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20563) );
  AOI22_X1 U22660 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n11170), .ZN(n20562) );
  OAI21_X1 U22661 ( .B1(n20563), .B2(n20597), .A(n20562), .ZN(U232) );
  INV_X1 U22662 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20565) );
  AOI22_X1 U22663 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n11170), .ZN(n20564) );
  OAI21_X1 U22664 ( .B1(n20565), .B2(n20597), .A(n20564), .ZN(U231) );
  INV_X1 U22665 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20567) );
  AOI22_X1 U22666 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n11170), .ZN(n20566) );
  OAI21_X1 U22667 ( .B1(n20567), .B2(n20597), .A(n20566), .ZN(U230) );
  AOI22_X1 U22668 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n11170), .ZN(n20568) );
  OAI21_X1 U22669 ( .B1(n20569), .B2(n20597), .A(n20568), .ZN(U229) );
  INV_X1 U22670 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20571) );
  AOI22_X1 U22671 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n11170), .ZN(n20570) );
  OAI21_X1 U22672 ( .B1(n20571), .B2(n20597), .A(n20570), .ZN(U228) );
  AOI22_X1 U22673 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n11170), .ZN(n20572) );
  OAI21_X1 U22674 ( .B1(n20573), .B2(n20597), .A(n20572), .ZN(U227) );
  INV_X1 U22675 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20575) );
  AOI22_X1 U22676 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n11170), .ZN(n20574) );
  OAI21_X1 U22677 ( .B1(n20575), .B2(n20597), .A(n20574), .ZN(U226) );
  INV_X1 U22678 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20577) );
  AOI22_X1 U22679 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n11170), .ZN(n20576) );
  OAI21_X1 U22680 ( .B1(n20577), .B2(n20597), .A(n20576), .ZN(U225) );
  INV_X1 U22681 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20579) );
  AOI22_X1 U22682 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n11170), .ZN(n20578) );
  OAI21_X1 U22683 ( .B1(n20579), .B2(n20597), .A(n20578), .ZN(U224) );
  INV_X1 U22684 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20581) );
  AOI22_X1 U22685 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n11170), .ZN(n20580) );
  OAI21_X1 U22686 ( .B1(n20581), .B2(n20597), .A(n20580), .ZN(U223) );
  INV_X1 U22687 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20583) );
  AOI22_X1 U22688 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n11170), .ZN(n20582) );
  OAI21_X1 U22689 ( .B1(n20583), .B2(n20597), .A(n20582), .ZN(U222) );
  INV_X1 U22690 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20586) );
  AOI22_X1 U22691 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n11170), .ZN(n20585) );
  OAI21_X1 U22692 ( .B1(n20586), .B2(n20597), .A(n20585), .ZN(U221) );
  INV_X1 U22693 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20588) );
  AOI22_X1 U22694 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n11170), .ZN(n20587) );
  OAI21_X1 U22695 ( .B1(n20588), .B2(n20597), .A(n20587), .ZN(U220) );
  INV_X1 U22696 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20590) );
  AOI22_X1 U22697 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n11170), .ZN(n20589) );
  OAI21_X1 U22698 ( .B1(n20590), .B2(n20597), .A(n20589), .ZN(U219) );
  AOI22_X1 U22699 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n11170), .ZN(n20591) );
  OAI21_X1 U22700 ( .B1(n20592), .B2(n20597), .A(n20591), .ZN(U218) );
  INV_X1 U22701 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20594) );
  AOI22_X1 U22702 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20584), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n11170), .ZN(n20593) );
  OAI21_X1 U22703 ( .B1(n20594), .B2(n20597), .A(n20593), .ZN(U217) );
  OAI222_X1 U22704 ( .A1(U212), .A2(n20598), .B1(n20597), .B2(n20596), .C1(
        U214), .C2(n20595), .ZN(U216) );
  AOI22_X1 U22705 ( .A1(n22596), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20599), 
        .B2(n22593), .ZN(P1_U3483) );
  AOI21_X1 U22706 ( .B1(n22224), .B2(n21770), .A(n20670), .ZN(n20600) );
  INV_X1 U22707 ( .A(n20600), .ZN(n20601) );
  AOI21_X1 U22708 ( .B1(n20602), .B2(n21807), .A(n20601), .ZN(n20608) );
  AOI21_X1 U22709 ( .B1(n20665), .B2(n20675), .A(n21339), .ZN(n20603) );
  OAI211_X1 U22710 ( .C1(n20604), .C2(n20603), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n22224), .ZN(n20605) );
  AOI21_X1 U22711 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20605), .A(n21823), 
        .ZN(n20607) );
  NAND2_X1 U22712 ( .A1(n20608), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20606) );
  OAI21_X1 U22713 ( .B1(n20608), .B2(n20607), .A(n20606), .ZN(P3_U3296) );
  INV_X1 U22714 ( .A(n20609), .ZN(n20610) );
  NAND2_X1 U22715 ( .A1(n21808), .A2(n20610), .ZN(n20663) );
  INV_X1 U22716 ( .A(n20663), .ZN(n20617) );
  AOI22_X1 U22717 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20657), .ZN(n20612) );
  OAI21_X1 U22718 ( .B1(n20613), .B2(n20663), .A(n20612), .ZN(P3_U2768) );
  AOI22_X1 U22719 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20657), .ZN(n20614) );
  OAI21_X1 U22720 ( .B1(n21159), .B2(n20663), .A(n20614), .ZN(P3_U2769) );
  AOI22_X1 U22721 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20657), .ZN(n20615) );
  OAI21_X1 U22722 ( .B1(n20616), .B2(n20663), .A(n20615), .ZN(P3_U2770) );
  AOI22_X1 U22723 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20657), .ZN(n20618) );
  OAI21_X1 U22724 ( .B1(n21180), .B2(n20659), .A(n20618), .ZN(P3_U2771) );
  AOI22_X1 U22725 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20657), .ZN(n20619) );
  OAI21_X1 U22726 ( .B1(n21170), .B2(n20659), .A(n20619), .ZN(P3_U2772) );
  AOI22_X1 U22727 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20657), .ZN(n20620) );
  OAI21_X1 U22728 ( .B1(n21171), .B2(n20659), .A(n20620), .ZN(P3_U2773) );
  AOI22_X1 U22729 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20657), .ZN(n20621) );
  OAI21_X1 U22730 ( .B1(n21195), .B2(n20659), .A(n20621), .ZN(P3_U2774) );
  AOI22_X1 U22731 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20657), .ZN(n20622) );
  OAI21_X1 U22732 ( .B1(n20623), .B2(n20659), .A(n20622), .ZN(P3_U2775) );
  AOI22_X1 U22733 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20657), .ZN(n20624) );
  OAI21_X1 U22734 ( .B1(n11384), .B2(n20659), .A(n20624), .ZN(P3_U2776) );
  AOI22_X1 U22735 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20657), .ZN(n20625) );
  OAI21_X1 U22736 ( .B1(n20626), .B2(n20659), .A(n20625), .ZN(P3_U2777) );
  AOI22_X1 U22737 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20657), .ZN(n20627) );
  OAI21_X1 U22738 ( .B1(n21204), .B2(n20659), .A(n20627), .ZN(P3_U2778) );
  AOI22_X1 U22739 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20657), .ZN(n20628) );
  OAI21_X1 U22740 ( .B1(n20629), .B2(n20659), .A(n20628), .ZN(P3_U2779) );
  AOI22_X1 U22741 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20657), .ZN(n20630) );
  OAI21_X1 U22742 ( .B1(n21220), .B2(n20659), .A(n20630), .ZN(P3_U2780) );
  AOI22_X1 U22743 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20657), .ZN(n20631) );
  OAI21_X1 U22744 ( .B1(n20632), .B2(n20659), .A(n20631), .ZN(P3_U2781) );
  AOI22_X1 U22745 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20661), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20657), .ZN(n20633) );
  OAI21_X1 U22746 ( .B1(n20634), .B2(n20659), .A(n20633), .ZN(P3_U2782) );
  AOI22_X1 U22747 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20657), .ZN(n20635) );
  OAI21_X1 U22748 ( .B1(n21281), .B2(n20659), .A(n20635), .ZN(P3_U2783) );
  AOI22_X1 U22749 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20657), .ZN(n20636) );
  OAI21_X1 U22750 ( .B1(n20637), .B2(n20659), .A(n20636), .ZN(P3_U2784) );
  AOI22_X1 U22751 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20657), .ZN(n20638) );
  OAI21_X1 U22752 ( .B1(n20639), .B2(n20659), .A(n20638), .ZN(P3_U2785) );
  AOI22_X1 U22753 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20657), .ZN(n20640) );
  OAI21_X1 U22754 ( .B1(n21149), .B2(n20659), .A(n20640), .ZN(P3_U2786) );
  AOI22_X1 U22755 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20660), .ZN(n20641) );
  OAI21_X1 U22756 ( .B1(n21145), .B2(n20659), .A(n20641), .ZN(P3_U2787) );
  AOI22_X1 U22757 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20660), .ZN(n20642) );
  OAI21_X1 U22758 ( .B1(n20643), .B2(n20659), .A(n20642), .ZN(P3_U2788) );
  AOI22_X1 U22759 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20660), .ZN(n20644) );
  OAI21_X1 U22760 ( .B1(n20645), .B2(n20659), .A(n20644), .ZN(P3_U2789) );
  AOI22_X1 U22761 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20652), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20660), .ZN(n20646) );
  OAI21_X1 U22762 ( .B1(n21129), .B2(n20659), .A(n20646), .ZN(P3_U2790) );
  AOI22_X1 U22763 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20652), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20660), .ZN(n20647) );
  OAI21_X1 U22764 ( .B1(n21267), .B2(n20659), .A(n20647), .ZN(P3_U2791) );
  AOI22_X1 U22765 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20652), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20660), .ZN(n20648) );
  OAI21_X1 U22766 ( .B1(n21156), .B2(n20663), .A(n20648), .ZN(P3_U2792) );
  AOI22_X1 U22767 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20652), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20660), .ZN(n20649) );
  OAI21_X1 U22768 ( .B1(n20650), .B2(n20659), .A(n20649), .ZN(P3_U2793) );
  AOI22_X1 U22769 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20652), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20660), .ZN(n20651) );
  OAI21_X1 U22770 ( .B1(n21112), .B2(n20663), .A(n20651), .ZN(P3_U2794) );
  AOI22_X1 U22771 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20652), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20660), .ZN(n20653) );
  OAI21_X1 U22772 ( .B1(n20654), .B2(n20659), .A(n20653), .ZN(P3_U2795) );
  AOI22_X1 U22773 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20660), .ZN(n20655) );
  OAI21_X1 U22774 ( .B1(n20656), .B2(n20663), .A(n20655), .ZN(P3_U2796) );
  AOI22_X1 U22775 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20657), .ZN(n20658) );
  OAI21_X1 U22776 ( .B1(n21253), .B2(n20659), .A(n20658), .ZN(P3_U2797) );
  AOI22_X1 U22777 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20661), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20660), .ZN(n20662) );
  OAI21_X1 U22778 ( .B1(n21257), .B2(n20663), .A(n20662), .ZN(P3_U2798) );
  INV_X1 U22779 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21094) );
  NOR4_X1 U22780 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n20664), .ZN(n20865) );
  INV_X1 U22781 ( .A(n20865), .ZN(n21815) );
  OAI21_X1 U22782 ( .B1(n20864), .B2(n21094), .A(n21069), .ZN(n20834) );
  AOI211_X1 U22783 ( .C1(n20665), .C2(n21339), .A(n22226), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n21809) );
  INV_X1 U22784 ( .A(n20811), .ZN(n20796) );
  AOI211_X4 U22785 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n21341), .A(n21809), .B(
        n20674), .ZN(n21075) );
  AOI22_X1 U22786 ( .A1(n20796), .A2(n20668), .B1(P3_EBX_REG_1__SCAN_IN), .B2(
        n21075), .ZN(n20681) );
  AND2_X1 U22787 ( .A1(n21812), .A2(n20669), .ZN(n21825) );
  NOR4_X2 U22788 ( .A1(n21769), .A2(n20670), .A3(n21069), .A4(n21825), .ZN(
        n21095) );
  INV_X1 U22789 ( .A(n21095), .ZN(n20810) );
  NAND3_X1 U22790 ( .A1(n21065), .A2(n21069), .A3(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20672) );
  AOI21_X1 U22791 ( .B1(n21090), .B2(n20672), .A(n20671), .ZN(n20679) );
  NAND2_X1 U22792 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n21341), .ZN(n20673) );
  AOI211_X4 U22793 ( .C1(n22224), .C2(n20675), .A(n20674), .B(n20673), .ZN(
        n21050) );
  NAND2_X1 U22794 ( .A1(n20676), .A2(n21294), .ZN(n21286) );
  OAI22_X1 U22795 ( .A1(n21093), .A2(n20677), .B1(n21286), .B2(n21100), .ZN(
        n20678) );
  AOI211_X1 U22796 ( .C1(n21095), .C2(P3_REIP_REG_1__SCAN_IN), .A(n20679), .B(
        n20678), .ZN(n20680) );
  OAI211_X1 U22797 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20834), .A(
        n20681), .B(n20680), .ZN(P3_U2670) );
  NAND2_X1 U22798 ( .A1(n21069), .A2(n20864), .ZN(n20868) );
  NAND2_X1 U22799 ( .A1(n21091), .A2(n20682), .ZN(n20683) );
  NOR3_X1 U22800 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20706) );
  AOI211_X1 U22801 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20683), .A(n20706), .B(
        n21093), .ZN(n20690) );
  NAND2_X1 U22802 ( .A1(n21772), .A2(n21294), .ZN(n21324) );
  NAND2_X1 U22803 ( .A1(n20684), .A2(n21324), .ZN(n21299) );
  INV_X1 U22804 ( .A(n21299), .ZN(n20686) );
  AOI22_X1 U22805 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n21095), .B1(n20686), 
        .B2(n20685), .ZN(n20688) );
  NAND2_X1 U22806 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20696) );
  OAI211_X1 U22807 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20796), .B(n20696), .ZN(n20687) );
  OAI211_X1 U22808 ( .C1(n21090), .C2(n20691), .A(n20688), .B(n20687), .ZN(
        n20689) );
  AOI211_X1 U22809 ( .C1(n21075), .C2(P3_EBX_REG_2__SCAN_IN), .A(n20690), .B(
        n20689), .ZN(n20693) );
  NAND2_X1 U22810 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n21094), .ZN(
        n20904) );
  INV_X1 U22811 ( .A(n20904), .ZN(n20716) );
  NOR2_X1 U22812 ( .A1(n20864), .A2(n21815), .ZN(n21086) );
  OAI221_X1 U22813 ( .B1(n20716), .B2(n20694), .C1(n20904), .C2(n20691), .A(
        n21086), .ZN(n20692) );
  OAI211_X1 U22814 ( .C1(n20868), .C2(n20694), .A(n20693), .B(n20692), .ZN(
        P3_U2669) );
  NOR2_X1 U22815 ( .A1(n20695), .A2(n20696), .ZN(n20723) );
  OAI21_X1 U22816 ( .B1(n20723), .B2(n20811), .A(n20810), .ZN(n20715) );
  OAI21_X1 U22817 ( .B1(n20811), .B2(n20696), .A(n20695), .ZN(n20704) );
  AOI21_X1 U22818 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20716), .A(
        n20864), .ZN(n20698) );
  OAI21_X1 U22819 ( .B1(n20699), .B2(n20698), .A(n20865), .ZN(n20697) );
  AOI21_X1 U22820 ( .B1(n20699), .B2(n20698), .A(n20697), .ZN(n20703) );
  NAND2_X1 U22821 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21312) );
  OAI21_X1 U22822 ( .B1(n21310), .B2(n21312), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21318) );
  NAND2_X1 U22823 ( .A1(n20700), .A2(n21318), .ZN(n21330) );
  INV_X1 U22824 ( .A(n21330), .ZN(n20701) );
  OAI22_X1 U22825 ( .A1(n20701), .A2(n21100), .B1(n20705), .B2(n21092), .ZN(
        n20702) );
  AOI211_X1 U22826 ( .C1(n20715), .C2(n20704), .A(n20703), .B(n20702), .ZN(
        n20708) );
  NAND2_X1 U22827 ( .A1(n20706), .A2(n20705), .ZN(n20710) );
  OAI211_X1 U22828 ( .C1(n20706), .C2(n20705), .A(n21050), .B(n20710), .ZN(
        n20707) );
  OAI211_X1 U22829 ( .C1(n21090), .C2(n20709), .A(n20708), .B(n20707), .ZN(
        P3_U2668) );
  NOR2_X1 U22830 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20710), .ZN(n20734) );
  AOI211_X1 U22831 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20710), .A(n20734), .B(
        n21093), .ZN(n20711) );
  AOI21_X1 U22832 ( .B1(n21056), .B2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20711), .ZN(n20722) );
  AOI211_X1 U22833 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n21065), .A(
        n20718), .B(n20834), .ZN(n20712) );
  AOI21_X1 U22834 ( .B1(n21075), .B2(P3_EBX_REG_4__SCAN_IN), .A(n20712), .ZN(
        n20721) );
  NAND3_X1 U22835 ( .A1(n20796), .A2(n20723), .A3(n21418), .ZN(n20713) );
  OAI221_X1 U22836 ( .B1(n21100), .B2(n14351), .C1(n21100), .C2(n21798), .A(
        n20713), .ZN(n20714) );
  AOI211_X1 U22837 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n20715), .A(n21769), .B(
        n20714), .ZN(n20720) );
  AOI21_X1 U22838 ( .B1(n20717), .B2(n20716), .A(n20864), .ZN(n20727) );
  NAND3_X1 U22839 ( .A1(n21069), .A2(n20727), .A3(n20718), .ZN(n20719) );
  NAND4_X1 U22840 ( .A1(n20722), .A2(n20721), .A3(n20720), .A4(n20719), .ZN(
        P3_U2667) );
  NAND2_X1 U22841 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20723), .ZN(n20729) );
  NOR2_X1 U22842 ( .A1(n20724), .A2(n20729), .ZN(n20752) );
  OAI21_X1 U22843 ( .B1(n20752), .B2(n20811), .A(n20810), .ZN(n20759) );
  INV_X1 U22844 ( .A(n20728), .ZN(n20726) );
  INV_X1 U22845 ( .A(n20727), .ZN(n20725) );
  AOI221_X1 U22846 ( .B1(n20728), .B2(n20727), .C1(n20726), .C2(n20725), .A(
        n21815), .ZN(n20732) );
  INV_X1 U22847 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20733) );
  OR3_X1 U22848 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20811), .A3(n20729), .ZN(
        n20730) );
  OAI211_X1 U22849 ( .C1(n20733), .C2(n21092), .A(n11173), .B(n20730), .ZN(
        n20731) );
  AOI211_X1 U22850 ( .C1(n20759), .C2(P3_REIP_REG_5__SCAN_IN), .A(n20732), .B(
        n20731), .ZN(n20736) );
  NAND2_X1 U22851 ( .A1(n20734), .A2(n20733), .ZN(n20745) );
  OAI211_X1 U22852 ( .C1(n20734), .C2(n20733), .A(n21050), .B(n20745), .ZN(
        n20735) );
  OAI211_X1 U22853 ( .C1(n21090), .C2(n20737), .A(n20736), .B(n20735), .ZN(
        P3_U2666) );
  INV_X1 U22854 ( .A(n20752), .ZN(n20738) );
  NOR3_X1 U22855 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20811), .A3(n20738), .ZN(
        n20760) );
  NOR2_X1 U22856 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20739), .ZN(
        n20805) );
  INV_X1 U22857 ( .A(n20805), .ZN(n20740) );
  NAND3_X1 U22858 ( .A1(n21086), .A2(n20744), .A3(n20740), .ZN(n20741) );
  OAI211_X1 U22859 ( .C1(n20742), .C2(n21090), .A(n11173), .B(n20741), .ZN(
        n20743) );
  AOI211_X1 U22860 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n20759), .A(n20760), .B(
        n20743), .ZN(n20749) );
  AOI211_X1 U22861 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n20868), .A(
        n20744), .B(n20834), .ZN(n20747) );
  NOR2_X1 U22862 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20745), .ZN(n20754) );
  AOI211_X1 U22863 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20745), .A(n20754), .B(
        n21093), .ZN(n20746) );
  AOI211_X1 U22864 ( .C1(n21075), .C2(P3_EBX_REG_6__SCAN_IN), .A(n20747), .B(
        n20746), .ZN(n20748) );
  NAND2_X1 U22865 ( .A1(n20749), .A2(n20748), .ZN(P3_U2665) );
  NOR2_X1 U22866 ( .A1(n20805), .A2(n20864), .ZN(n20750) );
  XNOR2_X1 U22867 ( .A(n20751), .B(n20750), .ZN(n20763) );
  NAND2_X1 U22868 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20752), .ZN(n20765) );
  NOR3_X1 U22869 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20811), .A3(n20765), .ZN(
        n20758) );
  NAND2_X1 U22870 ( .A1(n20754), .A2(n20753), .ZN(n20764) );
  OAI211_X1 U22871 ( .C1(n20754), .C2(n20753), .A(n21050), .B(n20764), .ZN(
        n20755) );
  OAI211_X1 U22872 ( .C1(n20756), .C2(n21090), .A(n11173), .B(n20755), .ZN(
        n20757) );
  AOI211_X1 U22873 ( .C1(n21075), .C2(P3_EBX_REG_7__SCAN_IN), .A(n20758), .B(
        n20757), .ZN(n20762) );
  OAI21_X1 U22874 ( .B1(n20760), .B2(n20759), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n20761) );
  OAI211_X1 U22875 ( .C1(n20763), .C2(n21815), .A(n20762), .B(n20761), .ZN(
        P3_U2664) );
  INV_X1 U22876 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20775) );
  NOR2_X1 U22877 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20764), .ZN(n20781) );
  AOI211_X1 U22878 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20764), .A(n20781), .B(
        n21093), .ZN(n20773) );
  NOR2_X1 U22879 ( .A1(n21442), .A2(n20765), .ZN(n20766) );
  AOI21_X1 U22880 ( .B1(n20796), .B2(n20766), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n20771) );
  NAND2_X1 U22881 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20766), .ZN(n20794) );
  AOI21_X1 U22882 ( .B1(n20796), .B2(n20794), .A(n21095), .ZN(n20790) );
  OAI21_X1 U22883 ( .B1(n20904), .B2(n20767), .A(n21065), .ZN(n20768) );
  XNOR2_X1 U22884 ( .A(n20769), .B(n20768), .ZN(n20770) );
  OAI22_X1 U22885 ( .A1(n20771), .A2(n20790), .B1(n21815), .B2(n20770), .ZN(
        n20772) );
  AOI211_X1 U22886 ( .C1(n21056), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20773), .B(n20772), .ZN(n20774) );
  OAI211_X1 U22887 ( .C1(n20775), .C2(n21092), .A(n20774), .B(n11173), .ZN(
        P3_U2663) );
  AOI211_X1 U22888 ( .C1(n20776), .C2(n20868), .A(n20779), .B(n20834), .ZN(
        n20786) );
  NAND2_X1 U22889 ( .A1(n20796), .A2(n21767), .ZN(n20777) );
  OAI22_X1 U22890 ( .A1(n20778), .A2(n21090), .B1(n20794), .B2(n20777), .ZN(
        n20785) );
  AOI211_X1 U22891 ( .C1(n20791), .C2(n21094), .A(n20864), .B(n21815), .ZN(
        n20789) );
  AOI22_X1 U22892 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n21075), .B1(n20779), .B2(
        n20789), .ZN(n20783) );
  NAND2_X1 U22893 ( .A1(n20781), .A2(n20780), .ZN(n20787) );
  OAI211_X1 U22894 ( .C1(n20781), .C2(n20780), .A(n21050), .B(n20787), .ZN(
        n20782) );
  OAI211_X1 U22895 ( .C1(n20790), .C2(n21767), .A(n20783), .B(n20782), .ZN(
        n20784) );
  OR4_X1 U22896 ( .A1(n18279), .A2(n20786), .A3(n20785), .A4(n20784), .ZN(
        P3_U2662) );
  NOR2_X1 U22897 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20787), .ZN(n20814) );
  AOI211_X1 U22898 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20787), .A(n20814), .B(
        n21093), .ZN(n20788) );
  AOI21_X1 U22899 ( .B1(n20792), .B2(n20789), .A(n20788), .ZN(n20803) );
  OAI21_X1 U22900 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n20811), .A(n20790), .ZN(
        n20801) );
  INV_X1 U22901 ( .A(n20791), .ZN(n20793) );
  AOI211_X1 U22902 ( .C1(n20793), .C2(n20868), .A(n20792), .B(n20834), .ZN(
        n20800) );
  NOR2_X1 U22903 ( .A1(n21767), .A2(n20794), .ZN(n20809) );
  NAND3_X1 U22904 ( .A1(n20796), .A2(n20809), .A3(n20795), .ZN(n20797) );
  OAI211_X1 U22905 ( .C1(n20798), .C2(n21090), .A(n11173), .B(n20797), .ZN(
        n20799) );
  AOI211_X1 U22906 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n20801), .A(n20800), 
        .B(n20799), .ZN(n20802) );
  OAI211_X1 U22907 ( .C1(n20804), .C2(n21092), .A(n20803), .B(n20802), .ZN(
        P3_U2661) );
  NAND2_X1 U22908 ( .A1(n20806), .A2(n20805), .ZN(n20825) );
  NAND2_X1 U22909 ( .A1(n21065), .A2(n20825), .ZN(n20807) );
  XNOR2_X1 U22910 ( .A(n20808), .B(n20807), .ZN(n20818) );
  NAND2_X1 U22911 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20809), .ZN(n20812) );
  NAND2_X1 U22912 ( .A1(n20811), .A2(n20810), .ZN(n21098) );
  INV_X1 U22913 ( .A(n21098), .ZN(n20938) );
  NOR3_X1 U22914 ( .A1(n21095), .A2(n20812), .A3(n20824), .ZN(n20896) );
  NOR2_X1 U22915 ( .A1(n20938), .A2(n20896), .ZN(n20847) );
  INV_X1 U22916 ( .A(n20847), .ZN(n20813) );
  AOI21_X1 U22917 ( .B1(n20824), .B2(n20823), .A(n20813), .ZN(n20817) );
  NAND2_X1 U22918 ( .A1(n20814), .A2(n20820), .ZN(n20821) );
  OAI211_X1 U22919 ( .C1(n20814), .C2(n20820), .A(n21050), .B(n20821), .ZN(
        n20815) );
  OAI21_X1 U22920 ( .B1(n21090), .B2(n20826), .A(n20815), .ZN(n20816) );
  AOI211_X1 U22921 ( .C1(n21069), .C2(n20818), .A(n20817), .B(n20816), .ZN(
        n20819) );
  OAI211_X1 U22922 ( .C1(n20820), .C2(n21092), .A(n20819), .B(n11173), .ZN(
        P3_U2660) );
  NOR2_X1 U22923 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20821), .ZN(n20836) );
  AOI211_X1 U22924 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20821), .A(n20836), .B(
        n21093), .ZN(n20822) );
  AOI211_X1 U22925 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n21075), .A(n21769), .B(
        n20822), .ZN(n20832) );
  NOR2_X4 U22926 ( .A1(n20824), .A2(n20823), .ZN(n20914) );
  NOR2_X1 U22927 ( .A1(n20826), .A2(n20825), .ZN(n20862) );
  OR2_X1 U22928 ( .A1(n20862), .A2(n20864), .ZN(n20828) );
  OAI21_X1 U22929 ( .B1(n20829), .B2(n20828), .A(n20865), .ZN(n20827) );
  AOI21_X1 U22930 ( .B1(n20829), .B2(n20828), .A(n20827), .ZN(n20830) );
  AOI221_X1 U22931 ( .B1(n20847), .B2(P3_REIP_REG_12__SCAN_IN), .C1(n20914), 
        .C2(n20848), .A(n20830), .ZN(n20831) );
  OAI211_X1 U22932 ( .C1(n20833), .C2(n21090), .A(n20832), .B(n20831), .ZN(
        P3_U2659) );
  NAND2_X1 U22933 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20914), .ZN(n20846) );
  AOI21_X1 U22934 ( .B1(n20914), .B2(n20848), .A(n20847), .ZN(n20845) );
  AOI21_X1 U22935 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20868), .A(
        n20834), .ZN(n20842) );
  AOI21_X1 U22936 ( .B1(n20835), .B2(n21094), .A(n20864), .ZN(n20852) );
  NAND2_X1 U22937 ( .A1(n21069), .A2(n20852), .ZN(n20853) );
  NAND2_X1 U22938 ( .A1(n20836), .A2(n20838), .ZN(n20855) );
  OAI211_X1 U22939 ( .C1(n20836), .C2(n20838), .A(n21050), .B(n20855), .ZN(
        n20837) );
  OAI211_X1 U22940 ( .C1(n20843), .C2(n20853), .A(n11173), .B(n20837), .ZN(
        n20841) );
  OAI22_X1 U22941 ( .A1(n20839), .A2(n21090), .B1(n20838), .B2(n21092), .ZN(
        n20840) );
  AOI211_X1 U22942 ( .C1(n20843), .C2(n20842), .A(n20841), .B(n20840), .ZN(
        n20844) );
  OAI221_X1 U22943 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n20846), .C1(n20849), 
        .C2(n20845), .A(n20844), .ZN(P3_U2658) );
  NAND3_X1 U22944 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(P3_REIP_REG_12__SCAN_IN), .ZN(n20877) );
  AOI21_X1 U22945 ( .B1(n20877), .B2(n21098), .A(n20847), .ZN(n20889) );
  NOR2_X1 U22946 ( .A1(n20849), .A2(n20848), .ZN(n20850) );
  AOI21_X1 U22947 ( .B1(n20850), .B2(n20914), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n20861) );
  AOI22_X1 U22948 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n21056), .B1(
        P3_EBX_REG_14__SCAN_IN), .B2(n21075), .ZN(n20860) );
  INV_X1 U22949 ( .A(n20854), .ZN(n20851) );
  NOR3_X1 U22950 ( .A1(n20852), .A2(n20851), .A3(n21815), .ZN(n20858) );
  NOR2_X1 U22951 ( .A1(n20854), .A2(n20853), .ZN(n20857) );
  NOR2_X1 U22952 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20855), .ZN(n20871) );
  AOI211_X1 U22953 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20855), .A(n20871), .B(
        n21093), .ZN(n20856) );
  NOR4_X1 U22954 ( .A1(n21769), .A2(n20858), .A3(n20857), .A4(n20856), .ZN(
        n20859) );
  OAI211_X1 U22955 ( .C1(n20889), .C2(n20861), .A(n20860), .B(n20859), .ZN(
        P3_U2657) );
  AND2_X1 U22956 ( .A1(n20863), .A2(n20862), .ZN(n20866) );
  AOI21_X1 U22957 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20866), .A(
        n20864), .ZN(n20881) );
  INV_X1 U22958 ( .A(n20881), .ZN(n20879) );
  OAI21_X1 U22959 ( .B1(n20866), .B2(n20869), .A(n20865), .ZN(n20867) );
  AOI22_X1 U22960 ( .A1(n20869), .A2(n20879), .B1(n20868), .B2(n20867), .ZN(
        n20870) );
  AOI211_X1 U22961 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n21075), .A(n21769), .B(
        n20870), .ZN(n20876) );
  INV_X1 U22962 ( .A(n20914), .ZN(n20897) );
  NOR3_X1 U22963 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20877), .A3(n20897), 
        .ZN(n20891) );
  NAND2_X1 U22964 ( .A1(n20871), .A2(n20872), .ZN(n20883) );
  OAI211_X1 U22965 ( .C1(n20872), .C2(n20871), .A(n20883), .B(n21050), .ZN(
        n20873) );
  INV_X1 U22966 ( .A(n20873), .ZN(n20874) );
  AOI211_X1 U22967 ( .C1(n21056), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20891), .B(n20874), .ZN(n20875) );
  OAI211_X1 U22968 ( .C1(n20889), .C2(n20878), .A(n20876), .B(n20875), .ZN(
        P3_U2656) );
  NOR2_X1 U22969 ( .A1(n20878), .A2(n20877), .ZN(n20895) );
  NAND2_X1 U22970 ( .A1(n20895), .A2(n20914), .ZN(n20894) );
  INV_X1 U22971 ( .A(n20882), .ZN(n20880) );
  AOI221_X1 U22972 ( .B1(n20882), .B2(n20881), .C1(n20880), .C2(n20879), .A(
        n21815), .ZN(n20888) );
  NOR2_X1 U22973 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20883), .ZN(n20899) );
  AOI211_X1 U22974 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20883), .A(n20899), .B(
        n21093), .ZN(n20887) );
  INV_X1 U22975 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n20884) );
  OAI22_X1 U22976 ( .A1(n20885), .A2(n21090), .B1(n20884), .B2(n21092), .ZN(
        n20886) );
  NOR4_X1 U22977 ( .A1(n21769), .A2(n20888), .A3(n20887), .A4(n20886), .ZN(
        n20893) );
  INV_X1 U22978 ( .A(n20889), .ZN(n20890) );
  OAI21_X1 U22979 ( .B1(n20891), .B2(n20890), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n20892) );
  OAI211_X1 U22980 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n20894), .A(n20893), 
        .B(n20892), .ZN(P3_U2655) );
  NAND2_X1 U22981 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20895), .ZN(n20898) );
  NOR2_X1 U22982 ( .A1(n20910), .A2(n20898), .ZN(n20915) );
  NAND2_X1 U22983 ( .A1(n20915), .A2(n20896), .ZN(n20937) );
  NAND2_X1 U22984 ( .A1(n21098), .A2(n20937), .ZN(n20935) );
  NOR3_X1 U22985 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20898), .A3(n20897), 
        .ZN(n20903) );
  INV_X1 U22986 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20901) );
  NAND2_X1 U22987 ( .A1(n20899), .A2(n20901), .ZN(n20911) );
  OAI211_X1 U22988 ( .C1(n20899), .C2(n20901), .A(n21050), .B(n20911), .ZN(
        n20900) );
  OAI211_X1 U22989 ( .C1(n20901), .C2(n21092), .A(n11173), .B(n20900), .ZN(
        n20902) );
  AOI211_X1 U22990 ( .C1(n21056), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20903), .B(n20902), .ZN(n20909) );
  OAI21_X1 U22991 ( .B1(n20905), .B2(n20904), .A(n21065), .ZN(n20906) );
  NAND2_X1 U22992 ( .A1(n20907), .A2(n20906), .ZN(n20916) );
  OAI211_X1 U22993 ( .C1(n20907), .C2(n20906), .A(n21069), .B(n20916), .ZN(
        n20908) );
  OAI211_X1 U22994 ( .C1(n20935), .C2(n20910), .A(n20909), .B(n20908), .ZN(
        P3_U2654) );
  NOR2_X1 U22995 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20911), .ZN(n20924) );
  AOI211_X1 U22996 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20911), .A(n20924), .B(
        n21093), .ZN(n20922) );
  OAI22_X1 U22997 ( .A1(n20913), .A2(n21090), .B1(n20912), .B2(n21092), .ZN(
        n20921) );
  NAND2_X1 U22998 ( .A1(n21065), .A2(n20916), .ZN(n20917) );
  NAND2_X1 U22999 ( .A1(n20918), .A2(n20917), .ZN(n20929) );
  OAI211_X1 U23000 ( .C1(n20918), .C2(n20917), .A(n21069), .B(n20929), .ZN(
        n20919) );
  OAI221_X1 U23001 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n20951), .C1(n20923), 
        .C2(n20935), .A(n20919), .ZN(n20920) );
  OR4_X1 U23002 ( .A1(n18279), .A2(n20922), .A3(n20921), .A4(n20920), .ZN(
        P3_U2653) );
  AOI221_X1 U23003 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n20923), .C2(n20934), .A(n20951), .ZN(n20928) );
  NAND2_X1 U23004 ( .A1(n20924), .A2(n20926), .ZN(n20939) );
  OAI211_X1 U23005 ( .C1(n20924), .C2(n20926), .A(n21050), .B(n20939), .ZN(
        n20925) );
  OAI211_X1 U23006 ( .C1(n20926), .C2(n21092), .A(n11173), .B(n20925), .ZN(
        n20927) );
  AOI211_X1 U23007 ( .C1(n21056), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20928), .B(n20927), .ZN(n20933) );
  OAI211_X1 U23008 ( .C1(n20931), .C2(n20930), .A(n21069), .B(n20944), .ZN(
        n20932) );
  OAI211_X1 U23009 ( .C1(n20935), .C2(n20934), .A(n20933), .B(n20932), .ZN(
        P3_U2652) );
  NAND3_X1 U23010 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(n20936), .ZN(n20949) );
  NAND3_X1 U23011 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(P3_REIP_REG_19__SCAN_IN), .ZN(n20950) );
  NOR2_X1 U23012 ( .A1(n20950), .A2(n20937), .ZN(n20974) );
  NOR2_X1 U23013 ( .A1(n20938), .A2(n20974), .ZN(n20967) );
  NOR2_X1 U23014 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20939), .ZN(n20957) );
  AOI211_X1 U23015 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20939), .A(n20957), .B(
        n21093), .ZN(n20943) );
  INV_X1 U23016 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n20940) );
  OAI22_X1 U23017 ( .A1(n20941), .A2(n21090), .B1(n20940), .B2(n21092), .ZN(
        n20942) );
  AOI211_X1 U23018 ( .C1(n20967), .C2(P3_REIP_REG_20__SCAN_IN), .A(n20943), 
        .B(n20942), .ZN(n20948) );
  OAI211_X1 U23019 ( .C1(n20946), .C2(n20945), .A(n21069), .B(n20953), .ZN(
        n20947) );
  OAI211_X1 U23020 ( .C1(n20949), .C2(n20951), .A(n20948), .B(n20947), .ZN(
        P3_U2651) );
  AOI22_X1 U23021 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n21056), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n21075), .ZN(n20961) );
  AOI22_X1 U23022 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20967), .B1(n20986), 
        .B2(n20952), .ZN(n20960) );
  NAND2_X1 U23023 ( .A1(n21065), .A2(n20953), .ZN(n20954) );
  NAND2_X1 U23024 ( .A1(n20955), .A2(n20954), .ZN(n20968) );
  OAI211_X1 U23025 ( .C1(n20955), .C2(n20954), .A(n21069), .B(n20968), .ZN(
        n20959) );
  NAND2_X1 U23026 ( .A1(n20957), .A2(n20956), .ZN(n20962) );
  OAI211_X1 U23027 ( .C1(n20957), .C2(n20956), .A(n21050), .B(n20962), .ZN(
        n20958) );
  NAND4_X1 U23028 ( .A1(n20961), .A2(n20960), .A3(n20959), .A4(n20958), .ZN(
        P3_U2650) );
  NOR2_X1 U23029 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20962), .ZN(n20981) );
  AOI211_X1 U23030 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20962), .A(n20981), .B(
        n21093), .ZN(n20966) );
  OAI22_X1 U23031 ( .A1(n20964), .A2(n21090), .B1(n20963), .B2(n21092), .ZN(
        n20965) );
  AOI211_X1 U23032 ( .C1(n20967), .C2(P3_REIP_REG_22__SCAN_IN), .A(n20966), 
        .B(n20965), .ZN(n20973) );
  NAND2_X1 U23033 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n20975) );
  OAI211_X1 U23034 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n20986), .B(n20975), .ZN(n20972) );
  NAND2_X1 U23035 ( .A1(n21065), .A2(n20968), .ZN(n20969) );
  NAND2_X1 U23036 ( .A1(n20970), .A2(n20969), .ZN(n20977) );
  OAI211_X1 U23037 ( .C1(n20970), .C2(n20969), .A(n21069), .B(n20977), .ZN(
        n20971) );
  NAND3_X1 U23038 ( .A1(n20973), .A2(n20972), .A3(n20971), .ZN(P3_U2649) );
  AOI22_X1 U23039 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n21056), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n21075), .ZN(n20985) );
  NAND4_X1 U23040 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .A4(n20974), .ZN(n20998) );
  AND2_X1 U23041 ( .A1(n21098), .A2(n20998), .ZN(n20992) );
  NOR2_X1 U23042 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20975), .ZN(n20976) );
  AOI22_X1 U23043 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n20992), .B1(n20986), 
        .B2(n20976), .ZN(n20984) );
  NAND2_X1 U23044 ( .A1(n21065), .A2(n20977), .ZN(n20978) );
  NAND2_X1 U23045 ( .A1(n20979), .A2(n20978), .ZN(n20993) );
  OAI211_X1 U23046 ( .C1(n20979), .C2(n20978), .A(n21069), .B(n20993), .ZN(
        n20983) );
  INV_X1 U23047 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20980) );
  NAND2_X1 U23048 ( .A1(n20981), .A2(n20980), .ZN(n20987) );
  OAI211_X1 U23049 ( .C1(n20981), .C2(n20980), .A(n21050), .B(n20987), .ZN(
        n20982) );
  NAND4_X1 U23050 ( .A1(n20985), .A2(n20984), .A3(n20983), .A4(n20982), .ZN(
        P3_U2648) );
  NAND4_X1 U23051 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .A4(n20986), .ZN(n20999) );
  NOR2_X1 U23052 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20987), .ZN(n21007) );
  AOI211_X1 U23053 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20987), .A(n21007), .B(
        n21093), .ZN(n20991) );
  OAI22_X1 U23054 ( .A1(n20989), .A2(n21090), .B1(n20988), .B2(n21092), .ZN(
        n20990) );
  AOI211_X1 U23055 ( .C1(n20992), .C2(P3_REIP_REG_24__SCAN_IN), .A(n20991), 
        .B(n20990), .ZN(n20997) );
  NAND2_X1 U23056 ( .A1(n21065), .A2(n20993), .ZN(n20994) );
  NAND2_X1 U23057 ( .A1(n20995), .A2(n20994), .ZN(n21003) );
  OAI211_X1 U23058 ( .C1(n20995), .C2(n20994), .A(n21069), .B(n21003), .ZN(
        n20996) );
  OAI211_X1 U23059 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n20999), .A(n20997), 
        .B(n20996), .ZN(P3_U2647) );
  AOI22_X1 U23060 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n21056), .B1(
        P3_EBX_REG_25__SCAN_IN), .B2(n21075), .ZN(n21011) );
  NOR2_X1 U23061 ( .A1(n21000), .A2(n20998), .ZN(n21013) );
  NOR2_X1 U23062 ( .A1(n21013), .A2(n21001), .ZN(n21002) );
  NOR2_X1 U23063 ( .A1(n21000), .A2(n20999), .ZN(n21012) );
  AOI22_X1 U23064 ( .A1(n21002), .A2(n21098), .B1(n21012), .B2(n21001), .ZN(
        n21010) );
  OAI211_X1 U23065 ( .C1(n21005), .C2(n21004), .A(n21069), .B(n21019), .ZN(
        n21009) );
  NAND2_X1 U23066 ( .A1(n21007), .A2(n21006), .ZN(n21014) );
  OAI211_X1 U23067 ( .C1(n21007), .C2(n21006), .A(n21050), .B(n21014), .ZN(
        n21008) );
  NAND4_X1 U23068 ( .A1(n21011), .A2(n21010), .A3(n21009), .A4(n21008), .ZN(
        P3_U2646) );
  NAND2_X1 U23069 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n21012), .ZN(n21024) );
  NAND3_X1 U23070 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n21013), .ZN(n21046) );
  AND2_X1 U23071 ( .A1(n21098), .A2(n21046), .ZN(n21042) );
  NOR2_X1 U23072 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n21014), .ZN(n21031) );
  AOI211_X1 U23073 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n21014), .A(n21031), .B(
        n21093), .ZN(n21018) );
  OAI22_X1 U23074 ( .A1(n21016), .A2(n21090), .B1(n21015), .B2(n21092), .ZN(
        n21017) );
  AOI211_X1 U23075 ( .C1(n21042), .C2(P3_REIP_REG_26__SCAN_IN), .A(n21018), 
        .B(n21017), .ZN(n21023) );
  OAI211_X1 U23076 ( .C1(n21021), .C2(n21020), .A(n21069), .B(n21027), .ZN(
        n21022) );
  OAI211_X1 U23077 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n21024), .A(n21023), 
        .B(n21022), .ZN(P3_U2645) );
  AOI22_X1 U23078 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n21056), .B1(
        P3_EBX_REG_27__SCAN_IN), .B2(n21075), .ZN(n21035) );
  AOI22_X1 U23079 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21042), .B1(n21066), 
        .B2(n21026), .ZN(n21034) );
  NAND2_X1 U23080 ( .A1(n21065), .A2(n21027), .ZN(n21028) );
  NAND2_X1 U23081 ( .A1(n21029), .A2(n21028), .ZN(n21057) );
  OAI211_X1 U23082 ( .C1(n21029), .C2(n21028), .A(n21069), .B(n21057), .ZN(
        n21033) );
  NAND2_X1 U23083 ( .A1(n21031), .A2(n21030), .ZN(n21037) );
  OAI211_X1 U23084 ( .C1(n21031), .C2(n21030), .A(n21050), .B(n21037), .ZN(
        n21032) );
  NAND4_X1 U23085 ( .A1(n21035), .A2(n21034), .A3(n21033), .A4(n21032), .ZN(
        P3_U2644) );
  NAND2_X1 U23086 ( .A1(n21065), .A2(n21057), .ZN(n21036) );
  XOR2_X1 U23087 ( .A(n21058), .B(n21036), .Z(n21045) );
  NOR2_X1 U23088 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21037), .ZN(n21051) );
  AOI211_X1 U23089 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21037), .A(n21051), .B(
        n21093), .ZN(n21041) );
  OAI22_X1 U23090 ( .A1(n21039), .A2(n21090), .B1(n21038), .B2(n21092), .ZN(
        n21040) );
  AOI211_X1 U23091 ( .C1(n21042), .C2(P3_REIP_REG_28__SCAN_IN), .A(n21041), 
        .B(n21040), .ZN(n21044) );
  NAND2_X1 U23092 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n21048) );
  OAI211_X1 U23093 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n21066), .B(n21048), .ZN(n21043) );
  OAI211_X1 U23094 ( .C1(n21815), .C2(n21045), .A(n21044), .B(n21043), .ZN(
        P3_U2643) );
  NAND3_X1 U23095 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n21047) );
  OAI21_X1 U23096 ( .B1(n21047), .B2(n21046), .A(n21098), .ZN(n21082) );
  INV_X1 U23097 ( .A(n21066), .ZN(n21049) );
  NOR3_X1 U23098 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n21049), .A3(n21048), 
        .ZN(n21055) );
  NAND2_X1 U23099 ( .A1(n21051), .A2(n21052), .ZN(n21070) );
  NAND2_X1 U23100 ( .A1(n21050), .A2(n21070), .ZN(n21067) );
  NOR2_X1 U23101 ( .A1(n21051), .A2(n21052), .ZN(n21053) );
  OAI22_X1 U23102 ( .A1(n21067), .A2(n21053), .B1(n21092), .B2(n21052), .ZN(
        n21054) );
  AOI211_X1 U23103 ( .C1(n21056), .C2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n21055), .B(n21054), .ZN(n21062) );
  OAI21_X1 U23104 ( .B1(n21058), .B2(n21057), .A(n21065), .ZN(n21059) );
  OAI211_X1 U23105 ( .C1(n21060), .C2(n21059), .A(n21069), .B(n21064), .ZN(
        n21061) );
  OAI211_X1 U23106 ( .C1(n21082), .C2(n21063), .A(n21062), .B(n21061), .ZN(
        P3_U2642) );
  NAND4_X1 U23107 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n21066), .A3(
        P3_REIP_REG_29__SCAN_IN), .A4(P3_REIP_REG_27__SCAN_IN), .ZN(n21078) );
  NOR2_X1 U23108 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n21078), .ZN(n21080) );
  OAI22_X1 U23109 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n21067), .B1(n11550), 
        .B2(n21090), .ZN(n21068) );
  NOR2_X1 U23110 ( .A1(n21093), .A2(n21070), .ZN(n21074) );
  OAI21_X1 U23111 ( .B1(n21075), .B2(n21074), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n21071) );
  OAI211_X1 U23112 ( .C1(n21079), .C2(n21082), .A(n21072), .B(n21071), .ZN(
        P3_U2641) );
  AOI22_X1 U23113 ( .A1(n21075), .A2(P3_EBX_REG_31__SCAN_IN), .B1(n21074), 
        .B2(n21073), .ZN(n21089) );
  NOR2_X1 U23114 ( .A1(n21077), .A2(n21076), .ZN(n21087) );
  NOR3_X1 U23115 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21079), .A3(n21078), 
        .ZN(n21085) );
  INV_X1 U23116 ( .A(n21080), .ZN(n21083) );
  AOI21_X1 U23117 ( .B1(n21083), .B2(n21082), .A(n21081), .ZN(n21084) );
  AOI211_X1 U23118 ( .C1(n21087), .C2(n21086), .A(n21085), .B(n21084), .ZN(
        n21088) );
  OAI211_X1 U23119 ( .C1(n11549), .C2(n21090), .A(n21089), .B(n21088), .ZN(
        P3_U2640) );
  AOI21_X1 U23120 ( .B1(n21093), .B2(n21092), .A(n21091), .ZN(n21097) );
  NOR3_X1 U23121 ( .A1(n21095), .A2(n21329), .A3(n21094), .ZN(n21096) );
  AOI211_X1 U23122 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n21098), .A(n21097), .B(
        n21096), .ZN(n21099) );
  OAI21_X1 U23123 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21100), .A(
        n21099), .ZN(P3_U2671) );
  NAND2_X1 U23124 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n21157) );
  NAND2_X1 U23125 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n21270) );
  NOR2_X2 U23126 ( .A1(n21152), .A2(n21149), .ZN(n21131) );
  NAND4_X1 U23127 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(n21131), .ZN(n21130) );
  NOR2_X2 U23128 ( .A1(n21130), .A2(n21129), .ZN(n21262) );
  NAND3_X1 U23129 ( .A1(n21263), .A2(n21262), .A3(P3_EAX_REG_8__SCAN_IN), .ZN(
        n21122) );
  NAND2_X1 U23130 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21126), .ZN(n21119) );
  NOR2_X1 U23131 ( .A1(n21157), .A2(n21119), .ZN(n21248) );
  INV_X1 U23132 ( .A(n21248), .ZN(n21109) );
  NAND2_X1 U23133 ( .A1(n21109), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n21108) );
  NAND2_X1 U23134 ( .A1(n21280), .A2(n21197), .ZN(n21249) );
  INV_X1 U23135 ( .A(n11189), .ZN(n21256) );
  AOI22_X1 U23136 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21278), .B1(n21277), .B2(
        n21106), .ZN(n21107) );
  OAI221_X1 U23137 ( .B1(n21109), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n21108), 
        .C2(n21256), .A(n21107), .ZN(P3_U2722) );
  INV_X1 U23138 ( .A(n21278), .ZN(n21141) );
  INV_X1 U23139 ( .A(n21119), .ZN(n21113) );
  AOI22_X1 U23140 ( .A1(n21113), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n11189), .ZN(n21111) );
  OAI222_X1 U23141 ( .A1(n21141), .A2(n21224), .B1(n21248), .B2(n21111), .C1(
        n21274), .C2(n21110), .ZN(P3_U2723) );
  NOR2_X1 U23142 ( .A1(n21112), .A2(n21119), .ZN(n21116) );
  AOI21_X1 U23143 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n11189), .A(n21113), .ZN(
        n21115) );
  OAI222_X1 U23144 ( .A1(n21141), .A2(n21117), .B1(n21116), .B2(n21115), .C1(
        n21274), .C2(n21114), .ZN(P3_U2724) );
  AOI22_X1 U23145 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21278), .B1(n21277), .B2(
        n21118), .ZN(n21121) );
  OAI211_X1 U23146 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n21126), .A(n11189), .B(
        n21119), .ZN(n21120) );
  NAND2_X1 U23147 ( .A1(n21121), .A2(n21120), .ZN(P3_U2725) );
  INV_X1 U23148 ( .A(n21122), .ZN(n21123) );
  AOI21_X1 U23149 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n11189), .A(n21123), .ZN(
        n21125) );
  OAI222_X1 U23150 ( .A1(n21141), .A2(n21127), .B1(n21126), .B2(n21125), .C1(
        n21274), .C2(n21124), .ZN(P3_U2726) );
  OR2_X1 U23151 ( .A1(n21256), .A2(n21262), .ZN(n21266) );
  AOI22_X1 U23152 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21278), .B1(n21277), .B2(
        n21353), .ZN(n21128) );
  OAI221_X1 U23153 ( .B1(n21266), .B2(n21130), .C1(n21266), .C2(n21129), .A(
        n21128), .ZN(P3_U2728) );
  NAND2_X1 U23154 ( .A1(n21263), .A2(n21131), .ZN(n21146) );
  NOR2_X1 U23155 ( .A1(n21145), .A2(n21146), .ZN(n21137) );
  AND2_X1 U23156 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n21137), .ZN(n21140) );
  AOI21_X1 U23157 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n11189), .A(n21140), .ZN(
        n21135) );
  NAND3_X1 U23158 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .ZN(n21132) );
  NOR2_X1 U23159 ( .A1(n21132), .A2(n21146), .ZN(n21134) );
  OAI222_X1 U23160 ( .A1(n21136), .A2(n21141), .B1(n21135), .B2(n21134), .C1(
        n21274), .C2(n21133), .ZN(P3_U2729) );
  AOI21_X1 U23161 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n11189), .A(n21137), .ZN(
        n21139) );
  OAI222_X1 U23162 ( .A1(n21142), .A2(n21141), .B1(n21140), .B2(n21139), .C1(
        n21274), .C2(n21138), .ZN(P3_U2730) );
  NAND2_X1 U23163 ( .A1(n11189), .A2(n21146), .ZN(n21150) );
  AOI22_X1 U23164 ( .A1(n21278), .A2(BUF2_REG_4__SCAN_IN), .B1(n21277), .B2(
        n21143), .ZN(n21144) );
  OAI221_X1 U23165 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21146), .C1(n21145), 
        .C2(n21150), .A(n21144), .ZN(P3_U2731) );
  AOI22_X1 U23166 ( .A1(n21278), .A2(BUF2_REG_3__SCAN_IN), .B1(n21277), .B2(
        n21147), .ZN(n21148) );
  OAI221_X1 U23167 ( .B1(n21150), .B2(n21152), .C1(n21150), .C2(n21149), .A(
        n21148), .ZN(P3_U2732) );
  AOI22_X1 U23168 ( .A1(n21278), .A2(BUF2_REG_2__SCAN_IN), .B1(n21277), .B2(
        n21151), .ZN(n21155) );
  OAI211_X1 U23169 ( .C1(n21153), .C2(P3_EAX_REG_2__SCAN_IN), .A(n11189), .B(
        n21152), .ZN(n21154) );
  NAND2_X1 U23170 ( .A1(n21155), .A2(n21154), .ZN(P3_U2733) );
  NOR4_X1 U23171 ( .A1(n21267), .A2(n21253), .A3(n21157), .A4(n21156), .ZN(
        n21158) );
  NOR2_X2 U23172 ( .A1(n21258), .A2(n21257), .ZN(n21255) );
  NAND2_X1 U23173 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n21189), .ZN(n21185) );
  NAND2_X1 U23174 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n21179), .ZN(n21166) );
  NAND2_X1 U23175 ( .A1(n11189), .A2(n21166), .ZN(n21174) );
  NOR2_X2 U23176 ( .A1(n21160), .A2(n21249), .ZN(n21243) );
  OAI22_X1 U23178 ( .A1(n21163), .A2(n21274), .B1(n21162), .B2(n22600), .ZN(
        n21164) );
  AOI21_X1 U23179 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21243), .A(n21164), .ZN(
        n21165) );
  OAI221_X1 U23180 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21166), .C1(n21171), 
        .C2(n21174), .A(n21165), .ZN(P3_U2714) );
  AOI22_X1 U23181 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n11163), .ZN(n21168) );
  OAI211_X1 U23182 ( .C1(n21179), .C2(P3_EAX_REG_20__SCAN_IN), .A(n11189), .B(
        n21166), .ZN(n21167) );
  OAI211_X1 U23183 ( .C1(n21169), .C2(n21274), .A(n21168), .B(n21167), .ZN(
        P3_U2715) );
  NOR2_X1 U23184 ( .A1(n21171), .A2(n21170), .ZN(n21172) );
  NAND4_X1 U23185 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(n21172), .ZN(n21196) );
  NOR2_X1 U23186 ( .A1(n21197), .A2(n21244), .ZN(n21191) );
  NAND2_X1 U23187 ( .A1(n21191), .A2(n21195), .ZN(n21178) );
  AOI22_X1 U23188 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n11163), .B1(n21277), .B2(
        n21173), .ZN(n21177) );
  NAND2_X1 U23189 ( .A1(n21263), .A2(n21280), .ZN(n21282) );
  OAI21_X1 U23190 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21282), .A(n21174), .ZN(
        n21175) );
  AOI22_X1 U23191 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n21243), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n21175), .ZN(n21176) );
  OAI211_X1 U23192 ( .C1(n21196), .C2(n21178), .A(n21177), .B(n21176), .ZN(
        P3_U2713) );
  AOI22_X1 U23193 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n11163), .ZN(n21183) );
  AOI211_X1 U23194 ( .C1(n21180), .C2(n21185), .A(n21179), .B(n21256), .ZN(
        n21181) );
  INV_X1 U23195 ( .A(n21181), .ZN(n21182) );
  OAI211_X1 U23196 ( .C1(n21184), .C2(n21274), .A(n21183), .B(n21182), .ZN(
        P3_U2716) );
  AOI22_X1 U23197 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n11163), .ZN(n21187) );
  OAI211_X1 U23198 ( .C1(n21189), .C2(P3_EAX_REG_18__SCAN_IN), .A(n11189), .B(
        n21185), .ZN(n21186) );
  OAI211_X1 U23199 ( .C1(n21188), .C2(n21274), .A(n21187), .B(n21186), .ZN(
        P3_U2717) );
  AOI22_X1 U23200 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n11163), .ZN(n21193) );
  INV_X1 U23201 ( .A(n21189), .ZN(n21190) );
  OAI211_X1 U23202 ( .C1(n21191), .C2(P3_EAX_REG_17__SCAN_IN), .A(n11189), .B(
        n21190), .ZN(n21192) );
  OAI211_X1 U23203 ( .C1(n21194), .C2(n21274), .A(n21193), .B(n21192), .ZN(
        P3_U2718) );
  AOI22_X1 U23204 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n11163), .ZN(n21200) );
  NOR3_X2 U23205 ( .A1(n21244), .A2(n21196), .A3(n21195), .ZN(n21238) );
  NAND2_X1 U23206 ( .A1(n21238), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21237) );
  OAI211_X1 U23207 ( .C1(n21198), .C2(P3_EAX_REG_25__SCAN_IN), .A(n11189), .B(
        n11215), .ZN(n21199) );
  OAI211_X1 U23208 ( .C1(n21201), .C2(n21274), .A(n21200), .B(n21199), .ZN(
        P3_U2710) );
  AOI22_X1 U23209 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n11163), .B1(n21277), .B2(
        n21202), .ZN(n21203) );
  INV_X1 U23210 ( .A(n21203), .ZN(n21206) );
  NOR2_X2 U23211 ( .A1(n11215), .A2(n21204), .ZN(n21226) );
  AOI211_X1 U23212 ( .C1(n21204), .C2(n11215), .A(n21226), .B(n21256), .ZN(
        n21205) );
  AOI211_X1 U23213 ( .C1(n21243), .C2(BUF2_REG_10__SCAN_IN), .A(n21206), .B(
        n21205), .ZN(n21207) );
  INV_X1 U23214 ( .A(n21207), .ZN(P3_U2709) );
  NAND2_X1 U23215 ( .A1(n21211), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21210) );
  OAI22_X1 U23216 ( .A1(n21256), .A2(n21211), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n21282), .ZN(n21208) );
  AOI22_X1 U23217 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n11163), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n21208), .ZN(n21209) );
  OAI21_X1 U23218 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n21210), .A(n21209), .ZN(
        P3_U2704) );
  AOI22_X1 U23219 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n11163), .ZN(n21213) );
  OAI211_X1 U23220 ( .C1(n21211), .C2(P3_EAX_REG_30__SCAN_IN), .A(n11189), .B(
        n21210), .ZN(n21212) );
  OAI211_X1 U23221 ( .C1(n21214), .C2(n21274), .A(n21213), .B(n21212), .ZN(
        P3_U2705) );
  AOI22_X1 U23222 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n11163), .ZN(n21217) );
  OAI211_X1 U23223 ( .C1(n11217), .C2(P3_EAX_REG_29__SCAN_IN), .A(n11189), .B(
        n21215), .ZN(n21216) );
  OAI211_X1 U23224 ( .C1(n21218), .C2(n21274), .A(n21217), .B(n21216), .ZN(
        P3_U2706) );
  INV_X1 U23225 ( .A(n21243), .ZN(n21236) );
  AOI22_X1 U23226 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n11163), .B1(n21277), .B2(
        n21219), .ZN(n21223) );
  AOI211_X1 U23227 ( .C1(n21220), .C2(n21225), .A(n11217), .B(n21256), .ZN(
        n21221) );
  INV_X1 U23228 ( .A(n21221), .ZN(n21222) );
  OAI211_X1 U23229 ( .C1(n21236), .C2(n21224), .A(n21223), .B(n21222), .ZN(
        P3_U2707) );
  AOI22_X1 U23230 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n11163), .ZN(n21228) );
  OAI211_X1 U23231 ( .C1(n21226), .C2(P3_EAX_REG_27__SCAN_IN), .A(n11189), .B(
        n21225), .ZN(n21227) );
  OAI211_X1 U23232 ( .C1(n21229), .C2(n21274), .A(n21228), .B(n21227), .ZN(
        P3_U2708) );
  AOI22_X1 U23233 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n11163), .B1(n21277), .B2(
        n21230), .ZN(n21234) );
  OAI211_X1 U23234 ( .C1(n21232), .C2(P3_EAX_REG_24__SCAN_IN), .A(n11189), .B(
        n21231), .ZN(n21233) );
  OAI211_X1 U23235 ( .C1(n21236), .C2(n21235), .A(n21234), .B(n21233), .ZN(
        P3_U2711) );
  AOI22_X1 U23236 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n11163), .ZN(n21240) );
  OAI211_X1 U23237 ( .C1(n21238), .C2(P3_EAX_REG_23__SCAN_IN), .A(n11189), .B(
        n21237), .ZN(n21239) );
  OAI211_X1 U23238 ( .C1(n21241), .C2(n21274), .A(n21240), .B(n21239), .ZN(
        P3_U2712) );
  AOI22_X1 U23239 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21243), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n11163), .ZN(n21246) );
  OAI211_X1 U23240 ( .C1(n21255), .C2(P3_EAX_REG_16__SCAN_IN), .A(n11189), .B(
        n21244), .ZN(n21245) );
  OAI211_X1 U23241 ( .C1(n21247), .C2(n21274), .A(n21246), .B(n21245), .ZN(
        P3_U2719) );
  NAND2_X1 U23242 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21248), .ZN(n21254) );
  NAND2_X1 U23243 ( .A1(n11189), .A2(n21258), .ZN(n21252) );
  AOI22_X1 U23244 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21278), .B1(n21277), .B2(
        n21250), .ZN(n21251) );
  OAI221_X1 U23245 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n21254), .C1(n21253), 
        .C2(n21252), .A(n21251), .ZN(P3_U2721) );
  AOI211_X1 U23246 ( .C1(n21258), .C2(n21257), .A(n21256), .B(n21255), .ZN(
        n21259) );
  AOI21_X1 U23247 ( .B1(n21278), .B2(BUF2_REG_15__SCAN_IN), .A(n21259), .ZN(
        n21260) );
  OAI21_X1 U23248 ( .B1(n21261), .B2(n21274), .A(n21260), .ZN(P3_U2720) );
  NAND2_X1 U23249 ( .A1(n21263), .A2(n21262), .ZN(n21268) );
  AOI22_X1 U23250 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21278), .B1(n21277), .B2(
        n21264), .ZN(n21265) );
  OAI221_X1 U23251 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n21268), .C1(n21267), 
        .C2(n21266), .A(n21265), .ZN(P3_U2727) );
  AOI22_X1 U23252 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21278), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n21269), .ZN(n21273) );
  INV_X1 U23253 ( .A(n21282), .ZN(n21271) );
  OAI211_X1 U23254 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(P3_EAX_REG_1__SCAN_IN), 
        .A(n21271), .B(n21270), .ZN(n21272) );
  OAI211_X1 U23255 ( .C1(n21275), .C2(n21274), .A(n21273), .B(n21272), .ZN(
        P3_U2734) );
  AOI22_X1 U23256 ( .A1(n21278), .A2(BUF2_REG_0__SCAN_IN), .B1(n21277), .B2(
        n21276), .ZN(n21279) );
  OAI221_X1 U23257 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21282), .C1(n21281), 
        .C2(n21280), .A(n21279), .ZN(P3_U2735) );
  INV_X1 U23258 ( .A(n21331), .ZN(n21334) );
  NOR2_X1 U23259 ( .A1(n21283), .A2(n21754), .ZN(n21285) );
  AOI22_X1 U23260 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21759), .B1(
        n21285), .B2(n21310), .ZN(n21786) );
  AOI222_X1 U23261 ( .A1(n21468), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21786), 
        .B2(n21329), .C1(n21310), .C2(n21822), .ZN(n21284) );
  AOI22_X1 U23262 ( .A1(n21334), .A2(n21310), .B1(n21284), .B2(n21331), .ZN(
        P3_U3290) );
  AOI21_X1 U23263 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21754), .A(
        n21742), .ZN(n21295) );
  OAI22_X1 U23264 ( .A1(n21285), .A2(n21286), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21295), .ZN(n21785) );
  INV_X1 U23265 ( .A(n21286), .ZN(n21288) );
  AOI22_X1 U23266 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18421), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21390), .ZN(n21300) );
  NAND2_X1 U23267 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21301) );
  INV_X1 U23268 ( .A(n21301), .ZN(n21287) );
  AOI222_X1 U23269 ( .A1(n21785), .A2(n21329), .B1(n21288), .B2(n21822), .C1(
        n21300), .C2(n21287), .ZN(n21289) );
  AOI22_X1 U23270 ( .A1(n21334), .A2(n21296), .B1(n21289), .B2(n21331), .ZN(
        P3_U3289) );
  NAND2_X1 U23271 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21294), .ZN(
        n21308) );
  INV_X1 U23272 ( .A(n21601), .ZN(n21782) );
  AOI22_X1 U23273 ( .A1(n21293), .A2(n21292), .B1(n21291), .B2(n21290), .ZN(
        n21319) );
  INV_X1 U23274 ( .A(n21294), .ZN(n21303) );
  AOI211_X1 U23275 ( .C1(n21328), .C2(n21319), .A(n21303), .B(n21772), .ZN(
        n21298) );
  AOI221_X1 U23276 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C1(n21772), .C2(n21296), .A(
        n21295), .ZN(n21297) );
  AOI211_X1 U23277 ( .C1(n21782), .C2(n21299), .A(n21298), .B(n21297), .ZN(
        n21771) );
  OAI22_X1 U23278 ( .A1(n21771), .A2(n21302), .B1(n21301), .B2(n21300), .ZN(
        n21306) );
  NAND2_X1 U23279 ( .A1(n21303), .A2(n21822), .ZN(n21304) );
  OAI21_X1 U23280 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n21304), .A(
        n21331), .ZN(n21305) );
  OAI22_X1 U23281 ( .A1(n21306), .A2(n21305), .B1(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n21331), .ZN(n21307) );
  OAI21_X1 U23282 ( .B1(n21309), .B2(n21308), .A(n21307), .ZN(P3_U3288) );
  NAND2_X1 U23283 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21310), .ZN(
        n21327) );
  NOR2_X1 U23284 ( .A1(n21314), .A2(n21311), .ZN(n21356) );
  INV_X1 U23285 ( .A(n21356), .ZN(n21322) );
  NAND2_X1 U23286 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21312), .ZN(
        n21313) );
  OAI21_X1 U23287 ( .B1(n21314), .B2(n21316), .A(n21313), .ZN(n21321) );
  NOR2_X1 U23288 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21315), .ZN(
        n21317) );
  OAI22_X1 U23289 ( .A1(n21319), .A2(n21318), .B1(n21317), .B2(n21316), .ZN(
        n21320) );
  AOI21_X1 U23290 ( .B1(n21322), .B2(n21321), .A(n21320), .ZN(n21326) );
  INV_X1 U23291 ( .A(n21324), .ZN(n21323) );
  OAI221_X1 U23292 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21324), 
        .C1(n21333), .C2(n21323), .A(n21782), .ZN(n21325) );
  OAI211_X1 U23293 ( .C1(n21328), .C2(n21327), .A(n21326), .B(n21325), .ZN(
        n21775) );
  AOI22_X1 U23294 ( .A1(n21822), .A2(n21330), .B1(n21329), .B2(n21775), .ZN(
        n21332) );
  AOI22_X1 U23295 ( .A1(n21334), .A2(n21333), .B1(n21332), .B2(n21331), .ZN(
        P3_U3285) );
  INV_X1 U23296 ( .A(n21335), .ZN(n21372) );
  OAI21_X1 U23297 ( .B1(n21338), .B2(n21337), .A(n21336), .ZN(n21347) );
  OAI21_X1 U23298 ( .B1(n21342), .B2(n21341), .A(n21339), .ZN(n21340) );
  AOI21_X1 U23299 ( .B1(n21342), .B2(n21341), .A(n21340), .ZN(n21796) );
  NOR3_X1 U23300 ( .A1(n21344), .A2(n21796), .A3(n21343), .ZN(n21346) );
  AOI211_X1 U23301 ( .C1(n21348), .C2(n21347), .A(n21346), .B(n21345), .ZN(
        n21350) );
  AOI221_X4 U23302 ( .B1(n21351), .B2(n21350), .C1(n21349), .C2(n21350), .A(
        n21807), .ZN(n21757) );
  NAND2_X1 U23303 ( .A1(n21352), .A2(n21613), .ZN(n21778) );
  NOR2_X2 U23304 ( .A1(n21778), .A2(n21353), .ZN(n21679) );
  AOI22_X1 U23305 ( .A1(n21679), .A2(n21701), .B1(n21780), .B2(n21472), .ZN(
        n21479) );
  NAND2_X1 U23306 ( .A1(n21696), .A2(n21354), .ZN(n21358) );
  NAND3_X1 U23307 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21432) );
  NOR2_X1 U23308 ( .A1(n21440), .A2(n21432), .ZN(n21444) );
  OAI21_X1 U23309 ( .B1(n21390), .B2(n21468), .A(n21399), .ZN(n21403) );
  NAND2_X1 U23310 ( .A1(n21444), .A2(n21403), .ZN(n21446) );
  NOR2_X1 U23311 ( .A1(n21478), .A2(n21446), .ZN(n21470) );
  NAND2_X1 U23312 ( .A1(n21696), .A2(n21470), .ZN(n21574) );
  NOR2_X1 U23313 ( .A1(n21355), .A2(n21574), .ZN(n21548) );
  NAND2_X1 U23314 ( .A1(n21357), .A2(n21356), .ZN(n21753) );
  NOR2_X1 U23315 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21742), .ZN(
        n21379) );
  NOR2_X1 U23316 ( .A1(n21707), .A2(n21379), .ZN(n21388) );
  NAND2_X1 U23317 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21404) );
  NOR2_X1 U23318 ( .A1(n21432), .A2(n21404), .ZN(n21423) );
  NAND2_X1 U23319 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21423), .ZN(
        n21445) );
  NOR2_X1 U23320 ( .A1(n21456), .A2(n21445), .ZN(n21758) );
  NAND2_X1 U23321 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21758), .ZN(
        n21741) );
  NOR2_X1 U23322 ( .A1(n21358), .A2(n21741), .ZN(n21360) );
  AOI22_X1 U23323 ( .A1(n21782), .A2(n21548), .B1(n21388), .B2(n21360), .ZN(
        n21591) );
  OAI21_X1 U23324 ( .B1(n21479), .B2(n21358), .A(n21591), .ZN(n21583) );
  NAND2_X1 U23325 ( .A1(n21757), .A2(n21583), .ZN(n21695) );
  NOR2_X1 U23326 ( .A1(n21359), .A2(n21778), .ZN(n21636) );
  INV_X1 U23327 ( .A(n21754), .ZN(n21598) );
  OAI221_X1 U23328 ( .B1(n21598), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n21598), .C2(n21360), .A(n21757), .ZN(n21683) );
  INV_X1 U23329 ( .A(n21732), .ZN(n21745) );
  INV_X1 U23330 ( .A(n21360), .ZN(n21595) );
  NOR2_X1 U23331 ( .A1(n21548), .A2(n21601), .ZN(n21361) );
  AOI221_X1 U23332 ( .B1(n21595), .B2(n21742), .C1(n21686), .C2(n21742), .A(
        n21361), .ZN(n21681) );
  AOI22_X1 U23333 ( .A1(n21679), .A2(n21363), .B1(n21780), .B2(n21362), .ZN(
        n21364) );
  OAI211_X1 U23334 ( .C1(n21745), .C2(n21365), .A(n21681), .B(n21364), .ZN(
        n21532) );
  AOI211_X1 U23335 ( .C1(n21754), .C2(n21366), .A(n21683), .B(n21532), .ZN(
        n21367) );
  NOR3_X1 U23336 ( .A1(n18279), .A2(n21367), .A3(n21533), .ZN(n21368) );
  AOI211_X1 U23337 ( .C1(n21765), .C2(n21370), .A(n21369), .B(n21368), .ZN(
        n21371) );
  OAI21_X1 U23338 ( .B1(n21372), .B2(n21695), .A(n21371), .ZN(P3_U2841) );
  NAND2_X1 U23339 ( .A1(n21757), .A2(n21780), .ZN(n21633) );
  OR2_X1 U23340 ( .A1(n21747), .A2(n21778), .ZN(n21454) );
  NOR2_X2 U23341 ( .A1(n21769), .A2(n21757), .ZN(n21730) );
  NOR2_X1 U23342 ( .A1(n11173), .A2(n21373), .ZN(n21375) );
  NOR2_X1 U23343 ( .A1(n21782), .A2(n21754), .ZN(n21689) );
  AOI221_X1 U23344 ( .B1(n21689), .B2(n21468), .C1(n21759), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21747), .ZN(n21374) );
  AOI211_X1 U23345 ( .C1(n21730), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21375), .B(n21374), .ZN(n21376) );
  OAI221_X1 U23346 ( .B1(n21378), .B2(n21633), .C1(n21377), .C2(n21454), .A(
        n21376), .ZN(P3_U2862) );
  NOR2_X1 U23347 ( .A1(n21613), .A2(n21379), .ZN(n21381) );
  NOR2_X1 U23348 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21689), .ZN(
        n21380) );
  MUX2_X1 U23349 ( .A(n21381), .B(n21380), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21385) );
  OAI22_X1 U23350 ( .A1(n21383), .A2(n21633), .B1(n21382), .B2(n21454), .ZN(
        n21384) );
  AOI21_X1 U23351 ( .B1(n21757), .B2(n21385), .A(n21384), .ZN(n21387) );
  NAND2_X1 U23352 ( .A1(n21769), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n21386) );
  OAI211_X1 U23353 ( .C1(n21712), .C2(n21390), .A(n21387), .B(n21386), .ZN(
        P3_U2861) );
  NOR2_X1 U23354 ( .A1(n21468), .A2(n21404), .ZN(n21401) );
  NOR2_X1 U23355 ( .A1(n21601), .A2(n21403), .ZN(n21400) );
  INV_X1 U23356 ( .A(n21388), .ZN(n21405) );
  NOR3_X1 U23357 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21390), .A3(
        n21405), .ZN(n21389) );
  AOI211_X1 U23358 ( .C1(n21782), .C2(n21401), .A(n21400), .B(n21389), .ZN(
        n21392) );
  NOR2_X1 U23359 ( .A1(n21598), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21536) );
  OAI211_X1 U23360 ( .C1(n21536), .C2(n21390), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n21753), .ZN(n21391) );
  AOI21_X1 U23361 ( .B1(n21392), .B2(n21391), .A(n21747), .ZN(n21396) );
  OAI22_X1 U23362 ( .A1(n21633), .A2(n21394), .B1(n21393), .B2(n21454), .ZN(
        n21395) );
  NOR2_X1 U23363 ( .A1(n21396), .A2(n21395), .ZN(n21398) );
  OAI211_X1 U23364 ( .C1(n21712), .C2(n21399), .A(n21398), .B(n21397), .ZN(
        P3_U2860) );
  AOI211_X1 U23365 ( .C1(n21742), .C2(n21404), .A(n21400), .B(n21420), .ZN(
        n21402) );
  AOI221_X1 U23366 ( .B1(n21598), .B2(n21402), .C1(n21401), .C2(n21402), .A(
        n21747), .ZN(n21411) );
  INV_X1 U23367 ( .A(n21403), .ZN(n21421) );
  OAI22_X1 U23368 ( .A1(n21421), .A2(n21601), .B1(n21405), .B2(n21404), .ZN(
        n21443) );
  OAI22_X1 U23369 ( .A1(n21633), .A2(n21407), .B1(n21406), .B2(n21454), .ZN(
        n21408) );
  AOI221_X1 U23370 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21411), .C1(
        n21443), .C2(n21411), .A(n21408), .ZN(n21410) );
  OAI211_X1 U23371 ( .C1(n21712), .C2(n21420), .A(n21410), .B(n21409), .ZN(
        P3_U2859) );
  OAI221_X1 U23372 ( .B1(n21730), .B2(n21411), .C1(n21730), .C2(n21721), .A(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21417) );
  NAND2_X1 U23373 ( .A1(n21757), .A2(n21443), .ZN(n21433) );
  NOR2_X1 U23374 ( .A1(n21433), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n21415) );
  OAI22_X1 U23375 ( .A1(n21633), .A2(n21413), .B1(n21412), .B2(n21454), .ZN(
        n21414) );
  AOI21_X1 U23376 ( .B1(n21415), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n21414), .ZN(n21416) );
  OAI211_X1 U23377 ( .C1(n11173), .C2(n21418), .A(n21417), .B(n21416), .ZN(
        P3_U2858) );
  NOR4_X1 U23378 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21420), .A3(
        n21419), .A4(n21433), .ZN(n21428) );
  OAI21_X1 U23379 ( .B1(n21421), .B2(n21432), .A(n21782), .ZN(n21422) );
  INV_X1 U23380 ( .A(n21536), .ZN(n21447) );
  OAI211_X1 U23381 ( .C1(n21707), .C2(n21423), .A(n21422), .B(n21447), .ZN(
        n21424) );
  AOI21_X1 U23382 ( .B1(n21757), .B2(n21424), .A(n21730), .ZN(n21441) );
  OAI22_X1 U23383 ( .A1(n21441), .A2(n21426), .B1(n21633), .B2(n21425), .ZN(
        n21427) );
  NOR2_X1 U23384 ( .A1(n21428), .A2(n21427), .ZN(n21430) );
  NAND2_X1 U23385 ( .A1(n21769), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21429) );
  OAI211_X1 U23386 ( .C1(n21431), .C2(n21454), .A(n21430), .B(n21429), .ZN(
        P3_U2857) );
  NOR3_X1 U23387 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21433), .A3(
        n21432), .ZN(n21437) );
  OAI22_X1 U23388 ( .A1(n21633), .A2(n21435), .B1(n21434), .B2(n21454), .ZN(
        n21436) );
  NOR2_X1 U23389 ( .A1(n21437), .A2(n21436), .ZN(n21439) );
  NAND2_X1 U23390 ( .A1(n21769), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n21438) );
  OAI211_X1 U23391 ( .C1(n21441), .C2(n21440), .A(n21439), .B(n21438), .ZN(
        P3_U2856) );
  INV_X1 U23392 ( .A(n21633), .ZN(n21581) );
  NOR2_X1 U23393 ( .A1(n11173), .A2(n21442), .ZN(n21451) );
  NAND2_X1 U23394 ( .A1(n21444), .A2(n21443), .ZN(n21477) );
  AOI22_X1 U23395 ( .A1(n21782), .A2(n21446), .B1(n21753), .B2(n21445), .ZN(
        n21448) );
  NAND3_X1 U23396 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21448), .A3(
        n21447), .ZN(n21457) );
  AOI22_X1 U23397 ( .A1(n21757), .A2(n21457), .B1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21730), .ZN(n21449) );
  AOI21_X1 U23398 ( .B1(n21456), .B2(n21477), .A(n21449), .ZN(n21450) );
  AOI211_X1 U23399 ( .C1(n21452), .C2(n21581), .A(n21451), .B(n21450), .ZN(
        n21453) );
  OAI21_X1 U23400 ( .B1(n21455), .B2(n21454), .A(n21453), .ZN(P3_U2855) );
  NOR2_X1 U23401 ( .A1(n21456), .A2(n21477), .ZN(n21459) );
  AND2_X1 U23402 ( .A1(n21721), .A2(n21457), .ZN(n21458) );
  MUX2_X1 U23403 ( .A(n21459), .B(n21458), .S(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n21460) );
  AOI21_X1 U23404 ( .B1(n21679), .B2(n21462), .A(n21460), .ZN(n21461) );
  OAI21_X1 U23405 ( .B1(n21463), .B2(n21462), .A(n21461), .ZN(n21464) );
  AOI22_X1 U23406 ( .A1(n21757), .A2(n21464), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21730), .ZN(n21466) );
  OAI211_X1 U23407 ( .C1(n21633), .C2(n21467), .A(n21466), .B(n21465), .ZN(
        P3_U2854) );
  NAND2_X1 U23408 ( .A1(n21700), .A2(n21644), .ZN(n21706) );
  NOR2_X1 U23409 ( .A1(n21468), .A2(n21741), .ZN(n21488) );
  AOI21_X1 U23410 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21488), .A(
        n21598), .ZN(n21473) );
  NAND2_X1 U23411 ( .A1(n21679), .A2(n21469), .ZN(n21471) );
  INV_X1 U23412 ( .A(n21470), .ZN(n21501) );
  NAND2_X1 U23413 ( .A1(n21782), .A2(n21501), .ZN(n21489) );
  OAI211_X1 U23414 ( .C1(n21472), .C2(n21644), .A(n21471), .B(n21489), .ZN(
        n21761) );
  AOI211_X1 U23415 ( .C1(n21475), .C2(n21706), .A(n21473), .B(n21761), .ZN(
        n21744) );
  NOR2_X1 U23416 ( .A1(n21492), .A2(n21601), .ZN(n21474) );
  AOI221_X1 U23417 ( .B1(n21475), .B2(n21742), .C1(n21741), .C2(n21742), .A(
        n21474), .ZN(n21491) );
  OAI211_X1 U23418 ( .C1(n21598), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n21744), .B(n21491), .ZN(n21476) );
  AOI21_X1 U23419 ( .B1(n21757), .B2(n21476), .A(n21730), .ZN(n21485) );
  NOR2_X1 U23420 ( .A1(n21478), .A2(n21477), .ZN(n21522) );
  INV_X1 U23421 ( .A(n21522), .ZN(n21500) );
  AOI22_X1 U23422 ( .A1(n21765), .A2(n21481), .B1(n21763), .B2(n21480), .ZN(
        n21483) );
  OAI211_X1 U23423 ( .C1(n21485), .C2(n21484), .A(n21483), .B(n21482), .ZN(
        P3_U2851) );
  AOI22_X1 U23424 ( .A1(n21679), .A2(n21487), .B1(n21780), .B2(n21486), .ZN(
        n21490) );
  INV_X1 U23425 ( .A(n21488), .ZN(n21752) );
  OAI21_X1 U23426 ( .B1(n21502), .B2(n21752), .A(n21754), .ZN(n21503) );
  NAND4_X1 U23427 ( .A1(n21491), .A2(n21490), .A3(n21489), .A4(n21503), .ZN(
        n21729) );
  OAI21_X1 U23428 ( .B1(n21759), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21731) );
  NOR2_X1 U23429 ( .A1(n21729), .A2(n21731), .ZN(n21498) );
  AOI22_X1 U23430 ( .A1(n21757), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n21492), .B2(n21763), .ZN(n21497) );
  AOI22_X1 U23431 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21730), .B1(
        n21765), .B2(n21493), .ZN(n21496) );
  INV_X1 U23432 ( .A(n21494), .ZN(n21495) );
  OAI211_X1 U23433 ( .C1(n21498), .C2(n21497), .A(n21496), .B(n21495), .ZN(
        P3_U2850) );
  AOI22_X1 U23434 ( .A1(n21769), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n21765), 
        .B2(n21499), .ZN(n21515) );
  NOR2_X1 U23435 ( .A1(n21506), .A2(n21500), .ZN(n21509) );
  OAI21_X1 U23436 ( .B1(n21502), .B2(n21501), .A(n21782), .ZN(n21504) );
  OAI211_X1 U23437 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n21689), .A(
        n21504), .B(n21503), .ZN(n21505) );
  AOI221_X1 U23438 ( .B1(n21506), .B2(n21742), .C1(n21741), .C2(n21742), .A(
        n21505), .ZN(n21507) );
  INV_X1 U23439 ( .A(n21507), .ZN(n21508) );
  MUX2_X1 U23440 ( .A(n21509), .B(n21508), .S(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n21513) );
  OAI22_X1 U23441 ( .A1(n21700), .A2(n21511), .B1(n21644), .B2(n21510), .ZN(
        n21512) );
  OAI21_X1 U23442 ( .B1(n21513), .B2(n21512), .A(n21757), .ZN(n21514) );
  OAI211_X1 U23443 ( .C1(n21712), .C2(n21516), .A(n21515), .B(n21514), .ZN(
        P3_U2848) );
  OAI22_X1 U23444 ( .A1(n21517), .A2(n21700), .B1(n21698), .B2(n21644), .ZN(
        n21719) );
  NOR3_X1 U23445 ( .A1(n21536), .A2(n21741), .A3(n21535), .ZN(n21519) );
  OAI21_X1 U23446 ( .B1(n21782), .B2(n21534), .A(n21574), .ZN(n21518) );
  OAI21_X1 U23447 ( .B1(n21707), .B2(n21519), .A(n21518), .ZN(n21720) );
  AOI221_X1 U23448 ( .B1(n21719), .B2(n21757), .C1(n21720), .C2(n21757), .A(
        n21730), .ZN(n21531) );
  NOR3_X1 U23449 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21520), .A3(
        n21633), .ZN(n21521) );
  AOI21_X1 U23450 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n21769), .A(n21521), 
        .ZN(n21530) );
  NAND2_X1 U23451 ( .A1(n21522), .A2(n21720), .ZN(n21526) );
  NAND2_X1 U23452 ( .A1(n21679), .A2(n21523), .ZN(n21524) );
  OAI22_X1 U23453 ( .A1(n21535), .A2(n21526), .B1(n21525), .B2(n21524), .ZN(
        n21528) );
  AOI22_X1 U23454 ( .A1(n21757), .A2(n21528), .B1(n21765), .B2(n21527), .ZN(
        n21529) );
  OAI211_X1 U23455 ( .C1(n21531), .C2(n21534), .A(n21530), .B(n21529), .ZN(
        P3_U2847) );
  AOI21_X1 U23456 ( .B1(n21732), .B2(n21533), .A(n21532), .ZN(n21541) );
  INV_X1 U23457 ( .A(n21576), .ZN(n21537) );
  NOR4_X1 U23458 ( .A1(n21536), .A2(n21535), .A3(n21534), .A4(n21741), .ZN(
        n21702) );
  NAND2_X1 U23459 ( .A1(n21537), .A2(n21702), .ZN(n21547) );
  OAI21_X1 U23460 ( .B1(n21546), .B2(n21754), .A(n21547), .ZN(n21540) );
  AOI21_X1 U23461 ( .B1(n21538), .B2(n21583), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21539) );
  AOI211_X1 U23462 ( .C1(n21541), .C2(n21540), .A(n21539), .B(n21747), .ZN(
        n21542) );
  AOI211_X1 U23463 ( .C1(n21544), .C2(n21765), .A(n21543), .B(n21542), .ZN(
        n21545) );
  OAI21_X1 U23464 ( .B1(n21546), .B2(n21712), .A(n21545), .ZN(P3_U2840) );
  NAND2_X1 U23465 ( .A1(n21753), .A2(n21547), .ZN(n21659) );
  INV_X1 U23466 ( .A(n21659), .ZN(n21549) );
  AOI21_X1 U23467 ( .B1(n21548), .B2(n21564), .A(n21601), .ZN(n21656) );
  NOR3_X1 U23468 ( .A1(n21549), .A2(n21572), .A3(n21656), .ZN(n21560) );
  NOR3_X1 U23469 ( .A1(n21613), .A2(n21560), .A3(n21565), .ZN(n21552) );
  NOR3_X1 U23470 ( .A1(n21591), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n21550), .ZN(n21551) );
  AOI211_X1 U23471 ( .C1(n21553), .C2(n21679), .A(n21552), .B(n21551), .ZN(
        n21558) );
  AOI22_X1 U23472 ( .A1(n21769), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21730), .ZN(n21557) );
  AOI22_X1 U23473 ( .A1(n21765), .A2(n21555), .B1(n21581), .B2(n21554), .ZN(
        n21556) );
  OAI211_X1 U23474 ( .C1(n21558), .C2(n21747), .A(n21557), .B(n21556), .ZN(
        P3_U2837) );
  NAND2_X1 U23475 ( .A1(n21769), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21570) );
  NOR2_X1 U23476 ( .A1(n21559), .A2(n21633), .ZN(n21568) );
  AOI21_X1 U23477 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21560), .A(
        n21613), .ZN(n21561) );
  AOI211_X1 U23478 ( .C1(n21679), .C2(n21603), .A(n21561), .B(n21562), .ZN(
        n21563) );
  OAI22_X1 U23479 ( .A1(n21563), .A2(n21747), .B1(n21562), .B2(n21712), .ZN(
        n21567) );
  NAND2_X1 U23480 ( .A1(n21564), .A2(n21583), .ZN(n21664) );
  NOR3_X1 U23481 ( .A1(n21565), .A2(n21572), .A3(n21664), .ZN(n21566) );
  OAI22_X1 U23482 ( .A1(n21568), .A2(n21567), .B1(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21566), .ZN(n21569) );
  OAI211_X1 U23483 ( .C1(n21571), .C2(n21750), .A(n21570), .B(n21569), .ZN(
        P3_U2836) );
  NOR2_X1 U23484 ( .A1(n21573), .A2(n21572), .ZN(n21579) );
  OR2_X1 U23485 ( .A1(n21575), .A2(n21574), .ZN(n21704) );
  NOR2_X1 U23486 ( .A1(n21704), .A2(n21576), .ZN(n21577) );
  AOI21_X1 U23487 ( .B1(n21579), .B2(n21577), .A(n21601), .ZN(n21600) );
  AOI211_X1 U23488 ( .C1(n21679), .C2(n21603), .A(n21600), .B(n21596), .ZN(
        n21578) );
  OAI211_X1 U23489 ( .C1(n21707), .C2(n21579), .A(n21578), .B(n21659), .ZN(
        n21582) );
  AOI22_X1 U23490 ( .A1(n21757), .A2(n21582), .B1(n21581), .B2(n21580), .ZN(
        n21584) );
  NAND2_X1 U23491 ( .A1(n21589), .A2(n21583), .ZN(n21638) );
  AOI222_X1 U23492 ( .A1(n21584), .A2(n21596), .B1(n21584), .B2(n21712), .C1(
        n21596), .C2(n21638), .ZN(n21585) );
  AOI211_X1 U23493 ( .C1(n21765), .C2(n21587), .A(n21586), .B(n21585), .ZN(
        n21588) );
  INV_X1 U23494 ( .A(n21588), .ZN(P3_U2835) );
  INV_X1 U23495 ( .A(n21646), .ZN(n21593) );
  INV_X1 U23496 ( .A(n21589), .ZN(n21594) );
  NOR3_X1 U23497 ( .A1(n21591), .A2(n21594), .A3(n21590), .ZN(n21624) );
  AOI21_X1 U23498 ( .B1(n21645), .B2(n21780), .A(n21624), .ZN(n21592) );
  OAI21_X1 U23499 ( .B1(n21700), .B2(n21593), .A(n21592), .ZN(n21618) );
  NOR3_X1 U23500 ( .A1(n21596), .A2(n21595), .A3(n21594), .ZN(n21597) );
  AOI222_X1 U23501 ( .A1(n21598), .A2(n21597), .B1(n21598), .B2(n21759), .C1(
        n21597), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21599) );
  NOR2_X1 U23502 ( .A1(n21600), .A2(n21599), .ZN(n21611) );
  OAI21_X1 U23503 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21601), .A(
        n21611), .ZN(n21648) );
  NOR2_X1 U23504 ( .A1(n21603), .A2(n21602), .ZN(n21605) );
  OAI222_X1 U23505 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21757), 
        .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21618), .C1(n18415), 
        .C2(n21607), .ZN(n21609) );
  OAI211_X1 U23506 ( .C1(n21610), .C2(n21750), .A(n21609), .B(n21608), .ZN(
        P3_U2833) );
  OAI211_X1 U23507 ( .C1(n21613), .C2(n21612), .A(n21611), .B(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21623) );
  OAI22_X1 U23508 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n21614), .B2(n21623), .ZN(
        n21616) );
  OAI22_X1 U23509 ( .A1(n21747), .A2(n21616), .B1(n21712), .B2(n21615), .ZN(
        n21617) );
  OAI21_X1 U23510 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n21618), .A(
        n21617), .ZN(n21619) );
  OAI211_X1 U23511 ( .C1(n21621), .C2(n21750), .A(n21620), .B(n21619), .ZN(
        P3_U2832) );
  AOI21_X1 U23512 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21730), .A(
        n21622), .ZN(n21632) );
  NAND3_X1 U23513 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21721), .A3(
        n21623), .ZN(n21627) );
  NAND3_X1 U23514 ( .A1(n21625), .A2(n21624), .A3(n18421), .ZN(n21626) );
  OAI211_X1 U23515 ( .C1(n21628), .C2(n21700), .A(n21627), .B(n21626), .ZN(
        n21630) );
  AOI22_X1 U23516 ( .A1(n21757), .A2(n21630), .B1(n21765), .B2(n21629), .ZN(
        n21631) );
  OAI211_X1 U23517 ( .C1(n21634), .C2(n21633), .A(n21632), .B(n21631), .ZN(
        P3_U2831) );
  NAND2_X1 U23518 ( .A1(n21636), .A2(n21635), .ZN(n21643) );
  OAI22_X1 U23519 ( .A1(n21639), .A2(n21638), .B1(n21637), .B2(n21643), .ZN(
        n21640) );
  AOI22_X1 U23520 ( .A1(n21757), .A2(n21640), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11173), .ZN(n21655) );
  INV_X1 U23521 ( .A(n21641), .ZN(n21642) );
  AOI21_X1 U23522 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21643), .A(
        n21642), .ZN(n21649) );
  OAI22_X1 U23523 ( .A1(n21646), .A2(n21700), .B1(n21645), .B2(n21644), .ZN(
        n21647) );
  OR3_X1 U23524 ( .A1(n21651), .A2(n21750), .A3(n21650), .ZN(n21653) );
  OAI211_X1 U23525 ( .C1(n21655), .C2(n21654), .A(n21653), .B(n21652), .ZN(
        P3_U2834) );
  INV_X1 U23526 ( .A(n21656), .ZN(n21662) );
  AOI22_X1 U23527 ( .A1(n21679), .A2(n21658), .B1(n21780), .B2(n21657), .ZN(
        n21660) );
  NAND3_X1 U23528 ( .A1(n21660), .A2(n21712), .A3(n21659), .ZN(n21673) );
  INV_X1 U23529 ( .A(n21673), .ZN(n21661) );
  NAND3_X1 U23530 ( .A1(n21662), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n21661), .ZN(n21663) );
  NAND2_X1 U23531 ( .A1(n11173), .A2(n21663), .ZN(n21671) );
  AOI221_X1 U23532 ( .B1(n21730), .B2(n21665), .C1(n21664), .C2(n21665), .A(
        n21671), .ZN(n21666) );
  AOI211_X1 U23533 ( .C1(n21668), .C2(n21765), .A(n21667), .B(n21666), .ZN(
        n21669) );
  INV_X1 U23534 ( .A(n21669), .ZN(P3_U2839) );
  AOI22_X1 U23535 ( .A1(n21769), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n21765), 
        .B2(n21670), .ZN(n21675) );
  INV_X1 U23536 ( .A(n21671), .ZN(n21672) );
  OAI211_X1 U23537 ( .C1(n21721), .C2(n21673), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21672), .ZN(n21674) );
  OAI211_X1 U23538 ( .C1(n21676), .C2(n21695), .A(n21675), .B(n21674), .ZN(
        P3_U2838) );
  AOI22_X1 U23539 ( .A1(n21679), .A2(n21678), .B1(n21780), .B2(n21677), .ZN(
        n21680) );
  NAND2_X1 U23540 ( .A1(n21681), .A2(n21680), .ZN(n21682) );
  OAI21_X1 U23541 ( .B1(n21683), .B2(n21682), .A(n11173), .ZN(n21687) );
  AOI22_X1 U23542 ( .A1(n21769), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n21765), 
        .B2(n21684), .ZN(n21685) );
  OAI221_X1 U23543 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21695), 
        .C1(n21686), .C2(n21687), .A(n21685), .ZN(P3_U2843) );
  NAND2_X1 U23544 ( .A1(n21686), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21688) );
  OAI21_X1 U23545 ( .B1(n21689), .B2(n21688), .A(n21687), .ZN(n21691) );
  AOI22_X1 U23546 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21691), .B1(
        n21765), .B2(n21690), .ZN(n21693) );
  OAI211_X1 U23547 ( .C1(n21695), .C2(n21694), .A(n21693), .B(n21692), .ZN(
        P3_U2842) );
  NAND2_X1 U23548 ( .A1(n21696), .A2(n21763), .ZN(n21728) );
  AOI22_X1 U23549 ( .A1(n21769), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n21765), 
        .B2(n21697), .ZN(n21710) );
  OAI211_X1 U23550 ( .C1(n21701), .C2(n21700), .A(n21699), .B(n21698), .ZN(
        n21705) );
  NAND2_X1 U23551 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21702), .ZN(
        n21703) );
  AOI222_X1 U23552 ( .A1(n21706), .A2(n21705), .B1(n21704), .B2(n21782), .C1(
        n21703), .C2(n21753), .ZN(n21713) );
  OAI211_X1 U23553 ( .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n21707), .A(
        n21757), .B(n21713), .ZN(n21708) );
  NAND3_X1 U23554 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11173), .A3(
        n21708), .ZN(n21709) );
  OAI211_X1 U23555 ( .C1(n21728), .C2(n21711), .A(n21710), .B(n21709), .ZN(
        P3_U2844) );
  OAI21_X1 U23556 ( .B1(n21713), .B2(n21747), .A(n21712), .ZN(n21715) );
  AOI22_X1 U23557 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21715), .B1(
        n21765), .B2(n21714), .ZN(n21717) );
  OAI211_X1 U23558 ( .C1(n21728), .C2(n21718), .A(n21717), .B(n21716), .ZN(
        P3_U2845) );
  AOI211_X1 U23559 ( .C1(n21721), .C2(n21720), .A(n21747), .B(n21719), .ZN(
        n21723) );
  NOR3_X1 U23560 ( .A1(n18279), .A2(n21723), .A3(n21722), .ZN(n21724) );
  AOI21_X1 U23561 ( .B1(n21765), .B2(n21725), .A(n21724), .ZN(n21727) );
  OAI211_X1 U23562 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n21728), .A(
        n21727), .B(n21726), .ZN(P3_U2846) );
  AOI211_X1 U23563 ( .C1(n21732), .C2(n21731), .A(n21730), .B(n21729), .ZN(
        n21734) );
  NOR3_X1 U23564 ( .A1(n21769), .A2(n21734), .A3(n21733), .ZN(n21735) );
  AOI21_X1 U23565 ( .B1(n21736), .B2(n21763), .A(n21735), .ZN(n21738) );
  OAI211_X1 U23566 ( .C1(n21739), .C2(n21750), .A(n21738), .B(n21737), .ZN(
        P3_U2849) );
  NOR2_X1 U23567 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21762), .ZN(
        n21740) );
  AOI22_X1 U23568 ( .A1(n21769), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21763), 
        .B2(n21740), .ZN(n21749) );
  NAND2_X1 U23569 ( .A1(n21742), .A2(n21741), .ZN(n21743) );
  OAI211_X1 U23570 ( .C1(n21745), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n21744), .B(n21743), .ZN(n21746) );
  OAI211_X1 U23571 ( .C1(n21747), .C2(n21746), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n11173), .ZN(n21748) );
  OAI211_X1 U23572 ( .C1(n21751), .C2(n21750), .A(n21749), .B(n21748), .ZN(
        P3_U2852) );
  OAI211_X1 U23573 ( .C1(n21755), .C2(n21754), .A(n21753), .B(n21752), .ZN(
        n21756) );
  OAI211_X1 U23574 ( .C1(n21759), .C2(n21758), .A(n21757), .B(n21756), .ZN(
        n21760) );
  OAI21_X1 U23575 ( .B1(n21761), .B2(n21760), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21768) );
  AOI22_X1 U23576 ( .A1(n21765), .A2(n21764), .B1(n21763), .B2(n21762), .ZN(
        n21766) );
  OAI221_X1 U23577 ( .B1(n21769), .B2(n21768), .C1(n11173), .C2(n21767), .A(
        n21766), .ZN(P3_U2853) );
  NAND2_X1 U23578 ( .A1(n22226), .A2(n21770), .ZN(n21820) );
  INV_X1 U23579 ( .A(n21789), .ZN(n21797) );
  AOI22_X1 U23580 ( .A1(n21789), .A2(n21772), .B1(n21771), .B2(n21797), .ZN(
        n21792) );
  AOI21_X1 U23581 ( .B1(n21774), .B2(n21773), .A(n21792), .ZN(n21806) );
  AOI22_X1 U23582 ( .A1(n21789), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21775), .B2(n21797), .ZN(n21805) );
  AOI221_X1 U23583 ( .B1(n21795), .B2(n21778), .C1(n21777), .C2(n21778), .A(
        n21776), .ZN(n21779) );
  AOI221_X1 U23584 ( .B1(n21782), .B2(n21781), .C1(n21780), .C2(n21781), .A(
        n21779), .ZN(n21834) );
  AOI222_X1 U23585 ( .A1(n21786), .A2(n21785), .B1(n21786), .B2(n21784), .C1(
        n21785), .C2(n21783), .ZN(n21788) );
  OAI21_X1 U23586 ( .B1(n21789), .B2(n21788), .A(n21787), .ZN(n21790) );
  AOI222_X1 U23587 ( .A1(n21792), .A2(n21791), .B1(n21792), .B2(n21790), .C1(
        n21791), .C2(n21790), .ZN(n21793) );
  AOI211_X1 U23588 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n21805), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n21793), .ZN(n21802) );
  NOR2_X1 U23589 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(P3_MORE_REG_SCAN_IN), .ZN(
        n21799) );
  OAI211_X1 U23590 ( .C1(n21796), .C2(n22226), .A(n21795), .B(n21794), .ZN(
        n21831) );
  OAI22_X1 U23591 ( .A1(n21799), .A2(n21831), .B1(n21798), .B2(n21797), .ZN(
        n21800) );
  NOR4_X1 U23592 ( .A1(n21803), .A2(n21802), .A3(n21801), .A4(n21800), .ZN(
        n21804) );
  OAI211_X1 U23593 ( .C1(n21806), .C2(n21805), .A(n21834), .B(n21804), .ZN(
        n21826) );
  AOI211_X1 U23594 ( .C1(n21809), .C2(n21808), .A(n21807), .B(n21826), .ZN(
        n21816) );
  AOI21_X1 U23595 ( .B1(n22226), .B2(n21810), .A(n21816), .ZN(n21829) );
  NAND3_X1 U23596 ( .A1(n21812), .A2(n21829), .A3(n21811), .ZN(n21813) );
  NAND4_X1 U23597 ( .A1(n21815), .A2(n21820), .A3(n21814), .A4(n21813), .ZN(
        P3_U2997) );
  NOR2_X1 U23598 ( .A1(n21816), .A2(n21830), .ZN(n21819) );
  OAI21_X1 U23599 ( .B1(n21819), .B2(n21818), .A(n21817), .ZN(P3_U3282) );
  INV_X1 U23600 ( .A(n21820), .ZN(n21821) );
  AOI211_X1 U23601 ( .C1(n21823), .C2(n21822), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n21821), .ZN(n21824) );
  AOI211_X1 U23602 ( .C1(n21832), .C2(n21826), .A(n21825), .B(n21824), .ZN(
        n21827) );
  OAI221_X1 U23603 ( .B1(n21830), .B2(n21829), .C1(n21830), .C2(n21828), .A(
        n21827), .ZN(P3_U2996) );
  NAND2_X1 U23604 ( .A1(n21832), .A2(n21831), .ZN(n21836) );
  NAND2_X1 U23605 ( .A1(n21836), .A2(P3_MORE_REG_SCAN_IN), .ZN(n21833) );
  OAI21_X1 U23606 ( .B1(n21836), .B2(n21834), .A(n21833), .ZN(P3_U3295) );
  AOI21_X1 U23607 ( .B1(n21836), .B2(P3_FLUSH_REG_SCAN_IN), .A(n21835), .ZN(
        n21837) );
  INV_X1 U23608 ( .A(n21837), .ZN(P3_U2637) );
  INV_X1 U23609 ( .A(n21838), .ZN(n21839) );
  AOI211_X1 U23610 ( .C1(n21842), .C2(n21841), .A(n21840), .B(n21839), .ZN(
        n21848) );
  OAI211_X1 U23611 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21844), .A(n21843), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21845) );
  AOI21_X1 U23612 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21845), .A(n22157), 
        .ZN(n21847) );
  NAND2_X1 U23613 ( .A1(n21848), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21846) );
  OAI21_X1 U23614 ( .B1(n21848), .B2(n21847), .A(n21846), .ZN(P1_U3485) );
  NOR2_X1 U23615 ( .A1(n21850), .A2(n21849), .ZN(n21860) );
  AOI211_X1 U23616 ( .C1(n21852), .C2(n21854), .A(n21860), .B(n21851), .ZN(
        n21868) );
  NOR2_X1 U23617 ( .A1(n21853), .A2(n22001), .ZN(n21859) );
  NOR2_X1 U23618 ( .A1(n21855), .A2(n21854), .ZN(n21857) );
  AOI22_X1 U23619 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21857), .B1(
        n21952), .B2(n21856), .ZN(n21858) );
  NOR2_X1 U23620 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21858), .ZN(
        n21866) );
  AOI211_X1 U23621 ( .C1(n21861), .C2(n21860), .A(n21859), .B(n21866), .ZN(
        n21865) );
  AOI22_X1 U23622 ( .A1(n21863), .A2(n22018), .B1(n22017), .B2(n21862), .ZN(
        n21864) );
  OAI211_X1 U23623 ( .C1(n21868), .C2(n21873), .A(n21865), .B(n21864), .ZN(
        P1_U3018) );
  INV_X1 U23624 ( .A(n21866), .ZN(n21869) );
  AOI21_X1 U23625 ( .B1(n21869), .B2(n21868), .A(n21867), .ZN(n21870) );
  AOI211_X1 U23626 ( .C1(n21872), .C2(n22018), .A(n21871), .B(n21870), .ZN(
        n21875) );
  OR3_X1 U23627 ( .A1(n21873), .A2(n21973), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21874) );
  OAI211_X1 U23628 ( .C1(n22014), .C2(n21876), .A(n21875), .B(n21874), .ZN(
        P1_U3017) );
  NAND2_X1 U23629 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21877), .ZN(
        n21892) );
  NOR2_X1 U23630 ( .A1(n21878), .A2(n21879), .ZN(n21882) );
  NOR2_X1 U23631 ( .A1(n21893), .A2(n21879), .ZN(n21881) );
  OAI21_X1 U23632 ( .B1(n21881), .B2(n21932), .A(n21880), .ZN(n21912) );
  AOI21_X1 U23633 ( .B1(n21952), .B2(n21882), .A(n21912), .ZN(n21891) );
  INV_X1 U23634 ( .A(n21883), .ZN(n21889) );
  INV_X1 U23635 ( .A(n21895), .ZN(n21894) );
  NOR2_X1 U23636 ( .A1(n21884), .A2(n21894), .ZN(n21888) );
  OAI22_X1 U23637 ( .A1(n22014), .A2(n21886), .B1(n21885), .B2(n22001), .ZN(
        n21887) );
  AOI211_X1 U23638 ( .C1(n21889), .C2(n22018), .A(n21888), .B(n21887), .ZN(
        n21890) );
  OAI221_X1 U23639 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21892), .C1(
        n21893), .C2(n21891), .A(n21890), .ZN(P1_U3029) );
  NOR2_X1 U23640 ( .A1(n21893), .A2(n21892), .ZN(n21917) );
  AOI21_X1 U23641 ( .B1(n21952), .B2(n21894), .A(n21917), .ZN(n21929) );
  NOR3_X1 U23642 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21929), .A3(
        n21909), .ZN(n21898) );
  AOI21_X1 U23643 ( .B1(n21952), .B2(n21895), .A(n21912), .ZN(n21910) );
  OR2_X1 U23644 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21929), .ZN(
        n21907) );
  AOI21_X1 U23645 ( .B1(n21910), .B2(n21907), .A(n21896), .ZN(n21897) );
  AOI211_X1 U23646 ( .C1(n21899), .C2(n22018), .A(n21898), .B(n21897), .ZN(
        n21901) );
  NAND2_X1 U23647 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22016), .ZN(n21900) );
  OAI211_X1 U23648 ( .C1(n22014), .C2(n21902), .A(n21901), .B(n21900), .ZN(
        P1_U3027) );
  INV_X1 U23649 ( .A(n21903), .ZN(n21905) );
  AOI222_X1 U23650 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n21906), .B1(n22018), 
        .B2(n21905), .C1(n21904), .C2(n22017), .ZN(n21908) );
  OAI211_X1 U23651 ( .C1(n21910), .C2(n21909), .A(n21908), .B(n21907), .ZN(
        P1_U3028) );
  NAND2_X1 U23652 ( .A1(n21911), .A2(n21915), .ZN(n21928) );
  INV_X1 U23653 ( .A(n21928), .ZN(n21916) );
  INV_X1 U23654 ( .A(n21931), .ZN(n21913) );
  AOI21_X1 U23655 ( .B1(n21952), .B2(n21913), .A(n21912), .ZN(n21914) );
  OAI21_X1 U23656 ( .B1(n21932), .B2(n21915), .A(n21914), .ZN(n21924) );
  AOI21_X1 U23657 ( .B1(n21917), .B2(n21916), .A(n21924), .ZN(n21923) );
  AOI22_X1 U23658 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22016), .B1(n22017), 
        .B2(n22035), .ZN(n21921) );
  NOR2_X1 U23659 ( .A1(n21929), .A2(n21918), .ZN(n21930) );
  AOI22_X1 U23660 ( .A1(n21919), .A2(n22018), .B1(n21930), .B2(n21922), .ZN(
        n21920) );
  OAI211_X1 U23661 ( .C1(n21923), .C2(n21922), .A(n21921), .B(n21920), .ZN(
        P1_U3025) );
  AOI22_X1 U23662 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22016), .B1(n22017), 
        .B2(n22025), .ZN(n21927) );
  AOI22_X1 U23663 ( .A1(n21925), .A2(n22018), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n21924), .ZN(n21926) );
  OAI211_X1 U23664 ( .C1(n21929), .C2(n21928), .A(n21927), .B(n21926), .ZN(
        P1_U3026) );
  NAND2_X1 U23665 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21930), .ZN(
        n21955) );
  OAI211_X1 U23666 ( .C1(n21933), .C2(n21932), .A(n21931), .B(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21935) );
  AOI21_X1 U23667 ( .B1(n21936), .B2(n21935), .A(n21934), .ZN(n21942) );
  AOI222_X1 U23668 ( .A1(n22046), .A2(n22017), .B1(n22016), .B2(
        P1_REIP_REG_7__SCAN_IN), .C1(n22018), .C2(n21937), .ZN(n21938) );
  OAI221_X1 U23669 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21955), .C1(
        n21939), .C2(n21942), .A(n21938), .ZN(P1_U3024) );
  INV_X1 U23670 ( .A(n21940), .ZN(n21945) );
  OAI21_X1 U23671 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n21956), .ZN(n21941) );
  OAI22_X1 U23672 ( .A1(n21943), .A2(n21942), .B1(n21955), .B2(n21941), .ZN(
        n21944) );
  AOI21_X1 U23673 ( .B1(n21945), .B2(n22018), .A(n21944), .ZN(n21947) );
  NAND2_X1 U23674 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22016), .ZN(n21946) );
  OAI211_X1 U23675 ( .C1(n22014), .C2(n21948), .A(n21947), .B(n21946), .ZN(
        P1_U3023) );
  INV_X1 U23676 ( .A(n21949), .ZN(n21950) );
  AOI21_X1 U23677 ( .B1(n21952), .B2(n21951), .A(n21950), .ZN(n21969) );
  AOI22_X1 U23678 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n22016), .B1(n22017), 
        .B2(n21953), .ZN(n21959) );
  INV_X1 U23679 ( .A(n21954), .ZN(n21957) );
  NOR2_X1 U23680 ( .A1(n21956), .A2(n21955), .ZN(n21966) );
  AOI22_X1 U23681 ( .A1(n21957), .A2(n22018), .B1(n21966), .B2(n21960), .ZN(
        n21958) );
  OAI211_X1 U23682 ( .C1(n21969), .C2(n21960), .A(n21959), .B(n21958), .ZN(
        P1_U3022) );
  OAI21_X1 U23683 ( .B1(n22014), .B2(n21962), .A(n21961), .ZN(n21963) );
  AOI21_X1 U23684 ( .B1(n21964), .B2(n22018), .A(n21963), .ZN(n21968) );
  OAI211_X1 U23685 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n21966), .B(n21965), .ZN(
        n21967) );
  OAI211_X1 U23686 ( .C1(n21969), .C2(n15658), .A(n21968), .B(n21967), .ZN(
        P1_U3021) );
  AOI22_X1 U23687 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n22016), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21970), .ZN(n21979) );
  AND3_X1 U23688 ( .A1(n21972), .A2(n21971), .A3(n22018), .ZN(n21977) );
  NOR4_X1 U23689 ( .A1(n21975), .A2(n21974), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n21973), .ZN(n21976) );
  NOR2_X1 U23690 ( .A1(n21977), .A2(n21976), .ZN(n21978) );
  OAI211_X1 U23691 ( .C1(n22014), .C2(n21980), .A(n21979), .B(n21978), .ZN(
        P1_U3013) );
  INV_X1 U23692 ( .A(n21981), .ZN(n21988) );
  INV_X1 U23693 ( .A(n21982), .ZN(n21985) );
  NOR3_X1 U23694 ( .A1(n21985), .A2(n21984), .A3(n21983), .ZN(n21986) );
  AOI211_X1 U23695 ( .C1(n21988), .C2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n21987), .B(n21986), .ZN(n21989) );
  OAI21_X1 U23696 ( .B1(n21990), .B2(n22004), .A(n21989), .ZN(n21991) );
  INV_X1 U23697 ( .A(n21991), .ZN(n21992) );
  OAI21_X1 U23698 ( .B1(n22014), .B2(n21993), .A(n21992), .ZN(P1_U3015) );
  AOI22_X1 U23699 ( .A1(n21994), .A2(n22018), .B1(n22017), .B2(n22101), .ZN(
        n21999) );
  AOI22_X1 U23700 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21997), .B1(
        n21996), .B2(n21995), .ZN(n21998) );
  OAI211_X1 U23701 ( .C1(n22001), .C2(n22000), .A(n21999), .B(n21998), .ZN(
        P1_U3012) );
  NOR3_X1 U23702 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n22003), .A3(
        n22002), .ZN(n22007) );
  NOR2_X1 U23703 ( .A1(n22005), .A2(n22004), .ZN(n22006) );
  AOI211_X1 U23704 ( .C1(n22016), .C2(P1_REIP_REG_22__SCAN_IN), .A(n22007), 
        .B(n22006), .ZN(n22012) );
  INV_X1 U23705 ( .A(n22008), .ZN(n22010) );
  OAI21_X1 U23706 ( .B1(n22010), .B2(n22009), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n22011) );
  OAI211_X1 U23707 ( .C1(n22014), .C2(n22013), .A(n22012), .B(n22011), .ZN(
        P1_U3009) );
  AOI22_X1 U23708 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n22016), .B1(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n22015), .ZN(n22021) );
  AOI22_X1 U23709 ( .A1(n22019), .A2(n22018), .B1(n22017), .B2(n22135), .ZN(
        n22020) );
  OAI211_X1 U23710 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n22022), .A(
        n22021), .B(n22020), .ZN(P1_U3008) );
  NAND2_X1 U23711 ( .A1(n22024), .A2(n22023), .ZN(n22027) );
  AOI22_X1 U23712 ( .A1(n22136), .A2(n22025), .B1(n22118), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n22026) );
  OAI21_X1 U23713 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n22027), .A(n22026), .ZN(
        n22028) );
  AOI211_X1 U23714 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n22100), .B(n22028), .ZN(n22033) );
  AOI22_X1 U23715 ( .A1(n22031), .A2(n22030), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n22029), .ZN(n22032) );
  OAI211_X1 U23716 ( .C1(n22034), .C2(n22128), .A(n22033), .B(n22032), .ZN(
        P1_U2835) );
  AOI22_X1 U23717 ( .A1(n22136), .A2(n22035), .B1(n22118), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n22037) );
  OR3_X1 U23718 ( .A1(n22073), .A2(P1_REIP_REG_6__SCAN_IN), .A3(n22040), .ZN(
        n22036) );
  NAND2_X1 U23719 ( .A1(n22037), .A2(n22036), .ZN(n22038) );
  AOI211_X1 U23720 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n22100), .B(n22038), .ZN(n22044) );
  OR3_X1 U23721 ( .A1(n22073), .A2(n22040), .A3(n22039), .ZN(n22048) );
  NAND2_X1 U23722 ( .A1(n22096), .A2(n22048), .ZN(n22051) );
  INV_X1 U23723 ( .A(n22051), .ZN(n22041) );
  AOI22_X1 U23724 ( .A1(n22042), .A2(n22137), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n22041), .ZN(n22043) );
  OAI211_X1 U23725 ( .C1(n22045), .C2(n22128), .A(n22044), .B(n22043), .ZN(
        P1_U2834) );
  AOI22_X1 U23726 ( .A1(n22136), .A2(n22046), .B1(n22118), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n22047) );
  OAI21_X1 U23727 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n22048), .A(n22047), .ZN(
        n22049) );
  AOI211_X1 U23728 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n22100), .B(n22049), .ZN(n22055) );
  NOR2_X1 U23729 ( .A1(n22051), .A2(n22050), .ZN(n22052) );
  AOI21_X1 U23730 ( .B1(n22053), .B2(n22137), .A(n22052), .ZN(n22054) );
  OAI211_X1 U23731 ( .C1(n22056), .C2(n22128), .A(n22055), .B(n22054), .ZN(
        P1_U2833) );
  INV_X1 U23732 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n22060) );
  INV_X1 U23733 ( .A(n22057), .ZN(n22058) );
  OAI22_X1 U23734 ( .A1(n22131), .A2(n22060), .B1(n22059), .B2(n22058), .ZN(
        n22061) );
  AOI211_X1 U23735 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n22100), .B(n22061), .ZN(n22068) );
  OAI21_X1 U23736 ( .B1(n22064), .B2(n22063), .A(n22062), .ZN(n22065) );
  AOI22_X1 U23737 ( .A1(n22137), .A2(n22066), .B1(n22076), .B2(n22065), .ZN(
        n22067) );
  OAI211_X1 U23738 ( .C1(n22069), .C2(n22128), .A(n22068), .B(n22067), .ZN(
        P1_U2829) );
  INV_X1 U23739 ( .A(n22070), .ZN(n22075) );
  INV_X1 U23740 ( .A(n22071), .ZN(n22072) );
  NOR3_X1 U23741 ( .A1(n22073), .A2(P1_REIP_REG_12__SCAN_IN), .A3(n22072), 
        .ZN(n22074) );
  AOI21_X1 U23742 ( .B1(n22075), .B2(n22136), .A(n22074), .ZN(n22082) );
  AOI22_X1 U23743 ( .A1(n22134), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n22076), .ZN(n22077) );
  OAI21_X1 U23744 ( .B1(n22131), .B2(n22078), .A(n22077), .ZN(n22079) );
  AOI211_X1 U23745 ( .C1(n22110), .C2(n22080), .A(n22100), .B(n22079), .ZN(
        n22081) );
  OAI211_X1 U23746 ( .C1(n22114), .C2(n22083), .A(n22082), .B(n22081), .ZN(
        P1_U2828) );
  AOI22_X1 U23747 ( .A1(n22085), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n22136), 
        .B2(n22084), .ZN(n22093) );
  INV_X1 U23748 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n22086) );
  OAI22_X1 U23749 ( .A1(n22087), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n22131), 
        .B2(n22086), .ZN(n22088) );
  AOI211_X1 U23750 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n22100), .B(n22088), .ZN(n22092) );
  AOI22_X1 U23751 ( .A1(n22090), .A2(n22137), .B1(n22110), .B2(n22089), .ZN(
        n22091) );
  NAND3_X1 U23752 ( .A1(n22093), .A2(n22092), .A3(n22091), .ZN(P1_U2825) );
  INV_X1 U23753 ( .A(n22094), .ZN(n22095) );
  AOI21_X1 U23754 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n22096), .A(n22095), 
        .ZN(n22105) );
  OAI22_X1 U23755 ( .A1(n22131), .A2(n22098), .B1(n22097), .B2(n22128), .ZN(
        n22099) );
  AOI211_X1 U23756 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n22100), .B(n22099), .ZN(n22104) );
  AOI22_X1 U23757 ( .A1(n22102), .A2(n22137), .B1(n22136), .B2(n22101), .ZN(
        n22103) );
  OAI211_X1 U23758 ( .C1(n22106), .C2(n22105), .A(n22104), .B(n22103), .ZN(
        P1_U2821) );
  INV_X1 U23759 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n22112) );
  INV_X1 U23760 ( .A(n22107), .ZN(n22108) );
  AOI22_X1 U23761 ( .A1(n22110), .A2(n22109), .B1(n22123), .B2(n22108), .ZN(
        n22111) );
  OAI21_X1 U23762 ( .B1(n22113), .B2(n22112), .A(n22111), .ZN(n22117) );
  NOR2_X1 U23763 ( .A1(n22115), .A2(n22114), .ZN(n22116) );
  AOI211_X1 U23764 ( .C1(n22118), .C2(P1_EBX_REG_21__SCAN_IN), .A(n22117), .B(
        n22116), .ZN(n22121) );
  NAND2_X1 U23765 ( .A1(n22136), .A2(n22119), .ZN(n22120) );
  OAI211_X1 U23766 ( .C1(n22123), .C2(n22122), .A(n22121), .B(n22120), .ZN(
        P1_U2819) );
  AOI211_X1 U23767 ( .C1(n22127), .C2(n22126), .A(n22125), .B(n22124), .ZN(
        n22133) );
  OAI22_X1 U23768 ( .A1(n22131), .A2(n22130), .B1(n22129), .B2(n22128), .ZN(
        n22132) );
  AOI211_X1 U23769 ( .C1(n22134), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n22133), .B(n22132), .ZN(n22140) );
  AOI22_X1 U23770 ( .A1(n22138), .A2(n22137), .B1(n22136), .B2(n22135), .ZN(
        n22139) );
  NAND2_X1 U23771 ( .A1(n22140), .A2(n22139), .ZN(P1_U2817) );
  OAI21_X1 U23772 ( .B1(n22143), .B2(n22142), .A(n22141), .ZN(P1_U2806) );
  INV_X1 U23773 ( .A(n22144), .ZN(n22147) );
  NAND4_X1 U23774 ( .A1(n22147), .A2(n22146), .A3(n22145), .A4(n22149), .ZN(
        n22148) );
  OAI21_X1 U23775 ( .B1(n22149), .B2(n12584), .A(n22148), .ZN(P1_U3468) );
  OAI211_X1 U23776 ( .C1(n22154), .C2(n12293), .A(n22151), .B(n22150), .ZN(
        P1_U3163) );
  OAI22_X1 U23777 ( .A1(n22154), .A2(n22280), .B1(n22153), .B2(n22152), .ZN(
        P1_U3466) );
  AOI21_X1 U23778 ( .B1(n22157), .B2(n22156), .A(n22155), .ZN(n22158) );
  OAI22_X1 U23779 ( .A1(n22160), .A2(n22159), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22158), .ZN(n22161) );
  OAI21_X1 U23780 ( .B1(n22163), .B2(n22162), .A(n22161), .ZN(P1_U3161) );
  INV_X1 U23781 ( .A(n22164), .ZN(n22165) );
  OAI21_X1 U23782 ( .B1(n22167), .B2(n22256), .A(n22165), .ZN(P1_U2805) );
  INV_X1 U23783 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22166) );
  OAI21_X1 U23784 ( .B1(n22167), .B2(n22166), .A(n22165), .ZN(P1_U3465) );
  INV_X1 U23785 ( .A(n22168), .ZN(n22170) );
  OAI21_X1 U23786 ( .B1(n22172), .B2(n22169), .A(n22170), .ZN(P2_U2818) );
  OAI21_X1 U23787 ( .B1(n22172), .B2(n22171), .A(n22170), .ZN(P2_U3592) );
  AOI21_X1 U23788 ( .B1(n17479), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n22174), 
        .ZN(n22173) );
  INV_X1 U23789 ( .A(n22173), .ZN(P3_U2636) );
  AOI21_X1 U23790 ( .B1(n17479), .B2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n22174), 
        .ZN(n22175) );
  INV_X1 U23791 ( .A(n22175), .ZN(P3_U3281) );
  INV_X1 U23792 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22217) );
  AOI21_X1 U23793 ( .B1(HOLD), .B2(n22176), .A(n22217), .ZN(n22178) );
  AOI21_X1 U23794 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n22226), .A(n22216), 
        .ZN(n22233) );
  INV_X1 U23795 ( .A(NA), .ZN(n22198) );
  OAI21_X1 U23796 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n22198), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n22232) );
  INV_X1 U23797 ( .A(n22232), .ZN(n22177) );
  OAI22_X1 U23798 ( .A1(n22179), .A2(n22178), .B1(n22233), .B2(n22177), .ZN(
        P3_U3029) );
  INV_X1 U23799 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22183) );
  NAND2_X1 U23800 ( .A1(n22181), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22191) );
  INV_X1 U23801 ( .A(HOLD), .ZN(n22215) );
  AOI21_X1 U23802 ( .B1(HOLD), .B2(P1_STATE_REG_2__SCAN_IN), .A(n22183), .ZN(
        n22192) );
  AOI21_X1 U23803 ( .B1(n22181), .B2(n22198), .A(n22180), .ZN(n22182) );
  OAI33_X1 U23804 ( .A1(n22183), .A2(NA), .A3(n22191), .B1(n22215), .B2(n22192), .B3(n22182), .ZN(n22186) );
  AOI22_X1 U23805 ( .A1(NA), .A2(n22184), .B1(P1_STATE_REG_0__SCAN_IN), .B2(
        n22191), .ZN(n22185) );
  AOI22_X1 U23806 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22186), .B1(
        P1_STATE_REG_2__SCAN_IN), .B2(n22185), .ZN(n22187) );
  INV_X1 U23807 ( .A(n22187), .ZN(P1_U3196) );
  AOI22_X1 U23808 ( .A1(HOLD), .A2(n22188), .B1(P1_STATE_REG_0__SCAN_IN), .B2(
        n22192), .ZN(n22190) );
  NAND3_X1 U23809 ( .A1(n22190), .A2(n22189), .A3(n22191), .ZN(P1_U3195) );
  AND2_X1 U23810 ( .A1(n22191), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22195) );
  OAI21_X1 U23811 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n22198), .A(n22192), 
        .ZN(n22193) );
  AOI21_X1 U23812 ( .B1(HOLD), .B2(P1_STATE_REG_1__SCAN_IN), .A(n22193), .ZN(
        n22194) );
  OAI22_X1 U23813 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22195), .B1(n22596), 
        .B2(n22194), .ZN(P1_U3194) );
  NAND2_X1 U23814 ( .A1(n22196), .A2(HOLD), .ZN(n22202) );
  NAND2_X1 U23815 ( .A1(n22197), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22209) );
  NAND2_X1 U23816 ( .A1(n22209), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n22208) );
  OAI21_X1 U23817 ( .B1(n22199), .B2(n22198), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n22213) );
  AOI22_X1 U23818 ( .A1(n22200), .A2(n17744), .B1(n22208), .B2(n22213), .ZN(
        n22201) );
  OAI21_X1 U23819 ( .B1(n22203), .B2(n22202), .A(n22201), .ZN(P2_U3209) );
  OAI211_X1 U23820 ( .C1(n22205), .C2(n22215), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22206) );
  NAND4_X1 U23821 ( .A1(n22207), .A2(n11687), .A3(n22209), .A4(n22206), .ZN(
        P2_U3210) );
  INV_X1 U23822 ( .A(n22208), .ZN(n22212) );
  OAI22_X1 U23823 ( .A1(NA), .A2(n22209), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22210) );
  OAI211_X1 U23824 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n22210), .ZN(n22211) );
  OAI221_X1 U23825 ( .B1(n22213), .B2(n22212), .C1(n22213), .C2(n22215), .A(
        n22211), .ZN(P2_U3211) );
  NOR2_X1 U23826 ( .A1(n22215), .A2(n22214), .ZN(n22229) );
  NOR3_X1 U23827 ( .A1(n22229), .A2(n22217), .A3(n22216), .ZN(n22218) );
  NOR2_X1 U23828 ( .A1(n22219), .A2(n22218), .ZN(n22222) );
  NOR2_X1 U23829 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22231)
         );
  AOI221_X1 U23830 ( .B1(n22229), .B2(n22224), .C1(n22231), .C2(n22224), .A(
        n22219), .ZN(n22220) );
  INV_X1 U23831 ( .A(n22220), .ZN(n22221) );
  MUX2_X1 U23832 ( .A(n22222), .B(n22221), .S(P3_STATE_REG_1__SCAN_IN), .Z(
        n22223) );
  OAI221_X1 U23833 ( .B1(n22225), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n22225), 
        .C2(n22224), .A(n22223), .ZN(P3_U3030) );
  NAND2_X1 U23834 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n22226), .ZN(n22227) );
  OAI22_X1 U23835 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n22227), .ZN(n22228) );
  OAI21_X1 U23836 ( .B1(n22229), .B2(n22228), .A(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n22230) );
  OAI22_X1 U23837 ( .A1(n22233), .A2(n22232), .B1(n22231), .B2(n22230), .ZN(
        P3_U3031) );
  NOR2_X1 U23838 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22234), .ZN(
        n22478) );
  AOI22_X1 U23839 ( .A1(n22587), .A2(n22299), .B1(n22478), .B2(n22292), .ZN(
        n22247) );
  NAND3_X1 U23840 ( .A1(n22491), .A2(n22253), .A3(n22235), .ZN(n22238) );
  INV_X1 U23841 ( .A(n22236), .ZN(n22237) );
  NAND2_X1 U23842 ( .A1(n22238), .A2(n22237), .ZN(n22243) );
  OR2_X1 U23843 ( .A1(n22239), .A2(n22286), .ZN(n22244) );
  NAND2_X1 U23844 ( .A1(n22241), .A2(n22240), .ZN(n22255) );
  AOI22_X1 U23845 ( .A1(n22243), .A2(n22244), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n22255), .ZN(n22242) );
  OAI211_X1 U23846 ( .C1(n22478), .C2(n22280), .A(n22278), .B(n22242), .ZN(
        n22482) );
  INV_X1 U23847 ( .A(n22243), .ZN(n22245) );
  AOI22_X1 U23848 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22482), .B1(
        n22291), .B2(n22481), .ZN(n22246) );
  OAI211_X1 U23849 ( .C1(n22302), .C2(n22491), .A(n22247), .B(n22246), .ZN(
        P1_U3033) );
  INV_X1 U23850 ( .A(n22248), .ZN(n22499) );
  OAI22_X1 U23851 ( .A1(n22500), .A2(n22267), .B1(n22266), .B2(n22499), .ZN(
        n22249) );
  INV_X1 U23852 ( .A(n22249), .ZN(n22251) );
  AOI22_X1 U23853 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22503), .B1(
        n22291), .B2(n22502), .ZN(n22250) );
  OAI211_X1 U23854 ( .C1(n22302), .C2(n22506), .A(n22251), .B(n22250), .ZN(
        P1_U3057) );
  NOR2_X1 U23855 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22252), .ZN(
        n22508) );
  NAND3_X1 U23856 ( .A1(n22258), .A2(n22253), .A3(n15410), .ZN(n22254) );
  OAI21_X1 U23857 ( .B1(n22255), .B2(n22289), .A(n22254), .ZN(n22507) );
  AOI22_X1 U23858 ( .A1(n22292), .A2(n22508), .B1(n22291), .B2(n22507), .ZN(
        n22262) );
  AOI21_X1 U23859 ( .B1(n22506), .B2(n22513), .A(n22256), .ZN(n22257) );
  AOI21_X1 U23860 ( .B1(n22258), .B2(n15410), .A(n22257), .ZN(n22259) );
  NOR2_X1 U23861 ( .A1(n22259), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22260) );
  AOI22_X1 U23862 ( .A1(n22510), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n22509), .B2(n22299), .ZN(n22261) );
  OAI211_X1 U23863 ( .C1(n22302), .C2(n22513), .A(n22262), .B(n22261), .ZN(
        P1_U3065) );
  INV_X1 U23864 ( .A(n22263), .ZN(n22515) );
  AOI22_X1 U23865 ( .A1(n22515), .A2(n22291), .B1(n22292), .B2(n22514), .ZN(
        n22265) );
  INV_X1 U23866 ( .A(n22513), .ZN(n22516) );
  AOI22_X1 U23867 ( .A1(n22517), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n22516), .B2(n22299), .ZN(n22264) );
  OAI211_X1 U23868 ( .C1(n22302), .C2(n22521), .A(n22265), .B(n22264), .ZN(
        P1_U3073) );
  OAI22_X1 U23869 ( .A1(n22521), .A2(n22267), .B1(n22520), .B2(n22266), .ZN(
        n22268) );
  INV_X1 U23870 ( .A(n22268), .ZN(n22270) );
  AOI22_X1 U23871 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22524), .B1(
        n22291), .B2(n22523), .ZN(n22269) );
  OAI211_X1 U23872 ( .C1(n22302), .C2(n22527), .A(n22270), .B(n22269), .ZN(
        P1_U3081) );
  NOR2_X1 U23873 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22271), .ZN(
        n22535) );
  AOI21_X1 U23874 ( .B1(n22272), .B2(n15410), .A(n22535), .ZN(n22276) );
  OAI22_X1 U23875 ( .A1(n22276), .A2(n22290), .B1(n22274), .B2(n22273), .ZN(
        n22536) );
  AOI22_X1 U23876 ( .A1(n22536), .A2(n22291), .B1(n22292), .B2(n22535), .ZN(
        n22282) );
  INV_X1 U23877 ( .A(n22546), .ZN(n22275) );
  OAI21_X1 U23878 ( .B1(n22275), .B2(n22537), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22277) );
  NAND2_X1 U23879 ( .A1(n22277), .A2(n22276), .ZN(n22279) );
  AOI22_X1 U23880 ( .A1(n22538), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n22537), .B2(n22299), .ZN(n22281) );
  OAI211_X1 U23881 ( .C1(n22302), .C2(n22546), .A(n22282), .B(n22281), .ZN(
        P1_U3097) );
  AOI22_X1 U23882 ( .A1(n22548), .A2(n22299), .B1(n22547), .B2(n22292), .ZN(
        n22284) );
  AOI22_X1 U23883 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22550), .B1(
        n22291), .B2(n22549), .ZN(n22283) );
  OAI211_X1 U23884 ( .C1(n22302), .C2(n22553), .A(n22284), .B(n22283), .ZN(
        P1_U3113) );
  NOR2_X1 U23885 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22285), .ZN(
        n22575) );
  NAND2_X1 U23886 ( .A1(n22287), .A2(n22286), .ZN(n22294) );
  OAI22_X1 U23887 ( .A1(n22294), .A2(n22290), .B1(n22289), .B2(n22288), .ZN(
        n22574) );
  AOI22_X1 U23888 ( .A1(n22292), .A2(n22575), .B1(n22291), .B2(n22574), .ZN(
        n22301) );
  INV_X1 U23889 ( .A(n22591), .ZN(n22293) );
  OAI21_X1 U23890 ( .B1(n22577), .B2(n22293), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22295) );
  AOI21_X1 U23891 ( .B1(n22295), .B2(n22294), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n22298) );
  AOI22_X1 U23892 ( .A1(n22578), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n22577), .B2(n22299), .ZN(n22300) );
  OAI211_X1 U23893 ( .C1(n22302), .C2(n22591), .A(n22301), .B(n22300), .ZN(
        P1_U3145) );
  AOI22_X1 U23894 ( .A1(n22587), .A2(n22327), .B1(n22478), .B2(n22326), .ZN(
        n22304) );
  AOI22_X1 U23895 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22482), .B1(
        n22325), .B2(n22481), .ZN(n22303) );
  OAI211_X1 U23896 ( .C1(n22330), .C2(n22491), .A(n22304), .B(n22303), .ZN(
        P1_U3034) );
  INV_X1 U23897 ( .A(n22305), .ZN(n22486) );
  AOI22_X1 U23898 ( .A1(n22486), .A2(n22325), .B1(n22326), .B2(n22485), .ZN(
        n22307) );
  INV_X1 U23899 ( .A(n22491), .ZN(n22435) );
  AOI22_X1 U23900 ( .A1(n22488), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n22435), .B2(n22327), .ZN(n22306) );
  OAI211_X1 U23901 ( .C1(n22330), .C2(n22493), .A(n22307), .B(n22306), .ZN(
        P1_U3042) );
  OAI22_X1 U23902 ( .A1(n22500), .A2(n22309), .B1(n22308), .B2(n22499), .ZN(
        n22310) );
  INV_X1 U23903 ( .A(n22310), .ZN(n22312) );
  AOI22_X1 U23904 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22503), .B1(
        n22325), .B2(n22502), .ZN(n22311) );
  OAI211_X1 U23905 ( .C1(n22330), .C2(n22506), .A(n22312), .B(n22311), .ZN(
        P1_U3058) );
  AOI22_X1 U23906 ( .A1(n22326), .A2(n22508), .B1(n22325), .B2(n22507), .ZN(
        n22314) );
  AOI22_X1 U23907 ( .A1(n22510), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n22509), .B2(n22327), .ZN(n22313) );
  OAI211_X1 U23908 ( .C1(n22330), .C2(n22513), .A(n22314), .B(n22313), .ZN(
        P1_U3066) );
  INV_X1 U23909 ( .A(n22315), .ZN(n22529) );
  AOI22_X1 U23910 ( .A1(n22529), .A2(n22325), .B1(n22528), .B2(n22326), .ZN(
        n22317) );
  AOI22_X1 U23911 ( .A1(n22531), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n22530), .B2(n22327), .ZN(n22316) );
  OAI211_X1 U23912 ( .C1(n22330), .C2(n22534), .A(n22317), .B(n22316), .ZN(
        P1_U3090) );
  AOI22_X1 U23913 ( .A1(n22536), .A2(n22325), .B1(n22326), .B2(n22535), .ZN(
        n22319) );
  AOI22_X1 U23914 ( .A1(n22538), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n22537), .B2(n22327), .ZN(n22318) );
  OAI211_X1 U23915 ( .C1(n22330), .C2(n22546), .A(n22319), .B(n22318), .ZN(
        P1_U3098) );
  AOI22_X1 U23916 ( .A1(n22548), .A2(n22327), .B1(n22547), .B2(n22326), .ZN(
        n22321) );
  AOI22_X1 U23917 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22550), .B1(
        n22325), .B2(n22549), .ZN(n22320) );
  OAI211_X1 U23918 ( .C1(n22330), .C2(n22553), .A(n22321), .B(n22320), .ZN(
        P1_U3114) );
  INV_X1 U23919 ( .A(n22322), .ZN(n22555) );
  AOI22_X1 U23920 ( .A1(n22555), .A2(n22325), .B1(n22326), .B2(n22554), .ZN(
        n22324) );
  AOI22_X1 U23921 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n22556), .B2(n22327), .ZN(n22323) );
  OAI211_X1 U23922 ( .C1(n22330), .C2(n22567), .A(n22324), .B(n22323), .ZN(
        P1_U3122) );
  AOI22_X1 U23923 ( .A1(n22326), .A2(n22575), .B1(n22325), .B2(n22574), .ZN(
        n22329) );
  AOI22_X1 U23924 ( .A1(n22578), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n22577), .B2(n22327), .ZN(n22328) );
  OAI211_X1 U23925 ( .C1(n22330), .C2(n22591), .A(n22329), .B(n22328), .ZN(
        P1_U3146) );
  AOI22_X1 U23926 ( .A1(n22587), .A2(n22356), .B1(n22478), .B2(n22355), .ZN(
        n22332) );
  AOI22_X1 U23927 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22482), .B1(
        n22354), .B2(n22481), .ZN(n22331) );
  OAI211_X1 U23928 ( .C1(n22359), .C2(n22491), .A(n22332), .B(n22331), .ZN(
        P1_U3035) );
  OAI22_X1 U23929 ( .A1(n22493), .A2(n22342), .B1(n22492), .B2(n22341), .ZN(
        n22333) );
  INV_X1 U23930 ( .A(n22333), .ZN(n22335) );
  AOI22_X1 U23931 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22496), .B1(
        n22354), .B2(n22495), .ZN(n22334) );
  OAI211_X1 U23932 ( .C1(n22359), .C2(n22500), .A(n22335), .B(n22334), .ZN(
        P1_U3051) );
  OAI22_X1 U23933 ( .A1(n22500), .A2(n22342), .B1(n22499), .B2(n22341), .ZN(
        n22336) );
  INV_X1 U23934 ( .A(n22336), .ZN(n22338) );
  AOI22_X1 U23935 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22503), .B1(
        n22354), .B2(n22502), .ZN(n22337) );
  OAI211_X1 U23936 ( .C1(n22359), .C2(n22506), .A(n22338), .B(n22337), .ZN(
        P1_U3059) );
  AOI22_X1 U23937 ( .A1(n22355), .A2(n22508), .B1(n22354), .B2(n22507), .ZN(
        n22340) );
  AOI22_X1 U23938 ( .A1(n22510), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n22509), .B2(n22356), .ZN(n22339) );
  OAI211_X1 U23939 ( .C1(n22359), .C2(n22513), .A(n22340), .B(n22339), .ZN(
        P1_U3067) );
  OAI22_X1 U23940 ( .A1(n22521), .A2(n22342), .B1(n22520), .B2(n22341), .ZN(
        n22343) );
  INV_X1 U23941 ( .A(n22343), .ZN(n22345) );
  AOI22_X1 U23942 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22524), .B1(
        n22354), .B2(n22523), .ZN(n22344) );
  OAI211_X1 U23943 ( .C1(n22359), .C2(n22527), .A(n22345), .B(n22344), .ZN(
        P1_U3083) );
  AOI22_X1 U23944 ( .A1(n22529), .A2(n22354), .B1(n22528), .B2(n22355), .ZN(
        n22347) );
  AOI22_X1 U23945 ( .A1(n22531), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n22530), .B2(n22356), .ZN(n22346) );
  OAI211_X1 U23946 ( .C1(n22359), .C2(n22534), .A(n22347), .B(n22346), .ZN(
        P1_U3091) );
  AOI22_X1 U23947 ( .A1(n22536), .A2(n22354), .B1(n22355), .B2(n22535), .ZN(
        n22349) );
  AOI22_X1 U23948 ( .A1(n22538), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22537), .B2(n22356), .ZN(n22348) );
  OAI211_X1 U23949 ( .C1(n22359), .C2(n22546), .A(n22349), .B(n22348), .ZN(
        P1_U3099) );
  AOI22_X1 U23950 ( .A1(n22548), .A2(n22356), .B1(n22355), .B2(n22547), .ZN(
        n22351) );
  AOI22_X1 U23951 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22550), .B1(
        n22354), .B2(n22549), .ZN(n22350) );
  OAI211_X1 U23952 ( .C1(n22359), .C2(n22553), .A(n22351), .B(n22350), .ZN(
        P1_U3115) );
  AOI22_X1 U23953 ( .A1(n22555), .A2(n22354), .B1(n22355), .B2(n22554), .ZN(
        n22353) );
  AOI22_X1 U23954 ( .A1(n22557), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n22556), .B2(n22356), .ZN(n22352) );
  OAI211_X1 U23955 ( .C1(n22359), .C2(n22567), .A(n22353), .B(n22352), .ZN(
        P1_U3123) );
  AOI22_X1 U23956 ( .A1(n22355), .A2(n22575), .B1(n22354), .B2(n22574), .ZN(
        n22358) );
  AOI22_X1 U23957 ( .A1(n22578), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n22577), .B2(n22356), .ZN(n22357) );
  OAI211_X1 U23958 ( .C1(n22359), .C2(n22591), .A(n22358), .B(n22357), .ZN(
        P1_U3147) );
  AOI22_X1 U23959 ( .A1(n22587), .A2(n22379), .B1(n22478), .B2(n22378), .ZN(
        n22361) );
  AOI22_X1 U23960 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22482), .B1(
        n22377), .B2(n22481), .ZN(n22360) );
  OAI211_X1 U23961 ( .C1(n22382), .C2(n22491), .A(n22361), .B(n22360), .ZN(
        P1_U3036) );
  OAI22_X1 U23962 ( .A1(n22493), .A2(n22371), .B1(n22492), .B2(n22370), .ZN(
        n22362) );
  INV_X1 U23963 ( .A(n22362), .ZN(n22364) );
  AOI22_X1 U23964 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22496), .B1(
        n22377), .B2(n22495), .ZN(n22363) );
  OAI211_X1 U23965 ( .C1(n22382), .C2(n22500), .A(n22364), .B(n22363), .ZN(
        P1_U3052) );
  OAI22_X1 U23966 ( .A1(n22500), .A2(n22371), .B1(n22499), .B2(n22370), .ZN(
        n22365) );
  INV_X1 U23967 ( .A(n22365), .ZN(n22367) );
  AOI22_X1 U23968 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22503), .B1(
        n22377), .B2(n22502), .ZN(n22366) );
  OAI211_X1 U23969 ( .C1(n22382), .C2(n22506), .A(n22367), .B(n22366), .ZN(
        P1_U3060) );
  AOI22_X1 U23970 ( .A1(n22378), .A2(n22508), .B1(n22377), .B2(n22507), .ZN(
        n22369) );
  AOI22_X1 U23971 ( .A1(n22510), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n22509), .B2(n22379), .ZN(n22368) );
  OAI211_X1 U23972 ( .C1(n22382), .C2(n22513), .A(n22369), .B(n22368), .ZN(
        P1_U3068) );
  OAI22_X1 U23973 ( .A1(n22521), .A2(n22371), .B1(n22520), .B2(n22370), .ZN(
        n22372) );
  INV_X1 U23974 ( .A(n22372), .ZN(n22374) );
  AOI22_X1 U23975 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22524), .B1(
        n22377), .B2(n22523), .ZN(n22373) );
  OAI211_X1 U23976 ( .C1(n22382), .C2(n22527), .A(n22374), .B(n22373), .ZN(
        P1_U3084) );
  AOI22_X1 U23977 ( .A1(n22536), .A2(n22377), .B1(n22378), .B2(n22535), .ZN(
        n22376) );
  AOI22_X1 U23978 ( .A1(n22538), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22537), .B2(n22379), .ZN(n22375) );
  OAI211_X1 U23979 ( .C1(n22382), .C2(n22546), .A(n22376), .B(n22375), .ZN(
        P1_U3100) );
  AOI22_X1 U23980 ( .A1(n22378), .A2(n22575), .B1(n22377), .B2(n22574), .ZN(
        n22381) );
  AOI22_X1 U23981 ( .A1(n22578), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n22577), .B2(n22379), .ZN(n22380) );
  OAI211_X1 U23982 ( .C1(n22382), .C2(n22591), .A(n22381), .B(n22380), .ZN(
        P1_U3148) );
  AOI22_X1 U23983 ( .A1(DATAI_20_), .A2(n11152), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n22474), .ZN(n22424) );
  INV_X1 U23984 ( .A(n22432), .ZN(n22421) );
  NOR2_X2 U23985 ( .A1(n22477), .A2(n11838), .ZN(n22428) );
  AOI22_X1 U23986 ( .A1(n22587), .A2(n22421), .B1(n22428), .B2(n22478), .ZN(
        n22385) );
  NOR2_X2 U23987 ( .A1(n22383), .A2(n22479), .ZN(n22427) );
  AOI22_X1 U23988 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22482), .B1(
        n22427), .B2(n22481), .ZN(n22384) );
  OAI211_X1 U23989 ( .C1(n22424), .C2(n22491), .A(n22385), .B(n22384), .ZN(
        P1_U3037) );
  AOI22_X1 U23990 ( .A1(n22486), .A2(n22427), .B1(n22485), .B2(n22428), .ZN(
        n22387) );
  INV_X1 U23991 ( .A(n22424), .ZN(n22429) );
  AOI22_X1 U23992 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22488), .B1(
        n22487), .B2(n22429), .ZN(n22386) );
  OAI211_X1 U23993 ( .C1(n22432), .C2(n22491), .A(n22387), .B(n22386), .ZN(
        P1_U3045) );
  INV_X1 U23994 ( .A(n22428), .ZN(n22414) );
  OAI22_X1 U23995 ( .A1(n22493), .A2(n22432), .B1(n22492), .B2(n22414), .ZN(
        n22388) );
  INV_X1 U23996 ( .A(n22388), .ZN(n22390) );
  AOI22_X1 U23997 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22496), .B1(
        n22427), .B2(n22495), .ZN(n22389) );
  OAI211_X1 U23998 ( .C1(n22424), .C2(n22500), .A(n22390), .B(n22389), .ZN(
        P1_U3053) );
  OAI22_X1 U23999 ( .A1(n22500), .A2(n22432), .B1(n22499), .B2(n22414), .ZN(
        n22391) );
  INV_X1 U24000 ( .A(n22391), .ZN(n22393) );
  AOI22_X1 U24001 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22503), .B1(
        n22427), .B2(n22502), .ZN(n22392) );
  OAI211_X1 U24002 ( .C1(n22424), .C2(n22506), .A(n22393), .B(n22392), .ZN(
        P1_U3061) );
  AOI22_X1 U24003 ( .A1(n22428), .A2(n22508), .B1(n22427), .B2(n22507), .ZN(
        n22395) );
  AOI22_X1 U24004 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n22510), .B1(
        n22509), .B2(n22421), .ZN(n22394) );
  OAI211_X1 U24005 ( .C1(n22424), .C2(n22513), .A(n22395), .B(n22394), .ZN(
        P1_U3069) );
  AOI22_X1 U24006 ( .A1(n22515), .A2(n22427), .B1(n22428), .B2(n22514), .ZN(
        n22398) );
  AOI22_X1 U24007 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n22517), .B1(
        n22396), .B2(n22429), .ZN(n22397) );
  OAI211_X1 U24008 ( .C1(n22432), .C2(n22513), .A(n22398), .B(n22397), .ZN(
        P1_U3077) );
  OAI22_X1 U24009 ( .A1(n22527), .A2(n22424), .B1(n22520), .B2(n22414), .ZN(
        n22399) );
  INV_X1 U24010 ( .A(n22399), .ZN(n22401) );
  AOI22_X1 U24011 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22524), .B1(
        n22427), .B2(n22523), .ZN(n22400) );
  OAI211_X1 U24012 ( .C1(n22432), .C2(n22521), .A(n22401), .B(n22400), .ZN(
        P1_U3085) );
  AOI22_X1 U24013 ( .A1(n22529), .A2(n22427), .B1(n22528), .B2(n22428), .ZN(
        n22403) );
  AOI22_X1 U24014 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n22531), .B1(
        n22537), .B2(n22429), .ZN(n22402) );
  OAI211_X1 U24015 ( .C1(n22432), .C2(n22527), .A(n22403), .B(n22402), .ZN(
        P1_U3093) );
  AOI22_X1 U24016 ( .A1(n22536), .A2(n22427), .B1(n22428), .B2(n22535), .ZN(
        n22405) );
  AOI22_X1 U24017 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n22538), .B1(
        n22537), .B2(n22421), .ZN(n22404) );
  OAI211_X1 U24018 ( .C1(n22424), .C2(n22546), .A(n22405), .B(n22404), .ZN(
        P1_U3101) );
  INV_X1 U24019 ( .A(n22406), .ZN(n22542) );
  AOI22_X1 U24020 ( .A1(n22542), .A2(n22427), .B1(n22541), .B2(n22428), .ZN(
        n22408) );
  AOI22_X1 U24021 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22543), .B1(
        n22548), .B2(n22429), .ZN(n22407) );
  OAI211_X1 U24022 ( .C1(n22432), .C2(n22546), .A(n22408), .B(n22407), .ZN(
        P1_U3109) );
  AOI22_X1 U24023 ( .A1(n22548), .A2(n22421), .B1(n22547), .B2(n22428), .ZN(
        n22410) );
  AOI22_X1 U24024 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22550), .B1(
        n22427), .B2(n22549), .ZN(n22409) );
  OAI211_X1 U24025 ( .C1(n22424), .C2(n22553), .A(n22410), .B(n22409), .ZN(
        P1_U3117) );
  AOI22_X1 U24026 ( .A1(n22555), .A2(n22427), .B1(n22554), .B2(n22428), .ZN(
        n22413) );
  AOI22_X1 U24027 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n22557), .B1(
        n22411), .B2(n22429), .ZN(n22412) );
  OAI211_X1 U24028 ( .C1(n22432), .C2(n22553), .A(n22413), .B(n22412), .ZN(
        P1_U3125) );
  OAI22_X1 U24029 ( .A1(n22573), .A2(n22424), .B1(n22561), .B2(n22414), .ZN(
        n22415) );
  INV_X1 U24030 ( .A(n22415), .ZN(n22417) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22564), .B1(
        n22427), .B2(n22563), .ZN(n22416) );
  OAI211_X1 U24032 ( .C1(n22432), .C2(n22567), .A(n22417), .B(n22416), .ZN(
        P1_U3133) );
  INV_X1 U24033 ( .A(n22418), .ZN(n22569) );
  AOI22_X1 U24034 ( .A1(n22427), .A2(n22569), .B1(n22428), .B2(n22568), .ZN(
        n22420) );
  AOI22_X1 U24035 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22570), .B1(
        n22577), .B2(n22429), .ZN(n22419) );
  OAI211_X1 U24036 ( .C1(n22432), .C2(n22573), .A(n22420), .B(n22419), .ZN(
        P1_U3141) );
  AOI22_X1 U24037 ( .A1(n22428), .A2(n22575), .B1(n22427), .B2(n22574), .ZN(
        n22423) );
  AOI22_X1 U24038 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22578), .B1(
        n22577), .B2(n22421), .ZN(n22422) );
  OAI211_X1 U24039 ( .C1(n22424), .C2(n22591), .A(n22423), .B(n22422), .ZN(
        P1_U3149) );
  INV_X1 U24040 ( .A(n22425), .ZN(n22584) );
  INV_X1 U24041 ( .A(n22426), .ZN(n22582) );
  AOI22_X1 U24042 ( .A1(n22428), .A2(n22584), .B1(n22427), .B2(n22582), .ZN(
        n22431) );
  AOI22_X1 U24043 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n22588), .B1(
        n22587), .B2(n22429), .ZN(n22430) );
  OAI211_X1 U24044 ( .C1(n22432), .C2(n22591), .A(n22431), .B(n22430), .ZN(
        P1_U3157) );
  AOI22_X1 U24045 ( .A1(n22587), .A2(n22456), .B1(n22455), .B2(n22478), .ZN(
        n22434) );
  AOI22_X1 U24046 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22482), .B1(
        n22454), .B2(n22481), .ZN(n22433) );
  OAI211_X1 U24047 ( .C1(n22459), .C2(n22491), .A(n22434), .B(n22433), .ZN(
        P1_U3038) );
  AOI22_X1 U24048 ( .A1(n22486), .A2(n22454), .B1(n22455), .B2(n22485), .ZN(
        n22437) );
  AOI22_X1 U24049 ( .A1(n22488), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n22435), .B2(n22456), .ZN(n22436) );
  OAI211_X1 U24050 ( .C1(n22459), .C2(n22493), .A(n22437), .B(n22436), .ZN(
        P1_U3046) );
  OAI22_X1 U24051 ( .A1(n22493), .A2(n22442), .B1(n22492), .B2(n22441), .ZN(
        n22438) );
  INV_X1 U24052 ( .A(n22438), .ZN(n22440) );
  AOI22_X1 U24053 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22496), .B1(
        n22454), .B2(n22495), .ZN(n22439) );
  OAI211_X1 U24054 ( .C1(n22459), .C2(n22500), .A(n22440), .B(n22439), .ZN(
        P1_U3054) );
  OAI22_X1 U24055 ( .A1(n22500), .A2(n22442), .B1(n22441), .B2(n22499), .ZN(
        n22443) );
  INV_X1 U24056 ( .A(n22443), .ZN(n22445) );
  AOI22_X1 U24057 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22503), .B1(
        n22454), .B2(n22502), .ZN(n22444) );
  OAI211_X1 U24058 ( .C1(n22459), .C2(n22506), .A(n22445), .B(n22444), .ZN(
        P1_U3062) );
  AOI22_X1 U24059 ( .A1(n22455), .A2(n22508), .B1(n22454), .B2(n22507), .ZN(
        n22447) );
  AOI22_X1 U24060 ( .A1(n22510), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n22509), .B2(n22456), .ZN(n22446) );
  OAI211_X1 U24061 ( .C1(n22459), .C2(n22513), .A(n22447), .B(n22446), .ZN(
        P1_U3070) );
  AOI22_X1 U24062 ( .A1(n22529), .A2(n22454), .B1(n22528), .B2(n22455), .ZN(
        n22449) );
  AOI22_X1 U24063 ( .A1(n22531), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n22530), .B2(n22456), .ZN(n22448) );
  OAI211_X1 U24064 ( .C1(n22459), .C2(n22534), .A(n22449), .B(n22448), .ZN(
        P1_U3094) );
  AOI22_X1 U24065 ( .A1(n22536), .A2(n22454), .B1(n22455), .B2(n22535), .ZN(
        n22451) );
  AOI22_X1 U24066 ( .A1(n22538), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n22537), .B2(n22456), .ZN(n22450) );
  OAI211_X1 U24067 ( .C1(n22459), .C2(n22546), .A(n22451), .B(n22450), .ZN(
        P1_U3102) );
  AOI22_X1 U24068 ( .A1(n22548), .A2(n22456), .B1(n22455), .B2(n22547), .ZN(
        n22453) );
  AOI22_X1 U24069 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22550), .B1(
        n22454), .B2(n22549), .ZN(n22452) );
  OAI211_X1 U24070 ( .C1(n22459), .C2(n22553), .A(n22453), .B(n22452), .ZN(
        P1_U3118) );
  AOI22_X1 U24071 ( .A1(n22455), .A2(n22575), .B1(n22454), .B2(n22574), .ZN(
        n22458) );
  AOI22_X1 U24072 ( .A1(n22578), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n22577), .B2(n22456), .ZN(n22457) );
  OAI211_X1 U24073 ( .C1(n22459), .C2(n22591), .A(n22458), .B(n22457), .ZN(
        P1_U3150) );
  AOI22_X1 U24074 ( .A1(n22587), .A2(n22470), .B1(n22478), .B2(n22468), .ZN(
        n22461) );
  AOI22_X1 U24075 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22482), .B1(
        n22469), .B2(n22481), .ZN(n22460) );
  OAI211_X1 U24076 ( .C1(n22473), .C2(n22491), .A(n22461), .B(n22460), .ZN(
        P1_U3039) );
  AOI22_X1 U24077 ( .A1(n22469), .A2(n22507), .B1(n22468), .B2(n22508), .ZN(
        n22463) );
  AOI22_X1 U24078 ( .A1(n22510), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n22509), .B2(n22470), .ZN(n22462) );
  OAI211_X1 U24079 ( .C1(n22473), .C2(n22513), .A(n22463), .B(n22462), .ZN(
        P1_U3071) );
  AOI22_X1 U24080 ( .A1(n22469), .A2(n22536), .B1(n22468), .B2(n22535), .ZN(
        n22465) );
  AOI22_X1 U24081 ( .A1(n22538), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22537), .B2(n22470), .ZN(n22464) );
  OAI211_X1 U24082 ( .C1(n22473), .C2(n22546), .A(n22465), .B(n22464), .ZN(
        P1_U3103) );
  AOI22_X1 U24083 ( .A1(n22548), .A2(n22470), .B1(n22547), .B2(n22468), .ZN(
        n22467) );
  AOI22_X1 U24084 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22550), .B1(
        n22469), .B2(n22549), .ZN(n22466) );
  OAI211_X1 U24085 ( .C1(n22473), .C2(n22553), .A(n22467), .B(n22466), .ZN(
        P1_U3119) );
  AOI22_X1 U24086 ( .A1(n22469), .A2(n22574), .B1(n22468), .B2(n22575), .ZN(
        n22472) );
  AOI22_X1 U24087 ( .A1(n22578), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n22577), .B2(n22470), .ZN(n22471) );
  OAI211_X1 U24088 ( .C1(n22473), .C2(n22591), .A(n22472), .B(n22471), .ZN(
        P1_U3151) );
  AOI22_X1 U24089 ( .A1(DATAI_31_), .A2(n11152), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n22474), .ZN(n22592) );
  INV_X1 U24090 ( .A(n22592), .ZN(n22576) );
  NOR2_X2 U24091 ( .A1(n22477), .A2(n22476), .ZN(n22585) );
  AOI22_X1 U24092 ( .A1(n22587), .A2(n22576), .B1(n22585), .B2(n22478), .ZN(
        n22484) );
  NOR2_X2 U24093 ( .A1(n22480), .A2(n22479), .ZN(n22583) );
  AOI22_X1 U24094 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22482), .B1(
        n22583), .B2(n22481), .ZN(n22483) );
  OAI211_X1 U24095 ( .C1(n22581), .C2(n22491), .A(n22484), .B(n22483), .ZN(
        P1_U3040) );
  AOI22_X1 U24096 ( .A1(n22486), .A2(n22583), .B1(n22485), .B2(n22585), .ZN(
        n22490) );
  INV_X1 U24097 ( .A(n22581), .ZN(n22586) );
  AOI22_X1 U24098 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22488), .B1(
        n22487), .B2(n22586), .ZN(n22489) );
  OAI211_X1 U24099 ( .C1(n22592), .C2(n22491), .A(n22490), .B(n22489), .ZN(
        P1_U3048) );
  INV_X1 U24100 ( .A(n22585), .ZN(n22560) );
  OAI22_X1 U24101 ( .A1(n22493), .A2(n22592), .B1(n22492), .B2(n22560), .ZN(
        n22494) );
  INV_X1 U24102 ( .A(n22494), .ZN(n22498) );
  AOI22_X1 U24103 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22496), .B1(
        n22583), .B2(n22495), .ZN(n22497) );
  OAI211_X1 U24104 ( .C1(n22581), .C2(n22500), .A(n22498), .B(n22497), .ZN(
        P1_U3056) );
  OAI22_X1 U24105 ( .A1(n22500), .A2(n22592), .B1(n22499), .B2(n22560), .ZN(
        n22501) );
  INV_X1 U24106 ( .A(n22501), .ZN(n22505) );
  AOI22_X1 U24107 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22503), .B1(
        n22583), .B2(n22502), .ZN(n22504) );
  OAI211_X1 U24108 ( .C1(n22581), .C2(n22506), .A(n22505), .B(n22504), .ZN(
        P1_U3064) );
  AOI22_X1 U24109 ( .A1(n22585), .A2(n22508), .B1(n22583), .B2(n22507), .ZN(
        n22512) );
  AOI22_X1 U24110 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n22510), .B1(
        n22509), .B2(n22576), .ZN(n22511) );
  OAI211_X1 U24111 ( .C1(n22581), .C2(n22513), .A(n22512), .B(n22511), .ZN(
        P1_U3072) );
  AOI22_X1 U24112 ( .A1(n22515), .A2(n22583), .B1(n22585), .B2(n22514), .ZN(
        n22519) );
  AOI22_X1 U24113 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22517), .B1(
        n22516), .B2(n22576), .ZN(n22518) );
  OAI211_X1 U24114 ( .C1(n22581), .C2(n22521), .A(n22519), .B(n22518), .ZN(
        P1_U3080) );
  OAI22_X1 U24115 ( .A1(n22521), .A2(n22592), .B1(n22520), .B2(n22560), .ZN(
        n22522) );
  INV_X1 U24116 ( .A(n22522), .ZN(n22526) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22524), .B1(
        n22583), .B2(n22523), .ZN(n22525) );
  OAI211_X1 U24118 ( .C1(n22581), .C2(n22527), .A(n22526), .B(n22525), .ZN(
        P1_U3088) );
  AOI22_X1 U24119 ( .A1(n22529), .A2(n22583), .B1(n22528), .B2(n22585), .ZN(
        n22533) );
  AOI22_X1 U24120 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22531), .B1(
        n22530), .B2(n22576), .ZN(n22532) );
  OAI211_X1 U24121 ( .C1(n22581), .C2(n22534), .A(n22533), .B(n22532), .ZN(
        P1_U3096) );
  AOI22_X1 U24122 ( .A1(n22536), .A2(n22583), .B1(n22585), .B2(n22535), .ZN(
        n22540) );
  AOI22_X1 U24123 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22538), .B1(
        n22537), .B2(n22576), .ZN(n22539) );
  OAI211_X1 U24124 ( .C1(n22581), .C2(n22546), .A(n22540), .B(n22539), .ZN(
        P1_U3104) );
  AOI22_X1 U24125 ( .A1(n22542), .A2(n22583), .B1(n22541), .B2(n22585), .ZN(
        n22545) );
  AOI22_X1 U24126 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22543), .B1(
        n22548), .B2(n22586), .ZN(n22544) );
  OAI211_X1 U24127 ( .C1(n22592), .C2(n22546), .A(n22545), .B(n22544), .ZN(
        P1_U3112) );
  AOI22_X1 U24128 ( .A1(n22548), .A2(n22576), .B1(n22547), .B2(n22585), .ZN(
        n22552) );
  AOI22_X1 U24129 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22550), .B1(
        n22583), .B2(n22549), .ZN(n22551) );
  OAI211_X1 U24130 ( .C1(n22581), .C2(n22553), .A(n22552), .B(n22551), .ZN(
        P1_U3120) );
  AOI22_X1 U24131 ( .A1(n22555), .A2(n22583), .B1(n22554), .B2(n22585), .ZN(
        n22559) );
  AOI22_X1 U24132 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n22557), .B1(
        n22556), .B2(n22576), .ZN(n22558) );
  OAI211_X1 U24133 ( .C1(n22581), .C2(n22567), .A(n22559), .B(n22558), .ZN(
        P1_U3128) );
  OAI22_X1 U24134 ( .A1(n22573), .A2(n22581), .B1(n22561), .B2(n22560), .ZN(
        n22562) );
  INV_X1 U24135 ( .A(n22562), .ZN(n22566) );
  AOI22_X1 U24136 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22564), .B1(
        n22583), .B2(n22563), .ZN(n22565) );
  OAI211_X1 U24137 ( .C1(n22592), .C2(n22567), .A(n22566), .B(n22565), .ZN(
        P1_U3136) );
  AOI22_X1 U24138 ( .A1(n22583), .A2(n22569), .B1(n22585), .B2(n22568), .ZN(
        n22572) );
  AOI22_X1 U24139 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22570), .B1(
        n22577), .B2(n22586), .ZN(n22571) );
  OAI211_X1 U24140 ( .C1(n22592), .C2(n22573), .A(n22572), .B(n22571), .ZN(
        P1_U3144) );
  AOI22_X1 U24141 ( .A1(n22585), .A2(n22575), .B1(n22583), .B2(n22574), .ZN(
        n22580) );
  AOI22_X1 U24142 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22578), .B1(
        n22577), .B2(n22576), .ZN(n22579) );
  OAI211_X1 U24143 ( .C1(n22581), .C2(n22591), .A(n22580), .B(n22579), .ZN(
        P1_U3152) );
  AOI22_X1 U24144 ( .A1(n22585), .A2(n22584), .B1(n22583), .B2(n22582), .ZN(
        n22590) );
  AOI22_X1 U24145 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22588), .B1(
        n22587), .B2(n22586), .ZN(n22589) );
  OAI211_X1 U24146 ( .C1(n22592), .C2(n22591), .A(n22590), .B(n22589), .ZN(
        P1_U3160) );
  AOI22_X1 U24147 ( .A1(n22596), .A2(n22595), .B1(n22594), .B2(n22593), .ZN(
        P1_U3486) );
  BUF_X1 U11568 ( .A(n14414), .Z(n18105) );
  CLKBUF_X3 U11598 ( .A(n18109), .Z(n11176) );
  AND2_X1 U14469 ( .A1(n12907), .A2(n12893), .ZN(n19682) );
  AOI221_X1 U11259 ( .B1(n19733), .B2(n19715), .C1(n19733), .C2(n20218), .A(
        n20211), .ZN(n19711) );
  CLKBUF_X1 U11306 ( .A(n12991), .Z(n19759) );
  CLKBUF_X1 U11308 ( .A(n18108), .Z(n17900) );
  NAND2_X1 U11312 ( .A1(n12476), .A2(n12475), .ZN(n12477) );
  CLKBUF_X1 U11314 ( .A(n11839), .Z(n14043) );
  AND2_X1 U11316 ( .A1(n18340), .A2(n18339), .ZN(n18352) );
  CLKBUF_X1 U11323 ( .A(n17722), .Z(n17732) );
  CLKBUF_X1 U11344 ( .A(n20660), .Z(n20657) );
  OR3_X1 U11362 ( .A1(n16549), .A2(n22476), .A3(n11832), .ZN(n22598) );
  OR3_X1 U11363 ( .A1(n22169), .A2(n15750), .A3(n19799), .ZN(n22599) );
  OR2_X1 U11392 ( .A1(n21351), .A2(n21249), .ZN(n22600) );
  OR2_X1 U11637 ( .A1(n21351), .A2(n19534), .ZN(n22601) );
endmodule

