

module b20_C_SARLock_k_64_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102;

  INV_X4 U4782 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U4783 ( .A1(n6710), .A2(n6707), .ZN(n7679) );
  INV_X1 U4785 ( .A(n4960), .ZN(n5094) );
  AND2_X2 U4787 ( .A1(n5775), .A2(n5976), .ZN(n6248) );
  NAND2_X1 U4788 ( .A1(n8192), .A2(n5977), .ZN(n5983) );
  NAND2_X1 U4789 ( .A1(n6827), .A2(n6794), .ZN(n4277) );
  NOR2_X1 U4790 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4801) );
  INV_X1 U4791 ( .A(n6286), .ZN(n6793) );
  OR2_X1 U4792 ( .A1(n9303), .A2(n4551), .ZN(n4545) );
  INV_X1 U4793 ( .A(n8547), .ZN(n8540) );
  AND2_X1 U4794 ( .A1(n8371), .A2(n8559), .ZN(n8547) );
  INV_X1 U4795 ( .A(n6794), .ZN(n6823) );
  INV_X2 U4796 ( .A(n5846), .ZN(n8225) );
  INV_X1 U4797 ( .A(n5846), .ZN(n5906) );
  INV_X1 U4798 ( .A(n6002), .ZN(n6188) );
  INV_X1 U4799 ( .A(n5983), .ZN(n5993) );
  NAND2_X1 U4800 ( .A1(n7679), .A2(n7683), .ZN(n7678) );
  NAND2_X1 U4801 ( .A1(n5779), .A2(n5778), .ZN(n5621) );
  CLKBUF_X2 U4802 ( .A(n5371), .Z(n8072) );
  AOI21_X2 U4803 ( .B1(n7956), .B2(n8030), .A(n8029), .ZN(n8028) );
  NOR2_X2 U4804 ( .A1(n6750), .A2(n6242), .ZN(n9350) );
  OAI211_X2 U4805 ( .C1(n6869), .C2(n4932), .A(n4598), .B(n4597), .ZN(n7264)
         );
  OAI22_X2 U4806 ( .A1(n8262), .A2(n8263), .B1(n8766), .B2(n5903), .ZN(n8241)
         );
  AOI22_X2 U4807 ( .A1(n8204), .A2(n8743), .B1(n5901), .B2(n5900), .ZN(n8262)
         );
  OAI21_X2 U4808 ( .B1(n8301), .B2(n8303), .A(n5908), .ZN(n5911) );
  AOI21_X2 U4809 ( .B1(n8241), .B2(n8242), .A(n4336), .ZN(n8301) );
  AND2_X1 U4810 ( .A1(n9126), .A2(n6804), .ZN(n6842) );
  NAND2_X1 U4811 ( .A1(n7459), .A2(n7463), .ZN(n7460) );
  NAND2_X1 U4812 ( .A1(n6304), .A2(n4306), .ZN(n7487) );
  NAND2_X4 U4813 ( .A1(n6827), .A2(n6794), .ZN(n6286) );
  NAND2_X1 U4814 ( .A1(n4836), .A2(n4835), .ZN(n4981) );
  CLKBUF_X1 U4815 ( .A(n6267), .Z(n4278) );
  CLKBUF_X2 U4816 ( .A(n5983), .Z(n6197) );
  CLKBUF_X1 U4817 ( .A(n5620), .Z(n5735) );
  NAND2_X1 U4818 ( .A1(n4807), .A2(n4806), .ZN(n8155) );
  AOI211_X1 U4819 ( .C1(n8181), .C2(n9836), .A(n8180), .B(n8179), .ZN(n8182)
         );
  AOI21_X1 U4820 ( .B1(n6842), .B2(n6841), .A(n6840), .ZN(n6843) );
  AOI211_X1 U4821 ( .C1(n10026), .C2(n8375), .A(n8201), .B(n8200), .ZN(n8202)
         );
  NOR2_X1 U4822 ( .A1(n9103), .A2(n9038), .ZN(n9043) );
  OAI21_X1 U4823 ( .B1(n5970), .B2(n5969), .A(n8523), .ZN(n6486) );
  OAI21_X1 U4824 ( .B1(n9301), .B2(n4448), .A(n4446), .ZN(n4445) );
  NAND2_X1 U4825 ( .A1(n8741), .A2(n4783), .ZN(n8731) );
  NAND2_X1 U4826 ( .A1(n6515), .A2(n6514), .ZN(n8188) );
  NAND2_X1 U4827 ( .A1(n5758), .A2(n5757), .ZN(n6672) );
  AND2_X1 U4828 ( .A1(n4453), .A2(n4282), .ZN(n9282) );
  XNOR2_X1 U4829 ( .A(n6507), .B(n6506), .ZN(n8326) );
  AOI21_X1 U4830 ( .B1(n9347), .B2(n6156), .A(n4771), .ZN(n9333) );
  AND2_X1 U4831 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  INV_X1 U4832 ( .A(n4454), .ZN(n9347) );
  NAND2_X1 U4833 ( .A1(n5257), .A2(n5256), .ZN(n8970) );
  NAND2_X1 U4834 ( .A1(n4589), .A2(n4587), .ZN(n8938) );
  AND2_X1 U4835 ( .A1(n4365), .A2(n4364), .ZN(n4363) );
  OAI21_X1 U4836 ( .B1(n8138), .B2(n8145), .A(n6113), .ZN(n9422) );
  OAI21_X1 U4837 ( .B1(n8002), .B2(n4468), .A(n4466), .ZN(n8138) );
  OAI21_X1 U4838 ( .B1(n7817), .B2(n4498), .A(n4497), .ZN(n5465) );
  NAND2_X1 U4839 ( .A1(n6320), .A2(n6319), .ZN(n7461) );
  NAND2_X1 U4840 ( .A1(n4496), .A2(n5459), .ZN(n7738) );
  OR2_X1 U4841 ( .A1(n9142), .A2(n8121), .ZN(n6722) );
  OR2_X1 U4842 ( .A1(n7670), .A2(n5457), .ZN(n4496) );
  NAND2_X1 U4843 ( .A1(n5693), .A2(n5692), .ZN(n9033) );
  OAI21_X1 U4844 ( .B1(n7526), .B2(n4540), .A(n4539), .ZN(n4538) );
  XNOR2_X1 U4845 ( .A(n5105), .B(n4780), .ZN(n7252) );
  NAND2_X1 U4846 ( .A1(n5689), .A2(n5688), .ZN(n8089) );
  OR2_X1 U4847 ( .A1(n9976), .A2(n7680), .ZN(n6569) );
  INV_X2 U4848 ( .A(n10034), .ZN(n4275) );
  OR2_X1 U4849 ( .A1(n7588), .A2(n9967), .ZN(n9818) );
  XNOR2_X1 U4850 ( .A(n4408), .B(n5027), .ZN(n6905) );
  NAND2_X1 U4851 ( .A1(n5822), .A2(n7240), .ZN(n5827) );
  NAND2_X2 U4852 ( .A1(n7358), .A2(n9878), .ZN(n9836) );
  CLKBUF_X1 U4853 ( .A(n5393), .Z(n5579) );
  INV_X2 U4854 ( .A(n6883), .ZN(n6943) );
  INV_X4 U4855 ( .A(n4952), .ZN(n8316) );
  AND4_X1 U4856 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n7680)
         );
  NAND4_X1 U4857 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n9176)
         );
  AND4_X1 U4858 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n7588)
         );
  OAI21_X1 U4859 ( .B1(n4979), .B2(n4981), .A(n4841), .ZN(n4994) );
  AND2_X1 U4860 ( .A1(n7353), .A2(n6847), .ZN(n6259) );
  OAI21_X1 U4861 ( .B1(n5169), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5171) );
  OR2_X1 U4862 ( .A1(n7074), .A2(n5530), .ZN(n7072) );
  NAND2_X1 U4863 ( .A1(n5804), .A2(n6745), .ZN(n6768) );
  AND3_X1 U4864 ( .A1(n5629), .A2(n5628), .A3(n5627), .ZN(n9924) );
  INV_X2 U4865 ( .A(n4932), .ZN(n8325) );
  CLKBUF_X1 U4866 ( .A(n4945), .Z(n5135) );
  INV_X1 U4867 ( .A(n5620), .ZN(n5720) );
  NOR2_X1 U4868 ( .A1(n5130), .A2(n5129), .ZN(n5133) );
  INV_X1 U4869 ( .A(n7772), .ZN(n6220) );
  MUX2_X1 U4870 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4805), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4807) );
  OAI211_X1 U4871 ( .C1(n4879), .C2(n4878), .A(n4877), .B(n4876), .ZN(n5371)
         );
  NAND2_X1 U4872 ( .A1(n5801), .A2(n5762), .ZN(n7772) );
  OAI21_X1 U4873 ( .B1(n5703), .B2(n4366), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5712) );
  XNOR2_X1 U4874 ( .A(n5773), .B(n5770), .ZN(n5778) );
  NAND2_X2 U4875 ( .A1(n6853), .A2(P1_U3086), .ZN(n9675) );
  OR2_X1 U4876 ( .A1(n5354), .A2(n4724), .ZN(n4876) );
  OR2_X1 U4877 ( .A1(n5609), .A2(n9670), .ZN(n4603) );
  AND2_X1 U4878 ( .A1(n5691), .A2(n5690), .ZN(n5701) );
  NOR2_X2 U4879 ( .A1(n4949), .A2(n4948), .ZN(n5534) );
  OR2_X1 U4880 ( .A1(n4724), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4508) );
  AND2_X1 U4881 ( .A1(n4793), .A2(n4295), .ZN(n4372) );
  AND4_X1 U4882 ( .A1(n4374), .A2(n4928), .A3(n4796), .A4(n4691), .ZN(n4373)
         );
  INV_X1 U4883 ( .A(n5600), .ZN(n4607) );
  AND2_X1 U4884 ( .A1(n4375), .A2(n4801), .ZN(n4374) );
  AND4_X1 U4885 ( .A1(n5604), .A2(n5603), .A3(n5602), .A4(n5601), .ZN(n5605)
         );
  AND3_X1 U4886 ( .A1(n5170), .A2(n5131), .A3(n4561), .ZN(n4793) );
  NAND2_X1 U4887 ( .A1(n9678), .A2(n4819), .ZN(n4820) );
  AND2_X1 U4888 ( .A1(n4692), .A2(n4799), .ZN(n4691) );
  NOR2_X1 U4889 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5601) );
  NOR2_X1 U4890 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5602) );
  NOR2_X1 U4891 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5603) );
  NOR2_X1 U4892 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5604) );
  INV_X4 U4893 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4894 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5170) );
  NOR2_X1 U4895 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5597) );
  NOR2_X1 U4896 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5596) );
  NOR2_X1 U4897 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5595) );
  INV_X1 U4898 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4882) );
  NOR2_X1 U4899 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5660) );
  AND2_X1 U4900 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9678) );
  NAND3_X2 U4901 ( .A1(n4872), .A2(n4871), .A3(n4764), .ZN(n5370) );
  NAND2_X2 U4902 ( .A1(n5669), .A2(n5668), .ZN(n9976) );
  OAI22_X2 U4903 ( .A1(n5059), .A2(n8572), .B1(n7934), .B2(n7946), .ZN(n8042)
         );
  XNOR2_X2 U4904 ( .A(n5771), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U4905 ( .A1(n5621), .A2(n5611), .ZN(n4276) );
  OAI21_X2 U4906 ( .B1(n9882), .B2(n6224), .A(n6699), .ZN(n6538) );
  AOI21_X2 U4907 ( .B1(n9852), .B2(n6228), .A(n6227), .ZN(n7470) );
  NAND2_X2 U4908 ( .A1(n6226), .A2(n4792), .ZN(n9852) );
  OAI211_X1 U4909 ( .C1(n5621), .C2(n6930), .A(n5617), .B(n5616), .ZN(n6267)
         );
  XNOR2_X2 U4910 ( .A(n4603), .B(n5610), .ZN(n5779) );
  XNOR2_X2 U4911 ( .A(n6268), .B(n6267), .ZN(n9892) );
  OAI21_X1 U4912 ( .B1(n8527), .B2(n8534), .A(n8533), .ZN(n4668) );
  NAND2_X1 U4913 ( .A1(n4409), .A2(n4300), .ZN(n6640) );
  NAND2_X1 U4914 ( .A1(n4410), .A2(n6636), .ZN(n4409) );
  OAI21_X1 U4915 ( .B1(n6633), .B2(n6632), .A(n6631), .ZN(n4410) );
  AND2_X1 U4916 ( .A1(n4642), .A2(n5027), .ZN(n4647) );
  NAND2_X1 U4917 ( .A1(n4895), .A2(n4855), .ZN(n4642) );
  NAND2_X1 U4918 ( .A1(n8731), .A2(n5327), .ZN(n5954) );
  AND2_X1 U4919 ( .A1(n8716), .A2(n5326), .ZN(n5327) );
  INV_X1 U4920 ( .A(n8131), .ZN(n4524) );
  NAND2_X1 U4921 ( .A1(n4526), .A2(n4530), .ZN(n5058) );
  INV_X1 U4922 ( .A(n4531), .ZN(n4530) );
  OAI21_X1 U4923 ( .B1(n7840), .B2(n4532), .A(n7841), .ZN(n4531) );
  OR2_X1 U4924 ( .A1(n8468), .A2(n8866), .ZN(n8475) );
  OAI22_X1 U4925 ( .A1(n9653), .A2(n6796), .B1(n9106), .B2(n6827), .ZN(n6430)
         );
  AND2_X1 U4926 ( .A1(n6344), .A2(n6338), .ZN(n4353) );
  NAND2_X1 U4927 ( .A1(n4390), .A2(n4389), .ZN(n8533) );
  AND2_X1 U4928 ( .A1(n8526), .A2(n8525), .ZN(n4389) );
  OR2_X1 U4929 ( .A1(n9004), .A2(n8868), .ZN(n8473) );
  AOI21_X2 U4930 ( .B1(n6231), .B2(n6551), .A(n6229), .ZN(n6661) );
  NAND2_X1 U4931 ( .A1(n4863), .A2(n9573), .ZN(n4866) );
  INV_X1 U4932 ( .A(n4512), .ZN(n4511) );
  OAI21_X1 U4933 ( .B1(n8835), .B2(n4513), .A(n5179), .ZN(n4512) );
  OR2_X1 U4934 ( .A1(n8914), .A2(n8838), .ZN(n5179) );
  AND2_X1 U4935 ( .A1(n8877), .A2(n8064), .ZN(n8131) );
  OR2_X1 U4936 ( .A1(n8711), .A2(n8721), .ZN(n8524) );
  NAND2_X1 U4937 ( .A1(n8711), .A2(n8721), .ZN(n8523) );
  OR2_X1 U4938 ( .A1(n8982), .A2(n8801), .ZN(n8502) );
  OR2_X1 U4939 ( .A1(n8275), .A2(n8568), .ZN(n8493) );
  OR2_X1 U4940 ( .A1(n8914), .A2(n8257), .ZN(n8484) );
  AND3_X1 U4941 ( .A1(n4800), .A2(n4898), .A3(n4899), .ZN(n4378) );
  NOR2_X1 U4942 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4800) );
  AND2_X1 U4943 ( .A1(n6441), .A2(n4732), .ZN(n4731) );
  OR2_X1 U4944 ( .A1(n9052), .A2(n4338), .ZN(n4732) );
  AOI21_X1 U4945 ( .B1(n4418), .B2(n6651), .A(n4416), .ZN(n4415) );
  NAND2_X1 U4946 ( .A1(n6647), .A2(n5759), .ZN(n4418) );
  NOR2_X1 U4947 ( .A1(n6650), .A2(n8188), .ZN(n4416) );
  OR2_X1 U4948 ( .A1(n8188), .A2(n6915), .ZN(n6760) );
  NAND2_X1 U4949 ( .A1(n8188), .A2(n6915), .ZN(n6770) );
  INV_X1 U4950 ( .A(n6248), .ZN(n6125) );
  OR2_X1 U4951 ( .A1(n6216), .A2(n6835), .ZN(n6676) );
  OAI21_X1 U4952 ( .B1(n4449), .B2(n9275), .A(n4318), .ZN(n4447) );
  INV_X1 U4953 ( .A(n4550), .ZN(n4549) );
  OAI21_X1 U4954 ( .B1(n6244), .B2(n4551), .A(n9275), .ZN(n4550) );
  INV_X1 U4955 ( .A(n4458), .ZN(n4456) );
  INV_X1 U4956 ( .A(n7683), .ZN(n4437) );
  NOR2_X1 U4957 ( .A1(n7683), .A2(n4443), .ZN(n4432) );
  INV_X1 U4958 ( .A(n9820), .ZN(n4443) );
  INV_X1 U4959 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5608) );
  INV_X1 U4960 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4475) );
  AND2_X1 U4961 ( .A1(n5120), .A2(n4780), .ZN(n5121) );
  OAI21_X1 U4962 ( .B1(n5045), .B2(n5044), .A(n4866), .ZN(n5063) );
  AND2_X1 U4963 ( .A1(n4860), .A2(n4859), .ZN(n5027) );
  NAND2_X1 U4964 ( .A1(n4853), .A2(n4852), .ZN(n4896) );
  NAND2_X1 U4965 ( .A1(n4851), .A2(SI_7_), .ZN(n4852) );
  OAI21_X1 U4966 ( .B1(n4994), .B2(n4993), .A(n4845), .ZN(n5010) );
  NAND2_X1 U4967 ( .A1(n7916), .A2(n5868), .ZN(n4715) );
  NAND2_X1 U4968 ( .A1(n4713), .A2(n4705), .ZN(n4704) );
  INV_X1 U4969 ( .A(n8270), .ZN(n4705) );
  INV_X1 U4970 ( .A(n8577), .ZN(n7417) );
  INV_X1 U4971 ( .A(n7309), .ZN(n5836) );
  AOI21_X1 U4972 ( .B1(n4712), .B2(n4711), .A(n4710), .ZN(n4709) );
  INV_X1 U4973 ( .A(n8211), .ZN(n4710) );
  INV_X1 U4974 ( .A(n8291), .ZN(n4711) );
  INV_X1 U4975 ( .A(n5053), .ZN(n5960) );
  NAND2_X1 U4976 ( .A1(n4809), .A2(n8155), .ZN(n8318) );
  NAND2_X1 U4977 ( .A1(n4685), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U4978 ( .A1(n7665), .A2(n7666), .ZN(n7664) );
  XNOR2_X1 U4979 ( .A(n5465), .B(n8025), .ZN(n8021) );
  OR2_X1 U4980 ( .A1(n8012), .A2(n4677), .ZN(n4674) );
  OR2_X1 U4981 ( .A1(n8618), .A2(n5068), .ZN(n4677) );
  NAND2_X1 U4982 ( .A1(n5503), .A2(n4676), .ZN(n4675) );
  INV_X1 U4983 ( .A(n8618), .ZN(n4676) );
  NAND2_X1 U4984 ( .A1(n5281), .A2(n5280), .ZN(n5301) );
  INV_X1 U4985 ( .A(n5282), .ZN(n5281) );
  NAND2_X1 U4986 ( .A1(n4514), .A2(n4516), .ZN(n8929) );
  AND2_X1 U4987 ( .A1(n8930), .A2(n4517), .ZN(n4516) );
  NAND2_X1 U4988 ( .A1(n4518), .A2(n4520), .ZN(n4517) );
  INV_X1 U4989 ( .A(n4538), .ZN(n7635) );
  AND2_X1 U4990 ( .A1(n7538), .A2(n8576), .ZN(n4540) );
  NAND2_X1 U4991 ( .A1(n7530), .A2(n7637), .ZN(n4539) );
  OAI21_X1 U4992 ( .B1(n8715), .B2(n8332), .A(n8520), .ZN(n5970) );
  NAND2_X1 U4993 ( .A1(n5898), .A2(n8743), .ZN(n5270) );
  NAND2_X1 U4994 ( .A1(n8970), .A2(n8743), .ZN(n8748) );
  INV_X1 U4995 ( .A(n6497), .ZN(n5190) );
  INV_X1 U4996 ( .A(n8928), .ZN(n8862) );
  NAND2_X1 U4997 ( .A1(n4876), .A2(n4870), .ZN(n4872) );
  NOR2_X1 U4998 ( .A1(n4869), .A2(n4868), .ZN(n4870) );
  AOI21_X1 U4999 ( .B1(n9052), .B2(n4360), .A(n4338), .ZN(n4359) );
  INV_X1 U5000 ( .A(n9052), .ZN(n4361) );
  INV_X1 U5001 ( .A(n6426), .ZN(n4360) );
  AND2_X1 U5002 ( .A1(n6193), .A2(n6192), .ZN(n6787) );
  OR2_X1 U5003 ( .A1(n9232), .A2(n9231), .ZN(n9234) );
  NAND2_X1 U5004 ( .A1(n6676), .A2(n6737), .ZN(n6669) );
  NOR2_X1 U5005 ( .A1(n9326), .A2(n9156), .ZN(n6172) );
  AOI21_X1 U5006 ( .B1(n4470), .B2(n4467), .A(n4311), .ZN(n4466) );
  INV_X1 U5007 ( .A(n4470), .ZN(n4468) );
  NAND2_X1 U5008 ( .A1(n5955), .A2(n5756), .ZN(n5744) );
  INV_X1 U5009 ( .A(n5621), .ZN(n5719) );
  NAND2_X1 U5010 ( .A1(n5610), .A2(n4735), .ZN(n4734) );
  INV_X1 U5011 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4735) );
  OAI21_X1 U5012 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(n6512) );
  AOI21_X1 U5013 ( .B1(n5966), .B2(n8928), .A(n5965), .ZN(n8162) );
  NOR2_X1 U5014 ( .A1(n6517), .A2(n9425), .ZN(n8184) );
  NOR2_X1 U5015 ( .A1(n6504), .A2(n6672), .ZN(n6516) );
  NAND2_X1 U5016 ( .A1(n4396), .A2(n8547), .ZN(n4395) );
  NAND2_X1 U5017 ( .A1(n8448), .A2(n4305), .ZN(n4396) );
  NAND2_X1 U5018 ( .A1(n8474), .A2(n4404), .ZN(n4403) );
  AND2_X1 U5019 ( .A1(n8473), .A2(n8540), .ZN(n4404) );
  NAND2_X1 U5020 ( .A1(n6600), .A2(n6641), .ZN(n6603) );
  AND2_X1 U5021 ( .A1(n9349), .A2(n6623), .ZN(n4424) );
  AND2_X1 U5022 ( .A1(n6685), .A2(n6649), .ZN(n4425) );
  INV_X1 U5023 ( .A(n6557), .ZN(n6231) );
  INV_X1 U5024 ( .A(n5593), .ZN(n4625) );
  INV_X1 U5025 ( .A(n8651), .ZN(n4673) );
  INV_X1 U5026 ( .A(n4591), .ZN(n4590) );
  OAI21_X1 U5027 ( .B1(n8458), .B2(n8456), .A(n8464), .ZN(n4591) );
  AOI21_X1 U5028 ( .B1(n4353), .B2(n6335), .A(n4351), .ZN(n4350) );
  INV_X1 U5029 ( .A(n6349), .ZN(n4351) );
  OR2_X1 U5030 ( .A1(n6199), .A2(n9130), .ZN(n6637) );
  AND2_X1 U5031 ( .A1(n9082), .A2(n9163), .ZN(n6594) );
  NAND2_X1 U5032 ( .A1(n6231), .A2(n6550), .ZN(n6659) );
  NOR2_X1 U5033 ( .A1(n9375), .A2(n9391), .ZN(n4621) );
  NAND2_X1 U5034 ( .A1(n4857), .A2(n4856), .ZN(n4860) );
  NOR2_X1 U5035 ( .A1(n8528), .A2(n8547), .ZN(n4662) );
  NAND2_X1 U5036 ( .A1(n4690), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U5037 ( .A1(n8660), .A2(n5512), .ZN(n8682) );
  AND2_X1 U5038 ( .A1(n8662), .A2(n4388), .ZN(n5556) );
  NAND2_X1 U5039 ( .A1(n5554), .A2(n8673), .ZN(n4388) );
  NAND2_X1 U5040 ( .A1(n5344), .A2(n5343), .ZN(n5363) );
  OR2_X1 U5041 ( .A1(n8909), .A2(n8826), .ZN(n8492) );
  AND2_X1 U5042 ( .A1(n7954), .A2(n8573), .ZN(n7840) );
  OR2_X1 U5043 ( .A1(n5329), .A2(n8333), .ZN(n8717) );
  AND2_X1 U5044 ( .A1(n8954), .A2(n8736), .ZN(n8332) );
  OR2_X1 U5045 ( .A1(n8267), .A2(n8735), .ZN(n8513) );
  OR2_X1 U5046 ( .A1(n8759), .A2(n8763), .ZN(n5265) );
  OR2_X1 U5047 ( .A1(n8773), .A2(n4290), .ZN(n8759) );
  OR2_X1 U5048 ( .A1(n4290), .A2(n5267), .ZN(n8760) );
  AND2_X1 U5049 ( .A1(n8776), .A2(n8774), .ZN(n5267) );
  OR2_X1 U5050 ( .A1(n8789), .A2(n8788), .ZN(n8774) );
  OR2_X1 U5051 ( .A1(n8803), .A2(n8789), .ZN(n8773) );
  NOR2_X1 U5052 ( .A1(n5427), .A2(n4570), .ZN(n4569) );
  INV_X1 U5053 ( .A(n8480), .ZN(n4570) );
  OR2_X1 U5054 ( .A1(n8998), .A2(n8851), .ZN(n8387) );
  XNOR2_X1 U5055 ( .A(n5189), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U5056 ( .A1(n5188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5189) );
  INV_X1 U5057 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4899) );
  INV_X1 U5058 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4898) );
  INV_X1 U5059 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4799) );
  OR2_X1 U5060 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  INV_X1 U5061 ( .A(n6651), .ZN(n4417) );
  NOR2_X1 U5062 ( .A1(n6669), .A2(n6643), .ZN(n6644) );
  NOR2_X1 U5063 ( .A1(n4413), .A2(n4415), .ZN(n4412) );
  NOR2_X1 U5064 ( .A1(n4299), .A2(n4414), .ZN(n4413) );
  INV_X1 U5065 ( .A(n6647), .ZN(n4414) );
  NAND2_X1 U5066 ( .A1(n9261), .A2(n7251), .ZN(n6642) );
  NOR2_X1 U5067 ( .A1(n6199), .A2(n4616), .ZN(n4615) );
  INV_X1 U5068 ( .A(n4617), .ZN(n4616) );
  AND2_X1 U5069 ( .A1(n4621), .A2(n9649), .ZN(n4620) );
  AND2_X1 U5070 ( .A1(n9375), .A2(n9159), .ZN(n6148) );
  OR2_X1 U5071 ( .A1(n9375), .A2(n9106), .ZN(n6616) );
  NAND2_X1 U5072 ( .A1(n8144), .A2(n8145), .ZN(n4558) );
  INV_X1 U5073 ( .A(n6594), .ZN(n6598) );
  NOR2_X1 U5074 ( .A1(n8003), .A2(n6104), .ZN(n8125) );
  OR2_X1 U5075 ( .A1(n8004), .A2(n9142), .ZN(n8003) );
  NOR2_X1 U5076 ( .A1(n8089), .A2(n4613), .ZN(n4612) );
  NAND2_X1 U5077 ( .A1(n8038), .A2(n9992), .ZN(n4613) );
  NAND2_X1 U5078 ( .A1(n9959), .A2(n6039), .ZN(n4606) );
  NOR2_X1 U5079 ( .A1(n9336), .A2(n9326), .ZN(n9325) );
  INV_X1 U5080 ( .A(n9829), .ZN(n5675) );
  INV_X1 U5081 ( .A(n4649), .ZN(n5290) );
  NAND2_X1 U5082 ( .A1(n4653), .A2(n4651), .ZN(n4650) );
  INV_X1 U5083 ( .A(n4656), .ZN(n4655) );
  NOR2_X1 U5084 ( .A1(n5249), .A2(n4659), .ZN(n4658) );
  INV_X1 U5085 ( .A(n5232), .ZN(n4659) );
  NAND2_X1 U5086 ( .A1(n4634), .A2(n4632), .ZN(n5216) );
  AOI21_X1 U5087 ( .B1(n4636), .B2(n4303), .A(n4633), .ZN(n4632) );
  INV_X1 U5088 ( .A(n5201), .ZN(n4633) );
  OAI21_X1 U5089 ( .B1(n5063), .B2(n5062), .A(n5061), .ZN(n5078) );
  NAND2_X1 U5090 ( .A1(n4323), .A2(n4643), .ZN(n4427) );
  NAND2_X1 U5091 ( .A1(n4429), .A2(n4854), .ZN(n4855) );
  OAI21_X1 U5092 ( .B1(n4429), .B2(n4854), .A(n4855), .ZN(n4895) );
  NAND2_X1 U5093 ( .A1(n4847), .A2(SI_6_), .ZN(n4848) );
  NAND2_X1 U5094 ( .A1(n5010), .A2(n5008), .ZN(n4849) );
  NAND2_X1 U5095 ( .A1(n4838), .A2(n4837), .ZN(n4841) );
  NOR2_X1 U5096 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5624) );
  AND2_X1 U5097 ( .A1(n8222), .A2(n5910), .ZN(n4698) );
  AND2_X1 U5098 ( .A1(n7512), .A2(n5845), .ZN(n4728) );
  INV_X1 U5099 ( .A(n4709), .ZN(n4708) );
  NOR2_X1 U5100 ( .A1(n4708), .A2(n8270), .ZN(n4707) );
  INV_X1 U5101 ( .A(n5886), .ZN(n4714) );
  OAI211_X1 U5102 ( .C1(n6867), .C2(n4932), .A(n4951), .B(n4950), .ZN(n7269)
         );
  OAI21_X1 U5103 ( .B1(n8365), .B2(n8532), .A(n8370), .ZN(n4595) );
  NOR2_X1 U5104 ( .A1(n8368), .A2(n8528), .ZN(n8370) );
  AOI21_X1 U5105 ( .B1(n8369), .B2(n8945), .A(n8390), .ZN(n4594) );
  NOR2_X1 U5106 ( .A1(n8544), .A2(n4400), .ZN(n4399) );
  OR2_X1 U5107 ( .A1(n8541), .A2(n8540), .ZN(n4774) );
  NAND2_X1 U5108 ( .A1(n8884), .A2(n8563), .ZN(n8548) );
  NAND2_X1 U5109 ( .A1(n8545), .A2(n8547), .ZN(n4401) );
  AND2_X1 U5110 ( .A1(n5247), .A2(n5246), .ZN(n8235) );
  NAND2_X1 U5111 ( .A1(n5480), .A2(n5479), .ZN(n4685) );
  XNOR2_X1 U5112 ( .A(n5531), .B(n5480), .ZN(n7017) );
  NAND2_X1 U5113 ( .A1(n6952), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U5114 ( .A1(n7017), .A2(n7016), .ZN(n7015) );
  XNOR2_X1 U5115 ( .A(n5534), .B(n5482), .ZN(n7035) );
  NAND2_X1 U5116 ( .A1(n5449), .A2(n7118), .ZN(n5450) );
  NAND2_X1 U5117 ( .A1(n4493), .A2(n4495), .ZN(n4494) );
  NAND3_X1 U5118 ( .A1(n4494), .A2(P2_REG2_REG_5__SCAN_IN), .A3(n5450), .ZN(
        n7122) );
  NOR2_X1 U5119 ( .A1(n7232), .A2(n4689), .ZN(n7230) );
  AND2_X1 U5120 ( .A1(n8587), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5491) );
  XNOR2_X1 U5121 ( .A(n5456), .B(n6909), .ZN(n7671) );
  NAND2_X1 U5122 ( .A1(n8583), .A2(n5545), .ZN(n7665) );
  NOR2_X1 U5123 ( .A1(n7671), .A2(n5019), .ZN(n7670) );
  OR2_X1 U5124 ( .A1(n7750), .A2(n7749), .ZN(n7752) );
  NAND2_X1 U5125 ( .A1(n7811), .A2(n5548), .ZN(n7881) );
  NAND2_X1 U5126 ( .A1(n7881), .A2(n7882), .ZN(n7880) );
  NAND2_X1 U5127 ( .A1(n7878), .A2(n5464), .ZN(n4497) );
  NAND2_X1 U5128 ( .A1(n4499), .A2(n5464), .ZN(n4498) );
  INV_X1 U5129 ( .A(n5462), .ZN(n4499) );
  NOR2_X1 U5130 ( .A1(n8021), .A2(n5069), .ZN(n8020) );
  XNOR2_X1 U5131 ( .A(n5506), .B(n5505), .ZN(n8633) );
  NAND2_X1 U5132 ( .A1(n8611), .A2(n5551), .ZN(n8628) );
  NAND2_X1 U5133 ( .A1(n8628), .A2(n8629), .ZN(n8627) );
  NOR2_X1 U5134 ( .A1(n8633), .A2(n8923), .ZN(n8632) );
  INV_X1 U5135 ( .A(n5506), .ZN(n5507) );
  XNOR2_X1 U5136 ( .A(n5471), .B(n8673), .ZN(n8670) );
  XNOR2_X1 U5137 ( .A(n5510), .B(n7405), .ZN(n8661) );
  NOR2_X1 U5138 ( .A1(n8661), .A2(n8917), .ZN(n8660) );
  NAND2_X1 U5139 ( .A1(n5300), .A2(n5299), .ZN(n5319) );
  AND2_X1 U5140 ( .A1(n8493), .A2(n8496), .ZN(n8803) );
  NAND2_X1 U5141 ( .A1(n8815), .A2(n8492), .ZN(n8804) );
  NAND2_X1 U5142 ( .A1(n4562), .A2(n4565), .ZN(n8817) );
  INV_X1 U5143 ( .A(n4566), .ZN(n4565) );
  OAI21_X1 U5144 ( .B1(n4567), .B2(n8824), .A(n8484), .ZN(n4566) );
  AOI21_X1 U5145 ( .B1(n4511), .B2(n4513), .A(n4333), .ZN(n4510) );
  NAND2_X1 U5146 ( .A1(n5159), .A2(n5158), .ZN(n5175) );
  INV_X1 U5147 ( .A(n5160), .ZN(n5159) );
  NAND2_X1 U5148 ( .A1(n4522), .A2(n4519), .ZN(n4515) );
  NAND2_X1 U5149 ( .A1(n8475), .A2(n5425), .ZN(n8930) );
  AND4_X1 U5150 ( .A1(n5076), .A2(n5075), .A3(n5074), .A4(n5073), .ZN(n8064)
         );
  NAND2_X1 U5151 ( .A1(n7547), .A2(n5016), .ZN(n4541) );
  OR2_X1 U5152 ( .A1(n8577), .A2(n7581), .ZN(n5016) );
  AND4_X2 U5153 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n7272)
         );
  OR2_X1 U5154 ( .A1(n8318), .A2(n4921), .ZN(n4922) );
  OR2_X1 U5155 ( .A1(n4960), .A2(n7262), .ZN(n4925) );
  XNOR2_X1 U5156 ( .A(n5967), .B(n8529), .ZN(n8330) );
  INV_X1 U5157 ( .A(n5951), .ZN(n8522) );
  AOI21_X1 U5158 ( .B1(n4575), .B2(n4573), .A(n4572), .ZN(n4571) );
  INV_X1 U5159 ( .A(n4575), .ZN(n4574) );
  INV_X1 U5160 ( .A(n8515), .ZN(n4572) );
  INV_X1 U5161 ( .A(n4578), .ZN(n4577) );
  OAI21_X1 U5162 ( .B1(n4581), .B2(n8507), .A(n8513), .ZN(n4578) );
  NOR2_X1 U5163 ( .A1(n8507), .A2(n4580), .ZN(n4579) );
  INV_X1 U5164 ( .A(n8381), .ZN(n4580) );
  INV_X1 U5165 ( .A(n8333), .ZN(n8732) );
  NOR2_X1 U5166 ( .A1(n8383), .A2(n4582), .ZN(n4581) );
  INV_X1 U5167 ( .A(n8756), .ZN(n8763) );
  NAND2_X1 U5168 ( .A1(n8506), .A2(n8748), .ZN(n8756) );
  NAND2_X1 U5169 ( .A1(n8772), .A2(n8381), .ZN(n4583) );
  INV_X1 U5170 ( .A(n8786), .ZN(n8789) );
  NAND2_X1 U5171 ( .A1(n8835), .A2(n8352), .ZN(n4567) );
  NAND2_X1 U5172 ( .A1(n5426), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U5173 ( .A1(n8836), .A2(n8835), .ZN(n8834) );
  OR2_X1 U5174 ( .A1(n9011), .A2(n8850), .ZN(n8845) );
  AND4_X1 U5175 ( .A1(n5144), .A2(n5143), .A3(n5142), .A4(n5141), .ZN(n8868)
         );
  NAND2_X1 U5176 ( .A1(n8845), .A2(n8471), .ZN(n8859) );
  NAND2_X1 U5177 ( .A1(n5424), .A2(n8475), .ZN(n4596) );
  INV_X1 U5178 ( .A(n7538), .ZN(n7530) );
  NOR2_X1 U5179 ( .A1(n5354), .A2(n4508), .ZN(n4804) );
  NAND2_X1 U5180 ( .A1(n4294), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U5181 ( .A1(n5386), .A2(n5380), .ZN(n5382) );
  INV_X1 U5182 ( .A(n8082), .ZN(n4742) );
  AOI21_X1 U5183 ( .B1(n4731), .B2(n4338), .A(n6447), .ZN(n4729) );
  AND2_X1 U5184 ( .A1(n6403), .A2(n4753), .ZN(n4747) );
  OR2_X1 U5185 ( .A1(n6411), .A2(n9115), .ZN(n4753) );
  INV_X1 U5186 ( .A(n8166), .ZN(n4358) );
  INV_X1 U5187 ( .A(n9115), .ZN(n4752) );
  NAND2_X1 U5188 ( .A1(n6411), .A2(n4751), .ZN(n4750) );
  AND2_X1 U5189 ( .A1(n9061), .A2(n6397), .ZN(n6396) );
  INV_X1 U5190 ( .A(n7503), .ZN(n6325) );
  AND3_X1 U5191 ( .A1(n6155), .A2(n6154), .A3(n6153), .ZN(n9053) );
  AND4_X1 U5192 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n7897)
         );
  AND4_X1 U5193 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n7726)
         );
  NAND2_X1 U5194 ( .A1(n5994), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5987) );
  NOR2_X1 U5195 ( .A1(n9190), .A2(n9189), .ZN(n9193) );
  AND2_X1 U5196 ( .A1(n9202), .A2(n9200), .ZN(n4492) );
  OR2_X1 U5197 ( .A1(n9193), .A2(n9192), .ZN(n9201) );
  XNOR2_X1 U5198 ( .A(n5718), .B(n5717), .ZN(n5804) );
  INV_X1 U5199 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U5200 ( .A1(n5716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U5201 ( .A1(n4548), .A2(n4546), .ZN(n9252) );
  AOI21_X1 U5202 ( .B1(n4549), .B2(n4551), .A(n4547), .ZN(n4546) );
  INV_X1 U5203 ( .A(n6635), .ZN(n4547) );
  NAND2_X1 U5204 ( .A1(n4545), .A2(n4549), .ZN(n9273) );
  AOI21_X1 U5205 ( .B1(n4451), .B2(n4450), .A(n4315), .ZN(n4449) );
  INV_X1 U5206 ( .A(n6184), .ZN(n4450) );
  NAND2_X1 U5207 ( .A1(n9303), .A2(n6244), .ZN(n9286) );
  AND2_X1 U5208 ( .A1(n9463), .A2(n9157), .ZN(n6165) );
  AND2_X1 U5209 ( .A1(n9339), .A2(n6622), .ZN(n4557) );
  INV_X1 U5210 ( .A(n9348), .ZN(n4556) );
  INV_X1 U5211 ( .A(n6622), .ZN(n4555) );
  NAND2_X1 U5212 ( .A1(n9350), .A2(n9349), .ZN(n9348) );
  AOI21_X1 U5213 ( .B1(n4461), .B2(n4459), .A(n4310), .ZN(n4458) );
  INV_X1 U5214 ( .A(n6131), .ZN(n4459) );
  AND2_X1 U5215 ( .A1(n6616), .A2(n6615), .ZN(n9367) );
  OR2_X1 U5216 ( .A1(n9426), .A2(n9162), .ZN(n6121) );
  OR2_X1 U5217 ( .A1(n8139), .A2(n9426), .ZN(n9423) );
  AND2_X1 U5218 ( .A1(n4471), .A2(n8117), .ZN(n4470) );
  INV_X1 U5219 ( .A(n6097), .ZN(n4471) );
  OR2_X1 U5220 ( .A1(n9033), .A2(n9164), .ZN(n6088) );
  OAI211_X1 U5221 ( .C1(n4437), .C2(n4435), .A(n4288), .B(n4433), .ZN(n4439)
         );
  NAND2_X1 U5222 ( .A1(n4437), .A2(n4778), .ZN(n4436) );
  NAND2_X1 U5223 ( .A1(n9877), .A2(n9881), .ZN(n6001) );
  NAND2_X1 U5224 ( .A1(n5739), .A2(n5738), .ZN(n9293) );
  NAND2_X1 U5225 ( .A1(n6905), .A2(n5756), .ZN(n5669) );
  NAND2_X1 U5226 ( .A1(n4736), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U5227 ( .A1(n4472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  AND2_X1 U5228 ( .A1(n5605), .A2(n4474), .ZN(n4473) );
  INV_X1 U5229 ( .A(n4734), .ZN(n4474) );
  NAND2_X1 U5230 ( .A1(n4627), .A2(n5333), .ZN(n5339) );
  NAND2_X1 U5231 ( .A1(n5332), .A2(n5331), .ZN(n4627) );
  XNOR2_X1 U5232 ( .A(n5332), .B(n5331), .ZN(n8039) );
  XNOR2_X1 U5233 ( .A(n5310), .B(n5309), .ZN(n7966) );
  XNOR2_X1 U5234 ( .A(n5250), .B(n5249), .ZN(n7771) );
  NAND2_X1 U5235 ( .A1(n4660), .A2(n5232), .ZN(n5250) );
  OAI21_X1 U5236 ( .B1(n5150), .B2(n4293), .A(n4636), .ZN(n5203) );
  NAND2_X1 U5237 ( .A1(n5712), .A2(n5711), .ZN(n5716) );
  NAND2_X1 U5238 ( .A1(n4639), .A2(n5165), .ZN(n5183) );
  NOR2_X1 U5239 ( .A1(n5600), .A2(n5635), .ZN(n5686) );
  INV_X1 U5240 ( .A(n8575), .ZN(n7517) );
  NAND2_X1 U5241 ( .A1(n5093), .A2(n5092), .ZN(n8468) );
  XNOR2_X1 U5242 ( .A(n5899), .B(n5901), .ZN(n8204) );
  AND4_X1 U5243 ( .A1(n4975), .A2(n4974), .A3(n4973), .A4(n4972), .ZN(n8410)
         );
  AND2_X1 U5244 ( .A1(n5213), .A2(n5212), .ZN(n8568) );
  OR2_X1 U5245 ( .A1(n5907), .A2(n8567), .ZN(n5908) );
  AND2_X1 U5246 ( .A1(n4887), .A2(n4886), .ZN(n8449) );
  INV_X1 U5247 ( .A(n8964), .ZN(n8267) );
  NAND2_X1 U5248 ( .A1(n4720), .A2(n5836), .ZN(n7306) );
  AND2_X1 U5249 ( .A1(n5264), .A2(n5263), .ZN(n8743) );
  INV_X1 U5250 ( .A(n8064), .ZN(n8933) );
  INV_X1 U5251 ( .A(n8134), .ZN(n8571) );
  NAND4_X1 U5252 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n4989), .ZN(n8578)
         );
  OR2_X1 U5253 ( .A1(n4952), .A2(n4986), .ZN(n4991) );
  OR2_X1 U5254 ( .A1(n5053), .A2(n7413), .ZN(n4989) );
  NAND2_X1 U5255 ( .A1(n7063), .A2(n4381), .ZN(n7131) );
  OR2_X1 U5256 ( .A1(n5537), .A2(n5538), .ZN(n4381) );
  NAND2_X1 U5257 ( .A1(n7131), .A2(n7130), .ZN(n7129) );
  NOR2_X1 U5258 ( .A1(n7218), .A2(n7219), .ZN(n7217) );
  OR2_X1 U5259 ( .A1(n8012), .A2(n5068), .ZN(n4679) );
  NOR2_X1 U5260 ( .A1(n8670), .A2(n8671), .ZN(n8669) );
  NOR2_X1 U5261 ( .A1(n8686), .A2(n7405), .ZN(n4505) );
  AOI21_X1 U5262 ( .B1(n8692), .B2(n8691), .A(n4385), .ZN(n4384) );
  NAND2_X1 U5263 ( .A1(n4686), .A2(n4386), .ZN(n4385) );
  INV_X1 U5264 ( .A(n8696), .ZN(n4386) );
  OAI21_X1 U5265 ( .B1(n5375), .B2(n8862), .A(n5374), .ZN(n8706) );
  NOR2_X1 U5266 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NOR2_X1 U5267 ( .A1(n8736), .A2(n8865), .ZN(n5372) );
  NAND2_X1 U5268 ( .A1(n5190), .A2(n5480), .ZN(n4597) );
  NAND2_X1 U5269 ( .A1(n4926), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4598) );
  INV_X1 U5270 ( .A(n8945), .ZN(n8884) );
  NAND2_X1 U5271 ( .A1(n5967), .A2(n8915), .ZN(n5968) );
  INV_X1 U5272 ( .A(n5579), .ZN(n8373) );
  AND2_X1 U5273 ( .A1(n9036), .A2(n9037), .ZN(n9038) );
  OAI21_X1 U5274 ( .B1(n9243), .B2(n9784), .A(n4483), .ZN(n4482) );
  OR2_X1 U5275 ( .A1(n9241), .A2(n9242), .ZN(n4483) );
  OAI211_X1 U5276 ( .C1(n9240), .C2(n9784), .A(n9239), .B(n9798), .ZN(n4485)
         );
  NOR2_X1 U5277 ( .A1(n5719), .A2(n6513), .ZN(n6514) );
  OR2_X1 U5278 ( .A1(n9016), .A2(n5611), .ZN(n6515) );
  XNOR2_X1 U5279 ( .A(n4465), .B(n6669), .ZN(n8183) );
  NAND2_X1 U5280 ( .A1(n9259), .A2(n6211), .ZN(n4465) );
  NAND2_X1 U5281 ( .A1(n9261), .A2(n6210), .ZN(n6211) );
  OR2_X1 U5282 ( .A1(n5643), .A2(n6856), .ZN(n5641) );
  INV_X1 U5283 ( .A(n6216), .ZN(n8178) );
  NOR2_X1 U5284 ( .A1(n8184), .A2(n6518), .ZN(n6526) );
  NAND2_X1 U5285 ( .A1(n8326), .A2(n5756), .ZN(n5758) );
  OR2_X1 U5286 ( .A1(n9435), .A2(n9998), .ZN(n5815) );
  OAI21_X1 U5287 ( .B1(n8183), .B2(n9941), .A(n4464), .ZN(n6816) );
  AND2_X1 U5288 ( .A1(n8174), .A2(n8175), .ZN(n4464) );
  NAND2_X1 U5289 ( .A1(n4393), .A2(n8462), .ZN(n8466) );
  NAND2_X1 U5290 ( .A1(n8461), .A2(n4394), .ZN(n4393) );
  NAND2_X1 U5291 ( .A1(n4402), .A2(n8483), .ZN(n8491) );
  OR2_X1 U5292 ( .A1(n6678), .A2(n6649), .ZN(n4420) );
  NAND2_X1 U5293 ( .A1(n4425), .A2(n6623), .ZN(n4421) );
  NAND2_X1 U5294 ( .A1(n4424), .A2(n4423), .ZN(n4422) );
  OAI21_X1 U5295 ( .B1(n4392), .B2(n8518), .A(n4314), .ZN(n4391) );
  AOI21_X1 U5296 ( .B1(n8510), .B2(n8511), .A(n8509), .ZN(n4392) );
  INV_X1 U5297 ( .A(n5248), .ZN(n4657) );
  NAND2_X1 U5298 ( .A1(n4536), .A2(n4533), .ZN(n4532) );
  INV_X1 U5299 ( .A(n4537), .ZN(n4533) );
  NOR2_X1 U5300 ( .A1(n4534), .A2(n4528), .ZN(n4527) );
  INV_X1 U5301 ( .A(n4777), .ZN(n4528) );
  OR2_X1 U5302 ( .A1(n7840), .A2(n4535), .ZN(n4534) );
  INV_X1 U5303 ( .A(n4536), .ZN(n4535) );
  NAND2_X1 U5304 ( .A1(n8580), .A2(n7320), .ZN(n8414) );
  AND2_X1 U5305 ( .A1(n9315), .A2(n9155), .ZN(n6632) );
  NAND2_X1 U5306 ( .A1(n6616), .A2(n9366), .ZN(n6697) );
  NAND2_X1 U5307 ( .A1(n5593), .A2(n5333), .ZN(n4626) );
  INV_X1 U5308 ( .A(n4624), .ZN(n4623) );
  OAI21_X1 U5309 ( .B1(n4628), .B2(n4625), .A(n4339), .ZN(n4624) );
  INV_X1 U5310 ( .A(n4629), .ZN(n4628) );
  OAI21_X1 U5311 ( .B1(n5331), .B2(n4630), .A(n5338), .ZN(n4629) );
  INV_X1 U5312 ( .A(n5273), .ZN(n4652) );
  OAI21_X1 U5313 ( .B1(n4658), .B2(n4657), .A(n5271), .ZN(n4656) );
  NOR2_X1 U5314 ( .A1(n4652), .A2(n4657), .ZN(n4651) );
  INV_X1 U5315 ( .A(n5233), .ZN(n4653) );
  NOR2_X1 U5316 ( .A1(n4637), .A2(n5202), .ZN(n4631) );
  INV_X1 U5317 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4818) );
  INV_X1 U5318 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4819) );
  OAI21_X1 U5319 ( .B1(n5836), .B2(n4719), .A(n7411), .ZN(n4717) );
  AND2_X1 U5320 ( .A1(n8543), .A2(n4666), .ZN(n4665) );
  NOR2_X1 U5321 ( .A1(n8532), .A2(n8540), .ZN(n4666) );
  AOI21_X1 U5322 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n7045), .A(n7033), .ZN(
        n5483) );
  NOR2_X1 U5323 ( .A1(n5483), .A2(n7084), .ZN(n5485) );
  AND2_X1 U5324 ( .A1(n7738), .A2(n5460), .ZN(n5461) );
  NAND3_X1 U5325 ( .A1(n4675), .A2(n4344), .A3(n4674), .ZN(n5506) );
  NAND2_X1 U5326 ( .A1(n4671), .A2(n4670), .ZN(n5510) );
  AOI21_X1 U5327 ( .B1(n5508), .B2(n4673), .A(n4672), .ZN(n4671) );
  INV_X1 U5328 ( .A(n5509), .ZN(n4672) );
  NOR2_X1 U5329 ( .A1(n8824), .A2(n4564), .ZN(n4563) );
  INV_X1 U5330 ( .A(n4569), .ZN(n4564) );
  INV_X1 U5331 ( .A(n4770), .ZN(n4513) );
  NAND2_X1 U5332 ( .A1(n7696), .A2(n7825), .ZN(n4537) );
  NAND2_X1 U5333 ( .A1(n7702), .A2(n8574), .ZN(n4536) );
  INV_X1 U5334 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7123) );
  NOR2_X1 U5335 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n4987) );
  AOI21_X1 U5336 ( .B1(n7200), .B2(n7201), .A(n4942), .ZN(n7270) );
  AND2_X1 U5337 ( .A1(n4577), .A2(n8516), .ZN(n4575) );
  INV_X1 U5338 ( .A(n4579), .ZN(n4573) );
  AOI21_X1 U5339 ( .B1(n4590), .B2(n8456), .A(n4588), .ZN(n4587) );
  INV_X1 U5340 ( .A(n8463), .ZN(n4588) );
  XNOR2_X1 U5341 ( .A(n7269), .B(n8581), .ZN(n8399) );
  NAND2_X1 U5342 ( .A1(n4763), .A2(n4725), .ZN(n4724) );
  INV_X1 U5343 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4869) );
  INV_X1 U5344 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4375) );
  INV_X1 U5345 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4798) );
  INV_X1 U5346 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4561) );
  INV_X1 U5347 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4794) );
  AND2_X1 U5348 ( .A1(n4795), .A2(n5128), .ZN(n4377) );
  NOR2_X1 U5349 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4795) );
  NOR2_X1 U5350 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5128) );
  NAND2_X1 U5351 ( .A1(n5066), .A2(n4883), .ZN(n5130) );
  INV_X1 U5352 ( .A(n5065), .ZN(n5066) );
  INV_X1 U5353 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U5354 ( .A1(n4352), .A2(n4350), .ZN(n4754) );
  AND2_X1 U5355 ( .A1(n6134), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6141) );
  OR2_X1 U5356 ( .A1(n7583), .A2(n6335), .ZN(n4354) );
  OR2_X1 U5357 ( .A1(n6391), .A2(n9071), .ZN(n6397) );
  AND2_X1 U5358 ( .A1(n6062), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6073) );
  INV_X1 U5359 ( .A(n9924), .ZN(n4370) );
  OR2_X1 U5360 ( .A1(n9315), .A2(n6796), .ZN(n6266) );
  NAND2_X1 U5361 ( .A1(n4746), .A2(n4745), .ZN(n4744) );
  INV_X1 U5362 ( .A(n4785), .ZN(n4745) );
  NAND2_X1 U5363 ( .A1(n4291), .A2(n9027), .ZN(n4746) );
  OAI22_X1 U5364 ( .A1(n4744), .A2(n4739), .B1(n9027), .B2(n4291), .ZN(n4738)
         );
  INV_X1 U5365 ( .A(n8083), .ZN(n4739) );
  AND2_X1 U5366 ( .A1(n6760), .A2(n6755), .ZN(n6740) );
  OR2_X1 U5367 ( .A1(n9261), .A2(n7251), .ZN(n6675) );
  INV_X1 U5368 ( .A(n6634), .ZN(n4551) );
  NOR2_X1 U5369 ( .A1(n9293), .A2(n9454), .ZN(n4617) );
  INV_X1 U5370 ( .A(n6632), .ZN(n9283) );
  INV_X1 U5371 ( .A(n8001), .ZN(n4467) );
  NAND2_X1 U5372 ( .A1(n4434), .A2(n4442), .ZN(n4433) );
  NAND2_X1 U5373 ( .A1(n7678), .A2(n6711), .ZN(n7723) );
  OAI21_X1 U5374 ( .B1(n6232), .B2(n6659), .A(n6661), .ZN(n6707) );
  AND2_X1 U5375 ( .A1(n6550), .A2(n7555), .ZN(n7557) );
  NAND2_X1 U5376 ( .A1(n9325), .A2(n9315), .ZN(n9309) );
  NAND2_X1 U5377 ( .A1(n9399), .A2(n4621), .ZN(n9372) );
  AND2_X1 U5378 ( .A1(n9399), .A2(n9657), .ZN(n9389) );
  AND2_X1 U5379 ( .A1(n5607), .A2(n5606), .ZN(n4755) );
  INV_X1 U5380 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5606) );
  INV_X1 U5381 ( .A(n5165), .ZN(n4638) );
  NOR2_X1 U5382 ( .A1(n5166), .A2(n4641), .ZN(n4640) );
  INV_X1 U5383 ( .A(n5149), .ZN(n4641) );
  INV_X1 U5384 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U5385 ( .A1(n5078), .A2(n5077), .ZN(n4648) );
  XNOR2_X1 U5386 ( .A(n5060), .B(SI_12_), .ZN(n5062) );
  NAND2_X1 U5387 ( .A1(n4866), .A2(n4865), .ZN(n5044) );
  INV_X1 U5388 ( .A(n4647), .ZN(n4646) );
  INV_X1 U5389 ( .A(n4855), .ZN(n4645) );
  INV_X1 U5390 ( .A(n4860), .ZN(n4644) );
  XNOR2_X1 U5391 ( .A(n4850), .B(SI_7_), .ZN(n4906) );
  OAI21_X1 U5392 ( .B1(n6853), .B2(n4843), .A(n4842), .ZN(n4844) );
  NAND2_X1 U5393 ( .A1(n6853), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4842) );
  OAI21_X1 U5394 ( .B1(n5611), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n4406), .ZN(
        n4833) );
  NAND2_X1 U5395 ( .A1(n5611), .A2(n4407), .ZN(n4406) );
  OAI21_X1 U5396 ( .B1(n4828), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4827), .ZN(
        n4829) );
  NAND2_X1 U5397 ( .A1(n4828), .A2(n6868), .ZN(n4827) );
  AND2_X1 U5398 ( .A1(n5857), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U5399 ( .A1(n7653), .A2(n5855), .ZN(n4723) );
  NAND2_X1 U5400 ( .A1(n7654), .A2(n5855), .ZN(n7867) );
  NAND2_X1 U5401 ( .A1(n8290), .A2(n8291), .ZN(n8289) );
  OR2_X1 U5402 ( .A1(n5357), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5359) );
  OR2_X1 U5403 ( .A1(n7022), .A2(n7262), .ZN(n7020) );
  AND2_X1 U5404 ( .A1(n4684), .A2(n4682), .ZN(n7034) );
  NOR2_X1 U5405 ( .A1(n7034), .A2(n7035), .ZN(n7033) );
  NOR2_X1 U5406 ( .A1(n5484), .A2(n5485), .ZN(n7077) );
  AND2_X1 U5407 ( .A1(n5483), .A2(n7084), .ZN(n5484) );
  OR2_X1 U5408 ( .A1(n5444), .A2(n6859), .ZN(n5445) );
  NAND2_X1 U5409 ( .A1(n5444), .A2(n6859), .ZN(n7052) );
  INV_X1 U5410 ( .A(n7122), .ZN(n7223) );
  OAI21_X1 U5411 ( .B1(n7223), .B2(n7221), .A(n7222), .ZN(n7225) );
  OR2_X1 U5412 ( .A1(n8602), .A2(n5454), .ZN(n5456) );
  NAND2_X1 U5413 ( .A1(n7664), .A2(n5546), .ZN(n7744) );
  NAND2_X1 U5414 ( .A1(n7744), .A2(n7745), .ZN(n7743) );
  NAND2_X1 U5415 ( .A1(n7752), .A2(n5495), .ZN(n5497) );
  NAND2_X1 U5416 ( .A1(n7812), .A2(n7813), .ZN(n7811) );
  NAND2_X1 U5417 ( .A1(n7880), .A2(n5549), .ZN(n8015) );
  NAND2_X1 U5418 ( .A1(n8612), .A2(n8613), .ZN(n8611) );
  NAND2_X1 U5419 ( .A1(n8627), .A2(n5552), .ZN(n8646) );
  AND2_X1 U5420 ( .A1(n8640), .A2(n5470), .ZN(n5471) );
  OAI21_X1 U5421 ( .B1(n8680), .B2(n4307), .A(n8697), .ZN(n4686) );
  INV_X1 U5422 ( .A(n8683), .ZN(n8684) );
  NOR2_X1 U5423 ( .A1(n8682), .A2(n8681), .ZN(n8680) );
  NAND2_X1 U5424 ( .A1(n5556), .A2(n5555), .ZN(n8683) );
  AND2_X1 U5425 ( .A1(n5369), .A2(n5368), .ZN(n8529) );
  NAND2_X1 U5426 ( .A1(n8531), .A2(n8376), .ZN(n8331) );
  INV_X1 U5427 ( .A(n8330), .ZN(n5958) );
  NAND2_X1 U5428 ( .A1(n5954), .A2(n4542), .ZN(n5352) );
  NOR2_X1 U5429 ( .A1(n4544), .A2(n4543), .ZN(n4542) );
  INV_X1 U5430 ( .A(n5947), .ZN(n4543) );
  INV_X1 U5431 ( .A(n5948), .ZN(n4544) );
  NAND2_X1 U5432 ( .A1(n8524), .A2(n8523), .ZN(n5951) );
  NOR2_X1 U5433 ( .A1(n8529), .A2(n8867), .ZN(n5373) );
  OR2_X1 U5434 ( .A1(n5319), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5345) );
  OR2_X1 U5435 ( .A1(n5258), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5282) );
  OR2_X1 U5436 ( .A1(n5241), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U5437 ( .A1(n5223), .A2(n8234), .ZN(n5241) );
  INV_X1 U5438 ( .A(n5224), .ZN(n5223) );
  NAND2_X1 U5439 ( .A1(n5194), .A2(n5193), .ZN(n5207) );
  INV_X1 U5440 ( .A(n5195), .ZN(n5194) );
  NAND2_X1 U5441 ( .A1(n5111), .A2(n5110), .ZN(n5139) );
  OR2_X1 U5442 ( .A1(n5096), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U5443 ( .A1(n5071), .A2(n5070), .ZN(n5096) );
  NOR2_X1 U5444 ( .A1(n5052), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5071) );
  OR2_X1 U5445 ( .A1(n5050), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U5446 ( .A1(n4529), .A2(n4536), .ZN(n7844) );
  NAND2_X1 U5447 ( .A1(n7692), .A2(n4537), .ZN(n4529) );
  NAND2_X1 U5448 ( .A1(n5021), .A2(n5020), .ZN(n5038) );
  AND2_X1 U5449 ( .A1(n8421), .A2(n8446), .ZN(n8345) );
  NAND2_X1 U5450 ( .A1(n5017), .A2(n4777), .ZN(n7692) );
  NOR2_X1 U5451 ( .A1(n5003), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n4915) );
  NOR2_X1 U5452 ( .A1(n8411), .A2(n4585), .ZN(n4584) );
  INV_X1 U5453 ( .A(n4782), .ZN(n4585) );
  NAND2_X1 U5454 ( .A1(n4987), .A2(n7123), .ZN(n5001) );
  OR2_X1 U5455 ( .A1(n5001), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U5456 ( .A1(n7421), .A2(n8339), .ZN(n4586) );
  OAI21_X1 U5457 ( .B1(n7270), .B2(n8399), .A(n4958), .ZN(n7321) );
  OR2_X1 U5458 ( .A1(n7269), .A2(n8581), .ZN(n4958) );
  AND4_X1 U5459 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n7271)
         );
  NAND2_X1 U5460 ( .A1(n5417), .A2(n7257), .ZN(n8391) );
  AND2_X1 U5461 ( .A1(n5351), .A2(n5350), .ZN(n8721) );
  AND2_X1 U5462 ( .A1(n8718), .A2(n8717), .ZN(n8720) );
  AND2_X1 U5463 ( .A1(n8519), .A2(n8520), .ZN(n8719) );
  INV_X1 U5464 ( .A(n8567), .ZN(n8736) );
  AND2_X1 U5465 ( .A1(n8762), .A2(n8760), .ZN(n5268) );
  AND2_X1 U5466 ( .A1(n8761), .A2(n8760), .ZN(n8778) );
  AND2_X1 U5467 ( .A1(n8775), .A2(n8774), .ZN(n8791) );
  NAND2_X1 U5468 ( .A1(n9011), .A2(n5118), .ZN(n5119) );
  AND2_X1 U5469 ( .A1(n4984), .A2(n4983), .ZN(n7424) );
  AND2_X1 U5470 ( .A1(n7848), .A2(n7950), .ZN(n8940) );
  NAND2_X1 U5471 ( .A1(n4302), .A2(n4378), .ZN(n4379) );
  OAI22_X1 U5472 ( .A1(n4928), .A2(n4946), .B1(P2_IR_REG_2__SCAN_IN), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U5473 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4946) );
  NAND2_X1 U5474 ( .A1(n5611), .A2(n4822), .ZN(n4941) );
  OR2_X1 U5475 ( .A1(n6151), .A2(n6150), .ZN(n6157) );
  OR2_X1 U5476 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  NAND2_X1 U5477 ( .A1(n6274), .A2(n4758), .ZN(n7091) );
  INV_X1 U5478 ( .A(n6442), .ZN(n9037) );
  AND2_X1 U5479 ( .A1(n8030), .A2(n6367), .ZN(n7957) );
  XNOR2_X1 U5480 ( .A(n6271), .B(n6794), .ZN(n6281) );
  AOI22_X1 U5481 ( .A1(n6268), .A2(n6451), .B1(n4278), .B2(n6825), .ZN(n6282)
         );
  OR2_X1 U5482 ( .A1(n6115), .A2(n6114), .ZN(n6123) );
  NAND2_X1 U5483 ( .A1(n7487), .A2(n6317), .ZN(n6320) );
  OAI21_X1 U5484 ( .B1(n8028), .B2(n4371), .A(n4737), .ZN(n6393) );
  NAND2_X1 U5485 ( .A1(n4740), .A2(n6377), .ZN(n4371) );
  INV_X1 U5486 ( .A(n4738), .ZN(n4737) );
  INV_X1 U5487 ( .A(n4744), .ZN(n4740) );
  OR2_X1 U5488 ( .A1(n6090), .A2(n7985), .ZN(n6098) );
  OR2_X1 U5489 ( .A1(n6082), .A2(n6081), .ZN(n6090) );
  NAND2_X1 U5490 ( .A1(n4415), .A2(n4417), .ZN(n4411) );
  AND3_X1 U5491 ( .A1(n6147), .A2(n6146), .A3(n6145), .ZN(n9106) );
  AND4_X1 U5492 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n8168)
         );
  AND4_X1 U5493 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n9118)
         );
  AND4_X1 U5494 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(n7997)
         );
  AND4_X1 U5495 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n7960)
         );
  AND4_X1 U5496 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n7361)
         );
  NAND2_X1 U5497 ( .A1(n5994), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6005) );
  NOR2_X1 U5498 ( .A1(n7157), .A2(n4478), .ZN(n7159) );
  NOR2_X1 U5499 ( .A1(n4480), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U5500 ( .A1(n7159), .A2(n7160), .ZN(n7288) );
  NOR2_X1 U5501 ( .A1(n7979), .A2(n4486), .ZN(n9188) );
  AND2_X1 U5502 ( .A1(n7980), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U5503 ( .A1(n4491), .A2(n4490), .ZN(n9225) );
  AOI21_X1 U5504 ( .B1(n4492), .B2(n9192), .A(n4347), .ZN(n4490) );
  OR2_X1 U5505 ( .A1(n6216), .A2(n6256), .ZN(n6504) );
  INV_X1 U5506 ( .A(n4445), .ZN(n9258) );
  NAND2_X1 U5507 ( .A1(n4451), .A2(n6668), .ZN(n4448) );
  INV_X1 U5508 ( .A(n4447), .ZN(n4446) );
  NAND2_X1 U5509 ( .A1(n6642), .A2(n6675), .ZN(n9257) );
  NAND2_X1 U5510 ( .A1(n9325), .A2(n4615), .ZN(n9268) );
  OR2_X1 U5511 ( .A1(n6157), .A2(n9591), .ZN(n6176) );
  AOI22_X1 U5512 ( .A1(n9350), .A2(n4297), .B1(n6679), .B2(n4554), .ZN(n4553)
         );
  INV_X1 U5513 ( .A(n4557), .ZN(n4554) );
  NAND2_X1 U5514 ( .A1(n9399), .A2(n4308), .ZN(n9336) );
  NAND2_X1 U5515 ( .A1(n9399), .A2(n4620), .ZN(n9354) );
  OAI21_X1 U5516 ( .B1(n9398), .B2(n4457), .A(n4455), .ZN(n4454) );
  NAND2_X1 U5517 ( .A1(n6149), .A2(n4461), .ZN(n4457) );
  AOI21_X1 U5518 ( .B1(n4456), .B2(n6149), .A(n6148), .ZN(n4455) );
  NOR2_X1 U5519 ( .A1(n9423), .A2(n9483), .ZN(n9399) );
  NAND2_X1 U5520 ( .A1(n4558), .A2(n6598), .ZN(n9413) );
  NAND2_X1 U5521 ( .A1(n7776), .A2(n4559), .ZN(n7992) );
  AND2_X1 U5522 ( .A1(n6663), .A2(n6716), .ZN(n4559) );
  OR2_X1 U5523 ( .A1(n8089), .A2(n9165), .ZN(n6080) );
  NOR2_X1 U5524 ( .A1(n4610), .A2(n9033), .ZN(n4609) );
  INV_X1 U5525 ( .A(n4612), .ZN(n4610) );
  NAND2_X1 U5526 ( .A1(n4611), .A2(n4612), .ZN(n7903) );
  OR2_X1 U5527 ( .A1(n6050), .A2(n6049), .ZN(n6056) );
  NOR2_X1 U5528 ( .A1(n4606), .A2(n9976), .ZN(n4605) );
  AND2_X1 U5529 ( .A1(n9818), .A2(n6556), .ZN(n7558) );
  NOR2_X1 U5530 ( .A1(n7475), .A2(n9845), .ZN(n9846) );
  INV_X1 U5531 ( .A(n7557), .ZN(n9838) );
  INV_X1 U5532 ( .A(n6658), .ZN(n7474) );
  NAND2_X1 U5533 ( .A1(n4600), .A2(n4599), .ZN(n9862) );
  AND2_X1 U5534 ( .A1(n7485), .A2(n9945), .ZN(n4599) );
  INV_X1 U5535 ( .A(n4601), .ZN(n4600) );
  NOR2_X1 U5536 ( .A1(n4601), .A2(n9937), .ZN(n9863) );
  NAND2_X1 U5537 ( .A1(n4602), .A2(n9930), .ZN(n9872) );
  OAI21_X1 U5538 ( .B1(n9892), .B2(n9891), .A(n5992), .ZN(n9877) );
  INV_X1 U5539 ( .A(n6669), .ZN(n6245) );
  NAND2_X1 U5540 ( .A1(n5615), .A2(n5614), .ZN(n6199) );
  NAND2_X1 U5541 ( .A1(n5709), .A2(n5708), .ZN(n9624) );
  NAND2_X1 U5542 ( .A1(n5706), .A2(n5705), .ZN(n6104) );
  INV_X1 U5543 ( .A(n7687), .ZN(n5674) );
  XNOR2_X1 U5544 ( .A(n5742), .B(n5741), .ZN(n5955) );
  NAND2_X1 U5545 ( .A1(n5594), .A2(n5740), .ZN(n5742) );
  NAND2_X1 U5546 ( .A1(n4654), .A2(n5248), .ZN(n5272) );
  NAND2_X1 U5547 ( .A1(n4660), .A2(n4658), .ZN(n4654) );
  NAND2_X1 U5548 ( .A1(n5761), .A2(n5760), .ZN(n5801) );
  NAND2_X1 U5549 ( .A1(n5710), .A2(n4367), .ZN(n4366) );
  INV_X1 U5550 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5710) );
  INV_X1 U5551 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4367) );
  XNOR2_X1 U5552 ( .A(n4428), .B(n5103), .ZN(n7195) );
  NAND2_X1 U5553 ( .A1(n4648), .A2(n5081), .ZN(n4428) );
  OAI21_X1 U5554 ( .B1(n4896), .B2(n4895), .A(n4855), .ZN(n4408) );
  NAND2_X1 U5555 ( .A1(n4841), .A2(n4840), .ZN(n4979) );
  INV_X1 U5556 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5598) );
  AND2_X1 U5557 ( .A1(n5626), .A2(n5631), .ZN(n6932) );
  NAND2_X1 U5558 ( .A1(n7576), .A2(n4728), .ZN(n7511) );
  NAND2_X1 U5559 ( .A1(n4715), .A2(n5870), .ZN(n8061) );
  NAND2_X1 U5560 ( .A1(n8289), .A2(n5886), .ZN(n8214) );
  NOR2_X1 U5561 ( .A1(n8312), .A2(n8223), .ZN(n4695) );
  NAND2_X1 U5562 ( .A1(n4322), .A2(n5916), .ZN(n4694) );
  NAND2_X1 U5563 ( .A1(n8226), .A2(n4701), .ZN(n4700) );
  INV_X1 U5564 ( .A(n5910), .ZN(n4701) );
  AOI21_X1 U5565 ( .B1(n4728), .B2(n7578), .A(n4316), .ZN(n4726) );
  INV_X1 U5566 ( .A(n4728), .ZN(n4727) );
  INV_X1 U5567 ( .A(n4703), .ZN(n4702) );
  OAI21_X1 U5568 ( .B1(n4704), .B2(n4708), .A(n5890), .ZN(n4703) );
  AND2_X1 U5569 ( .A1(n5288), .A2(n5287), .ZN(n8735) );
  NAND2_X1 U5570 ( .A1(n5298), .A2(n5297), .ZN(n8246) );
  AND3_X1 U5571 ( .A1(n5164), .A2(n5163), .A3(n5162), .ZN(n8851) );
  OR2_X1 U5572 ( .A1(n7652), .A2(n7653), .ZN(n7654) );
  OAI21_X1 U5573 ( .B1(n8290), .B2(n4713), .A(n4709), .ZN(n8271) );
  NAND2_X1 U5574 ( .A1(n5206), .A2(n5205), .ZN(n8275) );
  INV_X1 U5575 ( .A(n8576), .ZN(n7637) );
  NAND2_X1 U5576 ( .A1(n5015), .A2(n5014), .ZN(n7581) );
  NAND2_X1 U5578 ( .A1(n4593), .A2(n4592), .ZN(n8374) );
  NAND2_X1 U5579 ( .A1(n8372), .A2(n8390), .ZN(n4592) );
  NAND2_X1 U5580 ( .A1(n4595), .A2(n4594), .ZN(n4593) );
  NAND2_X1 U5581 ( .A1(n8552), .A2(n8550), .ZN(n8551) );
  OAI211_X1 U5582 ( .C1(n4401), .C2(n8546), .A(n4398), .B(n8548), .ZN(n8552)
         );
  INV_X1 U5583 ( .A(n8721), .ZN(n8566) );
  AND2_X1 U5584 ( .A1(n5308), .A2(n5307), .ZN(n8744) );
  NAND4_X1 U5585 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), .ZN(n8575)
         );
  NAND4_X1 U5586 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n8577)
         );
  OR2_X1 U5587 ( .A1(n4952), .A2(n7552), .ZN(n5006) );
  OR2_X1 U5588 ( .A1(n4960), .A2(n5451), .ZN(n5005) );
  OR2_X1 U5589 ( .A1(n5053), .A2(n10018), .ZN(n5004) );
  INV_X1 U5590 ( .A(n8410), .ZN(n8579) );
  INV_X1 U5591 ( .A(n7271), .ZN(n8580) );
  INV_X1 U5592 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6959) );
  XNOR2_X1 U5593 ( .A(n6952), .B(P2_IR_REG_0__SCAN_IN), .ZN(n6953) );
  NOR2_X1 U5594 ( .A1(n5481), .A2(n4684), .ZN(n7019) );
  INV_X1 U5595 ( .A(n4685), .ZN(n4683) );
  NAND2_X1 U5596 ( .A1(n7015), .A2(n4382), .ZN(n7042) );
  OR2_X1 U5597 ( .A1(n5532), .A2(n5480), .ZN(n4382) );
  NAND2_X1 U5598 ( .A1(n7042), .A2(n7041), .ZN(n7040) );
  NAND2_X1 U5599 ( .A1(n4494), .A2(n5450), .ZN(n7120) );
  NAND2_X1 U5600 ( .A1(n4687), .A2(n4690), .ZN(n7117) );
  NAND2_X1 U5601 ( .A1(n7129), .A2(n4380), .ZN(n7218) );
  OR2_X1 U5602 ( .A1(n5540), .A2(n4495), .ZN(n4380) );
  NAND2_X1 U5603 ( .A1(n5489), .A2(n8592), .ZN(n7397) );
  NAND2_X1 U5604 ( .A1(n4348), .A2(n8592), .ZN(n8594) );
  NAND2_X1 U5605 ( .A1(n8597), .A2(n4501), .ZN(n7390) );
  NOR2_X1 U5606 ( .A1(n8593), .A2(n4913), .ZN(n4681) );
  NOR2_X1 U5607 ( .A1(n7817), .A2(n5462), .ZN(n7879) );
  NOR2_X1 U5608 ( .A1(n8020), .A2(n5466), .ZN(n8610) );
  NAND2_X1 U5609 ( .A1(n4675), .A2(n4674), .ZN(n8617) );
  OR2_X1 U5610 ( .A1(n8643), .A2(n8642), .ZN(n8640) );
  OR2_X1 U5611 ( .A1(n8652), .A2(n8651), .ZN(n8654) );
  NOR2_X1 U5612 ( .A1(n8632), .A2(n5508), .ZN(n8652) );
  NAND2_X1 U5613 ( .A1(n5342), .A2(n5341), .ZN(n8711) );
  NAND2_X1 U5614 ( .A1(n5192), .A2(n5191), .ZN(n8909) );
  NAND2_X1 U5615 ( .A1(n5174), .A2(n5173), .ZN(n8914) );
  INV_X1 U5616 ( .A(n8468), .ZN(n9739) );
  NAND2_X1 U5617 ( .A1(n4515), .A2(n4518), .ZN(n8931) );
  AOI21_X1 U5618 ( .B1(n7138), .B2(n8325), .A(n5067), .ZN(n8877) );
  NAND2_X1 U5619 ( .A1(n8045), .A2(n8455), .ZN(n8135) );
  AND2_X1 U5620 ( .A1(n4521), .A2(n4525), .ZN(n8132) );
  NAND2_X1 U5621 ( .A1(n4522), .A2(n4280), .ZN(n4521) );
  INV_X1 U5622 ( .A(n8449), .ZN(n8052) );
  NAND2_X1 U5623 ( .A1(n5037), .A2(n5036), .ZN(n7954) );
  NAND2_X1 U5624 ( .A1(n4904), .A2(n4903), .ZN(n7646) );
  NAND2_X1 U5625 ( .A1(n4912), .A2(n4911), .ZN(n7538) );
  INV_X1 U5626 ( .A(n7581), .ZN(n10019) );
  INV_X1 U5627 ( .A(n7424), .ZN(n10027) );
  AND2_X1 U5628 ( .A1(n7245), .A2(n10017), .ZN(n10034) );
  INV_X1 U5629 ( .A(n10020), .ZN(n10026) );
  OAI21_X1 U5630 ( .B1(n8724), .B2(n8862), .A(n8723), .ZN(n8887) );
  INV_X1 U5631 ( .A(n8722), .ZN(n8723) );
  XNOR2_X1 U5632 ( .A(n8720), .B(n8719), .ZN(n8724) );
  OAI22_X1 U5633 ( .A1(n8721), .A2(n8867), .B1(n8865), .B2(n8744), .ZN(n8722)
         );
  NAND2_X1 U5634 ( .A1(n8315), .A2(n8314), .ZN(n8945) );
  NAND2_X1 U5635 ( .A1(n5318), .A2(n5317), .ZN(n8954) );
  INV_X1 U5636 ( .A(n8246), .ZN(n8959) );
  NAND2_X1 U5637 ( .A1(n4576), .A2(n4577), .ZN(n8729) );
  NAND2_X1 U5638 ( .A1(n8772), .A2(n4579), .ZN(n4576) );
  AND2_X1 U5639 ( .A1(n5279), .A2(n5278), .ZN(n8964) );
  XNOR2_X1 U5640 ( .A(n8752), .B(n8751), .ZN(n8965) );
  OR2_X1 U5641 ( .A1(n8750), .A2(n8749), .ZN(n8752) );
  AND2_X1 U5642 ( .A1(n4583), .A2(n4581), .ZN(n8750) );
  AND2_X1 U5643 ( .A1(n4583), .A2(n5431), .ZN(n8757) );
  NAND2_X1 U5644 ( .A1(n5240), .A2(n5239), .ZN(n8976) );
  NAND2_X1 U5645 ( .A1(n5222), .A2(n5221), .ZN(n8982) );
  NAND2_X1 U5646 ( .A1(n8822), .A2(n5428), .ZN(n8821) );
  NAND2_X1 U5647 ( .A1(n4568), .A2(n4567), .ZN(n8822) );
  NAND2_X1 U5648 ( .A1(n5157), .A2(n5156), .ZN(n8998) );
  AND2_X1 U5649 ( .A1(n8840), .A2(n8839), .ZN(n8996) );
  NAND2_X1 U5650 ( .A1(n5138), .A2(n5137), .ZN(n9004) );
  NAND2_X1 U5651 ( .A1(n4596), .A2(n5425), .ZN(n8860) );
  NAND2_X1 U5652 ( .A1(n4806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4803) );
  XNOR2_X1 U5653 ( .A(n5379), .B(n5378), .ZN(n7970) );
  NAND2_X1 U5654 ( .A1(n5382), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U5655 ( .A1(n5382), .A2(n5381), .ZN(n7933) );
  NAND2_X1 U5656 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4927) );
  NAND2_X1 U5657 ( .A1(n4742), .A2(n4741), .ZN(n9026) );
  NOR2_X1 U5658 ( .A1(n4291), .A2(n4785), .ZN(n4741) );
  NAND2_X1 U5659 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  OAI21_X1 U5660 ( .B1(n4749), .B2(n4337), .A(n4358), .ZN(n4355) );
  AND2_X1 U5661 ( .A1(n4747), .A2(n4358), .ZN(n4357) );
  NOR2_X1 U5662 ( .A1(n8028), .A2(n6378), .ZN(n8084) );
  XNOR2_X1 U5663 ( .A(n9036), .B(n9037), .ZN(n9105) );
  NAND2_X1 U5664 ( .A1(n6433), .A2(n6432), .ZN(n9104) );
  NAND2_X1 U5665 ( .A1(n5715), .A2(n5714), .ZN(n9426) );
  AND2_X1 U5666 ( .A1(n9127), .A2(n9124), .ZN(n6792) );
  CLKBUF_X1 U5667 ( .A(n9135), .Z(n9760) );
  INV_X1 U5668 ( .A(n7997), .ZN(n9164) );
  INV_X1 U5669 ( .A(n7897), .ZN(n9165) );
  NAND4_X1 U5670 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n9174)
         );
  INV_X1 U5671 ( .A(n6930), .ZN(n9775) );
  AOI21_X1 U5672 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6932), .A(n7186), .ZN(
        n6972) );
  AOI21_X1 U5673 ( .B1(n6934), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6970), .ZN(
        n9787) );
  AOI21_X1 U5674 ( .B1(n6986), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6982), .ZN(
        n6985) );
  NOR2_X1 U5675 ( .A1(n7095), .A2(n4332), .ZN(n7098) );
  NOR2_X1 U5676 ( .A1(n7098), .A2(n7097), .ZN(n7157) );
  NOR2_X1 U5677 ( .A1(n7428), .A2(n4489), .ZN(n7432) );
  AND2_X1 U5678 ( .A1(n7429), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4489) );
  NOR2_X1 U5679 ( .A1(n7432), .A2(n7431), .ZN(n7602) );
  NOR2_X1 U5680 ( .A1(n7602), .A2(n4488), .ZN(n7606) );
  AND2_X1 U5681 ( .A1(n7603), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U5682 ( .A1(n7606), .A2(n7605), .ZN(n7617) );
  NOR2_X1 U5683 ( .A1(n7706), .A2(n4487), .ZN(n7710) );
  AND2_X1 U5684 ( .A1(n7707), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4487) );
  NOR2_X1 U5685 ( .A1(n7710), .A2(n7709), .ZN(n7979) );
  XNOR2_X1 U5686 ( .A(n9188), .B(n9187), .ZN(n7981) );
  NAND2_X1 U5687 ( .A1(n9201), .A2(n4492), .ZN(n9223) );
  NAND2_X1 U5688 ( .A1(n9286), .A2(n6634), .ZN(n9274) );
  OAI21_X1 U5689 ( .B1(n9301), .B2(n4452), .A(n4449), .ZN(n9267) );
  NAND2_X1 U5690 ( .A1(n9301), .A2(n6184), .ZN(n4453) );
  NOR2_X1 U5691 ( .A1(n4556), .A2(n4555), .ZN(n4788) );
  NAND2_X1 U5692 ( .A1(n9348), .A2(n4557), .ZN(n9338) );
  OAI21_X1 U5693 ( .B1(n9398), .B2(n4460), .A(n4458), .ZN(n9363) );
  NAND2_X1 U5694 ( .A1(n9398), .A2(n6131), .ZN(n4462) );
  INV_X1 U5695 ( .A(n9624), .ZN(n9082) );
  NAND2_X1 U5696 ( .A1(n4469), .A2(n4470), .ZN(n8116) );
  NOR2_X1 U5697 ( .A1(n8000), .A2(n6097), .ZN(n8118) );
  NAND2_X1 U5698 ( .A1(n4345), .A2(n4441), .ZN(n4438) );
  INV_X1 U5699 ( .A(n9293), .ZN(n9639) );
  INV_X1 U5700 ( .A(n9426), .ZN(n9662) );
  INV_X1 U5701 ( .A(n6104), .ZN(n9668) );
  NAND2_X1 U5702 ( .A1(n5684), .A2(n5683), .ZN(n7768) );
  NOR2_X1 U5703 ( .A1(n5788), .A2(n4734), .ZN(n4733) );
  INV_X1 U5704 ( .A(n6932), .ZN(n7193) );
  INV_X1 U5705 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6870) );
  XNOR2_X1 U5706 ( .A(n4477), .B(n4476), .ZN(n6930) );
  NAND2_X1 U5707 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4477) );
  NAND2_X1 U5708 ( .A1(n7306), .A2(n5838), .ZN(n7412) );
  INV_X1 U5709 ( .A(n4496), .ZN(n7741) );
  NOR2_X1 U5710 ( .A1(n8672), .A2(n4505), .ZN(n4504) );
  OR2_X1 U5711 ( .A1(n8676), .A2(n8675), .ZN(n4503) );
  OAI21_X1 U5712 ( .B1(n8669), .B2(n4507), .A(n8601), .ZN(n4506) );
  OAI21_X1 U5713 ( .B1(n8699), .B2(n8698), .A(n4383), .ZN(P2_U3200) );
  AND2_X1 U5714 ( .A1(n4387), .A2(n4384), .ZN(n4383) );
  NAND2_X1 U5715 ( .A1(n8693), .A2(n5557), .ZN(n4387) );
  NOR2_X1 U5716 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  AND2_X1 U5717 ( .A1(n4757), .A2(n5971), .ZN(n5972) );
  NAND2_X1 U5718 ( .A1(n5974), .A2(n8942), .ZN(n5973) );
  OAI21_X1 U5719 ( .B1(n8714), .B2(n8927), .A(n5435), .ZN(n5436) );
  OR2_X1 U5720 ( .A1(n8714), .A2(n9014), .ZN(n5586) );
  NAND2_X1 U5721 ( .A1(n4484), .A2(n4481), .ZN(P1_U3262) );
  AOI21_X1 U5722 ( .B1(n4485), .B2(n6219), .A(n9246), .ZN(n4484) );
  NAND2_X1 U5723 ( .A1(n4482), .A2(n8189), .ZN(n4481) );
  OR2_X1 U5724 ( .A1(n9435), .A2(n10013), .ZN(n9436) );
  OAI21_X1 U5725 ( .B1(n8178), .B2(n9633), .A(n6817), .ZN(n6818) );
  AOI21_X1 U5726 ( .B1(n6521), .B2(n5816), .A(n6520), .ZN(n6522) );
  NAND2_X1 U5727 ( .A1(n6672), .A2(n5816), .ZN(n5817) );
  NAND2_X1 U5728 ( .A1(n4560), .A2(n6258), .ZN(P1_U3519) );
  NAND2_X1 U5729 ( .A1(n6816), .A2(n10000), .ZN(n4560) );
  OR2_X1 U5730 ( .A1(n8976), .A2(n8235), .ZN(n5431) );
  AND2_X1 U5731 ( .A1(n7638), .A2(n8440), .ZN(n4279) );
  INV_X2 U5732 ( .A(n4945), .ZN(n4926) );
  NAND2_X1 U5733 ( .A1(n5957), .A2(n5956), .ZN(n5967) );
  NAND2_X1 U5734 ( .A1(n8449), .A2(n8134), .ZN(n4280) );
  NAND2_X1 U5735 ( .A1(n9139), .A2(n9140), .ZN(n9060) );
  INV_X1 U5736 ( .A(n5431), .ZN(n8383) );
  AND2_X1 U5737 ( .A1(n4462), .A2(n4463), .ZN(n9383) );
  OAI21_X1 U5738 ( .B1(n6409), .B2(n4752), .A(n4750), .ZN(n4749) );
  XOR2_X1 U5739 ( .A(n4861), .B(SI_10_), .Z(n4281) );
  NAND2_X1 U5740 ( .A1(n5727), .A2(n5726), .ZN(n9375) );
  NAND2_X1 U5741 ( .A1(n4748), .A2(n6411), .ZN(n9114) );
  NAND2_X1 U5742 ( .A1(n9454), .A2(n9155), .ZN(n4282) );
  AND3_X1 U5743 ( .A1(n4793), .A2(n4377), .A3(n4796), .ZN(n4283) );
  INV_X1 U5744 ( .A(n4637), .ZN(n4636) );
  OAI21_X1 U5745 ( .B1(n4640), .B2(n4293), .A(n5181), .ZN(n4637) );
  AND2_X1 U5746 ( .A1(n5737), .A2(n5736), .ZN(n9315) );
  INV_X1 U5747 ( .A(n9315), .ZN(n9454) );
  AND2_X1 U5748 ( .A1(n5770), .A2(n5769), .ZN(n4284) );
  OR2_X1 U5749 ( .A1(n4700), .A2(n8312), .ZN(n4285) );
  AND2_X1 U5750 ( .A1(n8471), .A2(n5425), .ZN(n4286) );
  AND2_X1 U5751 ( .A1(n4615), .A2(n4614), .ZN(n4287) );
  AND2_X1 U5752 ( .A1(n4440), .A2(n4779), .ZN(n4288) );
  OR2_X1 U5753 ( .A1(n4325), .A2(n4523), .ZN(n4289) );
  NAND2_X1 U5754 ( .A1(n9817), .A2(n4432), .ZN(n4441) );
  NOR2_X1 U5755 ( .A1(n9813), .A2(n4613), .ZN(n7731) );
  NAND2_X1 U5756 ( .A1(n4340), .A2(n4441), .ZN(n9802) );
  NAND2_X1 U5757 ( .A1(n5681), .A2(n5680), .ZN(n9811) );
  INV_X1 U5758 ( .A(n6358), .ZN(n4362) );
  AND2_X1 U5759 ( .A1(n5630), .A2(n9924), .ZN(n4602) );
  NAND2_X1 U5760 ( .A1(n7460), .A2(n7461), .ZN(n7458) );
  AND2_X1 U5761 ( .A1(n5431), .A2(n8381), .ZN(n4290) );
  INV_X1 U5762 ( .A(n7392), .ZN(n4502) );
  XNOR2_X1 U5763 ( .A(n6794), .B(n6385), .ZN(n4291) );
  INV_X1 U5764 ( .A(n7118), .ZN(n4495) );
  OR2_X1 U5765 ( .A1(n6768), .A2(n6220), .ZN(n4292) );
  NAND2_X1 U5766 ( .A1(n6497), .A2(n5611), .ZN(n4932) );
  OR2_X1 U5767 ( .A1(n5182), .A2(n4638), .ZN(n4293) );
  OR2_X1 U5768 ( .A1(n5354), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4294) );
  NAND2_X1 U5769 ( .A1(n4691), .A2(n4928), .ZN(n4897) );
  INV_X1 U5770 ( .A(n5994), .ZN(n6180) );
  AND4_X1 U5771 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n6297)
         );
  NAND2_X1 U5772 ( .A1(n8328), .A2(n8327), .ZN(n8366) );
  NAND4_X1 U5773 ( .A1(n4373), .A2(n4378), .A3(n4372), .A4(n4377), .ZN(n5354)
         );
  AND3_X1 U5774 ( .A1(n4881), .A2(n4798), .A3(n4797), .ZN(n4295) );
  AOI21_X1 U5775 ( .B1(n6905), .B2(n8325), .A(n5030), .ZN(n7696) );
  AOI21_X1 U5776 ( .B1(n4647), .B2(n4645), .A(n4644), .ZN(n4643) );
  NAND2_X1 U5777 ( .A1(n4321), .A2(n4282), .ZN(n4452) );
  INV_X1 U5778 ( .A(n4713), .ZN(n4712) );
  OR2_X1 U5779 ( .A1(n8210), .A2(n4714), .ZN(n4713) );
  NAND4_X1 U5780 ( .A1(n5991), .A2(n5990), .A3(n5989), .A4(n5988), .ZN(n6275)
         );
  NAND2_X1 U5781 ( .A1(n6488), .A2(n6487), .ZN(n8375) );
  AOI21_X1 U5782 ( .B1(n9318), .B2(n6173), .A(n6172), .ZN(n9301) );
  NAND2_X1 U5783 ( .A1(n9095), .A2(n6426), .ZN(n9051) );
  AOI21_X1 U5784 ( .B1(n9333), .B2(n6166), .A(n6165), .ZN(n9318) );
  NAND4_X1 U5785 ( .A1(n4937), .A2(n4936), .A3(n4935), .A4(n4934), .ZN(n7113)
         );
  AOI21_X1 U5786 ( .B1(n5954), .B2(n5953), .A(n4790), .ZN(n6490) );
  NAND2_X1 U5787 ( .A1(n8834), .A2(n4770), .ZN(n8823) );
  XNOR2_X1 U5788 ( .A(n4823), .B(SI_1_), .ZN(n4930) );
  AND2_X1 U5789 ( .A1(n8458), .A2(n8453), .ZN(n4296) );
  AND2_X1 U5790 ( .A1(n6679), .A2(n9349), .ZN(n4297) );
  OR2_X1 U5791 ( .A1(n6679), .A2(n6649), .ZN(n4298) );
  OR2_X1 U5792 ( .A1(n6651), .A2(n5759), .ZN(n4299) );
  OAI21_X1 U5793 ( .B1(n9095), .B2(n4361), .A(n4359), .ZN(n9036) );
  NAND4_X1 U5794 ( .A1(n4476), .A2(n5599), .A3(n5625), .A4(n5598), .ZN(n5635)
         );
  NAND2_X1 U5795 ( .A1(n5613), .A2(n5612), .ZN(n6216) );
  INV_X1 U5796 ( .A(n8545), .ZN(n4400) );
  NAND2_X1 U5797 ( .A1(n5722), .A2(n5721), .ZN(n9483) );
  INV_X1 U5798 ( .A(n9142), .ZN(n8102) );
  NAND2_X1 U5799 ( .A1(n5699), .A2(n5698), .ZN(n9142) );
  NAND2_X1 U5800 ( .A1(n4730), .A2(n4729), .ZN(n6460) );
  NAND2_X1 U5801 ( .A1(n5732), .A2(n5731), .ZN(n9463) );
  INV_X1 U5802 ( .A(n9463), .ZN(n4619) );
  NAND2_X1 U5803 ( .A1(n9125), .A2(n6792), .ZN(n9126) );
  AND2_X1 U5804 ( .A1(n6635), .A2(n6634), .ZN(n4300) );
  OR2_X1 U5805 ( .A1(n9811), .A2(n9167), .ZN(n4301) );
  NAND2_X1 U5806 ( .A1(n5686), .A2(n5605), .ZN(n5766) );
  AND3_X1 U5807 ( .A1(n4691), .A2(n4928), .A3(n4801), .ZN(n4302) );
  OR2_X1 U5808 ( .A1(n8970), .A2(n8743), .ZN(n8506) );
  INV_X1 U5809 ( .A(n8506), .ZN(n4582) );
  INV_X1 U5810 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9670) );
  AND2_X1 U5811 ( .A1(n4293), .A2(n4635), .ZN(n4303) );
  AND2_X1 U5812 ( .A1(n9657), .A2(n8169), .ZN(n4304) );
  NAND2_X1 U5813 ( .A1(n4356), .A2(n4355), .ZN(n9094) );
  INV_X1 U5814 ( .A(n4461), .ZN(n4460) );
  NOR2_X1 U5815 ( .A1(n6130), .A2(n4304), .ZN(n4461) );
  AND2_X1 U5816 ( .A1(n8447), .A2(n8446), .ZN(n4305) );
  NAND2_X1 U5817 ( .A1(n9325), .A2(n4617), .ZN(n4618) );
  OR2_X1 U5818 ( .A1(n8375), .A2(n8378), .ZN(n8531) );
  NAND2_X1 U5819 ( .A1(n8396), .A2(n8400), .ZN(n7200) );
  OR2_X1 U5820 ( .A1(n7796), .A2(n7800), .ZN(n6344) );
  AND2_X1 U5821 ( .A1(n6312), .A2(n6303), .ZN(n4306) );
  AND2_X1 U5822 ( .A1(n8682), .A2(n8681), .ZN(n4307) );
  AND2_X1 U5823 ( .A1(n4880), .A2(n4881), .ZN(n5033) );
  AND2_X1 U5824 ( .A1(n4620), .A2(n4619), .ZN(n4308) );
  INV_X1 U5825 ( .A(n4778), .ZN(n4442) );
  INV_X1 U5826 ( .A(n6199), .ZN(n9272) );
  AND2_X1 U5827 ( .A1(n5608), .A2(n4475), .ZN(n4309) );
  NOR2_X1 U5828 ( .A1(n9657), .A2(n8169), .ZN(n4310) );
  NOR2_X1 U5829 ( .A1(n9668), .A2(n8146), .ZN(n4311) );
  INV_X1 U5830 ( .A(n4520), .ZN(n4519) );
  NAND2_X1 U5831 ( .A1(n4524), .A2(n4280), .ZN(n4520) );
  AND3_X1 U5832 ( .A1(n6646), .A2(n6645), .A3(n6644), .ZN(n4312) );
  INV_X1 U5833 ( .A(n4622), .ZN(n5747) );
  OAI21_X1 U5834 ( .B1(n5332), .B2(n4626), .A(n4623), .ZN(n4622) );
  AND2_X1 U5835 ( .A1(n4755), .A2(n4309), .ZN(n4313) );
  AND2_X1 U5836 ( .A1(n8719), .A2(n8517), .ZN(n4314) );
  AND2_X1 U5837 ( .A1(n9639), .A2(n6787), .ZN(n4315) );
  AND2_X1 U5838 ( .A1(n5848), .A2(n7637), .ZN(n4316) );
  NOR2_X1 U5839 ( .A1(n6458), .A2(n6457), .ZN(n4317) );
  NAND2_X1 U5840 ( .A1(n9272), .A2(n9130), .ZN(n4318) );
  AND3_X1 U5841 ( .A1(n4607), .A2(n4608), .A3(n5605), .ZN(n5763) );
  OR2_X1 U5842 ( .A1(n4379), .A2(n4376), .ZN(n4319) );
  NAND2_X1 U5843 ( .A1(n5763), .A2(n5606), .ZN(n4320) );
  NAND2_X1 U5844 ( .A1(n8387), .A2(n8352), .ZN(n8835) );
  OAI21_X1 U5845 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(n6447) );
  OR2_X1 U5846 ( .A1(n9639), .A2(n6787), .ZN(n4321) );
  AND2_X1 U5847 ( .A1(n4697), .A2(n4696), .ZN(n4322) );
  AND2_X1 U5848 ( .A1(n4646), .A2(n4281), .ZN(n4323) );
  INV_X1 U5849 ( .A(n4435), .ZN(n4434) );
  NAND2_X1 U5850 ( .A1(n4444), .A2(n4301), .ZN(n4435) );
  NAND2_X1 U5851 ( .A1(n9258), .A2(n9257), .ZN(n9259) );
  INV_X1 U5852 ( .A(n4452), .ZN(n4451) );
  OR2_X1 U5853 ( .A1(n5783), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4324) );
  OAI21_X1 U5854 ( .B1(n4896), .B2(n4646), .A(n4643), .ZN(n5031) );
  INV_X1 U5855 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4476) );
  AND2_X1 U5856 ( .A1(n7920), .A2(n8933), .ZN(n4325) );
  AOI21_X1 U5857 ( .B1(n6460), .B2(n6459), .A(n4317), .ZN(n9125) );
  NAND2_X1 U5858 ( .A1(n5729), .A2(n5728), .ZN(n9356) );
  AND2_X1 U5859 ( .A1(n4694), .A2(n8231), .ZN(n4326) );
  INV_X1 U5860 ( .A(n5838), .ZN(n4719) );
  AND2_X1 U5861 ( .A1(n5104), .A2(n5081), .ZN(n4327) );
  AND2_X1 U5862 ( .A1(n5871), .A2(n5870), .ZN(n4328) );
  OR2_X1 U5863 ( .A1(n4862), .A2(n9540), .ZN(n4329) );
  AND2_X1 U5864 ( .A1(n6238), .A2(n6598), .ZN(n4330) );
  NAND2_X1 U5865 ( .A1(n4289), .A2(n4524), .ZN(n4518) );
  OR2_X1 U5866 ( .A1(n8246), .A2(n8744), .ZN(n8516) );
  INV_X1 U5867 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U5868 ( .A1(n4929), .A2(n5478), .ZN(n7028) );
  AND2_X1 U5869 ( .A1(n6847), .A2(n6263), .ZN(n6288) );
  INV_X1 U5870 ( .A(n8042), .ZN(n4522) );
  INV_X1 U5871 ( .A(n8574), .ZN(n7825) );
  AND2_X1 U5872 ( .A1(n4363), .A2(n6358), .ZN(n4331) );
  XNOR2_X1 U5873 ( .A(n5745), .B(SI_29_), .ZN(n8153) );
  OAI21_X1 U5874 ( .B1(n4363), .B2(n4362), .A(n7957), .ZN(n7956) );
  INV_X1 U5875 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U5876 ( .A1(n5426), .A2(n8480), .ZN(n8833) );
  AND3_X1 U5877 ( .A1(n5641), .A2(n5640), .A3(n5639), .ZN(n7485) );
  NAND2_X1 U5878 ( .A1(n9420), .A2(n6121), .ZN(n9398) );
  AND2_X1 U5879 ( .A1(n7099), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4332) );
  NAND2_X1 U5880 ( .A1(n4706), .A2(n4702), .ZN(n8232) );
  AND2_X1 U5881 ( .A1(n8914), .A2(n8838), .ZN(n4333) );
  INV_X1 U5882 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5131) );
  INV_X1 U5883 ( .A(n4379), .ZN(n4880) );
  NOR2_X1 U5884 ( .A1(n8084), .A2(n8083), .ZN(n8082) );
  NOR2_X1 U5885 ( .A1(n6395), .A2(n6394), .ZN(n9139) );
  OR2_X1 U5886 ( .A1(n5703), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4334) );
  NAND2_X1 U5887 ( .A1(n6404), .A2(n6403), .ZN(n9073) );
  NAND2_X1 U5888 ( .A1(n5744), .A2(n5743), .ZN(n9261) );
  INV_X1 U5889 ( .A(n9261), .ZN(n4614) );
  INV_X1 U5890 ( .A(n9953), .ZN(n7477) );
  AND3_X1 U5891 ( .A1(n5654), .A2(n5653), .A3(n5652), .ZN(n9953) );
  NOR2_X1 U5892 ( .A1(n7879), .A2(n7878), .ZN(n4335) );
  INV_X1 U5893 ( .A(n9326), .ZN(n9644) );
  NAND2_X1 U5894 ( .A1(n5734), .A2(n5733), .ZN(n9326) );
  INV_X1 U5895 ( .A(n4469), .ZN(n8000) );
  NAND2_X1 U5896 ( .A1(n8002), .A2(n8001), .ZN(n4469) );
  INV_X1 U5897 ( .A(n9391), .ZN(n9657) );
  NAND2_X1 U5898 ( .A1(n5724), .A2(n5723), .ZN(n9391) );
  AND2_X1 U5899 ( .A1(n5905), .A2(n8744), .ZN(n4336) );
  AND2_X1 U5900 ( .A1(n6418), .A2(n6417), .ZN(n4337) );
  INV_X1 U5901 ( .A(n5202), .ZN(n4635) );
  NOR2_X1 U5902 ( .A1(n6431), .A2(n6430), .ZN(n4338) );
  NAND2_X1 U5903 ( .A1(n6354), .A2(n6355), .ZN(n6358) );
  OAI21_X1 U5904 ( .B1(n8082), .B2(n4785), .A(n4291), .ZN(n4743) );
  INV_X1 U5905 ( .A(n9959), .ZN(n9845) );
  AND2_X1 U5906 ( .A1(n5659), .A2(n5658), .ZN(n9959) );
  NAND2_X1 U5907 ( .A1(n5109), .A2(n5108), .ZN(n9011) );
  OR2_X1 U5908 ( .A1(n5592), .A2(n5741), .ZN(n4339) );
  AND2_X1 U5909 ( .A1(n4436), .A2(n4444), .ZN(n4340) );
  INV_X1 U5910 ( .A(n5967), .ZN(n8530) );
  AOI21_X1 U5911 ( .B1(n6404), .B2(n4747), .A(n4749), .ZN(n8165) );
  AND2_X1 U5912 ( .A1(n4354), .A2(n6338), .ZN(n7795) );
  AND2_X1 U5913 ( .A1(n9201), .A2(n9200), .ZN(n4341) );
  AND2_X1 U5914 ( .A1(n4679), .A2(n4678), .ZN(n4342) );
  AND2_X1 U5915 ( .A1(n5583), .A2(n5582), .ZN(n10060) );
  NOR2_X1 U5916 ( .A1(n7475), .A2(n4606), .ZN(n7563) );
  OR2_X1 U5917 ( .A1(n9813), .A2(n9811), .ZN(n4343) );
  OAI21_X1 U5918 ( .B1(n7554), .B2(n7558), .A(n6040), .ZN(n9817) );
  AOI21_X1 U5919 ( .B1(n9860), .B2(n9861), .A(n6019), .ZN(n7473) );
  OAI22_X1 U5920 ( .A1(n7473), .A2(n7474), .B1(n9172), .B2(n7477), .ZN(n9837)
         );
  AOI21_X1 U5921 ( .B1(n9817), .B2(n9820), .A(n4778), .ZN(n7682) );
  INV_X1 U5922 ( .A(n9813), .ZN(n4611) );
  NAND2_X1 U5923 ( .A1(n4541), .A2(n4759), .ZN(n7526) );
  NAND2_X1 U5924 ( .A1(n4586), .A2(n8415), .ZN(n7446) );
  NAND2_X1 U5925 ( .A1(n4438), .A2(n4779), .ZN(n7729) );
  AND2_X1 U5926 ( .A1(n6575), .A2(n6715), .ZN(n7730) );
  INV_X1 U5927 ( .A(n7730), .ZN(n4440) );
  AND2_X1 U5928 ( .A1(n5389), .A2(n6862), .ZN(n5395) );
  NAND2_X1 U5929 ( .A1(n7487), .A2(n6315), .ZN(n7459) );
  NAND2_X1 U5930 ( .A1(n6304), .A2(n6303), .ZN(n7486) );
  INV_X1 U5931 ( .A(n5333), .ZN(n4630) );
  NAND2_X1 U5932 ( .A1(n5843), .A2(n5842), .ZN(n7576) );
  NAND2_X1 U5933 ( .A1(n7197), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4344) );
  AND2_X1 U5934 ( .A1(n4436), .A2(n4434), .ZN(n4345) );
  AND2_X1 U5935 ( .A1(n7576), .A2(n5845), .ZN(n4346) );
  INV_X1 U5936 ( .A(n4525), .ZN(n4523) );
  NAND2_X1 U5937 ( .A1(n8052), .A2(n8571), .ZN(n4525) );
  INV_X2 U5938 ( .A(n4828), .ZN(n5611) );
  NAND2_X1 U5939 ( .A1(n5452), .A2(n7392), .ZN(n8597) );
  INV_X1 U5940 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4725) );
  NOR2_X1 U5941 ( .A1(n5486), .A2(n4495), .ZN(n7232) );
  NOR2_X1 U5942 ( .A1(n9222), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4347) );
  INV_X1 U5943 ( .A(n4602), .ZN(n9886) );
  AND2_X1 U5944 ( .A1(n5489), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4348) );
  INV_X1 U5945 ( .A(n7158), .ZN(n4480) );
  OR2_X1 U5946 ( .A1(n5481), .A2(n4683), .ZN(n4349) );
  NOR2_X1 U5947 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9677) );
  INV_X1 U5948 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4407) );
  AOI21_X1 U5949 ( .B1(n6255), .B2(n9868), .A(n6254), .ZN(n8174) );
  NOR2_X4 U5950 ( .A1(n5927), .A2(n6863), .ZN(P2_U3893) );
  OR2_X2 U5951 ( .A1(n6847), .A2(n6846), .ZN(n9177) );
  NAND2_X1 U5952 ( .A1(n4791), .A2(n5807), .ZN(n6847) );
  NAND2_X1 U5953 ( .A1(n7583), .A2(n4353), .ZN(n4352) );
  NAND2_X1 U5954 ( .A1(n6404), .A2(n4357), .ZN(n4356) );
  NAND2_X1 U5955 ( .A1(n6358), .A2(n4365), .ZN(n9747) );
  INV_X1 U5956 ( .A(n9748), .ZN(n4364) );
  NAND2_X1 U5957 ( .A1(n6357), .A2(n6356), .ZN(n4365) );
  XNOR2_X1 U5958 ( .A(n6823), .B(n4368), .ZN(n6293) );
  NAND2_X1 U5959 ( .A1(n4369), .A2(n6287), .ZN(n4368) );
  NAND2_X1 U5960 ( .A1(n6286), .A2(n4370), .ZN(n4369) );
  NAND4_X1 U5961 ( .A1(n4377), .A2(n4295), .A3(n4793), .A4(n4796), .ZN(n4376)
         );
  NAND3_X1 U5962 ( .A1(n4391), .A2(n8521), .A3(n8522), .ZN(n4390) );
  NAND3_X1 U5963 ( .A1(n4397), .A2(n4395), .A3(n4296), .ZN(n4394) );
  NAND3_X1 U5964 ( .A1(n8429), .A2(n8447), .A3(n8540), .ZN(n4397) );
  NAND2_X1 U5965 ( .A1(n8546), .A2(n4399), .ZN(n4398) );
  NAND3_X1 U5966 ( .A1(n4405), .A2(n4403), .A3(n8482), .ZN(n4402) );
  NAND3_X1 U5967 ( .A1(n8481), .A2(n8547), .A3(n8480), .ZN(n4405) );
  MUX2_X1 U5968 ( .A(n6852), .B(n6855), .S(n5611), .Z(n4838) );
  NAND2_X1 U5969 ( .A1(n6627), .A2(n6626), .ZN(n6633) );
  OAI21_X1 U5970 ( .B1(n4412), .B2(n4312), .A(n4411), .ZN(n6652) );
  NAND2_X1 U5971 ( .A1(n4419), .A2(n4298), .ZN(n6624) );
  NAND3_X1 U5972 ( .A1(n4422), .A2(n4421), .A3(n4420), .ZN(n4419) );
  INV_X1 U5973 ( .A(n6621), .ZN(n4423) );
  NAND3_X1 U5974 ( .A1(n4427), .A2(n4426), .A3(n4329), .ZN(n5045) );
  NAND3_X1 U5975 ( .A1(n4896), .A2(n4643), .A3(n4281), .ZN(n4426) );
  INV_X4 U5976 ( .A(n5611), .ZN(n6853) );
  OAI21_X1 U5977 ( .B1(n5611), .B2(P2_DATAO_REG_8__SCAN_IN), .A(n4430), .ZN(
        n4429) );
  NAND2_X1 U5978 ( .A1(n5611), .A2(n6902), .ZN(n4430) );
  NAND3_X1 U5979 ( .A1(n4439), .A2(n6070), .A3(n4431), .ZN(n7787) );
  NAND3_X1 U5980 ( .A1(n4288), .A2(n4432), .A3(n9817), .ZN(n4431) );
  OR2_X1 U5981 ( .A1(n7687), .A2(n9168), .ZN(n4444) );
  NAND3_X1 U5982 ( .A1(n5976), .A2(n5775), .A3(P1_REG2_REG_0__SCAN_IN), .ZN(
        n5991) );
  NAND3_X1 U5983 ( .A1(n5976), .A2(n5775), .A3(P1_REG2_REG_1__SCAN_IN), .ZN(
        n5985) );
  NAND2_X1 U5984 ( .A1(n6248), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U5985 ( .A1(n6248), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6006) );
  INV_X1 U5986 ( .A(n6130), .ZN(n4463) );
  NAND4_X1 U5987 ( .A1(n4313), .A2(n4607), .A3(n5605), .A4(n4608), .ZN(n5788)
         );
  NAND4_X1 U5988 ( .A1(n4473), .A2(n4313), .A3(n4607), .A4(n4608), .ZN(n4472)
         );
  NAND4_X1 U5989 ( .A1(n4607), .A2(n4608), .A3(n5605), .A4(n4755), .ZN(n5783)
         );
  NAND2_X1 U5990 ( .A1(n9193), .A2(n4492), .ZN(n4491) );
  NAND2_X1 U5991 ( .A1(n4928), .A2(n4692), .ZN(n4947) );
  NOR2_X4 U5992 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4928) );
  INV_X1 U5993 ( .A(n5449), .ZN(n4493) );
  NAND2_X1 U5994 ( .A1(n4500), .A2(n4502), .ZN(n4501) );
  INV_X1 U5995 ( .A(n5452), .ZN(n4500) );
  NAND3_X1 U5996 ( .A1(n4501), .A2(P2_REG2_REG_7__SCAN_IN), .A3(n8597), .ZN(
        n7389) );
  NAND3_X1 U5997 ( .A1(n4506), .A2(n4504), .A3(n4503), .ZN(P2_U3199) );
  AND2_X1 U5998 ( .A1(n8670), .A2(n8671), .ZN(n4507) );
  NAND2_X1 U5999 ( .A1(n4810), .A2(n4812), .ZN(n5053) );
  NAND3_X1 U6000 ( .A1(n4812), .A2(n4810), .A3(P2_REG3_REG_2__SCAN_IN), .ZN(
        n4954) );
  NAND3_X1 U6001 ( .A1(n4812), .A2(n4810), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n4923) );
  NAND2_X1 U6002 ( .A1(n4509), .A2(n4510), .ZN(n8809) );
  NAND2_X1 U6003 ( .A1(n8836), .A2(n4511), .ZN(n4509) );
  NAND2_X1 U6004 ( .A1(n8042), .A2(n4518), .ZN(n4514) );
  NAND2_X1 U6005 ( .A1(n5017), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U6006 ( .A1(n9303), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U6007 ( .A1(n4930), .A2(n4931), .ZN(n4826) );
  OAI21_X1 U6008 ( .B1(n5619), .B2(n5618), .A(n4941), .ZN(n4931) );
  NAND2_X1 U6009 ( .A1(n4828), .A2(SI_0_), .ZN(n5619) );
  NAND2_X1 U6010 ( .A1(n4552), .A2(n4669), .ZN(n4823) );
  NAND2_X1 U6011 ( .A1(n4828), .A2(n6870), .ZN(n4552) );
  INV_X1 U6012 ( .A(n4553), .ZN(n9322) );
  NAND2_X1 U6013 ( .A1(n4558), .A2(n4330), .ZN(n9415) );
  NAND2_X1 U6014 ( .A1(n7776), .A2(n6716), .ZN(n7896) );
  NAND2_X1 U6015 ( .A1(n7992), .A2(n6235), .ZN(n7994) );
  NAND2_X1 U6016 ( .A1(n5426), .A2(n4563), .ZN(n4562) );
  OAI21_X1 U6017 ( .B1(n8772), .B2(n4574), .A(n4571), .ZN(n8715) );
  NAND2_X1 U6018 ( .A1(n4586), .A2(n4584), .ZN(n7545) );
  NAND2_X1 U6019 ( .A1(n8046), .A2(n4590), .ZN(n4589) );
  NAND2_X1 U6020 ( .A1(n8046), .A2(n8458), .ZN(n8045) );
  NAND2_X1 U6021 ( .A1(n4596), .A2(n4286), .ZN(n8844) );
  INV_X1 U6022 ( .A(n7264), .ZN(n7170) );
  NAND2_X1 U6023 ( .A1(n7272), .A2(n7264), .ZN(n8400) );
  NAND2_X1 U6024 ( .A1(n4602), .A2(n9930), .ZN(n4601) );
  INV_X1 U6025 ( .A(n7475), .ZN(n4604) );
  NAND2_X1 U6026 ( .A1(n4604), .A2(n4605), .ZN(n9829) );
  NOR2_X2 U6027 ( .A1(n5635), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U6028 ( .A1(n4611), .A2(n4609), .ZN(n8004) );
  NAND2_X1 U6029 ( .A1(n9325), .A2(n4287), .ZN(n6256) );
  INV_X1 U6030 ( .A(n4618), .ZN(n9292) );
  OAI21_X1 U6031 ( .B1(n5332), .B2(n4630), .A(n4628), .ZN(n5594) );
  NAND2_X1 U6032 ( .A1(n5150), .A2(n4631), .ZN(n4634) );
  NAND2_X1 U6033 ( .A1(n5150), .A2(n4640), .ZN(n4639) );
  NAND2_X1 U6034 ( .A1(n5150), .A2(n5149), .ZN(n5167) );
  NAND2_X1 U6035 ( .A1(n4648), .A2(n4327), .ZN(n5122) );
  OAI22_X1 U6036 ( .A1(n5234), .A2(n4650), .B1(n4652), .B2(n4655), .ZN(n4649)
         );
  OR2_X1 U6037 ( .A1(n5234), .A2(n5233), .ZN(n4660) );
  NAND2_X1 U6038 ( .A1(n4664), .A2(n4661), .ZN(n8538) );
  NAND2_X1 U6039 ( .A1(n4663), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U6040 ( .A1(n8539), .A2(n8376), .ZN(n8528) );
  NAND2_X1 U6041 ( .A1(n4668), .A2(n8529), .ZN(n4663) );
  NAND2_X1 U6042 ( .A1(n4667), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U6043 ( .A1(n4668), .A2(n8530), .ZN(n4667) );
  NAND2_X2 U6044 ( .A1(n4821), .A2(n4820), .ZN(n4828) );
  NAND3_X1 U6045 ( .A1(n4821), .A2(n4820), .A3(n6854), .ZN(n4669) );
  NAND2_X1 U6046 ( .A1(n8632), .A2(n4673), .ZN(n4670) );
  INV_X1 U6047 ( .A(n5503), .ZN(n4678) );
  INV_X1 U6048 ( .A(n4679), .ZN(n8011) );
  OAI21_X1 U6049 ( .B1(n8592), .B2(n8593), .A(n4680), .ZN(n8596) );
  NAND2_X1 U6050 ( .A1(n5489), .A2(n4681), .ZN(n4680) );
  INV_X1 U6051 ( .A(n5481), .ZN(n4682) );
  MUX2_X1 U6052 ( .A(n9025), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6053 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9025), .S(n6497), .Z(n7257) );
  NAND2_X1 U6054 ( .A1(n4687), .A2(n4689), .ZN(n4688) );
  NAND2_X1 U6055 ( .A1(n5486), .A2(n4495), .ZN(n4690) );
  INV_X1 U6056 ( .A(n7232), .ZN(n4687) );
  NAND2_X1 U6057 ( .A1(n4688), .A2(n7231), .ZN(n7229) );
  NAND2_X2 U6058 ( .A1(n8582), .A2(n7170), .ZN(n8396) );
  NOR2_X1 U6059 ( .A1(n8582), .A2(n7264), .ZN(n4942) );
  INV_X2 U6060 ( .A(n7272), .ZN(n8582) );
  INV_X1 U6061 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4692) );
  OAI211_X1 U6062 ( .C1(n5911), .C2(n4285), .A(n4326), .B(n4693), .ZN(P2_U3160) );
  NAND3_X1 U6063 ( .A1(n5911), .A2(n4695), .A3(n4699), .ZN(n4693) );
  NOR2_X1 U6064 ( .A1(n5911), .A2(n5910), .ZN(n8224) );
  NAND2_X1 U6065 ( .A1(n8226), .A2(n8222), .ZN(n4696) );
  OR2_X1 U6066 ( .A1(n8226), .A2(n4698), .ZN(n4697) );
  INV_X1 U6067 ( .A(n8226), .ZN(n4699) );
  NAND2_X1 U6068 ( .A1(n8290), .A2(n4707), .ZN(n4706) );
  NAND2_X1 U6069 ( .A1(n4715), .A2(n4328), .ZN(n8074) );
  NAND2_X1 U6070 ( .A1(n7308), .A2(n5838), .ZN(n4718) );
  INV_X1 U6071 ( .A(n7308), .ZN(n4720) );
  NAND2_X1 U6072 ( .A1(n4718), .A2(n4716), .ZN(n5841) );
  INV_X1 U6073 ( .A(n4717), .ZN(n4716) );
  NAND2_X1 U6074 ( .A1(n4721), .A2(n4722), .ZN(n5864) );
  NAND2_X1 U6075 ( .A1(n7652), .A2(n5855), .ZN(n4721) );
  OAI21_X2 U6076 ( .B1(n5843), .B2(n4727), .A(n4726), .ZN(n7611) );
  NAND2_X1 U6077 ( .A1(n9051), .A2(n4731), .ZN(n4730) );
  NOR2_X1 U6078 ( .A1(n5788), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6079 ( .A1(n4284), .A2(n4733), .ZN(n4736) );
  NAND2_X1 U6080 ( .A1(n9073), .A2(n6409), .ZN(n9113) );
  NAND2_X1 U6081 ( .A1(n9073), .A2(n6410), .ZN(n4748) );
  INV_X1 U6082 ( .A(n6410), .ZN(n4751) );
  NAND3_X1 U6083 ( .A1(n7460), .A2(n7461), .A3(n6325), .ZN(n7501) );
  NAND2_X1 U6084 ( .A1(n4754), .A2(n6352), .ZN(n6357) );
  NAND2_X1 U6085 ( .A1(n5675), .A2(n5674), .ZN(n9813) );
  NAND2_X1 U6086 ( .A1(n5655), .A2(n9953), .ZN(n7475) );
  NAND2_X1 U6087 ( .A1(n5768), .A2(n9901), .ZN(n9250) );
  XNOR2_X1 U6088 ( .A(n6504), .B(n5759), .ZN(n5768) );
  AOI21_X1 U6089 ( .B1(n8555), .B2(n8554), .A(n8553), .ZN(n8562) );
  INV_X1 U6090 ( .A(n9862), .ZN(n5655) );
  NAND2_X1 U6091 ( .A1(n5393), .A2(n7544), .ZN(n5819) );
  INV_X1 U6092 ( .A(n4278), .ZN(n6701) );
  NAND2_X1 U6093 ( .A1(n6001), .A2(n6000), .ZN(n7347) );
  XNOR2_X1 U6094 ( .A(n9043), .B(n9042), .ZN(n9050) );
  INV_X1 U6095 ( .A(n7348), .ZN(n6007) );
  OAI21_X1 U6096 ( .B1(n8224), .B2(n5946), .A(n4789), .ZN(P2_U3154) );
  NOR2_X1 U6097 ( .A1(n9105), .A2(n9104), .ZN(n9103) );
  OAI22_X2 U6098 ( .A1(n6486), .A2(n6485), .B1(n8529), .B2(n5967), .ZN(n8365)
         );
  OR2_X1 U6099 ( .A1(n9174), .A2(n7485), .ZN(n9851) );
  OAI21_X2 U6100 ( .B1(n7450), .B2(n7448), .A(n7447), .ZN(n7547) );
  INV_X1 U6101 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U6102 ( .A1(n5911), .A2(n5910), .ZN(n5917) );
  AND2_X1 U6103 ( .A1(n5686), .A2(n5685), .ZN(n5691) );
  OR2_X1 U6104 ( .A1(n8158), .A2(n9014), .ZN(n4756) );
  INV_X1 U6105 ( .A(n8312), .ZN(n5916) );
  OR2_X1 U6106 ( .A1(n8158), .A2(n8927), .ZN(n4757) );
  OR2_X1 U6107 ( .A1(n6847), .A2(n9777), .ZN(n4758) );
  OR2_X1 U6108 ( .A1(n7417), .A2(n10019), .ZN(n4759) );
  INV_X1 U6109 ( .A(n8824), .ZN(n5428) );
  AND2_X1 U6110 ( .A1(n7271), .A2(n7320), .ZN(n4760) );
  OR2_X1 U6111 ( .A1(n10057), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n4761) );
  OR2_X1 U6112 ( .A1(n10057), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4762) );
  INV_X1 U6113 ( .A(n9667), .ZN(n5816) );
  AND3_X1 U6114 ( .A1(n4873), .A2(n5387), .A3(n4875), .ZN(n4763) );
  AND3_X1 U6115 ( .A1(n6140), .A2(n6139), .A3(n6138), .ZN(n8169) );
  INV_X1 U6116 ( .A(n9633), .ZN(n6529) );
  OR2_X1 U6117 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4764) );
  AND2_X1 U6118 ( .A1(n7136), .A2(n6745), .ZN(n9901) );
  OR2_X1 U6119 ( .A1(n6533), .A2(n8989), .ZN(n4765) );
  AND4_X1 U6120 ( .A1(n8522), .A2(n8719), .A3(n8732), .A4(n8361), .ZN(n4766)
         );
  NOR2_X1 U6121 ( .A1(n8763), .A2(n5268), .ZN(n4767) );
  OR2_X1 U6122 ( .A1(n8826), .A2(n8217), .ZN(n4768) );
  OR2_X1 U6123 ( .A1(n9739), .A2(n8866), .ZN(n4769) );
  OR2_X1 U6124 ( .A1(n8261), .A2(n8851), .ZN(n4770) );
  AND2_X1 U6125 ( .A1(n9649), .A2(n9053), .ZN(n4771) );
  AND3_X1 U6126 ( .A1(n6831), .A2(n6830), .A3(n9148), .ZN(n4772) );
  OR2_X1 U6127 ( .A1(n6533), .A2(n8908), .ZN(n4773) );
  OR2_X1 U6128 ( .A1(n6769), .A2(n6768), .ZN(n4775) );
  AND2_X1 U6129 ( .A1(n9998), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4776) );
  OR2_X1 U6130 ( .A1(n7640), .A2(n7517), .ZN(n4777) );
  AND2_X1 U6131 ( .A1(n9830), .A2(n7680), .ZN(n4778) );
  OR2_X1 U6132 ( .A1(n9992), .A2(n7726), .ZN(n4779) );
  XOR2_X1 U6133 ( .A(n5123), .B(SI_15_), .Z(n4780) );
  AND4_X1 U6134 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(n9119)
         );
  OR2_X1 U6135 ( .A1(n7357), .A2(n6525), .ZN(n10013) );
  INV_X1 U6136 ( .A(n5522), .ZN(n5505) );
  AND4_X1 U6137 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n8121)
         );
  OR2_X1 U6138 ( .A1(n10015), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n4781) );
  OR2_X1 U6139 ( .A1(n7495), .A2(n8578), .ZN(n4782) );
  NAND2_X1 U6140 ( .A1(n6351), .A2(n7857), .ZN(n6352) );
  INV_X1 U6141 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4843) );
  OR2_X1 U6142 ( .A1(n8964), .A2(n8735), .ZN(n4783) );
  OR2_X1 U6143 ( .A1(n6739), .A2(n6757), .ZN(n4784) );
  NOR2_X1 U6144 ( .A1(n8366), .A2(n8329), .ZN(n8542) );
  INV_X1 U6145 ( .A(n6672), .ZN(n5759) );
  AND2_X1 U6146 ( .A1(n6384), .A2(n6383), .ZN(n4785) );
  OR2_X1 U6147 ( .A1(n8115), .A2(n8868), .ZN(n4786) );
  INV_X1 U6148 ( .A(n8188), .ZN(n6521) );
  INV_X1 U6149 ( .A(n9900), .ZN(n5630) );
  INV_X1 U6150 ( .A(n7588), .ZN(n9170) );
  NOR2_X1 U6151 ( .A1(n5021), .A2(n4890), .ZN(n4787) );
  AND4_X1 U6152 ( .A1(n5117), .A2(n5116), .A3(n5115), .A4(n5114), .ZN(n8850)
         );
  INV_X1 U6153 ( .A(n8850), .ZN(n5118) );
  AND2_X1 U6154 ( .A1(n5945), .A2(n5944), .ZN(n4789) );
  NOR2_X1 U6155 ( .A1(n5952), .A2(n5951), .ZN(n4790) );
  NAND2_X1 U6156 ( .A1(n5664), .A2(n5663), .ZN(n9967) );
  INV_X1 U6157 ( .A(n6219), .ZN(n8189) );
  AND2_X1 U6158 ( .A1(n7911), .A2(n5810), .ZN(n4791) );
  NAND2_X1 U6159 ( .A1(n7485), .A2(n9174), .ZN(n4792) );
  OR2_X1 U6160 ( .A1(n6568), .A2(n6567), .ZN(n6593) );
  NAND2_X1 U6161 ( .A1(n6597), .A2(n6596), .ZN(n6610) );
  NAND2_X1 U6162 ( .A1(n6601), .A2(n6649), .ZN(n6602) );
  NAND2_X1 U6163 ( .A1(n6603), .A2(n6602), .ZN(n6614) );
  AOI21_X1 U6164 ( .B1(n6620), .B2(n6619), .A(n6618), .ZN(n6621) );
  NOR2_X1 U6165 ( .A1(n6638), .A2(n6641), .ZN(n6639) );
  OR2_X1 U6166 ( .A1(n8375), .A2(n8547), .ZN(n8377) );
  OR2_X1 U6167 ( .A1(n8564), .A2(n8547), .ZN(n8379) );
  INV_X1 U6168 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4797) );
  INV_X1 U6169 ( .A(n8542), .ZN(n8543) );
  AND2_X1 U6170 ( .A1(n4794), .A2(n4882), .ZN(n4796) );
  INV_X1 U6171 ( .A(n9967), .ZN(n6039) );
  NAND2_X1 U6172 ( .A1(n4774), .A2(n8543), .ZN(n8544) );
  OAI21_X1 U6173 ( .B1(n8945), .B2(n8367), .A(n8548), .ZN(n8368) );
  INV_X1 U6174 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4868) );
  INV_X1 U6175 ( .A(n5345), .ZN(n5344) );
  INV_X1 U6176 ( .A(n9421), .ZN(n6238) );
  NAND2_X1 U6177 ( .A1(n7359), .A2(n6008), .ZN(n6009) );
  INV_X1 U6178 ( .A(n7578), .ZN(n5842) );
  OR2_X1 U6179 ( .A1(n7868), .A2(n8573), .ZN(n5856) );
  INV_X1 U6180 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5482) );
  AND2_X1 U6181 ( .A1(n4915), .A2(n4889), .ZN(n5021) );
  INV_X1 U6182 ( .A(n7489), .ZN(n6312) );
  INV_X1 U6183 ( .A(n6742), .ZN(n6745) );
  NOR2_X1 U6184 ( .A1(n9483), .A2(n9161), .ZN(n6130) );
  XNOR2_X1 U6185 ( .A(n7320), .B(n8225), .ZN(n5833) );
  AND2_X1 U6186 ( .A1(n7871), .A2(n5856), .ZN(n5857) );
  OR2_X1 U6187 ( .A1(n5363), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U6188 ( .A1(n5534), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5440) );
  OAI21_X1 U6189 ( .B1(n7228), .B2(n5451), .A(n7225), .ZN(n5452) );
  INV_X1 U6190 ( .A(n5301), .ZN(n5300) );
  INV_X1 U6191 ( .A(n5112), .ZN(n5111) );
  OR2_X1 U6192 ( .A1(n5038), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5050) );
  NOR2_X1 U6193 ( .A1(n8578), .A2(n7454), .ZN(n7448) );
  NAND2_X1 U6194 ( .A1(n8414), .A2(n8430), .ZN(n5421) );
  OAI21_X1 U6195 ( .B1(n6297), .B2(n6796), .A(n6296), .ZN(n6298) );
  OR2_X1 U6196 ( .A1(n9624), .A2(n9163), .ZN(n6113) );
  INV_X1 U6197 ( .A(n8121), .ZN(n6096) );
  OR2_X1 U6198 ( .A1(n7768), .A2(n9166), .ZN(n6070) );
  NOR2_X1 U6199 ( .A1(n6275), .A2(n9902), .ZN(n9893) );
  NAND2_X1 U6200 ( .A1(n6219), .A2(n7772), .ZN(n6649) );
  XNOR2_X1 U6201 ( .A(n5747), .B(n5748), .ZN(n5745) );
  INV_X1 U6202 ( .A(n5763), .ZN(n5764) );
  XNOR2_X1 U6203 ( .A(n4846), .B(SI_6_), .ZN(n5008) );
  INV_X1 U6204 ( .A(n8909), .ZN(n8217) );
  INV_X1 U6205 ( .A(n5959), .ZN(n8197) );
  OAI21_X1 U6206 ( .B1(n5534), .B2(P2_REG2_REG_2__SCAN_IN), .A(n5440), .ZN(
        n7031) );
  INV_X1 U6207 ( .A(n5518), .ZN(n5515) );
  OR2_X1 U6208 ( .A1(n5207), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5224) );
  OR2_X1 U6209 ( .A1(n5139), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5160) );
  OR2_X1 U6210 ( .A1(n7954), .A2(n8573), .ZN(n7841) );
  INV_X1 U6211 ( .A(n8436), .ZN(n5422) );
  INV_X1 U6212 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U6213 ( .A1(n8039), .A2(n8325), .ZN(n5318) );
  INV_X1 U6214 ( .A(n8352), .ZN(n5427) );
  INV_X1 U6215 ( .A(n7646), .ZN(n7640) );
  AOI21_X1 U6216 ( .B1(n9463), .B2(n6825), .A(n6440), .ZN(n9040) );
  AND2_X1 U6217 ( .A1(n6420), .A2(n6419), .ZN(n8166) );
  AND2_X1 U6218 ( .A1(n6343), .A2(n6342), .ZN(n7800) );
  AND2_X1 U6219 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6014) );
  NOR2_X1 U6220 ( .A1(n6853), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6513) );
  NOR2_X1 U6221 ( .A1(n9142), .A2(n6096), .ZN(n6097) );
  INV_X1 U6222 ( .A(n6663), .ZN(n7900) );
  INV_X1 U6223 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5813) );
  AND2_X1 U6224 ( .A1(n6708), .A2(n9803), .ZN(n7683) );
  AND2_X1 U6225 ( .A1(n8324), .A2(n5964), .ZN(n8378) );
  AND2_X1 U6226 ( .A1(n5230), .A2(n5229), .ZN(n8801) );
  AND4_X1 U6227 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n8134)
         );
  NAND2_X1 U6228 ( .A1(n8944), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5971) );
  INV_X1 U6229 ( .A(n8939), .ZN(n8915) );
  OAI21_X1 U6230 ( .B1(n9272), .B2(n9749), .A(n6812), .ZN(n6813) );
  AND2_X1 U6231 ( .A1(n6164), .A2(n6163), .ZN(n9107) );
  AND4_X1 U6232 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n7961)
         );
  AND2_X1 U6233 ( .A1(n6598), .A2(n6604), .ZN(n8145) );
  OR2_X1 U6234 ( .A1(n6913), .A2(n6467), .ZN(n9878) );
  NOR2_X1 U6235 ( .A1(n10000), .A2(n6519), .ZN(n6520) );
  OR2_X1 U6236 ( .A1(n5790), .A2(n8041), .ZN(n6897) );
  OR2_X1 U6237 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  XNOR2_X1 U6238 ( .A(n4844), .B(SI_5_), .ZN(n4993) );
  XNOR2_X1 U6239 ( .A(n4833), .B(SI_3_), .ZN(n4966) );
  AND2_X1 U6240 ( .A1(n5915), .A2(n5914), .ZN(n8312) );
  INV_X1 U6241 ( .A(n9011), .ZN(n8081) );
  NAND2_X1 U6242 ( .A1(n5325), .A2(n5324), .ZN(n8567) );
  AND4_X1 U6243 ( .A1(n5102), .A2(n5101), .A3(n5100), .A4(n5099), .ZN(n8866)
         );
  OR2_X1 U6244 ( .A1(n5819), .A2(n5920), .ZN(n10017) );
  INV_X1 U6245 ( .A(n8942), .ZN(n8944) );
  OAI21_X1 U6246 ( .B1(n5974), .B2(n10060), .A(n4761), .ZN(n5975) );
  INV_X1 U6247 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6876) );
  INV_X1 U6248 ( .A(n6813), .ZN(n6814) );
  INV_X1 U6249 ( .A(n6482), .ZN(n6483) );
  AND4_X1 U6250 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n8146)
         );
  AOI21_X1 U6251 ( .B1(n6521), .B2(n6529), .A(n6528), .ZN(n6530) );
  NOR2_X1 U6252 ( .A1(n4776), .A2(n6257), .ZN(n6258) );
  INV_X1 U6253 ( .A(n9375), .ZN(n9653) );
  OR2_X1 U6254 ( .A1(n6525), .A2(n6524), .ZN(n9998) );
  INV_X1 U6255 ( .A(n5976), .ZN(n8192) );
  INV_X1 U6256 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U6257 ( .A1(n5973), .A2(n5972), .ZN(P2_U3487) );
  NOR2_X1 U6258 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4873) );
  INV_X1 U6259 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5387) );
  INV_X1 U6260 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4875) );
  INV_X1 U6261 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U6262 ( .A1(n4804), .A2(n4802), .ZN(n4806) );
  INV_X1 U6263 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9017) );
  XNOR2_X2 U6264 ( .A(n4803), .B(n9017), .ZN(n4809) );
  INV_X1 U6265 ( .A(n4804), .ZN(n4871) );
  NAND2_X1 U6266 ( .A1(n4871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U6267 ( .A1(n4959), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n4817) );
  INV_X2 U6268 ( .A(n8155), .ZN(n4810) );
  NAND2_X2 U6269 ( .A1(n4809), .A2(n4810), .ZN(n4952) );
  INV_X1 U6270 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n4808) );
  OR2_X1 U6271 ( .A1(n4952), .A2(n4808), .ZN(n4816) );
  INV_X1 U6272 ( .A(n4809), .ZN(n4812) );
  INV_X1 U6273 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4889) );
  INV_X1 U6274 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5020) );
  AND2_X1 U6275 ( .A1(n5052), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n4811) );
  NOR2_X1 U6276 ( .A1(n5071), .A2(n4811), .ZN(n8049) );
  OR2_X1 U6277 ( .A1(n5053), .A2(n8049), .ZN(n4815) );
  NAND2_X4 U6278 ( .A1(n4812), .A2(n8155), .ZN(n4960) );
  INV_X1 U6279 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n4813) );
  OR2_X1 U6280 ( .A1(n4960), .A2(n4813), .ZN(n4814) );
  NAND2_X1 U6281 ( .A1(n9677), .A2(n4818), .ZN(n4821) );
  INV_X1 U6282 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6854) );
  INV_X1 U6283 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5618) );
  AND2_X1 U6284 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4822) );
  INV_X1 U6285 ( .A(n4823), .ZN(n4824) );
  NAND2_X1 U6286 ( .A1(n4824), .A2(SI_1_), .ZN(n4825) );
  NAND2_X1 U6287 ( .A1(n4826), .A2(n4825), .ZN(n4943) );
  INV_X1 U6288 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6857) );
  INV_X1 U6289 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6868) );
  XNOR2_X1 U6290 ( .A(n4829), .B(SI_2_), .ZN(n4944) );
  NAND2_X1 U6291 ( .A1(n4943), .A2(n4944), .ZN(n4832) );
  INV_X1 U6292 ( .A(n4829), .ZN(n4830) );
  NAND2_X1 U6293 ( .A1(n4830), .A2(SI_2_), .ZN(n4831) );
  NAND2_X1 U6294 ( .A1(n4832), .A2(n4831), .ZN(n4965) );
  INV_X1 U6295 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U6296 ( .A1(n4965), .A2(n4966), .ZN(n4836) );
  INV_X1 U6297 ( .A(n4833), .ZN(n4834) );
  NAND2_X1 U6298 ( .A1(n4834), .A2(SI_3_), .ZN(n4835) );
  INV_X1 U6299 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6855) );
  INV_X1 U6300 ( .A(SI_4_), .ZN(n4837) );
  INV_X1 U6301 ( .A(n4838), .ZN(n4839) );
  NAND2_X1 U6302 ( .A1(n4839), .A2(SI_4_), .ZN(n4840) );
  NAND2_X1 U6303 ( .A1(n4844), .A2(SI_5_), .ZN(n4845) );
  INV_X1 U6304 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6875) );
  MUX2_X1 U6305 ( .A(n6876), .B(n6875), .S(n6853), .Z(n4846) );
  INV_X1 U6306 ( .A(n4846), .ZN(n4847) );
  NAND2_X1 U6307 ( .A1(n4849), .A2(n4848), .ZN(n4905) );
  INV_X1 U6308 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6881) );
  INV_X1 U6309 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6880) );
  MUX2_X1 U6310 ( .A(n6881), .B(n6880), .S(n6853), .Z(n4850) );
  NAND2_X1 U6311 ( .A1(n4905), .A2(n4906), .ZN(n4853) );
  INV_X1 U6312 ( .A(n4850), .ZN(n4851) );
  INV_X1 U6313 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6902) );
  INV_X1 U6314 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6901) );
  INV_X1 U6315 ( .A(SI_8_), .ZN(n4854) );
  INV_X1 U6316 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6907) );
  INV_X1 U6317 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6906) );
  MUX2_X1 U6318 ( .A(n6907), .B(n6906), .S(n6853), .Z(n4857) );
  INV_X1 U6319 ( .A(SI_9_), .ZN(n4856) );
  INV_X1 U6320 ( .A(n4857), .ZN(n4858) );
  NAND2_X1 U6321 ( .A1(n4858), .A2(SI_9_), .ZN(n4859) );
  MUX2_X1 U6322 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6853), .Z(n4861) );
  INV_X1 U6323 ( .A(n4861), .ZN(n4862) );
  INV_X1 U6324 ( .A(SI_10_), .ZN(n9540) );
  INV_X1 U6325 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7048) );
  INV_X1 U6326 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7047) );
  MUX2_X1 U6327 ( .A(n7048), .B(n7047), .S(n6853), .Z(n4863) );
  INV_X1 U6328 ( .A(SI_11_), .ZN(n9573) );
  INV_X1 U6329 ( .A(n4863), .ZN(n4864) );
  NAND2_X1 U6330 ( .A1(n4864), .A2(SI_11_), .ZN(n4865) );
  MUX2_X1 U6331 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6853), .Z(n5060) );
  INV_X1 U6332 ( .A(n5062), .ZN(n4867) );
  XNOR2_X1 U6333 ( .A(n5063), .B(n4867), .ZN(n7087) );
  INV_X1 U6334 ( .A(n4873), .ZN(n5384) );
  NAND2_X1 U6335 ( .A1(n5387), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4874) );
  NOR2_X1 U6336 ( .A1(n5384), .A2(n4874), .ZN(n4879) );
  XNOR2_X1 U6337 ( .A(n4875), .B(P2_IR_REG_31__SCAN_IN), .ZN(n4878) );
  NAND3_X1 U6338 ( .A1(n4294), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n4877) );
  NAND2_X4 U6339 ( .A1(n5370), .A2(n5371), .ZN(n6497) );
  NAND2_X1 U6340 ( .A1(n7087), .A2(n8325), .ZN(n4887) );
  NAND2_X1 U6341 ( .A1(n6497), .A2(n6853), .ZN(n4945) );
  INV_X1 U6342 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U6343 ( .A1(n5033), .A2(n4882), .ZN(n5065) );
  NAND2_X1 U6344 ( .A1(n5065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4884) );
  INV_X1 U6345 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4883) );
  XNOR2_X1 U6346 ( .A(n4884), .B(n4883), .ZN(n7112) );
  OAI22_X1 U6347 ( .A1(n5135), .A2(n7110), .B1(n6497), .B2(n7112), .ZN(n4885)
         );
  INV_X1 U6348 ( .A(n4885), .ZN(n4886) );
  NAND2_X1 U6349 ( .A1(n4959), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n4894) );
  INV_X1 U6350 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5490) );
  OR2_X1 U6351 ( .A1(n4952), .A2(n5490), .ZN(n4893) );
  INV_X1 U6352 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n4888) );
  OR2_X1 U6353 ( .A1(n4960), .A2(n4888), .ZN(n4892) );
  NOR2_X1 U6354 ( .A1(n4915), .A2(n4889), .ZN(n4890) );
  OR2_X1 U6355 ( .A1(n5053), .A2(n4787), .ZN(n4891) );
  XNOR2_X1 U6356 ( .A(n4896), .B(n4895), .ZN(n6900) );
  NAND2_X1 U6357 ( .A1(n6900), .A2(n8325), .ZN(n4904) );
  OR2_X1 U6358 ( .A1(n4897), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4995) );
  NOR2_X1 U6359 ( .A1(n4995), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5011) );
  AND2_X1 U6360 ( .A1(n5011), .A2(n4898), .ZN(n4908) );
  NAND2_X1 U6361 ( .A1(n4908), .A2(n4899), .ZN(n5028) );
  NAND2_X1 U6362 ( .A1(n5028), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4901) );
  INV_X1 U6363 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4900) );
  XNOR2_X1 U6364 ( .A(n4901), .B(n4900), .ZN(n8587) );
  OAI22_X1 U6365 ( .A1(n5135), .A2(n6902), .B1(n6497), .B2(n8587), .ZN(n4902)
         );
  INV_X1 U6366 ( .A(n4902), .ZN(n4903) );
  INV_X1 U6367 ( .A(n4906), .ZN(n4907) );
  XNOR2_X1 U6368 ( .A(n4905), .B(n4907), .ZN(n6879) );
  NAND2_X1 U6369 ( .A1(n6879), .A2(n8325), .ZN(n4912) );
  NOR2_X1 U6370 ( .A1(n4908), .A2(n4868), .ZN(n4909) );
  XNOR2_X1 U6371 ( .A(n4909), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7392) );
  OAI22_X1 U6372 ( .A1(n5135), .A2(n6881), .B1(n6497), .B2(n7392), .ZN(n4910)
         );
  INV_X1 U6373 ( .A(n4910), .ZN(n4911) );
  NAND2_X1 U6374 ( .A1(n4959), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n4919) );
  INV_X1 U6375 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n4913) );
  OR2_X1 U6376 ( .A1(n4952), .A2(n4913), .ZN(n4918) );
  OR2_X1 U6377 ( .A1(n4960), .A2(n7536), .ZN(n4917) );
  AND2_X1 U6378 ( .A1(n5003), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n4914) );
  NOR2_X1 U6379 ( .A1(n4915), .A2(n4914), .ZN(n7535) );
  OR2_X1 U6380 ( .A1(n5053), .A2(n7535), .ZN(n4916) );
  NAND4_X1 U6381 ( .A1(n4919), .A2(n4918), .A3(n4917), .A4(n4916), .ZN(n8576)
         );
  INV_X1 U6382 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7262) );
  NAND2_X1 U6383 ( .A1(n8316), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4924) );
  INV_X1 U6384 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n4920) );
  INV_X1 U6385 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n4921) );
  MUX2_X1 U6386 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4927), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n4929) );
  INV_X1 U6387 ( .A(n4928), .ZN(n5478) );
  XNOR2_X1 U6388 ( .A(n4930), .B(n4931), .ZN(n6869) );
  NAND2_X1 U6389 ( .A1(n4959), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4937) );
  INV_X1 U6390 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5477) );
  OR2_X1 U6391 ( .A1(n4952), .A2(n5477), .ZN(n4936) );
  INV_X1 U6392 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n4933) );
  OR2_X1 U6393 ( .A1(n4960), .A2(n4933), .ZN(n4935) );
  INV_X1 U6394 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6956) );
  OR2_X1 U6395 ( .A1(n5053), .A2(n6956), .ZN(n4934) );
  INV_X1 U6396 ( .A(SI_0_), .ZN(n4939) );
  INV_X1 U6397 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4938) );
  OAI21_X1 U6398 ( .B1(n6853), .B2(n4939), .A(n4938), .ZN(n4940) );
  AND2_X1 U6399 ( .A1(n4941), .A2(n4940), .ZN(n9025) );
  NAND2_X1 U6400 ( .A1(n7113), .A2(n7257), .ZN(n7201) );
  XNOR2_X1 U6401 ( .A(n4943), .B(n4944), .ZN(n6867) );
  NAND2_X1 U6402 ( .A1(n4926), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4951) );
  INV_X1 U6403 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6404 ( .A1(n5190), .A2(n5534), .ZN(n4950) );
  NAND2_X1 U6405 ( .A1(n5094), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4957) );
  OR2_X1 U6406 ( .A1(n4952), .A2(n5482), .ZN(n4956) );
  INV_X1 U6407 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n4953) );
  OR2_X1 U6408 ( .A1(n8318), .A2(n4953), .ZN(n4955) );
  INV_X1 U6409 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7331) );
  NAND4_X2 U6410 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), .ZN(n8581)
         );
  NAND2_X1 U6411 ( .A1(n4959), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4964) );
  INV_X1 U6412 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5529) );
  OR2_X1 U6413 ( .A1(n4952), .A2(n5529), .ZN(n4963) );
  OR2_X1 U6414 ( .A1(n5053), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n4962) );
  INV_X1 U6415 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5530) );
  OR2_X1 U6416 ( .A1(n4960), .A2(n5530), .ZN(n4961) );
  XNOR2_X1 U6417 ( .A(n4965), .B(n4966), .ZN(n6858) );
  NAND2_X1 U6418 ( .A1(n4926), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6419 ( .A1(n4947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4967) );
  MUX2_X1 U6420 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4967), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n4968) );
  AND2_X1 U6421 ( .A1(n4968), .A2(n4897), .ZN(n7084) );
  NAND2_X1 U6422 ( .A1(n5190), .A2(n7084), .ZN(n4969) );
  OAI211_X1 U6423 ( .C1(n6858), .C2(n4932), .A(n4970), .B(n4969), .ZN(n7371)
         );
  INV_X1 U6424 ( .A(n7371), .ZN(n7320) );
  NAND2_X1 U6425 ( .A1(n7271), .A2(n7371), .ZN(n8430) );
  AOI21_X2 U6426 ( .B1(n7321), .B2(n5421), .A(n4760), .ZN(n7422) );
  NAND2_X1 U6427 ( .A1(n4959), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4975) );
  OR2_X1 U6428 ( .A1(n4952), .A2(n7426), .ZN(n4974) );
  AND2_X1 U6429 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n4971) );
  NOR2_X1 U6430 ( .A1(n4987), .A2(n4971), .ZN(n7310) );
  OR2_X1 U6431 ( .A1(n5053), .A2(n7310), .ZN(n4973) );
  INV_X1 U6432 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5446) );
  OR2_X1 U6433 ( .A1(n4960), .A2(n5446), .ZN(n4972) );
  NAND2_X1 U6434 ( .A1(n4897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4977) );
  INV_X1 U6435 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4976) );
  XNOR2_X1 U6436 ( .A(n4977), .B(n4976), .ZN(n7068) );
  OAI22_X1 U6437 ( .A1(n5135), .A2(n6855), .B1(n6497), .B2(n7068), .ZN(n4978)
         );
  INV_X1 U6438 ( .A(n4978), .ZN(n4984) );
  INV_X1 U6439 ( .A(n4979), .ZN(n4980) );
  XNOR2_X1 U6440 ( .A(n4981), .B(n4980), .ZN(n6856) );
  INV_X1 U6441 ( .A(n6856), .ZN(n4982) );
  NAND2_X1 U6442 ( .A1(n4982), .A2(n8325), .ZN(n4983) );
  NAND2_X1 U6443 ( .A1(n8410), .A2(n7424), .ZN(n4985) );
  AOI22_X1 U6444 ( .A1(n7422), .A2(n4985), .B1(n8579), .B2(n10027), .ZN(n7450)
         );
  NAND2_X1 U6445 ( .A1(n4959), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4992) );
  INV_X1 U6446 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4986) );
  INV_X1 U6447 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7452) );
  OR2_X1 U6448 ( .A1(n4960), .A2(n7452), .ZN(n4990) );
  OR2_X1 U6449 ( .A1(n4987), .A2(n7123), .ZN(n4988) );
  AND2_X1 U6450 ( .A1(n5001), .A2(n4988), .ZN(n7413) );
  XNOR2_X1 U6451 ( .A(n4994), .B(n4993), .ZN(n6873) );
  OR2_X1 U6452 ( .A1(n4932), .A2(n6873), .ZN(n5000) );
  NAND2_X1 U6453 ( .A1(n4995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4997) );
  INV_X1 U6454 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4996) );
  XNOR2_X1 U6455 ( .A(n4997), .B(n4996), .ZN(n7118) );
  OAI22_X1 U6456 ( .A1(n5135), .A2(n4843), .B1(n6497), .B2(n7118), .ZN(n4998)
         );
  INV_X1 U6457 ( .A(n4998), .ZN(n4999) );
  NAND2_X1 U6458 ( .A1(n5000), .A2(n4999), .ZN(n7454) );
  NAND2_X1 U6459 ( .A1(n8578), .A2(n7454), .ZN(n7447) );
  NAND2_X1 U6460 ( .A1(n4959), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5007) );
  INV_X1 U6461 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6462 ( .A1(n5001), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5002) );
  AND2_X1 U6463 ( .A1(n5003), .A2(n5002), .ZN(n10018) );
  INV_X1 U6464 ( .A(n5008), .ZN(n5009) );
  XNOR2_X1 U6465 ( .A(n5010), .B(n5009), .ZN(n6874) );
  NAND2_X1 U6466 ( .A1(n6874), .A2(n8325), .ZN(n5015) );
  NOR2_X1 U6467 ( .A1(n5011), .A2(n4868), .ZN(n5012) );
  XNOR2_X1 U6468 ( .A(n5012), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6878) );
  OAI22_X1 U6469 ( .A1(n5135), .A2(n6876), .B1(n6497), .B2(n6878), .ZN(n5013)
         );
  INV_X1 U6470 ( .A(n5013), .ZN(n5014) );
  OAI21_X1 U6471 ( .B1(n8575), .B2(n7646), .A(n7635), .ZN(n5017) );
  NAND2_X1 U6472 ( .A1(n4959), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5026) );
  INV_X1 U6473 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5018) );
  OR2_X1 U6474 ( .A1(n4952), .A2(n5018), .ZN(n5025) );
  INV_X1 U6475 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5019) );
  OR2_X1 U6476 ( .A1(n4960), .A2(n5019), .ZN(n5024) );
  OR2_X1 U6477 ( .A1(n5021), .A2(n5020), .ZN(n5022) );
  AND2_X1 U6478 ( .A1(n5038), .A2(n5022), .ZN(n7700) );
  OR2_X1 U6479 ( .A1(n5053), .A2(n7700), .ZN(n5023) );
  NAND4_X1 U6480 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n8574)
         );
  OAI21_X1 U6481 ( .B1(n5028), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5029) );
  XNOR2_X1 U6482 ( .A(n5029), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7675) );
  INV_X1 U6483 ( .A(n7675), .ZN(n6909) );
  OAI22_X1 U6484 ( .A1(n5135), .A2(n6907), .B1(n6497), .B2(n6909), .ZN(n5030)
         );
  XNOR2_X1 U6485 ( .A(n5031), .B(n4281), .ZN(n6918) );
  NAND2_X1 U6486 ( .A1(n6918), .A2(n8325), .ZN(n5037) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6920) );
  NOR2_X1 U6488 ( .A1(n4880), .A2(n4868), .ZN(n5032) );
  MUX2_X1 U6489 ( .A(n4868), .B(n5032), .S(P2_IR_REG_10__SCAN_IN), .Z(n5034)
         );
  OR2_X1 U6490 ( .A1(n5034), .A2(n5033), .ZN(n7742) );
  OAI22_X1 U6491 ( .A1(n5135), .A2(n6920), .B1(n6497), .B2(n7742), .ZN(n5035)
         );
  INV_X1 U6492 ( .A(n5035), .ZN(n5036) );
  NAND2_X1 U6493 ( .A1(n4959), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5043) );
  INV_X1 U6494 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5494) );
  OR2_X1 U6495 ( .A1(n4952), .A2(n5494), .ZN(n5042) );
  INV_X1 U6496 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5458) );
  OR2_X1 U6497 ( .A1(n4960), .A2(n5458), .ZN(n5041) );
  NAND2_X1 U6498 ( .A1(n5038), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5039) );
  AND2_X1 U6499 ( .A1(n5050), .A2(n5039), .ZN(n7849) );
  OR2_X1 U6500 ( .A1(n5053), .A2(n7849), .ZN(n5040) );
  NAND4_X1 U6501 ( .A1(n5043), .A2(n5042), .A3(n5041), .A4(n5040), .ZN(n8573)
         );
  XNOR2_X1 U6502 ( .A(n5045), .B(n5044), .ZN(n7046) );
  OR2_X1 U6503 ( .A1(n5033), .A2(n4868), .ZN(n5046) );
  XNOR2_X1 U6504 ( .A(n5046), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7822) );
  INV_X1 U6505 ( .A(n7822), .ZN(n7050) );
  OAI22_X1 U6506 ( .A1(n5135), .A2(n7048), .B1(n6497), .B2(n7050), .ZN(n5047)
         );
  AOI21_X1 U6507 ( .B1(n7046), .B2(n8325), .A(n5047), .ZN(n7940) );
  NOR2_X1 U6508 ( .A1(n5058), .A2(n7940), .ZN(n5059) );
  NAND2_X1 U6509 ( .A1(n4959), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5057) );
  INV_X1 U6510 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5048) );
  OR2_X1 U6511 ( .A1(n4952), .A2(n5048), .ZN(n5056) );
  INV_X1 U6512 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5049) );
  OR2_X1 U6513 ( .A1(n4960), .A2(n5049), .ZN(n5055) );
  NAND2_X1 U6514 ( .A1(n5050), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5051) );
  AND2_X1 U6515 ( .A1(n5052), .A2(n5051), .ZN(n7944) );
  OR2_X1 U6516 ( .A1(n5053), .A2(n7944), .ZN(n5054) );
  NAND4_X1 U6517 ( .A1(n5057), .A2(n5056), .A3(n5055), .A4(n5054), .ZN(n8572)
         );
  INV_X1 U6518 ( .A(n5058), .ZN(n7934) );
  INV_X1 U6519 ( .A(n7940), .ZN(n7946) );
  NAND2_X1 U6520 ( .A1(n5060), .A2(SI_12_), .ZN(n5061) );
  INV_X1 U6521 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9523) );
  INV_X1 U6522 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7139) );
  MUX2_X1 U6523 ( .A(n9523), .B(n7139), .S(n6853), .Z(n5079) );
  XNOR2_X1 U6524 ( .A(n5079), .B(SI_13_), .ZN(n5077) );
  INV_X1 U6525 ( .A(n5077), .ZN(n5064) );
  XNOR2_X1 U6526 ( .A(n5078), .B(n5064), .ZN(n7138) );
  NAND2_X1 U6527 ( .A1(n5130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5086) );
  XNOR2_X1 U6528 ( .A(n5086), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8025) );
  INV_X1 U6529 ( .A(n8025), .ZN(n7141) );
  OAI22_X1 U6530 ( .A1(n5135), .A2(n9523), .B1(n6497), .B2(n7141), .ZN(n5067)
         );
  INV_X1 U6531 ( .A(n8877), .ZN(n7920) );
  NAND2_X1 U6532 ( .A1(n4959), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5076) );
  INV_X1 U6533 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6534 ( .A1(n4952), .A2(n5068), .ZN(n5075) );
  INV_X1 U6535 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5069) );
  OR2_X1 U6536 ( .A1(n4960), .A2(n5069), .ZN(n5074) );
  INV_X1 U6537 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5070) );
  OR2_X1 U6538 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  AND2_X1 U6539 ( .A1(n5072), .A2(n5096), .ZN(n8876) );
  OR2_X1 U6540 ( .A1(n5053), .A2(n8876), .ZN(n5073) );
  INV_X1 U6541 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6542 ( .A1(n5080), .A2(SI_13_), .ZN(n5081) );
  INV_X1 U6543 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7196) );
  INV_X1 U6544 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7199) );
  MUX2_X1 U6545 ( .A(n7196), .B(n7199), .S(n6853), .Z(n5083) );
  INV_X1 U6546 ( .A(SI_14_), .ZN(n5082) );
  NAND2_X1 U6547 ( .A1(n5083), .A2(n5082), .ZN(n5120) );
  INV_X1 U6548 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6549 ( .A1(n5084), .A2(SI_14_), .ZN(n5085) );
  NAND2_X1 U6550 ( .A1(n5120), .A2(n5085), .ZN(n5103) );
  NAND2_X1 U6551 ( .A1(n7195), .A2(n8325), .ZN(n5093) );
  INV_X1 U6552 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6553 ( .A1(n5086), .A2(n5127), .ZN(n5087) );
  NAND2_X1 U6554 ( .A1(n5087), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5089) );
  INV_X1 U6555 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6556 ( .A1(n5089), .A2(n5088), .ZN(n5106) );
  OR2_X1 U6557 ( .A1(n5089), .A2(n5088), .ZN(n5090) );
  NAND2_X1 U6558 ( .A1(n5106), .A2(n5090), .ZN(n7197) );
  OAI22_X1 U6559 ( .A1(n5135), .A2(n7196), .B1(n6497), .B2(n7197), .ZN(n5091)
         );
  INV_X1 U6560 ( .A(n5091), .ZN(n5092) );
  NAND2_X1 U6561 ( .A1(n5094), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5102) );
  INV_X1 U6562 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5095) );
  OR2_X1 U6563 ( .A1(n4952), .A2(n5095), .ZN(n5101) );
  NAND2_X1 U6564 ( .A1(n5096), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5097) );
  AND2_X1 U6565 ( .A1(n5112), .A2(n5097), .ZN(n9743) );
  OR2_X1 U6566 ( .A1(n9743), .A2(n5053), .ZN(n5100) );
  INV_X1 U6567 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6568 ( .A1(n8318), .A2(n5098), .ZN(n5099) );
  NAND2_X1 U6569 ( .A1(n8468), .A2(n8866), .ZN(n5425) );
  NAND2_X1 U6570 ( .A1(n8929), .A2(n4769), .ZN(n8861) );
  NAND2_X1 U6571 ( .A1(n5122), .A2(n5120), .ZN(n5105) );
  MUX2_X1 U6572 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6853), .Z(n5123) );
  NAND2_X1 U6573 ( .A1(n7252), .A2(n8325), .ZN(n5109) );
  NAND2_X1 U6574 ( .A1(n5106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5107) );
  XNOR2_X1 U6575 ( .A(n5107), .B(P2_IR_REG_15__SCAN_IN), .ZN(n5522) );
  AOI22_X1 U6576 ( .A1(n4926), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5522), .B2(
        n5190), .ZN(n5108) );
  INV_X1 U6577 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6578 ( .A1(n5112), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6579 ( .A1(n5139), .A2(n5113), .ZN(n8873) );
  NAND2_X1 U6580 ( .A1(n5960), .A2(n8873), .ZN(n5117) );
  INV_X1 U6581 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9009) );
  OR2_X1 U6582 ( .A1(n8318), .A2(n9009), .ZN(n5116) );
  INV_X1 U6583 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8923) );
  OR2_X1 U6584 ( .A1(n4952), .A2(n8923), .ZN(n5115) );
  INV_X1 U6585 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8872) );
  OR2_X1 U6586 ( .A1(n4960), .A2(n8872), .ZN(n5114) );
  NAND2_X1 U6587 ( .A1(n9011), .A2(n8850), .ZN(n8471) );
  NAND2_X1 U6588 ( .A1(n8861), .A2(n8859), .ZN(n8870) );
  NAND2_X1 U6589 ( .A1(n8870), .A2(n5119), .ZN(n8847) );
  NAND2_X1 U6590 ( .A1(n5122), .A2(n5121), .ZN(n5125) );
  NAND2_X1 U6591 ( .A1(n5123), .A2(SI_15_), .ZN(n5124) );
  NAND2_X1 U6592 ( .A1(n5125), .A2(n5124), .ZN(n5146) );
  INV_X1 U6593 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7302) );
  INV_X1 U6594 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7305) );
  MUX2_X1 U6595 ( .A(n7302), .B(n7305), .S(n6853), .Z(n5147) );
  XNOR2_X1 U6596 ( .A(n5147), .B(SI_16_), .ZN(n5145) );
  INV_X1 U6597 ( .A(n5145), .ZN(n5126) );
  XNOR2_X1 U6598 ( .A(n5146), .B(n5126), .ZN(n7301) );
  NAND2_X1 U6599 ( .A1(n7301), .A2(n8325), .ZN(n5138) );
  NAND2_X1 U6600 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  OR2_X1 U6601 ( .A1(n5133), .A2(n4868), .ZN(n5132) );
  MUX2_X1 U6602 ( .A(n5132), .B(P2_IR_REG_31__SCAN_IN), .S(n5131), .Z(n5134)
         );
  NAND2_X1 U6603 ( .A1(n5133), .A2(n5131), .ZN(n5169) );
  NAND2_X1 U6604 ( .A1(n5134), .A2(n5169), .ZN(n7303) );
  OAI22_X1 U6605 ( .A1(n5135), .A2(n7302), .B1(n6497), .B2(n7303), .ZN(n5136)
         );
  INV_X1 U6606 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6607 ( .A1(n5139), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6608 ( .A1(n5160), .A2(n5140), .ZN(n8856) );
  NAND2_X1 U6609 ( .A1(n8856), .A2(n5960), .ZN(n5144) );
  NAND2_X1 U6610 ( .A1(n4959), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6611 ( .A1(n8316), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6612 ( .A1(n5094), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6613 ( .A1(n9004), .A2(n8868), .ZN(n8480) );
  NAND2_X1 U6614 ( .A1(n8473), .A2(n8480), .ZN(n8334) );
  NAND2_X1 U6615 ( .A1(n8847), .A2(n8334), .ZN(n8853) );
  INV_X1 U6616 ( .A(n9004), .ZN(n8115) );
  NAND2_X1 U6617 ( .A1(n8853), .A2(n4786), .ZN(n8836) );
  NAND2_X1 U6618 ( .A1(n5146), .A2(n5145), .ZN(n5150) );
  INV_X1 U6619 ( .A(n5147), .ZN(n5148) );
  NAND2_X1 U6620 ( .A1(n5148), .A2(SI_16_), .ZN(n5149) );
  INV_X1 U6621 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7404) );
  INV_X1 U6622 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7407) );
  MUX2_X1 U6623 ( .A(n7404), .B(n7407), .S(n6853), .Z(n5152) );
  INV_X1 U6624 ( .A(SI_17_), .ZN(n5151) );
  NAND2_X1 U6625 ( .A1(n5152), .A2(n5151), .ZN(n5165) );
  INV_X1 U6626 ( .A(n5152), .ZN(n5153) );
  NAND2_X1 U6627 ( .A1(n5153), .A2(SI_17_), .ZN(n5154) );
  NAND2_X1 U6628 ( .A1(n5165), .A2(n5154), .ZN(n5166) );
  XNOR2_X1 U6629 ( .A(n5167), .B(n5166), .ZN(n7403) );
  NAND2_X1 U6630 ( .A1(n7403), .A2(n8325), .ZN(n5157) );
  NAND2_X1 U6631 ( .A1(n5169), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5155) );
  XNOR2_X1 U6632 ( .A(n5155), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8673) );
  AOI22_X1 U6633 ( .A1(n4926), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5190), .B2(
        n8673), .ZN(n5156) );
  INV_X1 U6634 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6635 ( .A1(n5160), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6636 ( .A1(n5175), .A2(n5161), .ZN(n8841) );
  NAND2_X1 U6637 ( .A1(n8841), .A2(n5960), .ZN(n5164) );
  AOI22_X1 U6638 ( .A1(n5094), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8316), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6639 ( .A1(n4959), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6640 ( .A1(n8998), .A2(n8851), .ZN(n8352) );
  INV_X1 U6641 ( .A(n8998), .ZN(n8261) );
  MUX2_X1 U6642 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6853), .Z(n5180) );
  XNOR2_X1 U6643 ( .A(n5180), .B(SI_18_), .ZN(n5182) );
  INV_X1 U6644 ( .A(n5182), .ZN(n5168) );
  XNOR2_X1 U6645 ( .A(n5183), .B(n5168), .ZN(n7409) );
  NAND2_X1 U6646 ( .A1(n7409), .A2(n8325), .ZN(n5174) );
  NAND2_X1 U6647 ( .A1(n5171), .A2(n5170), .ZN(n5188) );
  OR2_X1 U6648 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  AND2_X1 U6649 ( .A1(n5188), .A2(n5172), .ZN(n5557) );
  AOI22_X1 U6650 ( .A1(n4926), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5557), .B2(
        n5190), .ZN(n5173) );
  INV_X1 U6651 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8829) );
  OR2_X2 U6652 ( .A1(n5175), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6653 ( .A1(n5175), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6654 ( .A1(n5195), .A2(n5176), .ZN(n8827) );
  NAND2_X1 U6655 ( .A1(n8827), .A2(n5960), .ZN(n5178) );
  AOI22_X1 U6656 ( .A1(n4959), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n8316), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n5177) );
  OAI211_X1 U6657 ( .C1(n4960), .C2(n8829), .A(n5178), .B(n5177), .ZN(n8838)
         );
  NAND2_X1 U6658 ( .A1(n5180), .A2(SI_18_), .ZN(n5181) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7500) );
  INV_X1 U6660 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8191) );
  MUX2_X1 U6661 ( .A(n7500), .B(n8191), .S(n6853), .Z(n5185) );
  INV_X1 U6662 ( .A(SI_19_), .ZN(n5184) );
  NAND2_X1 U6663 ( .A1(n5185), .A2(n5184), .ZN(n5201) );
  INV_X1 U6664 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6665 ( .A1(n5186), .A2(SI_19_), .ZN(n5187) );
  NAND2_X1 U6666 ( .A1(n5201), .A2(n5187), .ZN(n5202) );
  XNOR2_X1 U6667 ( .A(n5203), .B(n5202), .ZN(n7499) );
  NAND2_X1 U6668 ( .A1(n7499), .A2(n8325), .ZN(n5192) );
  AOI22_X1 U6669 ( .A1(n5579), .A2(n5190), .B1(n4926), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n5191) );
  INV_X1 U6670 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6671 ( .A1(n5195), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6672 ( .A1(n5207), .A2(n5196), .ZN(n8812) );
  INV_X1 U6673 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U6674 ( .A1(n8316), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6675 ( .A1(n4959), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5197) );
  OAI211_X1 U6676 ( .C1(n4960), .C2(n8814), .A(n5198), .B(n5197), .ZN(n5199)
         );
  AOI21_X1 U6677 ( .B1(n8812), .B2(n5960), .A(n5199), .ZN(n8826) );
  NAND2_X1 U6678 ( .A1(n8909), .A2(n8826), .ZN(n8488) );
  NAND2_X1 U6679 ( .A1(n8492), .A2(n8488), .ZN(n8357) );
  NAND2_X1 U6680 ( .A1(n8809), .A2(n8357), .ZN(n5200) );
  NAND2_X1 U6681 ( .A1(n5200), .A2(n4768), .ZN(n8758) );
  INV_X1 U6682 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7542) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7523) );
  MUX2_X1 U6684 ( .A(n7542), .B(n7523), .S(n6853), .Z(n5214) );
  XNOR2_X1 U6685 ( .A(n5214), .B(SI_20_), .ZN(n5204) );
  XNOR2_X1 U6686 ( .A(n5216), .B(n5204), .ZN(n7522) );
  NAND2_X1 U6687 ( .A1(n7522), .A2(n8325), .ZN(n5206) );
  NAND2_X1 U6688 ( .A1(n4926), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6689 ( .A1(n5207), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6690 ( .A1(n5224), .A2(n5208), .ZN(n8802) );
  NAND2_X1 U6691 ( .A1(n8802), .A2(n5960), .ZN(n5213) );
  INV_X1 U6692 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U6693 ( .A1(n4959), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6694 ( .A1(n8316), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5209) );
  OAI211_X1 U6695 ( .C1(n8805), .C2(n4960), .A(n5210), .B(n5209), .ZN(n5211)
         );
  INV_X1 U6696 ( .A(n5211), .ZN(n5212) );
  NAND2_X1 U6697 ( .A1(n8275), .A2(n8568), .ZN(n8496) );
  INV_X1 U6698 ( .A(SI_20_), .ZN(n5215) );
  OAI21_X1 U6699 ( .B1(n5216), .B2(n5215), .A(n5214), .ZN(n5218) );
  NAND2_X1 U6700 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6701 ( .A1(n5218), .A2(n5217), .ZN(n5234) );
  MUX2_X1 U6702 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6853), .Z(n5231) );
  INV_X1 U6703 ( .A(n5231), .ZN(n5219) );
  XNOR2_X1 U6704 ( .A(n5219), .B(SI_21_), .ZN(n5220) );
  XNOR2_X1 U6705 ( .A(n5234), .B(n5220), .ZN(n5725) );
  NAND2_X1 U6706 ( .A1(n5725), .A2(n8325), .ZN(n5222) );
  NAND2_X1 U6707 ( .A1(n4926), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5221) );
  INV_X1 U6708 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U6709 ( .A1(n5224), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6710 ( .A1(n5241), .A2(n5225), .ZN(n8795) );
  NAND2_X1 U6711 ( .A1(n8795), .A2(n5960), .ZN(n5230) );
  INV_X1 U6712 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U6713 ( .A1(n4959), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6714 ( .A1(n8316), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5226) );
  OAI211_X1 U6715 ( .C1(n8794), .C2(n4960), .A(n5227), .B(n5226), .ZN(n5228)
         );
  INV_X1 U6716 ( .A(n5228), .ZN(n5229) );
  NAND2_X1 U6717 ( .A1(n8982), .A2(n8801), .ZN(n8501) );
  NAND2_X1 U6718 ( .A1(n8502), .A2(n8501), .ZN(n8786) );
  NOR2_X1 U6719 ( .A1(n5231), .A2(SI_21_), .ZN(n5233) );
  NAND2_X1 U6720 ( .A1(n5231), .A2(SI_21_), .ZN(n5232) );
  INV_X1 U6721 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7773) );
  INV_X1 U6722 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9604) );
  MUX2_X1 U6723 ( .A(n7773), .B(n9604), .S(n6853), .Z(n5236) );
  INV_X1 U6724 ( .A(SI_22_), .ZN(n5235) );
  NAND2_X1 U6725 ( .A1(n5236), .A2(n5235), .ZN(n5248) );
  INV_X1 U6726 ( .A(n5236), .ZN(n5237) );
  NAND2_X1 U6727 ( .A1(n5237), .A2(SI_22_), .ZN(n5238) );
  NAND2_X1 U6728 ( .A1(n5248), .A2(n5238), .ZN(n5249) );
  NAND2_X1 U6729 ( .A1(n7771), .A2(n8325), .ZN(n5240) );
  NAND2_X1 U6730 ( .A1(n4926), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6731 ( .A1(n5241), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6732 ( .A1(n5258), .A2(n5242), .ZN(n8783) );
  NAND2_X1 U6733 ( .A1(n8783), .A2(n5960), .ZN(n5247) );
  INV_X1 U6734 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9534) );
  NAND2_X1 U6735 ( .A1(n4959), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6736 ( .A1(n5094), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5243) );
  OAI211_X1 U6737 ( .C1(n4952), .C2(n9534), .A(n5244), .B(n5243), .ZN(n5245)
         );
  INV_X1 U6738 ( .A(n5245), .ZN(n5246) );
  NAND2_X1 U6739 ( .A1(n8976), .A2(n8235), .ZN(n8381) );
  INV_X1 U6740 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5251) );
  INV_X1 U6741 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5730) );
  MUX2_X1 U6742 ( .A(n5251), .B(n5730), .S(n6853), .Z(n5253) );
  INV_X1 U6743 ( .A(SI_23_), .ZN(n5252) );
  NAND2_X1 U6744 ( .A1(n5253), .A2(n5252), .ZN(n5273) );
  INV_X1 U6745 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6746 ( .A1(n5254), .A2(SI_23_), .ZN(n5255) );
  AND2_X1 U6747 ( .A1(n5273), .A2(n5255), .ZN(n5271) );
  XNOR2_X1 U6748 ( .A(n5272), .B(n5271), .ZN(n7758) );
  NAND2_X1 U6749 ( .A1(n7758), .A2(n8325), .ZN(n5257) );
  NAND2_X1 U6750 ( .A1(n4926), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6751 ( .A1(n5258), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6752 ( .A1(n5282), .A2(n5259), .ZN(n8769) );
  NAND2_X1 U6753 ( .A1(n8769), .A2(n5960), .ZN(n5264) );
  INV_X1 U6754 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U6755 ( .A1(n8316), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6756 ( .A1(n4959), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5260) );
  OAI211_X1 U6757 ( .C1(n4960), .C2(n8768), .A(n5261), .B(n5260), .ZN(n5262)
         );
  INV_X1 U6758 ( .A(n5262), .ZN(n5263) );
  NOR2_X1 U6759 ( .A1(n8758), .A2(n5265), .ZN(n5269) );
  INV_X1 U6760 ( .A(n8976), .ZN(n8288) );
  NAND2_X1 U6761 ( .A1(n8288), .A2(n8235), .ZN(n8762) );
  INV_X1 U6762 ( .A(n8982), .ZN(n5266) );
  NAND2_X1 U6763 ( .A1(n5266), .A2(n8801), .ZN(n8776) );
  INV_X1 U6764 ( .A(n8275), .ZN(n8990) );
  NAND2_X1 U6765 ( .A1(n8990), .A2(n8568), .ZN(n8788) );
  NOR2_X1 U6766 ( .A1(n5269), .A2(n4767), .ZN(n8765) );
  INV_X1 U6767 ( .A(n8970), .ZN(n5898) );
  NAND2_X1 U6768 ( .A1(n8765), .A2(n5270), .ZN(n8741) );
  INV_X1 U6769 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7931) );
  INV_X1 U6770 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7912) );
  MUX2_X1 U6771 ( .A(n7931), .B(n7912), .S(n6853), .Z(n5275) );
  INV_X1 U6772 ( .A(SI_24_), .ZN(n5274) );
  NAND2_X1 U6773 ( .A1(n5275), .A2(n5274), .ZN(n5291) );
  INV_X1 U6774 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6775 ( .A1(n5276), .A2(SI_24_), .ZN(n5277) );
  AND2_X1 U6776 ( .A1(n5291), .A2(n5277), .ZN(n5289) );
  XNOR2_X1 U6777 ( .A(n5290), .B(n5289), .ZN(n7910) );
  NAND2_X1 U6778 ( .A1(n7910), .A2(n8325), .ZN(n5279) );
  NAND2_X1 U6779 ( .A1(n4926), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5278) );
  INV_X1 U6780 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6781 ( .A1(n5282), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6782 ( .A1(n5301), .A2(n5283), .ZN(n8745) );
  NAND2_X1 U6783 ( .A1(n8745), .A2(n5960), .ZN(n5288) );
  INV_X1 U6784 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U6785 ( .A1(n8316), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6786 ( .A1(n4959), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5284) );
  OAI211_X1 U6787 ( .C1(n4960), .C2(n8755), .A(n5285), .B(n5284), .ZN(n5286)
         );
  INV_X1 U6788 ( .A(n5286), .ZN(n5287) );
  NAND2_X1 U6789 ( .A1(n8964), .A2(n8735), .ZN(n8730) );
  NAND2_X1 U6790 ( .A1(n5290), .A2(n5289), .ZN(n5292) );
  NAND2_X1 U6791 ( .A1(n5292), .A2(n5291), .ZN(n5310) );
  INV_X1 U6792 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7968) );
  INV_X1 U6793 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9517) );
  MUX2_X1 U6794 ( .A(n7968), .B(n9517), .S(n6853), .Z(n5294) );
  INV_X1 U6795 ( .A(SI_25_), .ZN(n5293) );
  NAND2_X1 U6796 ( .A1(n5294), .A2(n5293), .ZN(n5311) );
  INV_X1 U6797 ( .A(n5294), .ZN(n5295) );
  NAND2_X1 U6798 ( .A1(n5295), .A2(SI_25_), .ZN(n5296) );
  AND2_X1 U6799 ( .A1(n5311), .A2(n5296), .ZN(n5309) );
  NAND2_X1 U6800 ( .A1(n7966), .A2(n8325), .ZN(n5298) );
  NAND2_X1 U6801 ( .A1(n4926), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5297) );
  INV_X1 U6802 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6803 ( .A1(n5301), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6804 ( .A1(n5319), .A2(n5302), .ZN(n8738) );
  NAND2_X1 U6805 ( .A1(n8738), .A2(n5960), .ZN(n5308) );
  INV_X1 U6806 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6807 ( .A1(n8316), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6808 ( .A1(n4959), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5303) );
  OAI211_X1 U6809 ( .C1(n5305), .C2(n4960), .A(n5304), .B(n5303), .ZN(n5306)
         );
  INV_X1 U6810 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6811 ( .A1(n8959), .A2(n8744), .ZN(n5328) );
  AND2_X1 U6812 ( .A1(n8730), .A2(n5328), .ZN(n8716) );
  NAND2_X1 U6813 ( .A1(n5310), .A2(n5309), .ZN(n5312) );
  NAND2_X1 U6814 ( .A1(n5312), .A2(n5311), .ZN(n5332) );
  INV_X1 U6815 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8059) );
  INV_X1 U6816 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8040) );
  MUX2_X1 U6817 ( .A(n8059), .B(n8040), .S(n6853), .Z(n5314) );
  INV_X1 U6818 ( .A(SI_26_), .ZN(n5313) );
  NAND2_X1 U6819 ( .A1(n5314), .A2(n5313), .ZN(n5333) );
  INV_X1 U6820 ( .A(n5314), .ZN(n5315) );
  NAND2_X1 U6821 ( .A1(n5315), .A2(SI_26_), .ZN(n5316) );
  AND2_X1 U6822 ( .A1(n5333), .A2(n5316), .ZN(n5331) );
  NAND2_X1 U6823 ( .A1(n4926), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6824 ( .A1(n5319), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6825 ( .A1(n5345), .A2(n5320), .ZN(n8726) );
  NAND2_X1 U6826 ( .A1(n8726), .A2(n5960), .ZN(n5325) );
  INV_X1 U6827 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U6828 ( .A1(n5094), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6829 ( .A1(n8316), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5321) );
  OAI211_X1 U6830 ( .C1(n8318), .C2(n8953), .A(n5322), .B(n5321), .ZN(n5323)
         );
  INV_X1 U6831 ( .A(n5323), .ZN(n5324) );
  NOR2_X1 U6832 ( .A1(n8954), .A2(n8567), .ZN(n5330) );
  INV_X1 U6833 ( .A(n5330), .ZN(n5326) );
  INV_X1 U6834 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6835 ( .A1(n8246), .A2(n8744), .ZN(n8515) );
  NAND2_X1 U6836 ( .A1(n8516), .A2(n8515), .ZN(n8333) );
  OR2_X1 U6837 ( .A1(n5330), .A2(n8717), .ZN(n5948) );
  NAND2_X1 U6838 ( .A1(n8954), .A2(n8567), .ZN(n5947) );
  INV_X1 U6839 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9576) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8164) );
  MUX2_X1 U6841 ( .A(n9576), .B(n8164), .S(n6853), .Z(n5335) );
  INV_X1 U6842 ( .A(SI_27_), .ZN(n5334) );
  NAND2_X1 U6843 ( .A1(n5335), .A2(n5334), .ZN(n5740) );
  INV_X1 U6844 ( .A(n5335), .ZN(n5336) );
  NAND2_X1 U6845 ( .A1(n5336), .A2(SI_27_), .ZN(n5337) );
  AND2_X1 U6846 ( .A1(n5740), .A2(n5337), .ZN(n5338) );
  OR2_X1 U6847 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  NAND2_X1 U6848 ( .A1(n5340), .A2(n5594), .ZN(n8071) );
  NAND2_X1 U6849 ( .A1(n8071), .A2(n8325), .ZN(n5342) );
  NAND2_X1 U6850 ( .A1(n4926), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5341) );
  INV_X1 U6851 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6852 ( .A1(n5345), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6853 ( .A1(n5363), .A2(n5346), .ZN(n8707) );
  NAND2_X1 U6854 ( .A1(n8707), .A2(n5960), .ZN(n5351) );
  INV_X1 U6855 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U6856 ( .A1(n8316), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6857 ( .A1(n4959), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5347) );
  OAI211_X1 U6858 ( .C1(n4960), .C2(n8708), .A(n5348), .B(n5347), .ZN(n5349)
         );
  INV_X1 U6859 ( .A(n5349), .ZN(n5350) );
  XNOR2_X1 U6860 ( .A(n5352), .B(n5951), .ZN(n5375) );
  NAND2_X1 U6861 ( .A1(n4319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5353) );
  MUX2_X1 U6862 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5353), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5355) );
  NAND2_X1 U6863 ( .A1(n5355), .A2(n5354), .ZN(n7775) );
  INV_X1 U6864 ( .A(n7775), .ZN(n8559) );
  NAND2_X1 U6865 ( .A1(n5579), .A2(n8559), .ZN(n5362) );
  NAND2_X1 U6866 ( .A1(n5033), .A2(n4283), .ZN(n5357) );
  NAND2_X1 U6867 ( .A1(n5359), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5356) );
  XNOR2_X1 U6868 ( .A(n5356), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U6869 ( .A1(n5357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5358) );
  MUX2_X1 U6870 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5358), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5360) );
  AND2_X1 U6871 ( .A1(n5360), .A2(n5359), .ZN(n8554) );
  NAND2_X1 U6872 ( .A1(n8371), .A2(n8554), .ZN(n5361) );
  NAND2_X1 U6873 ( .A1(n5362), .A2(n5361), .ZN(n8928) );
  NAND2_X1 U6874 ( .A1(n5363), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6875 ( .A1(n5959), .A2(n5364), .ZN(n8227) );
  NAND2_X1 U6876 ( .A1(n8227), .A2(n5960), .ZN(n5369) );
  INV_X1 U6877 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U6878 ( .A1(n4959), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6879 ( .A1(n8316), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5365) );
  OAI211_X1 U6880 ( .C1(n8156), .C2(n4960), .A(n5366), .B(n5365), .ZN(n5367)
         );
  INV_X1 U6881 ( .A(n5367), .ZN(n5368) );
  OAI21_X1 U6882 ( .B1(n5370), .B2(n8072), .A(n6497), .ZN(n5922) );
  NAND2_X1 U6883 ( .A1(n5922), .A2(n8547), .ZN(n8867) );
  INV_X1 U6884 ( .A(n5922), .ZN(n5923) );
  NAND2_X1 U6885 ( .A1(n5923), .A2(n8547), .ZN(n8865) );
  INV_X1 U6886 ( .A(n8711), .ZN(n5376) );
  INV_X1 U6887 ( .A(n8371), .ZN(n8390) );
  NAND2_X1 U6888 ( .A1(n8390), .A2(n7775), .ZN(n8939) );
  NOR2_X1 U6889 ( .A1(n5376), .A2(n8939), .ZN(n5377) );
  NOR2_X1 U6890 ( .A1(n8706), .A2(n5377), .ZN(n5584) );
  NAND2_X1 U6891 ( .A1(n8373), .A2(n8559), .ZN(n5432) );
  INV_X1 U6892 ( .A(n8554), .ZN(n7544) );
  OR2_X1 U6893 ( .A1(n5432), .A2(n7544), .ZN(n5394) );
  INV_X1 U6894 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5380) );
  INV_X1 U6895 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5378) );
  OR2_X1 U6896 ( .A1(n5386), .A2(n5380), .ZN(n5381) );
  XNOR2_X1 U6897 ( .A(n7933), .B(P2_B_REG_SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6898 ( .A1(n7970), .A2(n5383), .ZN(n5389) );
  NAND2_X1 U6899 ( .A1(n5384), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6900 ( .A1(n5386), .A2(n5385), .ZN(n5388) );
  XNOR2_X1 U6901 ( .A(n5388), .B(n5387), .ZN(n6862) );
  INV_X1 U6902 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U6903 ( .A1(n5395), .A2(n6866), .ZN(n5391) );
  INV_X1 U6904 ( .A(n6862), .ZN(n8058) );
  NAND2_X1 U6905 ( .A1(n8058), .A2(n7933), .ZN(n5390) );
  NAND2_X1 U6906 ( .A1(n5391), .A2(n5390), .ZN(n5575) );
  NOR2_X1 U6907 ( .A1(n5575), .A2(n8547), .ZN(n5392) );
  NAND2_X1 U6908 ( .A1(n5394), .A2(n5392), .ZN(n7242) );
  NOR2_X1 U6909 ( .A1(n5819), .A2(n8939), .ZN(n5398) );
  NAND2_X1 U6910 ( .A1(n5394), .A2(n8540), .ZN(n5397) );
  INV_X1 U6911 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6864) );
  AND2_X1 U6912 ( .A1(n7970), .A2(n8058), .ZN(n5396) );
  AOI21_X1 U6913 ( .B1(n5395), .B2(n6864), .A(n5396), .ZN(n7239) );
  NAND2_X1 U6914 ( .A1(n5397), .A2(n7239), .ZN(n7243) );
  OAI21_X1 U6915 ( .B1(n7242), .B2(n5398), .A(n7243), .ZN(n5416) );
  NAND2_X1 U6916 ( .A1(n8373), .A2(n7544), .ZN(n8549) );
  NAND2_X1 U6917 ( .A1(n8549), .A2(n8547), .ZN(n5928) );
  INV_X1 U6918 ( .A(n5395), .ZN(n6861) );
  NOR2_X1 U6919 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5402) );
  NOR4_X1 U6920 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5401) );
  NOR4_X1 U6921 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5400) );
  NOR4_X1 U6922 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5399) );
  NAND4_X1 U6923 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n5408)
         );
  NOR4_X1 U6924 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5406) );
  NOR4_X1 U6925 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5405) );
  NOR4_X1 U6926 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5404) );
  NOR4_X1 U6927 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5403) );
  NAND4_X1 U6928 ( .A1(n5406), .A2(n5405), .A3(n5404), .A4(n5403), .ZN(n5407)
         );
  NOR2_X1 U6929 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  OR2_X1 U6930 ( .A1(n6861), .A2(n5409), .ZN(n5574) );
  INV_X1 U6931 ( .A(n7933), .ZN(n5410) );
  AND2_X1 U6932 ( .A1(n6862), .A2(n5410), .ZN(n5412) );
  INV_X1 U6933 ( .A(n7970), .ZN(n5411) );
  NAND2_X1 U6934 ( .A1(n5412), .A2(n5411), .ZN(n5927) );
  NAND2_X1 U6935 ( .A1(n5354), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5413) );
  XNOR2_X1 U6936 ( .A(n5413), .B(n4725), .ZN(n5926) );
  AND2_X1 U6937 ( .A1(n5926), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6860) );
  AND2_X1 U6938 ( .A1(n5927), .A2(n6860), .ZN(n5919) );
  AND2_X1 U6939 ( .A1(n5574), .A2(n5919), .ZN(n5414) );
  NAND2_X1 U6940 ( .A1(n5928), .A2(n5414), .ZN(n7238) );
  INV_X1 U6941 ( .A(n5575), .ZN(n7240) );
  AND2_X1 U6942 ( .A1(n7240), .A2(n7239), .ZN(n5571) );
  NOR2_X1 U6943 ( .A1(n7238), .A2(n5571), .ZN(n5415) );
  AND2_X2 U6944 ( .A1(n5416), .A2(n5415), .ZN(n8942) );
  INV_X1 U6945 ( .A(n7200), .ZN(n5419) );
  INV_X1 U6946 ( .A(n7113), .ZN(n5417) );
  INV_X1 U6947 ( .A(n8391), .ZN(n5418) );
  NAND2_X1 U6948 ( .A1(n5419), .A2(n5418), .ZN(n7206) );
  NAND2_X1 U6949 ( .A1(n7206), .A2(n8400), .ZN(n7268) );
  NAND2_X1 U6950 ( .A1(n7268), .A2(n8399), .ZN(n5420) );
  INV_X1 U6951 ( .A(n8581), .ZN(n7323) );
  NAND2_X1 U6952 ( .A1(n7323), .A2(n7269), .ZN(n8404) );
  NAND2_X1 U6953 ( .A1(n5420), .A2(n8404), .ZN(n7319) );
  INV_X1 U6954 ( .A(n5421), .ZN(n8337) );
  NAND2_X1 U6955 ( .A1(n7319), .A2(n8337), .ZN(n7318) );
  NAND2_X1 U6956 ( .A1(n7318), .A2(n8430), .ZN(n7421) );
  XNOR2_X1 U6957 ( .A(n8579), .B(n10027), .ZN(n8339) );
  NAND2_X1 U6958 ( .A1(n8410), .A2(n10027), .ZN(n8415) );
  INV_X1 U6959 ( .A(n7454), .ZN(n7495) );
  NAND2_X1 U6960 ( .A1(n10019), .A2(n8577), .ZN(n8438) );
  NAND2_X1 U6961 ( .A1(n7495), .A2(n8578), .ZN(n8432) );
  AND2_X1 U6962 ( .A1(n8438), .A2(n8432), .ZN(n8417) );
  NAND2_X1 U6963 ( .A1(n7417), .A2(n7581), .ZN(n8436) );
  AOI21_X2 U6964 ( .B1(n7545), .B2(n8417), .A(n5422), .ZN(n7525) );
  OR2_X1 U6965 ( .A1(n7538), .A2(n7637), .ZN(n7638) );
  NAND2_X1 U6966 ( .A1(n7538), .A2(n7637), .ZN(n8440) );
  NAND2_X1 U6967 ( .A1(n7525), .A2(n4279), .ZN(n7524) );
  OR2_X1 U6968 ( .A1(n7646), .A2(n7517), .ZN(n8420) );
  AND2_X1 U6969 ( .A1(n8420), .A2(n7638), .ZN(n8424) );
  AND2_X1 U6970 ( .A1(n7646), .A2(n7517), .ZN(n8422) );
  AOI21_X2 U6971 ( .B1(n7524), .B2(n8424), .A(n8422), .ZN(n7691) );
  INV_X1 U6972 ( .A(n7696), .ZN(n7702) );
  OR2_X1 U6973 ( .A1(n7702), .A2(n7825), .ZN(n8421) );
  NAND2_X1 U6974 ( .A1(n7702), .A2(n7825), .ZN(n8446) );
  NAND2_X1 U6975 ( .A1(n7691), .A2(n8345), .ZN(n7690) );
  INV_X1 U6976 ( .A(n8573), .ZN(n7936) );
  OR2_X1 U6977 ( .A1(n7954), .A2(n7936), .ZN(n8450) );
  AND2_X1 U6978 ( .A1(n8450), .A2(n8421), .ZN(n8427) );
  NAND2_X1 U6979 ( .A1(n7690), .A2(n8427), .ZN(n7938) );
  INV_X1 U6980 ( .A(n8572), .ZN(n8044) );
  NAND2_X1 U6981 ( .A1(n7946), .A2(n8044), .ZN(n8452) );
  NAND2_X1 U6982 ( .A1(n7954), .A2(n7936), .ZN(n7937) );
  AND2_X1 U6983 ( .A1(n8452), .A2(n7937), .ZN(n8447) );
  NAND2_X1 U6984 ( .A1(n7938), .A2(n8447), .ZN(n5423) );
  OR2_X1 U6985 ( .A1(n7946), .A2(n8044), .ZN(n8453) );
  NAND2_X1 U6986 ( .A1(n5423), .A2(n8453), .ZN(n8046) );
  XNOR2_X1 U6987 ( .A(n8052), .B(n8571), .ZN(n8458) );
  OR2_X1 U6988 ( .A1(n8052), .A2(n8134), .ZN(n8455) );
  NAND2_X1 U6989 ( .A1(n7920), .A2(n8064), .ZN(n8464) );
  OR2_X1 U6990 ( .A1(n7920), .A2(n8064), .ZN(n8463) );
  INV_X1 U6991 ( .A(n8938), .ZN(n5424) );
  AND2_X1 U6992 ( .A1(n8473), .A2(n8845), .ZN(n8478) );
  NAND2_X1 U6993 ( .A1(n8844), .A2(n8478), .ZN(n5426) );
  INV_X1 U6994 ( .A(n8835), .ZN(n8482) );
  INV_X1 U6995 ( .A(n8838), .ZN(n8257) );
  NAND2_X1 U6996 ( .A1(n8914), .A2(n8257), .ZN(n8487) );
  NAND2_X1 U6997 ( .A1(n8484), .A2(n8487), .ZN(n8824) );
  INV_X1 U6998 ( .A(n8357), .ZN(n8816) );
  NAND2_X1 U6999 ( .A1(n8817), .A2(n8816), .ZN(n8815) );
  INV_X1 U7000 ( .A(n8493), .ZN(n5429) );
  OAI21_X1 U7001 ( .B1(n8804), .B2(n5429), .A(n8496), .ZN(n8787) );
  INV_X1 U7002 ( .A(n8501), .ZN(n5430) );
  OAI21_X2 U7003 ( .B1(n8787), .B2(n5430), .A(n8502), .ZN(n8772) );
  NAND2_X1 U7004 ( .A1(n8267), .A2(n8735), .ZN(n8512) );
  NAND2_X1 U7005 ( .A1(n8512), .A2(n8748), .ZN(n8507) );
  OR2_X2 U7006 ( .A1(n8954), .A2(n8736), .ZN(n8520) );
  XNOR2_X1 U7007 ( .A(n5970), .B(n8522), .ZN(n8714) );
  OR2_X1 U7008 ( .A1(n8549), .A2(n8540), .ZN(n5936) );
  NAND2_X1 U7009 ( .A1(n5936), .A2(n8939), .ZN(n7246) );
  AND2_X1 U7010 ( .A1(n8549), .A2(n5432), .ZN(n5433) );
  OR2_X1 U7011 ( .A1(n7246), .A2(n5433), .ZN(n7848) );
  OR2_X1 U7012 ( .A1(n5819), .A2(n8559), .ZN(n7950) );
  INV_X1 U7013 ( .A(n8940), .ZN(n8905) );
  NAND2_X1 U7014 ( .A1(n8905), .A2(n8942), .ZN(n8927) );
  INV_X1 U7015 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5434) );
  OR2_X1 U7016 ( .A1(n8942), .A2(n5434), .ZN(n5435) );
  INV_X1 U7017 ( .A(n5436), .ZN(n5437) );
  OAI21_X1 U7018 ( .B1(n5584), .B2(n8944), .A(n5437), .ZN(P2_U3486) );
  INV_X1 U7019 ( .A(n6860), .ZN(n6863) );
  NAND2_X1 U7020 ( .A1(n5927), .A2(n8540), .ZN(n5438) );
  NAND2_X1 U7021 ( .A1(n5438), .A2(n5926), .ZN(n5561) );
  NAND2_X1 U7022 ( .A1(n5561), .A2(n6497), .ZN(n5439) );
  NAND2_X1 U7023 ( .A1(n5439), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7024 ( .A(n6878), .ZN(n7228) );
  INV_X1 U7025 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9594) );
  AND2_X1 U7026 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n6959), .ZN(n5441) );
  NAND2_X1 U7027 ( .A1(n4928), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5442) );
  OAI21_X1 U7028 ( .B1(n7028), .B2(n5441), .A(n5442), .ZN(n7022) );
  NAND2_X1 U7029 ( .A1(n7020), .A2(n5442), .ZN(n7030) );
  NAND2_X1 U7030 ( .A1(n7031), .A2(n7030), .ZN(n7029) );
  OR2_X1 U7031 ( .A1(n5534), .A2(n9594), .ZN(n5443) );
  NAND2_X1 U7032 ( .A1(n7029), .A2(n5443), .ZN(n5444) );
  INV_X1 U7033 ( .A(n7084), .ZN(n6859) );
  NAND2_X1 U7034 ( .A1(n7052), .A2(n5445), .ZN(n7074) );
  NAND2_X1 U7035 ( .A1(n7072), .A2(n7052), .ZN(n5447) );
  XNOR2_X1 U7036 ( .A(n7068), .B(n5446), .ZN(n7051) );
  NAND2_X1 U7037 ( .A1(n5447), .A2(n7051), .ZN(n7055) );
  NAND2_X1 U7038 ( .A1(n7068), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7039 ( .A1(n7055), .A2(n5448), .ZN(n5449) );
  INV_X1 U7040 ( .A(n5450), .ZN(n7221) );
  MUX2_X1 U7041 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n5451), .S(n6878), .Z(n7222)
         );
  INV_X1 U7042 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7536) );
  MUX2_X1 U7043 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n4888), .S(n8587), .Z(n8599)
         );
  INV_X1 U7044 ( .A(n8599), .ZN(n5453) );
  AOI21_X1 U7045 ( .B1(n7389), .B2(n8597), .A(n5453), .ZN(n8602) );
  AND2_X1 U7046 ( .A1(n8587), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5454) );
  INV_X1 U7047 ( .A(n5456), .ZN(n5455) );
  NOR2_X1 U7048 ( .A1(n7675), .A2(n5455), .ZN(n5457) );
  MUX2_X1 U7049 ( .A(n5458), .B(P2_REG2_REG_10__SCAN_IN), .S(n7742), .Z(n7740)
         );
  INV_X1 U7050 ( .A(n7740), .ZN(n5459) );
  NAND2_X1 U7051 ( .A1(n7742), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U7052 ( .A(n7822), .B(n5461), .ZN(n7818) );
  NOR2_X1 U7053 ( .A1(n5049), .A2(n7818), .ZN(n7817) );
  NOR2_X1 U7054 ( .A1(n7822), .A2(n5461), .ZN(n5462) );
  NAND2_X1 U7055 ( .A1(n7112), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5464) );
  OR2_X1 U7056 ( .A1(n7112), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U7057 ( .A1(n5464), .A2(n5463), .ZN(n7878) );
  NOR2_X1 U7058 ( .A1(n8025), .A2(n5465), .ZN(n5466) );
  NAND2_X1 U7059 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7197), .ZN(n5467) );
  OAI21_X1 U7060 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7197), .A(n5467), .ZN(
        n8609) );
  NOR2_X1 U7061 ( .A1(n8610), .A2(n8609), .ZN(n8608) );
  AOI21_X1 U7062 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7197), .A(n8608), .ZN(
        n5468) );
  XNOR2_X1 U7063 ( .A(n5468), .B(n5522), .ZN(n8626) );
  NOR2_X1 U7064 ( .A1(n8626), .A2(n8872), .ZN(n8625) );
  NOR2_X1 U7065 ( .A1(n5522), .A2(n5468), .ZN(n5469) );
  NOR2_X1 U7066 ( .A1(n8625), .A2(n5469), .ZN(n8643) );
  INV_X1 U7067 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8855) );
  MUX2_X1 U7068 ( .A(n8855), .B(P2_REG2_REG_16__SCAN_IN), .S(n7303), .Z(n8642)
         );
  NAND2_X1 U7069 ( .A1(n7303), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5470) );
  NOR2_X1 U7070 ( .A1(n8673), .A2(n5471), .ZN(n5472) );
  INV_X1 U7071 ( .A(n8673), .ZN(n7405) );
  INV_X1 U7072 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8671) );
  NOR2_X1 U7073 ( .A1(n5472), .A2(n8669), .ZN(n8679) );
  INV_X1 U7074 ( .A(n5557), .ZN(n8691) );
  NAND2_X1 U7075 ( .A1(n8691), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5473) );
  OAI21_X1 U7076 ( .B1(n8691), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5473), .ZN(
        n8678) );
  NOR2_X1 U7077 ( .A1(n8679), .A2(n8678), .ZN(n8677) );
  INV_X1 U7078 ( .A(n5473), .ZN(n5474) );
  NOR2_X1 U7079 ( .A1(n8677), .A2(n5474), .ZN(n5475) );
  MUX2_X1 U7080 ( .A(n8814), .B(P2_REG2_REG_19__SCAN_IN), .S(n5579), .Z(n5519)
         );
  XNOR2_X1 U7081 ( .A(n5475), .B(n5519), .ZN(n5570) );
  NOR2_X1 U7082 ( .A1(n5370), .A2(P2_U3151), .ZN(n8092) );
  AND2_X1 U7083 ( .A1(n5561), .A2(n8092), .ZN(n6954) );
  INV_X1 U7084 ( .A(n6954), .ZN(n5476) );
  OR2_X1 U7085 ( .A1(n5476), .A2(n8072), .ZN(n8698) );
  INV_X1 U7086 ( .A(n5534), .ZN(n7045) );
  INV_X1 U7087 ( .A(n7028), .ZN(n5480) );
  NAND2_X1 U7088 ( .A1(n6959), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5479) );
  NOR2_X1 U7089 ( .A1(n5478), .A2(n5477), .ZN(n5481) );
  NAND2_X1 U7090 ( .A1(n7077), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7078) );
  INV_X1 U7091 ( .A(n5485), .ZN(n7056) );
  XNOR2_X1 U7092 ( .A(n7068), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7057) );
  AOI21_X1 U7093 ( .B1(n7078), .B2(n7056), .A(n7057), .ZN(n7059) );
  AOI21_X1 U7094 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7068), .A(n7059), .ZN(
        n5486) );
  INV_X1 U7095 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7552) );
  MUX2_X1 U7096 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7552), .S(n6878), .Z(n7231)
         );
  OAI21_X1 U7097 ( .B1(n7228), .B2(n7552), .A(n7229), .ZN(n5487) );
  NAND2_X1 U7098 ( .A1(n5487), .A2(n7392), .ZN(n8592) );
  NAND2_X1 U7099 ( .A1(n5488), .A2(n4502), .ZN(n5489) );
  MUX2_X1 U7100 ( .A(n5490), .B(P2_REG1_REG_8__SCAN_IN), .S(n8587), .Z(n8593)
         );
  NOR2_X1 U7101 ( .A1(n8596), .A2(n5491), .ZN(n5492) );
  XNOR2_X1 U7102 ( .A(n5492), .B(n7675), .ZN(n7662) );
  NOR2_X1 U7103 ( .A1(n7662), .A2(n5018), .ZN(n7661) );
  NOR2_X1 U7104 ( .A1(n7675), .A2(n5492), .ZN(n5493) );
  NOR2_X1 U7105 ( .A1(n7661), .A2(n5493), .ZN(n7750) );
  MUX2_X1 U7106 ( .A(n5494), .B(P2_REG1_REG_10__SCAN_IN), .S(n7742), .Z(n7749)
         );
  NAND2_X1 U7107 ( .A1(n7742), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5495) );
  INV_X1 U7108 ( .A(n5497), .ZN(n5496) );
  NOR2_X1 U7109 ( .A1(n7822), .A2(n5496), .ZN(n5498) );
  XNOR2_X1 U7110 ( .A(n5497), .B(n7050), .ZN(n7810) );
  NOR2_X1 U7111 ( .A1(n5048), .A2(n7810), .ZN(n7809) );
  NOR2_X1 U7112 ( .A1(n5498), .A2(n7809), .ZN(n7887) );
  NAND2_X1 U7113 ( .A1(n7112), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5500) );
  OR2_X1 U7114 ( .A1(n7112), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7115 ( .A1(n5500), .A2(n5499), .ZN(n7886) );
  OR2_X1 U7116 ( .A1(n7887), .A2(n7886), .ZN(n7889) );
  NAND2_X1 U7117 ( .A1(n7889), .A2(n5500), .ZN(n5501) );
  XNOR2_X1 U7118 ( .A(n5501), .B(n7141), .ZN(n8012) );
  INV_X1 U7119 ( .A(n5501), .ZN(n5502) );
  NOR2_X1 U7120 ( .A1(n8025), .A2(n5502), .ZN(n5503) );
  NAND2_X1 U7121 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7197), .ZN(n5504) );
  OAI21_X1 U7122 ( .B1(n7197), .B2(P2_REG1_REG_14__SCAN_IN), .A(n5504), .ZN(
        n8618) );
  NOR2_X1 U7123 ( .A1(n5522), .A2(n5507), .ZN(n5508) );
  NAND2_X1 U7124 ( .A1(n7303), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5509) );
  OAI21_X1 U7125 ( .B1(n7303), .B2(P2_REG1_REG_16__SCAN_IN), .A(n5509), .ZN(
        n8651) );
  INV_X1 U7126 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8917) );
  INV_X1 U7127 ( .A(n5510), .ZN(n5511) );
  NOR2_X1 U7128 ( .A1(n8673), .A2(n5511), .ZN(n5512) );
  NAND2_X1 U7129 ( .A1(n8691), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5513) );
  OAI21_X1 U7130 ( .B1(n8691), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5513), .ZN(
        n8681) );
  INV_X1 U7131 ( .A(n5513), .ZN(n5514) );
  NOR2_X1 U7132 ( .A1(n8680), .A2(n5514), .ZN(n5516) );
  XNOR2_X1 U7133 ( .A(n5579), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5518) );
  XNOR2_X1 U7134 ( .A(n5516), .B(n5515), .ZN(n5517) );
  AND2_X1 U7135 ( .A1(n6954), .A2(n8072), .ZN(n8697) );
  NAND2_X1 U7136 ( .A1(n5517), .A2(n8697), .ZN(n5569) );
  MUX2_X1 U7137 ( .A(n5519), .B(n5518), .S(n8072), .Z(n5559) );
  MUX2_X1 U7138 ( .A(n8671), .B(n8917), .S(n8072), .Z(n5554) );
  XNOR2_X1 U7139 ( .A(n7405), .B(n5554), .ZN(n8664) );
  INV_X1 U7140 ( .A(n7303), .ZN(n8657) );
  INV_X1 U7141 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8920) );
  MUX2_X1 U7142 ( .A(n8855), .B(n8920), .S(n8072), .Z(n5520) );
  NAND2_X1 U7143 ( .A1(n8657), .A2(n5520), .ZN(n5553) );
  XNOR2_X1 U7144 ( .A(n5520), .B(n7303), .ZN(n8647) );
  MUX2_X1 U7145 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8072), .Z(n5521) );
  OR2_X1 U7146 ( .A1(n5521), .A2(n5505), .ZN(n5552) );
  XNOR2_X1 U7147 ( .A(n5522), .B(n5521), .ZN(n8629) );
  MUX2_X1 U7148 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8072), .Z(n5523) );
  OR2_X1 U7149 ( .A1(n5523), .A2(n7197), .ZN(n5551) );
  INV_X1 U7150 ( .A(n7197), .ZN(n8622) );
  XNOR2_X1 U7151 ( .A(n5523), .B(n8622), .ZN(n8613) );
  MUX2_X1 U7152 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8072), .Z(n5524) );
  OR2_X1 U7153 ( .A1(n5524), .A2(n7141), .ZN(n5550) );
  XNOR2_X1 U7154 ( .A(n5524), .B(n8025), .ZN(n8016) );
  MUX2_X1 U7155 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8072), .Z(n5525) );
  OR2_X1 U7156 ( .A1(n5525), .A2(n7112), .ZN(n5549) );
  INV_X1 U7157 ( .A(n7112), .ZN(n7892) );
  XNOR2_X1 U7158 ( .A(n5525), .B(n7892), .ZN(n7882) );
  MUX2_X1 U7159 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8072), .Z(n5526) );
  OR2_X1 U7160 ( .A1(n5526), .A2(n7050), .ZN(n5548) );
  XNOR2_X1 U7161 ( .A(n5526), .B(n7822), .ZN(n7813) );
  MUX2_X1 U7162 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8072), .Z(n5527) );
  OR2_X1 U7163 ( .A1(n5527), .A2(n7742), .ZN(n5547) );
  XOR2_X1 U7164 ( .A(n7742), .B(n5527), .Z(n7745) );
  MUX2_X1 U7165 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8072), .Z(n5528) );
  OR2_X1 U7166 ( .A1(n5528), .A2(n6909), .ZN(n5546) );
  XNOR2_X1 U7167 ( .A(n5528), .B(n7675), .ZN(n7666) );
  MUX2_X1 U7168 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8072), .Z(n5544) );
  OR2_X1 U7169 ( .A1(n5544), .A2(n8587), .ZN(n5545) );
  MUX2_X1 U7170 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8072), .Z(n5541) );
  INV_X1 U7171 ( .A(n5541), .ZN(n5542) );
  MUX2_X1 U7172 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8072), .Z(n5539) );
  INV_X1 U7173 ( .A(n5539), .ZN(n5540) );
  INV_X1 U7174 ( .A(n7068), .ZN(n5538) );
  MUX2_X1 U7175 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8072), .Z(n5536) );
  INV_X1 U7176 ( .A(n5536), .ZN(n5537) );
  MUX2_X1 U7177 ( .A(n5530), .B(n5529), .S(n8072), .Z(n5535) );
  MUX2_X1 U7178 ( .A(n9594), .B(n5482), .S(n8072), .Z(n5533) );
  MUX2_X1 U7179 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8072), .Z(n5531) );
  INV_X1 U7180 ( .A(n5531), .ZN(n5532) );
  MUX2_X1 U7181 ( .A(n4933), .B(n5477), .S(n8072), .Z(n6952) );
  XNOR2_X1 U7182 ( .A(n5533), .B(n7045), .ZN(n7041) );
  OAI21_X1 U7183 ( .B1(n5534), .B2(n5533), .A(n7040), .ZN(n7070) );
  XNOR2_X1 U7184 ( .A(n5535), .B(n7084), .ZN(n7071) );
  NOR2_X1 U7185 ( .A1(n7070), .A2(n7071), .ZN(n7069) );
  AOI21_X1 U7186 ( .B1(n7084), .B2(n5535), .A(n7069), .ZN(n7065) );
  XOR2_X1 U7187 ( .A(n7068), .B(n5536), .Z(n7064) );
  NAND2_X1 U7188 ( .A1(n7065), .A2(n7064), .ZN(n7063) );
  XNOR2_X1 U7189 ( .A(n5539), .B(n4495), .ZN(n7130) );
  XNOR2_X1 U7190 ( .A(n5541), .B(n6878), .ZN(n7219) );
  AOI21_X1 U7191 ( .B1(n7228), .B2(n5542), .A(n7217), .ZN(n7388) );
  MUX2_X1 U7192 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8072), .Z(n5543) );
  XNOR2_X1 U7193 ( .A(n5543), .B(n7392), .ZN(n7387) );
  OAI22_X1 U7194 ( .A1(n7388), .A2(n7387), .B1(n5543), .B2(n7392), .ZN(n8585)
         );
  XOR2_X1 U7195 ( .A(n8587), .B(n5544), .Z(n8584) );
  NAND2_X1 U7196 ( .A1(n8585), .A2(n8584), .ZN(n8583) );
  NAND2_X1 U7197 ( .A1(n5547), .A2(n7743), .ZN(n7812) );
  NAND2_X1 U7198 ( .A1(n8016), .A2(n8015), .ZN(n8014) );
  NAND2_X1 U7199 ( .A1(n5550), .A2(n8014), .ZN(n8612) );
  NAND2_X1 U7200 ( .A1(n8647), .A2(n8646), .ZN(n8645) );
  NAND2_X1 U7201 ( .A1(n5553), .A2(n8645), .ZN(n8663) );
  NAND2_X1 U7202 ( .A1(n8664), .A2(n8663), .ZN(n8662) );
  MUX2_X1 U7203 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8072), .Z(n5555) );
  NOR2_X1 U7204 ( .A1(n5556), .A2(n5555), .ZN(n8685) );
  AOI21_X1 U7205 ( .B1(n5557), .B2(n8683), .A(n8685), .ZN(n5558) );
  XNOR2_X1 U7206 ( .A(n5559), .B(n5558), .ZN(n5560) );
  NAND2_X1 U7207 ( .A1(P2_U3893), .A2(n5370), .ZN(n8689) );
  NOR2_X1 U7208 ( .A1(n5560), .A2(n8689), .ZN(n5567) );
  AND2_X1 U7209 ( .A1(n5561), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5562) );
  INV_X1 U7210 ( .A(n5370), .ZN(n8556) );
  MUX2_X1 U7211 ( .A(n5562), .B(P2_U3893), .S(n8556), .Z(n5563) );
  NAND2_X1 U7212 ( .A1(n5563), .A2(n6497), .ZN(n8686) );
  NAND2_X1 U7213 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8215) );
  INV_X1 U7214 ( .A(n5926), .ZN(n7761) );
  NOR2_X1 U7215 ( .A1(n5927), .A2(n7761), .ZN(n5564) );
  OR2_X1 U7216 ( .A1(P2_U3150), .A2(n5564), .ZN(n8695) );
  INV_X1 U7217 ( .A(n8695), .ZN(n7394) );
  NAND2_X1 U7218 ( .A1(n7394), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5565) );
  OAI211_X1 U7219 ( .C1(n8686), .C2(n8373), .A(n8215), .B(n5565), .ZN(n5566)
         );
  OAI211_X1 U7220 ( .C1(n5570), .C2(n8698), .A(n5569), .B(n5568), .ZN(P2_U3201) );
  INV_X1 U7221 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7222 ( .A1(n5571), .A2(n5574), .ZN(n5925) );
  INV_X1 U7223 ( .A(n5919), .ZN(n5935) );
  NOR2_X1 U7224 ( .A1(n5925), .A2(n5935), .ZN(n5918) );
  NAND2_X1 U7225 ( .A1(n8554), .A2(n8559), .ZN(n5577) );
  NOR2_X1 U7226 ( .A1(n5577), .A2(n8371), .ZN(n5572) );
  NAND2_X1 U7227 ( .A1(n5579), .A2(n5572), .ZN(n5929) );
  NAND2_X1 U7228 ( .A1(n5936), .A2(n5929), .ZN(n5573) );
  NAND2_X1 U7229 ( .A1(n5918), .A2(n5573), .ZN(n5583) );
  NAND2_X1 U7230 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  NOR2_X1 U7231 ( .A1(n5576), .A2(n7239), .ZN(n5937) );
  NAND2_X1 U7232 ( .A1(n5937), .A2(n5919), .ZN(n5924) );
  NAND2_X1 U7233 ( .A1(n5819), .A2(n8915), .ZN(n9738) );
  INV_X1 U7234 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7235 ( .A1(n5579), .A2(n5578), .ZN(n5581) );
  NOR2_X1 U7236 ( .A1(n8915), .A2(n8547), .ZN(n5580) );
  NAND2_X1 U7237 ( .A1(n5581), .A2(n5580), .ZN(n5912) );
  AND2_X1 U7238 ( .A1(n9738), .A2(n5912), .ZN(n5932) );
  OR2_X1 U7239 ( .A1(n5924), .A2(n5932), .ZN(n5582) );
  INV_X2 U7240 ( .A(n10060), .ZN(n10057) );
  MUX2_X1 U7241 ( .A(n5585), .B(n5584), .S(n10057), .Z(n5587) );
  OR2_X1 U7242 ( .A1(n10060), .A2(n8940), .ZN(n9014) );
  NAND2_X1 U7243 ( .A1(n5587), .A2(n5586), .ZN(P2_U3454) );
  INV_X1 U7244 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5588) );
  INV_X1 U7245 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8151) );
  MUX2_X1 U7246 ( .A(n5588), .B(n8151), .S(n6853), .Z(n5591) );
  INV_X1 U7247 ( .A(SI_28_), .ZN(n5589) );
  NAND2_X1 U7248 ( .A1(n5591), .A2(n5589), .ZN(n5590) );
  AND2_X1 U7249 ( .A1(n5740), .A2(n5590), .ZN(n5593) );
  INV_X1 U7250 ( .A(n5590), .ZN(n5592) );
  XNOR2_X1 U7251 ( .A(n5591), .B(SI_28_), .ZN(n5741) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8154) );
  INV_X1 U7253 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9607) );
  MUX2_X1 U7254 ( .A(n8154), .B(n9607), .S(n6853), .Z(n5748) );
  NAND4_X1 U7255 ( .A1(n5660), .A2(n5597), .A3(n5596), .A4(n5595), .ZN(n5600)
         );
  NOR2_X1 U7256 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5607) );
  INV_X1 U7257 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5610) );
  INV_X1 U7258 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5770) );
  NAND2_X2 U7259 ( .A1(n5621), .A2(n6853), .ZN(n5643) );
  INV_X2 U7260 ( .A(n5643), .ZN(n5756) );
  NAND2_X1 U7261 ( .A1(n8153), .A2(n5756), .ZN(n5613) );
  NAND2_X1 U7262 ( .A1(n5621), .A2(n5611), .ZN(n5620) );
  OR2_X1 U7263 ( .A1(n5735), .A2(n9607), .ZN(n5612) );
  NAND2_X1 U7264 ( .A1(n8071), .A2(n5756), .ZN(n5615) );
  OR2_X1 U7265 ( .A1(n5735), .A2(n8164), .ZN(n5614) );
  OR2_X1 U7266 ( .A1(n5643), .A2(n6869), .ZN(n5617) );
  OR2_X1 U7267 ( .A1(n4276), .A2(n6870), .ZN(n5616) );
  XNOR2_X1 U7268 ( .A(n5619), .B(n5618), .ZN(n6849) );
  MUX2_X1 U7269 ( .A(n5599), .B(n6849), .S(n5621), .Z(n9902) );
  NAND2_X1 U7270 ( .A1(n6701), .A2(n9902), .ZN(n9900) );
  OR2_X1 U7271 ( .A1(n5643), .A2(n6867), .ZN(n5629) );
  OR2_X1 U7272 ( .A1(n5620), .A2(n6868), .ZN(n5628) );
  INV_X1 U7273 ( .A(n5624), .ZN(n5622) );
  NAND2_X1 U7274 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5622), .ZN(n5623) );
  INV_X1 U7275 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5625) );
  MUX2_X1 U7276 ( .A(n5623), .B(P1_IR_REG_31__SCAN_IN), .S(n5625), .Z(n5626)
         );
  NAND2_X1 U7277 ( .A1(n5625), .A2(n5624), .ZN(n5631) );
  OR2_X1 U7278 ( .A1(n5621), .A2(n7193), .ZN(n5627) );
  NAND2_X1 U7279 ( .A1(n5631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5632) );
  XNOR2_X1 U7280 ( .A(n5632), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6934) );
  INV_X1 U7281 ( .A(n6934), .ZN(n6979) );
  OR2_X1 U7282 ( .A1(n5643), .A2(n6858), .ZN(n5634) );
  OR2_X1 U7283 ( .A1(n5620), .A2(n6851), .ZN(n5633) );
  OAI211_X1 U7284 ( .C1(n5621), .C2(n6979), .A(n5634), .B(n5633), .ZN(n9870)
         );
  OR2_X1 U7285 ( .A1(n5620), .A2(n6852), .ZN(n5640) );
  NAND2_X1 U7286 ( .A1(n5635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5636) );
  MUX2_X1 U7287 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5636), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5638) );
  NOR2_X1 U7288 ( .A1(n5635), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5647) );
  INV_X1 U7289 ( .A(n5647), .ZN(n5637) );
  NAND2_X1 U7290 ( .A1(n5638), .A2(n5637), .ZN(n9797) );
  OR2_X1 U7291 ( .A1(n5621), .A2(n9797), .ZN(n5639) );
  INV_X1 U7292 ( .A(n7485), .ZN(n9937) );
  OR2_X1 U7293 ( .A1(n5647), .A2(n9670), .ZN(n5642) );
  XNOR2_X1 U7294 ( .A(n5642), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6986) );
  INV_X1 U7295 ( .A(n6986), .ZN(n6872) );
  OR2_X1 U7296 ( .A1(n5643), .A2(n6873), .ZN(n5645) );
  INV_X1 U7297 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6871) );
  OR2_X1 U7298 ( .A1(n5735), .A2(n6871), .ZN(n5644) );
  OAI211_X1 U7299 ( .C1(n5621), .C2(n6872), .A(n5645), .B(n5644), .ZN(n9859)
         );
  INV_X1 U7300 ( .A(n9859), .ZN(n9945) );
  NAND2_X1 U7301 ( .A1(n5756), .A2(n6874), .ZN(n5654) );
  INV_X1 U7302 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5646) );
  AND2_X1 U7303 ( .A1(n5647), .A2(n5646), .ZN(n5661) );
  OR2_X1 U7304 ( .A1(n5661), .A2(n9670), .ZN(n5650) );
  INV_X1 U7305 ( .A(n5650), .ZN(n5648) );
  NAND2_X1 U7306 ( .A1(n5648), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5651) );
  INV_X1 U7307 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7308 ( .A1(n5650), .A2(n5649), .ZN(n5656) );
  AND2_X1 U7309 ( .A1(n5651), .A2(n5656), .ZN(n7001) );
  INV_X1 U7310 ( .A(n7001), .ZN(n7005) );
  OR2_X1 U7311 ( .A1(n5621), .A2(n7005), .ZN(n5653) );
  OR2_X1 U7312 ( .A1(n5735), .A2(n6875), .ZN(n5652) );
  NAND2_X1 U7313 ( .A1(n5656), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5657) );
  XNOR2_X1 U7314 ( .A(n5657), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7099) );
  AOI22_X1 U7315 ( .A1(n5720), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5719), .B2(
        n7099), .ZN(n5659) );
  NAND2_X1 U7316 ( .A1(n6879), .A2(n5756), .ZN(n5658) );
  NAND2_X1 U7317 ( .A1(n6900), .A2(n5756), .ZN(n5664) );
  AND2_X1 U7318 ( .A1(n5661), .A2(n5660), .ZN(n5666) );
  OR2_X1 U7319 ( .A1(n5666), .A2(n9670), .ZN(n5662) );
  XNOR2_X1 U7320 ( .A(n5662), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7158) );
  AOI22_X1 U7321 ( .A1(n5720), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5719), .B2(
        n7158), .ZN(n5663) );
  INV_X1 U7322 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7323 ( .A1(n5666), .A2(n5665), .ZN(n5670) );
  NAND2_X1 U7324 ( .A1(n5670), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5667) );
  XNOR2_X1 U7325 ( .A(n5667), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7291) );
  AOI22_X1 U7326 ( .A1(n5720), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5719), .B2(
        n7291), .ZN(n5668) );
  INV_X1 U7327 ( .A(n9976), .ZN(n9830) );
  NAND2_X1 U7328 ( .A1(n6918), .A2(n5756), .ZN(n5673) );
  OR2_X1 U7329 ( .A1(n5670), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7330 ( .A1(n5671), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5677) );
  INV_X1 U7331 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U7332 ( .A(n5677), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7429) );
  AOI22_X1 U7333 ( .A1(n5720), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5719), .B2(
        n7429), .ZN(n5672) );
  NAND2_X1 U7334 ( .A1(n5673), .A2(n5672), .ZN(n7687) );
  NAND2_X1 U7335 ( .A1(n7046), .A2(n5756), .ZN(n5681) );
  NAND2_X1 U7336 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  NAND2_X1 U7337 ( .A1(n5678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U7338 ( .A(n5679), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7603) );
  AOI22_X1 U7339 ( .A1(n5720), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5719), .B2(
        n7603), .ZN(n5680) );
  NAND2_X1 U7340 ( .A1(n7087), .A2(n5756), .ZN(n5684) );
  OR2_X1 U7341 ( .A1(n5686), .A2(n9670), .ZN(n5682) );
  XNOR2_X1 U7342 ( .A(n5682), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7620) );
  AOI22_X1 U7343 ( .A1(n5720), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5719), .B2(
        n7620), .ZN(n5683) );
  INV_X1 U7344 ( .A(n7768), .ZN(n8038) );
  NAND2_X1 U7345 ( .A1(n7138), .A2(n5756), .ZN(n5689) );
  INV_X1 U7346 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5685) );
  OR2_X1 U7347 ( .A1(n5691), .A2(n9670), .ZN(n5687) );
  XNOR2_X1 U7348 ( .A(n5687), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7707) );
  AOI22_X1 U7349 ( .A1(n5720), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5719), .B2(
        n7707), .ZN(n5688) );
  INV_X1 U7350 ( .A(n8089), .ZN(n7930) );
  NAND2_X1 U7351 ( .A1(n7195), .A2(n5756), .ZN(n5693) );
  INV_X1 U7352 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5690) );
  OR2_X1 U7353 ( .A1(n5701), .A2(n9670), .ZN(n5695) );
  XNOR2_X1 U7354 ( .A(n5695), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7980) );
  AOI22_X1 U7355 ( .A1(n5720), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5719), .B2(
        n7980), .ZN(n5692) );
  NAND2_X1 U7356 ( .A1(n7252), .A2(n5756), .ZN(n5699) );
  INV_X1 U7357 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7358 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  NAND2_X1 U7359 ( .A1(n5696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5697) );
  XNOR2_X1 U7360 ( .A(n5697), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9182) );
  AOI22_X1 U7361 ( .A1(n5720), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5719), .B2(
        n9182), .ZN(n5698) );
  NAND2_X1 U7362 ( .A1(n7301), .A2(n5756), .ZN(n5706) );
  NOR2_X1 U7363 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5700) );
  NAND2_X1 U7364 ( .A1(n5701), .A2(n5700), .ZN(n5703) );
  NAND2_X1 U7365 ( .A1(n5703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5702) );
  MUX2_X1 U7366 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5702), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5704) );
  AND2_X1 U7367 ( .A1(n5704), .A2(n4334), .ZN(n9196) );
  AOI22_X1 U7368 ( .A1(n5720), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5719), .B2(
        n9196), .ZN(n5705) );
  NAND2_X1 U7369 ( .A1(n7403), .A2(n5756), .ZN(n5709) );
  NAND2_X1 U7370 ( .A1(n4334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5707) );
  XNOR2_X1 U7371 ( .A(n5707), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9222) );
  AOI22_X1 U7372 ( .A1(n5720), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5719), .B2(
        n9222), .ZN(n5708) );
  NAND2_X1 U7373 ( .A1(n8125), .A2(n9082), .ZN(n8139) );
  NAND2_X1 U7374 ( .A1(n7409), .A2(n5756), .ZN(n5715) );
  INV_X1 U7375 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5711) );
  OR2_X1 U7376 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  AND2_X1 U7377 ( .A1(n5716), .A2(n5713), .ZN(n9235) );
  AOI22_X1 U7378 ( .A1(n5720), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5719), .B2(
        n9235), .ZN(n5714) );
  NAND2_X1 U7379 ( .A1(n7499), .A2(n5756), .ZN(n5722) );
  INV_X1 U7380 ( .A(n5804), .ZN(n6219) );
  AOI22_X1 U7381 ( .A1(n5720), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6219), .B2(
        n5719), .ZN(n5721) );
  NAND2_X1 U7382 ( .A1(n7522), .A2(n5756), .ZN(n5724) );
  OR2_X1 U7383 ( .A1(n5735), .A2(n7523), .ZN(n5723) );
  NAND2_X1 U7384 ( .A1(n5725), .A2(n5756), .ZN(n5727) );
  INV_X1 U7385 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n9514) );
  OR2_X1 U7386 ( .A1(n5735), .A2(n9514), .ZN(n5726) );
  NAND2_X1 U7387 ( .A1(n7771), .A2(n5756), .ZN(n5729) );
  OR2_X1 U7388 ( .A1(n5735), .A2(n9604), .ZN(n5728) );
  NAND2_X1 U7389 ( .A1(n7758), .A2(n5756), .ZN(n5732) );
  OR2_X1 U7390 ( .A1(n5735), .A2(n5730), .ZN(n5731) );
  NAND2_X1 U7391 ( .A1(n7910), .A2(n5756), .ZN(n5734) );
  OR2_X1 U7392 ( .A1(n5735), .A2(n7912), .ZN(n5733) );
  NAND2_X1 U7393 ( .A1(n7966), .A2(n5756), .ZN(n5737) );
  OR2_X1 U7394 ( .A1(n5735), .A2(n9517), .ZN(n5736) );
  NAND2_X1 U7395 ( .A1(n8039), .A2(n5756), .ZN(n5739) );
  OR2_X1 U7396 ( .A1(n5735), .A2(n8040), .ZN(n5738) );
  OR2_X1 U7397 ( .A1(n5735), .A2(n8151), .ZN(n5743) );
  INV_X1 U7398 ( .A(n5745), .ZN(n5746) );
  NAND2_X1 U7399 ( .A1(n5746), .A2(SI_29_), .ZN(n5751) );
  INV_X1 U7400 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U7401 ( .A1(n4622), .A2(n5749), .ZN(n5750) );
  NAND2_X1 U7402 ( .A1(n5751), .A2(n5750), .ZN(n6507) );
  INV_X1 U7403 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9022) );
  INV_X1 U7404 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8193) );
  MUX2_X1 U7405 ( .A(n9022), .B(n8193), .S(n6853), .Z(n5753) );
  INV_X1 U7406 ( .A(SI_30_), .ZN(n5752) );
  NAND2_X1 U7407 ( .A1(n5753), .A2(n5752), .ZN(n6505) );
  INV_X1 U7408 ( .A(n5753), .ZN(n5754) );
  NAND2_X1 U7409 ( .A1(n5754), .A2(SI_30_), .ZN(n5755) );
  NAND2_X1 U7410 ( .A1(n6505), .A2(n5755), .ZN(n6506) );
  OR2_X1 U7411 ( .A1(n5735), .A2(n8193), .ZN(n5757) );
  NAND2_X1 U7412 ( .A1(n4320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5761) );
  INV_X1 U7413 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7414 ( .A1(n5764), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5765) );
  XNOR2_X1 U7415 ( .A(n5765), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6655) );
  INV_X1 U7416 ( .A(n6655), .ZN(n7643) );
  AND2_X1 U7417 ( .A1(n7772), .A2(n7643), .ZN(n7136) );
  NAND2_X1 U7418 ( .A1(n5766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5767) );
  XNOR2_X1 U7419 ( .A(n5767), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6742) );
  INV_X1 U7420 ( .A(n9901), .ZN(n9425) );
  INV_X1 U7421 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7422 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5772) );
  NAND2_X1 U7423 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  XNOR2_X2 U7424 ( .A(n5774), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5775) );
  INV_X1 U7425 ( .A(n5775), .ZN(n5977) );
  INV_X1 U7426 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U7427 ( .A1(n6248), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5777) );
  AND2_X2 U7428 ( .A1(n8192), .A2(n5775), .ZN(n5994) );
  NAND2_X1 U7429 ( .A1(n5994), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5776) );
  OAI211_X1 U7430 ( .C1(n6197), .C2(n6527), .A(n5777), .B(n5776), .ZN(n6915)
         );
  INV_X1 U7431 ( .A(n5778), .ZN(n7182) );
  NOR2_X1 U7432 ( .A1(n7772), .A2(n7643), .ZN(n6911) );
  NAND2_X1 U7433 ( .A1(n5778), .A2(n6911), .ZN(n9129) );
  INV_X1 U7434 ( .A(P1_B_REG_SCAN_IN), .ZN(n5786) );
  NOR2_X1 U7435 ( .A1(n5779), .A2(n5786), .ZN(n5780) );
  OR2_X1 U7436 ( .A1(n9129), .A2(n5780), .ZN(n6253) );
  INV_X1 U7437 ( .A(n6253), .ZN(n5781) );
  AND2_X1 U7438 ( .A1(n6915), .A2(n5781), .ZN(n6518) );
  INV_X1 U7439 ( .A(n6518), .ZN(n8185) );
  NAND2_X1 U7440 ( .A1(n9250), .A2(n8185), .ZN(n9435) );
  NAND2_X1 U7441 ( .A1(n4324), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5782) );
  XNOR2_X1 U7442 ( .A(n5782), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5807) );
  NOR2_X1 U7443 ( .A1(n5807), .A2(n5786), .ZN(n5787) );
  NAND2_X1 U7444 ( .A1(n5783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5784) );
  MUX2_X1 U7445 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5784), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5785) );
  AND2_X1 U7446 ( .A1(n5785), .A2(n4324), .ZN(n7911) );
  MUX2_X1 U7447 ( .A(n5787), .B(n5786), .S(n7911), .Z(n5790) );
  NAND2_X1 U7448 ( .A1(n5788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5789) );
  XNOR2_X1 U7449 ( .A(n5789), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5810) );
  INV_X1 U7450 ( .A(n5810), .ZN(n8041) );
  NOR4_X1 U7451 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5799) );
  NOR4_X1 U7452 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5798) );
  INV_X1 U7453 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9912) );
  INV_X1 U7454 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9911) );
  INV_X1 U7455 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9914) );
  INV_X1 U7456 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9910) );
  NAND4_X1 U7457 ( .A1(n9912), .A2(n9911), .A3(n9914), .A4(n9910), .ZN(n5796)
         );
  NOR4_X1 U7458 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5794) );
  NOR4_X1 U7459 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5793) );
  NOR4_X1 U7460 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5792) );
  NOR4_X1 U7461 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5791) );
  NAND4_X1 U7462 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(n5795)
         );
  NOR4_X1 U7463 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n5796), .A4(n5795), .ZN(n5797) );
  AND3_X1 U7464 ( .A1(n5799), .A2(n5798), .A3(n5797), .ZN(n5800) );
  NOR2_X1 U7465 ( .A1(n6897), .A2(n5800), .ZN(n6463) );
  INV_X1 U7466 ( .A(n6463), .ZN(n5809) );
  NAND2_X1 U7467 ( .A1(n5801), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5803) );
  INV_X1 U7468 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U7469 ( .A(n5803), .B(n5802), .ZN(n6910) );
  AND2_X1 U7470 ( .A1(n6910), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6845) );
  NAND2_X1 U7471 ( .A1(n6847), .A2(n6845), .ZN(n6913) );
  INV_X1 U7472 ( .A(n6913), .ZN(n6896) );
  NAND2_X1 U7473 ( .A1(n6768), .A2(n6911), .ZN(n5805) );
  NAND2_X1 U7474 ( .A1(n6896), .A2(n5805), .ZN(n7354) );
  NAND2_X1 U7475 ( .A1(n6219), .A2(n9901), .ZN(n6467) );
  INV_X1 U7476 ( .A(n6467), .ZN(n5806) );
  NOR2_X1 U7477 ( .A1(n7354), .A2(n5806), .ZN(n5808) );
  INV_X1 U7478 ( .A(n5807), .ZN(n7967) );
  NAND2_X1 U7479 ( .A1(n8041), .A2(n7967), .ZN(n9669) );
  OAI21_X1 U7480 ( .B1(n6897), .B2(P1_D_REG_1__SCAN_IN), .A(n9669), .ZN(n6464)
         );
  NAND3_X1 U7481 ( .A1(n5809), .A2(n5808), .A3(n6464), .ZN(n6525) );
  INV_X1 U7482 ( .A(n6897), .ZN(n5812) );
  INV_X1 U7483 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5811) );
  NOR2_X1 U7484 ( .A1(n5810), .A2(n7911), .ZN(n6899) );
  AOI21_X1 U7485 ( .B1(n5812), .B2(n5811), .A(n6899), .ZN(n6524) );
  NAND2_X1 U7486 ( .A1(n9998), .A2(n5813), .ZN(n5814) );
  NAND2_X1 U7487 ( .A1(n5815), .A2(n5814), .ZN(n5818) );
  INV_X2 U7488 ( .A(n9998), .ZN(n10000) );
  NAND2_X1 U7489 ( .A1(n6768), .A2(n7136), .ZN(n9991) );
  INV_X1 U7490 ( .A(n9991), .ZN(n9977) );
  NAND2_X1 U7491 ( .A1(n10000), .A2(n9977), .ZN(n9667) );
  NAND2_X1 U7492 ( .A1(n5818), .A2(n5817), .ZN(P1_U3520) );
  NAND2_X1 U7493 ( .A1(n5819), .A2(n8390), .ZN(n5821) );
  NAND2_X1 U7494 ( .A1(n7544), .A2(n8371), .ZN(n5820) );
  NAND2_X1 U7495 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  INV_X2 U7496 ( .A(n5827), .ZN(n5846) );
  INV_X1 U7497 ( .A(n7257), .ZN(n7114) );
  NAND2_X1 U7498 ( .A1(n8225), .A2(n7114), .ZN(n5823) );
  NAND2_X1 U7499 ( .A1(n5823), .A2(n8391), .ZN(n7167) );
  XNOR2_X1 U7500 ( .A(n5827), .B(n7170), .ZN(n5824) );
  XNOR2_X1 U7501 ( .A(n5824), .B(n8582), .ZN(n7168) );
  NAND2_X1 U7502 ( .A1(n7167), .A2(n7168), .ZN(n5826) );
  NAND2_X1 U7503 ( .A1(n5824), .A2(n7272), .ZN(n5825) );
  NAND2_X1 U7504 ( .A1(n5826), .A2(n5825), .ZN(n7147) );
  INV_X1 U7505 ( .A(n7269), .ZN(n8402) );
  XNOR2_X1 U7506 ( .A(n8402), .B(n5827), .ZN(n5828) );
  XNOR2_X1 U7507 ( .A(n5828), .B(n8581), .ZN(n7148) );
  NAND2_X1 U7508 ( .A1(n7147), .A2(n7148), .ZN(n5830) );
  NAND2_X1 U7509 ( .A1(n5828), .A2(n7323), .ZN(n5829) );
  NAND2_X1 U7510 ( .A1(n5830), .A2(n5829), .ZN(n7342) );
  INV_X1 U7511 ( .A(n7342), .ZN(n5832) );
  XNOR2_X1 U7512 ( .A(n5833), .B(n7271), .ZN(n7343) );
  INV_X1 U7513 ( .A(n7343), .ZN(n5831) );
  NAND2_X1 U7514 ( .A1(n5832), .A2(n5831), .ZN(n7340) );
  INV_X1 U7515 ( .A(n5833), .ZN(n5834) );
  NAND2_X1 U7516 ( .A1(n5834), .A2(n8580), .ZN(n5835) );
  NAND2_X1 U7517 ( .A1(n7340), .A2(n5835), .ZN(n7308) );
  XNOR2_X1 U7518 ( .A(n8225), .B(n7424), .ZN(n5837) );
  XNOR2_X1 U7519 ( .A(n5837), .B(n8410), .ZN(n7309) );
  NAND2_X1 U7520 ( .A1(n5837), .A2(n8410), .ZN(n5838) );
  XNOR2_X1 U7521 ( .A(n8225), .B(n7495), .ZN(n5839) );
  XNOR2_X1 U7522 ( .A(n5839), .B(n8578), .ZN(n7411) );
  INV_X1 U7523 ( .A(n8578), .ZN(n7549) );
  NAND2_X1 U7524 ( .A1(n5839), .A2(n7549), .ZN(n5840) );
  NAND2_X1 U7525 ( .A1(n5841), .A2(n5840), .ZN(n7575) );
  INV_X1 U7526 ( .A(n7575), .ZN(n5843) );
  XNOR2_X1 U7527 ( .A(n8225), .B(n7581), .ZN(n5844) );
  XNOR2_X1 U7528 ( .A(n5844), .B(n8577), .ZN(n7578) );
  NAND2_X1 U7529 ( .A1(n5844), .A2(n8577), .ZN(n5845) );
  XNOR2_X1 U7530 ( .A(n7538), .B(n5906), .ZN(n5847) );
  XNOR2_X1 U7531 ( .A(n5847), .B(n7637), .ZN(n7512) );
  INV_X1 U7532 ( .A(n5847), .ZN(n5848) );
  XNOR2_X1 U7533 ( .A(n7646), .B(n8225), .ZN(n5849) );
  XNOR2_X1 U7534 ( .A(n5849), .B(n7517), .ZN(n7610) );
  NAND2_X1 U7535 ( .A1(n7611), .A2(n7610), .ZN(n5852) );
  INV_X1 U7536 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U7537 ( .A1(n5850), .A2(n7517), .ZN(n5851) );
  NAND2_X1 U7538 ( .A1(n5852), .A2(n5851), .ZN(n7652) );
  XNOR2_X1 U7539 ( .A(n7696), .B(n5906), .ZN(n5853) );
  XNOR2_X1 U7540 ( .A(n5853), .B(n7825), .ZN(n7653) );
  INV_X1 U7541 ( .A(n5853), .ZN(n5854) );
  NAND2_X1 U7542 ( .A1(n5854), .A2(n8574), .ZN(n5855) );
  XNOR2_X1 U7543 ( .A(n7940), .B(n8572), .ZN(n8348) );
  XNOR2_X1 U7544 ( .A(n8348), .B(n5906), .ZN(n7871) );
  XNOR2_X1 U7545 ( .A(n7954), .B(n8225), .ZN(n7868) );
  NAND2_X1 U7546 ( .A1(n5846), .A2(n8573), .ZN(n5858) );
  OAI22_X1 U7547 ( .A1(n7954), .A2(n5858), .B1(n8044), .B2(n5846), .ZN(n5862)
         );
  NAND2_X1 U7548 ( .A1(n5846), .A2(n8572), .ZN(n5860) );
  NAND3_X1 U7549 ( .A1(n7954), .A2(n8573), .A3(n8225), .ZN(n5859) );
  NAND3_X1 U7550 ( .A1(n8348), .A2(n5860), .A3(n5859), .ZN(n5861) );
  OAI21_X1 U7551 ( .B1(n8348), .B2(n5862), .A(n5861), .ZN(n5863) );
  NAND2_X1 U7552 ( .A1(n5864), .A2(n5863), .ZN(n7834) );
  XNOR2_X1 U7553 ( .A(n8449), .B(n5906), .ZN(n5865) );
  XNOR2_X1 U7554 ( .A(n5865), .B(n8571), .ZN(n7833) );
  NAND2_X1 U7555 ( .A1(n7834), .A2(n7833), .ZN(n7832) );
  INV_X1 U7556 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U7557 ( .A1(n5866), .A2(n8571), .ZN(n5867) );
  NAND2_X1 U7558 ( .A1(n7832), .A2(n5867), .ZN(n7916) );
  XNOR2_X1 U7559 ( .A(n8877), .B(n5906), .ZN(n7914) );
  NAND2_X1 U7560 ( .A1(n7914), .A2(n8064), .ZN(n5868) );
  INV_X1 U7561 ( .A(n7914), .ZN(n5869) );
  NAND2_X1 U7562 ( .A1(n5869), .A2(n8933), .ZN(n5870) );
  XNOR2_X1 U7563 ( .A(n8468), .B(n5846), .ZN(n5872) );
  XNOR2_X1 U7564 ( .A(n5872), .B(n8866), .ZN(n8062) );
  INV_X1 U7565 ( .A(n8062), .ZN(n5871) );
  XNOR2_X1 U7566 ( .A(n9011), .B(n5906), .ZN(n5877) );
  XNOR2_X1 U7567 ( .A(n5877), .B(n8850), .ZN(n8075) );
  NAND2_X1 U7568 ( .A1(n5872), .A2(n8866), .ZN(n8073) );
  AND2_X1 U7569 ( .A1(n8075), .A2(n8073), .ZN(n5873) );
  NAND2_X1 U7570 ( .A1(n8074), .A2(n5873), .ZN(n8108) );
  XNOR2_X1 U7571 ( .A(n9004), .B(n5846), .ZN(n5874) );
  NAND2_X1 U7572 ( .A1(n5874), .A2(n8868), .ZN(n8249) );
  INV_X1 U7573 ( .A(n5874), .ZN(n5875) );
  INV_X1 U7574 ( .A(n8868), .ZN(n8837) );
  NAND2_X1 U7575 ( .A1(n5875), .A2(n8837), .ZN(n5876) );
  NAND2_X1 U7576 ( .A1(n8249), .A2(n5876), .ZN(n8105) );
  AND2_X1 U7577 ( .A1(n5877), .A2(n5118), .ZN(n8104) );
  NOR2_X1 U7578 ( .A1(n8105), .A2(n8104), .ZN(n5878) );
  NAND2_X1 U7579 ( .A1(n8108), .A2(n5878), .ZN(n8103) );
  NAND2_X1 U7580 ( .A1(n8103), .A2(n8249), .ZN(n5882) );
  XNOR2_X1 U7581 ( .A(n8998), .B(n5846), .ZN(n5879) );
  NAND2_X1 U7582 ( .A1(n5879), .A2(n8851), .ZN(n5883) );
  INV_X1 U7583 ( .A(n5879), .ZN(n5880) );
  INV_X1 U7584 ( .A(n8851), .ZN(n8570) );
  NAND2_X1 U7585 ( .A1(n5880), .A2(n8570), .ZN(n5881) );
  AND2_X1 U7586 ( .A1(n5883), .A2(n5881), .ZN(n8250) );
  NAND2_X1 U7587 ( .A1(n5882), .A2(n8250), .ZN(n8253) );
  NAND2_X1 U7588 ( .A1(n8253), .A2(n5883), .ZN(n8290) );
  XNOR2_X1 U7589 ( .A(n8914), .B(n5906), .ZN(n5884) );
  XNOR2_X1 U7590 ( .A(n5884), .B(n8257), .ZN(n8291) );
  INV_X1 U7591 ( .A(n5884), .ZN(n5885) );
  NAND2_X1 U7592 ( .A1(n5885), .A2(n8257), .ZN(n5886) );
  XNOR2_X1 U7593 ( .A(n8909), .B(n5846), .ZN(n5887) );
  AND2_X1 U7594 ( .A1(n5887), .A2(n8826), .ZN(n8210) );
  INV_X1 U7595 ( .A(n5887), .ZN(n5888) );
  INV_X1 U7596 ( .A(n8826), .ZN(n8569) );
  NAND2_X1 U7597 ( .A1(n5888), .A2(n8569), .ZN(n8211) );
  XNOR2_X1 U7598 ( .A(n8275), .B(n5846), .ZN(n5889) );
  XNOR2_X1 U7599 ( .A(n5889), .B(n8568), .ZN(n8270) );
  NAND2_X1 U7600 ( .A1(n5889), .A2(n8568), .ZN(n5890) );
  XNOR2_X1 U7601 ( .A(n8982), .B(n5906), .ZN(n5891) );
  XNOR2_X1 U7602 ( .A(n5891), .B(n8801), .ZN(n8233) );
  NAND2_X1 U7603 ( .A1(n8232), .A2(n8233), .ZN(n8279) );
  XNOR2_X1 U7604 ( .A(n8976), .B(n5846), .ZN(n5895) );
  XNOR2_X1 U7605 ( .A(n5895), .B(n8235), .ZN(n8280) );
  INV_X1 U7606 ( .A(n8280), .ZN(n5893) );
  INV_X1 U7607 ( .A(n5891), .ZN(n5892) );
  NAND2_X1 U7608 ( .A1(n5892), .A2(n8801), .ZN(n8278) );
  AND2_X1 U7609 ( .A1(n5893), .A2(n8278), .ZN(n5894) );
  NAND2_X1 U7610 ( .A1(n8279), .A2(n5894), .ZN(n8282) );
  INV_X1 U7611 ( .A(n5895), .ZN(n5896) );
  INV_X1 U7612 ( .A(n8235), .ZN(n8792) );
  NAND2_X1 U7613 ( .A1(n5896), .A2(n8792), .ZN(n5897) );
  NAND2_X1 U7614 ( .A1(n8282), .A2(n5897), .ZN(n5899) );
  XNOR2_X1 U7615 ( .A(n5898), .B(n5906), .ZN(n5901) );
  INV_X1 U7616 ( .A(n5899), .ZN(n5900) );
  XNOR2_X1 U7617 ( .A(n8964), .B(n5906), .ZN(n5902) );
  XNOR2_X1 U7618 ( .A(n5902), .B(n8735), .ZN(n8263) );
  INV_X1 U7619 ( .A(n8735), .ZN(n8766) );
  INV_X1 U7620 ( .A(n5902), .ZN(n5903) );
  XNOR2_X1 U7621 ( .A(n8246), .B(n5906), .ZN(n5904) );
  XNOR2_X1 U7622 ( .A(n5904), .B(n8744), .ZN(n8242) );
  INV_X1 U7623 ( .A(n5904), .ZN(n5905) );
  XNOR2_X1 U7624 ( .A(n8954), .B(n5906), .ZN(n5907) );
  XNOR2_X1 U7625 ( .A(n5907), .B(n8567), .ZN(n8303) );
  XNOR2_X1 U7626 ( .A(n8711), .B(n8225), .ZN(n5909) );
  NAND2_X1 U7627 ( .A1(n5909), .A2(n8566), .ZN(n8222) );
  OAI21_X1 U7628 ( .B1(n5909), .B2(n8566), .A(n8222), .ZN(n5910) );
  INV_X1 U7629 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U7630 ( .A1(n5918), .A2(n5913), .ZN(n5915) );
  OR2_X1 U7631 ( .A1(n5924), .A2(n5929), .ZN(n5914) );
  NAND2_X1 U7632 ( .A1(n5917), .A2(n5916), .ZN(n5946) );
  NAND2_X1 U7633 ( .A1(n5918), .A2(n8915), .ZN(n5921) );
  NAND2_X1 U7634 ( .A1(n5919), .A2(n8915), .ZN(n5920) );
  NAND2_X1 U7635 ( .A1(n5921), .A2(n10017), .ZN(n8310) );
  NAND2_X1 U7636 ( .A1(n8711), .A2(n8310), .ZN(n5945) );
  OR3_X1 U7637 ( .A1(n5924), .A2(n5936), .A3(n5922), .ZN(n8308) );
  INV_X1 U7638 ( .A(n8529), .ZN(n8565) );
  OR3_X1 U7639 ( .A1(n5924), .A2(n5923), .A3(n5936), .ZN(n8295) );
  INV_X1 U7640 ( .A(n8295), .ZN(n8304) );
  NAND2_X1 U7641 ( .A1(n8565), .A2(n8304), .ZN(n5942) );
  INV_X1 U7642 ( .A(n5925), .ZN(n5933) );
  AND3_X1 U7643 ( .A1(n5928), .A2(n5927), .A3(n5926), .ZN(n5931) );
  OR2_X1 U7644 ( .A1(n5937), .A2(n5929), .ZN(n5930) );
  OAI211_X1 U7645 ( .C1(n5933), .C2(n5932), .A(n5931), .B(n5930), .ZN(n5934)
         );
  NAND2_X1 U7646 ( .A1(n5934), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5940) );
  NOR2_X1 U7647 ( .A1(n5936), .A2(n5935), .ZN(n8557) );
  INV_X1 U7648 ( .A(n5937), .ZN(n5938) );
  NAND2_X1 U7649 ( .A1(n8557), .A2(n5938), .ZN(n5939) );
  NAND2_X1 U7650 ( .A1(n5940), .A2(n5939), .ZN(n8305) );
  AOI22_X1 U7651 ( .A1(n8707), .A2(n8305), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n5941) );
  OAI211_X1 U7652 ( .C1(n8736), .C2(n8308), .A(n5942), .B(n5941), .ZN(n5943)
         );
  INV_X1 U7653 ( .A(n5943), .ZN(n5944) );
  NAND2_X1 U7654 ( .A1(n8711), .A2(n8566), .ZN(n5950) );
  AND2_X1 U7655 ( .A1(n5947), .A2(n5950), .ZN(n5949) );
  AND2_X1 U7656 ( .A1(n5949), .A2(n5948), .ZN(n5953) );
  INV_X1 U7657 ( .A(n5950), .ZN(n5952) );
  NAND2_X1 U7658 ( .A1(n5955), .A2(n8325), .ZN(n5957) );
  NAND2_X1 U7659 ( .A1(n4926), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7660 ( .A(n6490), .B(n5958), .ZN(n5966) );
  NAND2_X1 U7661 ( .A1(n8197), .A2(n5960), .ZN(n8324) );
  INV_X1 U7662 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U7663 ( .A1(n4959), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7664 ( .A1(n8316), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5961) );
  OAI211_X1 U7665 ( .C1(n8198), .C2(n4960), .A(n5962), .B(n5961), .ZN(n5963)
         );
  INV_X1 U7666 ( .A(n5963), .ZN(n5964) );
  OAI22_X1 U7667 ( .A1(n8378), .A2(n8867), .B1(n8721), .B2(n8865), .ZN(n5965)
         );
  NAND2_X1 U7668 ( .A1(n8162), .A2(n5968), .ZN(n5974) );
  INV_X1 U7669 ( .A(n8524), .ZN(n5969) );
  XNOR2_X1 U7670 ( .A(n6486), .B(n8330), .ZN(n8158) );
  NAND2_X1 U7671 ( .A1(n5975), .A2(n4756), .ZN(P2_U3455) );
  NAND2_X1 U7672 ( .A1(n5994), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7673 ( .A1(n5993), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5981) );
  AND2_X2 U7674 ( .A1(n5977), .A2(n5976), .ZN(n6002) );
  NOR2_X1 U7675 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5978) );
  NOR2_X1 U7676 ( .A1(n6014), .A2(n5978), .ZN(n7492) );
  NAND2_X1 U7677 ( .A1(n6002), .A2(n7492), .ZN(n5980) );
  NAND2_X1 U7678 ( .A1(n6248), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7679 ( .A1(n4792), .A2(n9851), .ZN(n7359) );
  INV_X1 U7680 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6925) );
  OR2_X1 U7681 ( .A1(n5983), .A2(n6925), .ZN(n5986) );
  NAND2_X1 U7682 ( .A1(n6002), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5984) );
  NAND4_X2 U7683 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n6268)
         );
  INV_X1 U7684 ( .A(n9902), .ZN(n7135) );
  NAND2_X1 U7685 ( .A1(n5993), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7686 ( .A1(n6002), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7687 ( .A1(n5994), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5988) );
  AND2_X1 U7688 ( .A1(n7135), .A2(n6275), .ZN(n9891) );
  OR2_X1 U7689 ( .A1(n6268), .A2(n4278), .ZN(n5992) );
  NAND2_X1 U7690 ( .A1(n6002), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7691 ( .A1(n5993), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7692 ( .A1(n5994), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5995) );
  NOR2_X1 U7693 ( .A1(n9924), .A2(n9176), .ZN(n6224) );
  INV_X1 U7694 ( .A(n6224), .ZN(n5999) );
  NAND2_X1 U7695 ( .A1(n9924), .A2(n9176), .ZN(n6699) );
  NAND2_X1 U7696 ( .A1(n5999), .A2(n6699), .ZN(n9881) );
  INV_X1 U7697 ( .A(n9176), .ZN(n7282) );
  NAND2_X1 U7698 ( .A1(n7282), .A2(n9924), .ZN(n6000) );
  OR2_X1 U7699 ( .A1(n6188), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6004) );
  INV_X1 U7700 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6924) );
  OR2_X1 U7701 ( .A1(n6197), .A2(n6924), .ZN(n6003) );
  NAND2_X1 U7702 ( .A1(n6297), .A2(n9870), .ZN(n6539) );
  INV_X1 U7703 ( .A(n9870), .ZN(n9930) );
  INV_X1 U7704 ( .A(n6297), .ZN(n9175) );
  NAND2_X1 U7705 ( .A1(n9930), .A2(n9175), .ZN(n6700) );
  AND2_X1 U7706 ( .A1(n6539), .A2(n6700), .ZN(n7348) );
  NAND3_X1 U7707 ( .A1(n7359), .A2(n7347), .A3(n6007), .ZN(n6012) );
  INV_X1 U7708 ( .A(n9174), .ZN(n7283) );
  NAND2_X1 U7709 ( .A1(n7283), .A2(n7485), .ZN(n6010) );
  NAND2_X1 U7710 ( .A1(n6297), .A2(n9930), .ZN(n7349) );
  INV_X1 U7711 ( .A(n7349), .ZN(n6008) );
  AND2_X1 U7712 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  NAND2_X1 U7713 ( .A1(n6012), .A2(n6011), .ZN(n9860) );
  NAND2_X1 U7714 ( .A1(n6249), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7715 ( .A1(n6248), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6017) );
  INV_X1 U7716 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7717 ( .A1(n6197), .A2(n6013), .ZN(n6016) );
  NAND2_X1 U7718 ( .A1(n6014), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6026) );
  OAI21_X1 U7719 ( .B1(n6014), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6026), .ZN(
        n9857) );
  OR2_X1 U7720 ( .A1(n6188), .A2(n9857), .ZN(n6015) );
  NAND2_X1 U7721 ( .A1(n7361), .A2(n9859), .ZN(n6542) );
  INV_X1 U7722 ( .A(n7361), .ZN(n9173) );
  AND2_X1 U7723 ( .A1(n9945), .A2(n9173), .ZN(n6227) );
  INV_X1 U7724 ( .A(n6227), .ZN(n6704) );
  NAND2_X1 U7725 ( .A1(n6542), .A2(n6704), .ZN(n9861) );
  AND2_X1 U7726 ( .A1(n7361), .A2(n9945), .ZN(n6019) );
  NAND2_X1 U7727 ( .A1(n6249), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7728 ( .A1(n5993), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6022) );
  XNOR2_X1 U7729 ( .A(n6026), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U7730 ( .A1(n6002), .A2(n7508), .ZN(n6021) );
  NAND2_X1 U7731 ( .A1(n6248), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6020) );
  NAND4_X1 U7732 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n9172)
         );
  OR2_X1 U7733 ( .A1(n9172), .A2(n9953), .ZN(n6546) );
  NAND2_X1 U7734 ( .A1(n9953), .A2(n9172), .ZN(n6545) );
  NAND2_X1 U7735 ( .A1(n6546), .A2(n6545), .ZN(n6658) );
  INV_X1 U7736 ( .A(n6026), .ZN(n6024) );
  AOI21_X1 U7737 ( .B1(n6024), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7738 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6025) );
  NOR2_X1 U7739 ( .A1(n6026), .A2(n6025), .ZN(n6033) );
  OR2_X1 U7740 ( .A1(n6027), .A2(n6033), .ZN(n9843) );
  OR2_X1 U7741 ( .A1(n6188), .A2(n9843), .ZN(n6031) );
  NAND2_X1 U7742 ( .A1(n5993), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7743 ( .A1(n6249), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7744 ( .A1(n6248), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6028) );
  NAND4_X1 U7745 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n9171)
         );
  NAND2_X1 U7746 ( .A1(n9959), .A2(n9171), .ZN(n6550) );
  INV_X1 U7747 ( .A(n9171), .ZN(n6032) );
  NAND2_X1 U7748 ( .A1(n6032), .A2(n9845), .ZN(n7555) );
  AOI22_X1 U7749 ( .A1(n9837), .A2(n9838), .B1(n6032), .B2(n9959), .ZN(n7554)
         );
  NAND2_X1 U7750 ( .A1(n6249), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6038) );
  INV_X1 U7751 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7102) );
  OR2_X1 U7752 ( .A1(n6197), .A2(n7102), .ZN(n6037) );
  OR2_X1 U7753 ( .A1(n6125), .A2(n4479), .ZN(n6036) );
  NAND2_X1 U7754 ( .A1(n6033), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6050) );
  OR2_X1 U7755 ( .A1(n6033), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7756 ( .A1(n6050), .A2(n6034), .ZN(n7804) );
  OR2_X1 U7757 ( .A1(n6188), .A2(n7804), .ZN(n6035) );
  NAND2_X1 U7758 ( .A1(n9967), .A2(n7588), .ZN(n6556) );
  NAND2_X1 U7759 ( .A1(n7588), .A2(n6039), .ZN(n6040) );
  NAND2_X1 U7760 ( .A1(n6249), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6046) );
  INV_X1 U7761 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6041) );
  OR2_X1 U7762 ( .A1(n6197), .A2(n6041), .ZN(n6045) );
  INV_X1 U7763 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7764 ( .A1(n6125), .A2(n6042), .ZN(n6044) );
  INV_X1 U7765 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6048) );
  XNOR2_X1 U7766 ( .A(n6050), .B(n6048), .ZN(n9823) );
  OR2_X1 U7767 ( .A1(n6188), .A2(n9823), .ZN(n6043) );
  NAND2_X1 U7768 ( .A1(n9976), .A2(n7680), .ZN(n6563) );
  NAND2_X1 U7769 ( .A1(n6569), .A2(n6563), .ZN(n9820) );
  NAND2_X1 U7770 ( .A1(n6249), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6055) );
  INV_X1 U7771 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7294) );
  OR2_X1 U7772 ( .A1(n6197), .A2(n7294), .ZN(n6054) );
  INV_X1 U7773 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7684) );
  OR2_X1 U7774 ( .A1(n6125), .A2(n7684), .ZN(n6053) );
  INV_X1 U7775 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6047) );
  OAI21_X1 U7776 ( .B1(n6050), .B2(n6048), .A(n6047), .ZN(n6051) );
  NAND2_X1 U7777 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n6049) );
  NAND2_X1 U7778 ( .A1(n6051), .A2(n6056), .ZN(n9759) );
  OR2_X1 U7779 ( .A1(n6188), .A2(n9759), .ZN(n6052) );
  OR2_X1 U7780 ( .A1(n7687), .A2(n7960), .ZN(n6708) );
  NAND2_X1 U7781 ( .A1(n7687), .A2(n7960), .ZN(n9803) );
  INV_X1 U7782 ( .A(n7960), .ZN(n9168) );
  NAND2_X1 U7783 ( .A1(n6248), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7784 ( .A1(n6249), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6060) );
  INV_X1 U7785 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7438) );
  NOR2_X1 U7786 ( .A1(n6056), .A2(n7438), .ZN(n6062) );
  INV_X1 U7787 ( .A(n6062), .ZN(n6064) );
  NAND2_X1 U7788 ( .A1(n6056), .A2(n7438), .ZN(n6057) );
  NAND2_X1 U7789 ( .A1(n6064), .A2(n6057), .ZN(n9809) );
  OR2_X1 U7790 ( .A1(n6188), .A2(n9809), .ZN(n6059) );
  INV_X1 U7791 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7435) );
  OR2_X1 U7792 ( .A1(n6197), .A2(n7435), .ZN(n6058) );
  INV_X1 U7793 ( .A(n7726), .ZN(n9167) );
  INV_X1 U7794 ( .A(n9811), .ZN(n9992) );
  NAND2_X1 U7795 ( .A1(n6249), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6069) );
  INV_X1 U7796 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7596) );
  OR2_X1 U7797 ( .A1(n6197), .A2(n7596), .ZN(n6068) );
  INV_X1 U7798 ( .A(n6073), .ZN(n6074) );
  INV_X1 U7799 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7800 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  NAND2_X1 U7801 ( .A1(n6074), .A2(n6065), .ZN(n8032) );
  OR2_X1 U7802 ( .A1(n6188), .A2(n8032), .ZN(n6067) );
  INV_X1 U7803 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7732) );
  OR2_X1 U7804 ( .A1(n6125), .A2(n7732), .ZN(n6066) );
  OR2_X1 U7805 ( .A1(n7768), .A2(n7961), .ZN(n6575) );
  NAND2_X1 U7806 ( .A1(n7768), .A2(n7961), .ZN(n6715) );
  INV_X1 U7807 ( .A(n7961), .ZN(n9166) );
  NAND2_X1 U7808 ( .A1(n5994), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6079) );
  INV_X1 U7809 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6071) );
  OR2_X1 U7810 ( .A1(n6197), .A2(n6071), .ZN(n6078) );
  INV_X1 U7811 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6072) );
  OR2_X1 U7812 ( .A1(n6125), .A2(n6072), .ZN(n6077) );
  NAND2_X1 U7813 ( .A1(n6073), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6082) );
  INV_X1 U7814 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7628) );
  NAND2_X1 U7815 ( .A1(n6074), .A2(n7628), .ZN(n6075) );
  NAND2_X1 U7816 ( .A1(n6082), .A2(n6075), .ZN(n8087) );
  OR2_X1 U7817 ( .A1(n6188), .A2(n8087), .ZN(n6076) );
  OR2_X1 U7818 ( .A1(n8089), .A2(n7897), .ZN(n6718) );
  NAND2_X1 U7819 ( .A1(n8089), .A2(n7897), .ZN(n6716) );
  NAND2_X1 U7820 ( .A1(n6718), .A2(n6716), .ZN(n7786) );
  NAND2_X1 U7821 ( .A1(n7787), .A2(n7786), .ZN(n7785) );
  NAND2_X1 U7822 ( .A1(n7785), .A2(n6080), .ZN(n7901) );
  NAND2_X1 U7823 ( .A1(n5994), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6087) );
  INV_X1 U7824 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7711) );
  OR2_X1 U7825 ( .A1(n6197), .A2(n7711), .ZN(n6086) );
  INV_X1 U7826 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7827 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  NAND2_X1 U7828 ( .A1(n6090), .A2(n6083), .ZN(n9031) );
  OR2_X1 U7829 ( .A1(n6188), .A2(n9031), .ZN(n6085) );
  INV_X1 U7830 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7904) );
  OR2_X1 U7831 ( .A1(n6125), .A2(n7904), .ZN(n6084) );
  XNOR2_X1 U7832 ( .A(n9033), .B(n9164), .ZN(n6663) );
  NAND2_X1 U7833 ( .A1(n7901), .A2(n7900), .ZN(n7899) );
  NAND2_X1 U7834 ( .A1(n7899), .A2(n6088), .ZN(n8002) );
  NAND2_X1 U7835 ( .A1(n5994), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6095) );
  INV_X1 U7836 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6089) );
  OR2_X1 U7837 ( .A1(n6197), .A2(n6089), .ZN(n6094) );
  INV_X1 U7838 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U7839 ( .A1(n6090), .A2(n7985), .ZN(n6091) );
  NAND2_X1 U7840 ( .A1(n6098), .A2(n6091), .ZN(n9146) );
  OR2_X1 U7841 ( .A1(n6188), .A2(n9146), .ZN(n6093) );
  INV_X1 U7842 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8005) );
  OR2_X1 U7843 ( .A1(n6125), .A2(n8005), .ZN(n6092) );
  NAND2_X1 U7844 ( .A1(n9142), .A2(n8121), .ZN(n6589) );
  NAND2_X1 U7845 ( .A1(n6722), .A2(n6589), .ZN(n8001) );
  NAND2_X1 U7846 ( .A1(n5994), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7847 ( .A1(n6248), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6102) );
  INV_X1 U7848 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9179) );
  OR2_X1 U7849 ( .A1(n6197), .A2(n9179), .ZN(n6101) );
  INV_X1 U7850 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9065) );
  NOR2_X1 U7851 ( .A1(n6098), .A2(n9065), .ZN(n6105) );
  INV_X1 U7852 ( .A(n6105), .ZN(n6107) );
  NAND2_X1 U7853 ( .A1(n6098), .A2(n9065), .ZN(n6099) );
  NAND2_X1 U7854 ( .A1(n6107), .A2(n6099), .ZN(n9066) );
  OR2_X1 U7855 ( .A1(n6188), .A2(n9066), .ZN(n6100) );
  OR2_X1 U7856 ( .A1(n6104), .A2(n8146), .ZN(n6605) );
  NAND2_X1 U7857 ( .A1(n6104), .A2(n8146), .ZN(n6724) );
  NAND2_X1 U7858 ( .A1(n6605), .A2(n6724), .ZN(n8117) );
  NAND2_X1 U7859 ( .A1(n6248), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6112) );
  INV_X1 U7860 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9205) );
  OR2_X1 U7861 ( .A1(n6197), .A2(n9205), .ZN(n6111) );
  INV_X1 U7862 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9511) );
  OR2_X1 U7863 ( .A1(n6180), .A2(n9511), .ZN(n6110) );
  NAND2_X1 U7864 ( .A1(n6105), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6115) );
  INV_X1 U7865 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7866 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  NAND2_X1 U7867 ( .A1(n6115), .A2(n6108), .ZN(n9077) );
  OR2_X1 U7868 ( .A1(n6188), .A2(n9077), .ZN(n6109) );
  INV_X1 U7869 ( .A(n9118), .ZN(n9163) );
  NAND2_X1 U7870 ( .A1(n9624), .A2(n9118), .ZN(n6604) );
  NAND2_X1 U7871 ( .A1(n5994), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7872 ( .A1(n5993), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7873 ( .A1(n6248), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6118) );
  INV_X1 U7874 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7875 ( .A1(n6115), .A2(n6114), .ZN(n6116) );
  NAND2_X1 U7876 ( .A1(n6123), .A2(n6116), .ZN(n9428) );
  OR2_X1 U7877 ( .A1(n6188), .A2(n9428), .ZN(n6117) );
  OR2_X1 U7878 ( .A1(n9426), .A2(n8168), .ZN(n6606) );
  NAND2_X1 U7879 ( .A1(n9426), .A2(n8168), .ZN(n9404) );
  NAND2_X1 U7880 ( .A1(n6606), .A2(n9404), .ZN(n9421) );
  NAND2_X1 U7881 ( .A1(n9422), .A2(n9421), .ZN(n9420) );
  INV_X1 U7882 ( .A(n8168), .ZN(n9162) );
  NAND2_X1 U7883 ( .A1(n5994), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7884 ( .A1(n5993), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6128) );
  INV_X1 U7885 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6122) );
  NOR2_X1 U7886 ( .A1(n6123), .A2(n6122), .ZN(n6134) );
  INV_X1 U7887 ( .A(n6134), .ZN(n6136) );
  NAND2_X1 U7888 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  NAND2_X1 U7889 ( .A1(n6136), .A2(n6124), .ZN(n9400) );
  OR2_X1 U7890 ( .A1(n6188), .A2(n9400), .ZN(n6127) );
  INV_X1 U7891 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9233) );
  OR2_X1 U7892 ( .A1(n6125), .A2(n9233), .ZN(n6126) );
  INV_X1 U7893 ( .A(n9119), .ZN(n9161) );
  NAND2_X1 U7894 ( .A1(n9483), .A2(n9161), .ZN(n6131) );
  INV_X1 U7895 ( .A(n9483), .ZN(n9403) );
  NAND2_X1 U7896 ( .A1(n6249), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7897 ( .A1(n5993), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6132) );
  AND2_X1 U7898 ( .A1(n6133), .A2(n6132), .ZN(n6140) );
  INV_X1 U7899 ( .A(n6141), .ZN(n6143) );
  INV_X1 U7900 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7901 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  AND2_X1 U7902 ( .A1(n6143), .A2(n6137), .ZN(n9392) );
  NAND2_X1 U7903 ( .A1(n9392), .A2(n6002), .ZN(n6139) );
  NAND2_X1 U7904 ( .A1(n6248), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6138) );
  INV_X1 U7905 ( .A(n8169), .ZN(n9160) );
  NAND2_X1 U7906 ( .A1(n6141), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6151) );
  INV_X1 U7907 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7908 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  NAND2_X1 U7909 ( .A1(n6151), .A2(n6144), .ZN(n9376) );
  OR2_X1 U7910 ( .A1(n9376), .A2(n6188), .ZN(n6147) );
  AOI22_X1 U7911 ( .A1(n5993), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5994), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7912 ( .A1(n6248), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7913 ( .A1(n9375), .A2(n9106), .ZN(n6615) );
  INV_X1 U7914 ( .A(n9367), .ZN(n6149) );
  INV_X1 U7915 ( .A(n9106), .ZN(n9159) );
  INV_X1 U7916 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7917 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  AND2_X1 U7918 ( .A1(n6157), .A2(n6152), .ZN(n9357) );
  NAND2_X1 U7919 ( .A1(n9357), .A2(n6002), .ZN(n6155) );
  AOI22_X1 U7920 ( .A1(n5993), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n6249), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7921 ( .A1(n6248), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6153) );
  INV_X1 U7922 ( .A(n9053), .ZN(n9158) );
  NAND2_X1 U7923 ( .A1(n9356), .A2(n9158), .ZN(n6156) );
  INV_X1 U7924 ( .A(n9356), .ZN(n9649) );
  INV_X1 U7925 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U7926 ( .A1(n6157), .A2(n9591), .ZN(n6158) );
  NAND2_X1 U7927 ( .A1(n6176), .A2(n6158), .ZN(n9047) );
  INV_X1 U7928 ( .A(n9047), .ZN(n9342) );
  NAND2_X1 U7929 ( .A1(n9342), .A2(n6002), .ZN(n6164) );
  INV_X1 U7930 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7931 ( .A1(n6249), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7932 ( .A1(n6248), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U7933 ( .C1(n6197), .C2(n6161), .A(n6160), .B(n6159), .ZN(n6162)
         );
  INV_X1 U7934 ( .A(n6162), .ZN(n6163) );
  NAND2_X1 U7935 ( .A1(n4619), .A2(n9107), .ZN(n6166) );
  INV_X1 U7936 ( .A(n9107), .ZN(n9157) );
  XNOR2_X1 U7937 ( .A(n6176), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U7938 ( .A1(n9327), .A2(n6002), .ZN(n6171) );
  INV_X1 U7939 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U7940 ( .A1(n6248), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7941 ( .A1(n5993), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6167) );
  OAI211_X1 U7942 ( .C1(n6180), .C2(n9642), .A(n6168), .B(n6167), .ZN(n6169)
         );
  INV_X1 U7943 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7944 ( .A1(n6171), .A2(n6170), .ZN(n9156) );
  NAND2_X1 U7945 ( .A1(n9326), .A2(n9156), .ZN(n6173) );
  INV_X1 U7946 ( .A(n9156), .ZN(n6625) );
  NAND2_X1 U7947 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n6174) );
  NOR2_X1 U7948 ( .A1(n6176), .A2(n6174), .ZN(n6185) );
  INV_X1 U7949 ( .A(n6185), .ZN(n6186) );
  INV_X1 U7950 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9089) );
  INV_X1 U7951 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6175) );
  OAI21_X1 U7952 ( .B1(n6176), .B2(n9089), .A(n6175), .ZN(n6177) );
  AND2_X1 U7953 ( .A1(n6186), .A2(n6177), .ZN(n9312) );
  NAND2_X1 U7954 ( .A1(n9312), .A2(n6002), .ZN(n6183) );
  INV_X1 U7955 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U7956 ( .A1(n5993), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7957 ( .A1(n6248), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7958 ( .C1(n6180), .C2(n9536), .A(n6179), .B(n6178), .ZN(n6181)
         );
  INV_X1 U7959 ( .A(n6181), .ZN(n6182) );
  NAND2_X1 U7960 ( .A1(n6183), .A2(n6182), .ZN(n9155) );
  INV_X1 U7961 ( .A(n9155), .ZN(n6243) );
  NAND2_X1 U7962 ( .A1(n9315), .A2(n6243), .ZN(n6184) );
  AND2_X1 U7963 ( .A1(n6185), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6203) );
  INV_X1 U7964 ( .A(n6203), .ZN(n6201) );
  INV_X1 U7965 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U7966 ( .A1(n6186), .A2(n9134), .ZN(n6187) );
  NAND2_X1 U7967 ( .A1(n6201), .A2(n6187), .ZN(n9294) );
  OR2_X1 U7968 ( .A1(n9294), .A2(n6188), .ZN(n6193) );
  INV_X1 U7969 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9450) );
  NAND2_X1 U7970 ( .A1(n5994), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7971 ( .A1(n6248), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6189) );
  OAI211_X1 U7972 ( .C1(n6197), .C2(n9450), .A(n6190), .B(n6189), .ZN(n6191)
         );
  INV_X1 U7973 ( .A(n6191), .ZN(n6192) );
  XNOR2_X1 U7974 ( .A(n6201), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9270) );
  INV_X1 U7975 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7976 ( .A1(n5994), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7977 ( .A1(n6248), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6194) );
  OAI211_X1 U7978 ( .C1(n6197), .C2(n6196), .A(n6195), .B(n6194), .ZN(n6198)
         );
  AOI21_X1 U7979 ( .B1(n9270), .B2(n6002), .A(n6198), .ZN(n9130) );
  NAND2_X1 U7980 ( .A1(n6199), .A2(n9130), .ZN(n6635) );
  NAND2_X1 U7981 ( .A1(n6637), .A2(n6635), .ZN(n6668) );
  INV_X1 U7982 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6810) );
  INV_X1 U7983 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6200) );
  OAI21_X1 U7984 ( .B1(n6201), .B2(n6810), .A(n6200), .ZN(n6205) );
  AND2_X1 U7985 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6202) );
  AND2_X1 U7986 ( .A1(n6203), .A2(n6202), .ZN(n8176) );
  INV_X1 U7987 ( .A(n8176), .ZN(n6204) );
  AND2_X1 U7988 ( .A1(n6205), .A2(n6204), .ZN(n9262) );
  INV_X1 U7989 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7990 ( .A1(n5994), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7991 ( .A1(n6248), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6206) );
  OAI211_X1 U7992 ( .C1(n6197), .C2(n6208), .A(n6207), .B(n6206), .ZN(n6209)
         );
  AOI21_X1 U7993 ( .B1(n9262), .B2(n6002), .A(n6209), .ZN(n7251) );
  INV_X1 U7994 ( .A(n7251), .ZN(n6210) );
  INV_X1 U7995 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7996 ( .A1(n5994), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7997 ( .A1(n6248), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6212) );
  OAI211_X1 U7998 ( .C1(n6197), .C2(n6214), .A(n6213), .B(n6212), .ZN(n6215)
         );
  AOI21_X1 U7999 ( .B1(n8176), .B2(n6002), .A(n6215), .ZN(n6835) );
  NAND2_X1 U8000 ( .A1(n6216), .A2(n6835), .ZN(n6737) );
  INV_X1 U8001 ( .A(n6911), .ZN(n6470) );
  OR2_X1 U8002 ( .A1(n6768), .A2(n6470), .ZN(n6218) );
  INV_X1 U8003 ( .A(n7136), .ZN(n6217) );
  NAND2_X1 U8004 ( .A1(n6218), .A2(n6217), .ZN(n7379) );
  NAND2_X1 U8005 ( .A1(n5804), .A2(n6220), .ZN(n6260) );
  AND2_X1 U8006 ( .A1(n6260), .A2(n6768), .ZN(n6221) );
  OR2_X1 U8007 ( .A1(n7379), .A2(n6221), .ZN(n7352) );
  OR2_X1 U8008 ( .A1(n6649), .A2(n6742), .ZN(n9969) );
  AND2_X1 U8009 ( .A1(n7352), .A2(n9969), .ZN(n9941) );
  OR2_X1 U8010 ( .A1(n9391), .A2(n8169), .ZN(n9366) );
  NAND2_X1 U8011 ( .A1(n9893), .A2(n9892), .ZN(n6223) );
  INV_X1 U8012 ( .A(n6268), .ZN(n7092) );
  NAND2_X1 U8013 ( .A1(n7092), .A2(n4278), .ZN(n6222) );
  NAND2_X1 U8014 ( .A1(n6223), .A2(n6222), .ZN(n9882) );
  NAND2_X1 U8015 ( .A1(n6538), .A2(n6539), .ZN(n6225) );
  NAND2_X1 U8016 ( .A1(n6225), .A2(n6700), .ZN(n7360) );
  INV_X1 U8017 ( .A(n7360), .ZN(n6226) );
  AND2_X1 U8018 ( .A1(n9851), .A2(n6542), .ZN(n6228) );
  INV_X1 U8019 ( .A(n7470), .ZN(n6230) );
  NAND2_X1 U8020 ( .A1(n6569), .A2(n9818), .ZN(n6557) );
  NAND2_X1 U8021 ( .A1(n6556), .A2(n7555), .ZN(n6551) );
  INV_X1 U8022 ( .A(n6563), .ZN(n6229) );
  NAND3_X1 U8023 ( .A1(n6230), .A2(n6661), .A3(n6546), .ZN(n6710) );
  INV_X1 U8024 ( .A(n6545), .ZN(n6232) );
  NAND2_X1 U8025 ( .A1(n9811), .A2(n7726), .ZN(n6573) );
  NAND2_X1 U8026 ( .A1(n6573), .A2(n9803), .ZN(n6564) );
  INV_X1 U8027 ( .A(n6564), .ZN(n6711) );
  OR2_X1 U8028 ( .A1(n9811), .A2(n7726), .ZN(n7722) );
  AND2_X1 U8029 ( .A1(n6575), .A2(n7722), .ZN(n6713) );
  NAND2_X1 U8030 ( .A1(n7723), .A2(n6713), .ZN(n7779) );
  NAND2_X1 U8031 ( .A1(n7779), .A2(n6715), .ZN(n6233) );
  INV_X1 U8032 ( .A(n7786), .ZN(n7778) );
  NAND2_X1 U8033 ( .A1(n6233), .A2(n7778), .ZN(n7776) );
  OR2_X1 U8034 ( .A1(n9033), .A2(n7997), .ZN(n7991) );
  INV_X1 U8035 ( .A(n7991), .ZN(n6234) );
  NOR2_X1 U8036 ( .A1(n8001), .A2(n6234), .ZN(n6235) );
  NAND2_X1 U8037 ( .A1(n7994), .A2(n6589), .ZN(n8120) );
  INV_X1 U8038 ( .A(n6724), .ZN(n6236) );
  OR2_X2 U8039 ( .A1(n8120), .A2(n6236), .ZN(n6237) );
  NAND2_X1 U8040 ( .A1(n6237), .A2(n6605), .ZN(n8144) );
  OR2_X1 U8041 ( .A1(n9483), .A2(n9119), .ZN(n6608) );
  NAND2_X1 U8042 ( .A1(n9483), .A2(n9119), .ZN(n6729) );
  NAND2_X1 U8043 ( .A1(n6608), .A2(n6729), .ZN(n9405) );
  INV_X1 U8044 ( .A(n9404), .ZN(n6239) );
  NOR2_X1 U8045 ( .A1(n9405), .A2(n6239), .ZN(n6240) );
  NAND2_X1 U8046 ( .A1(n9415), .A2(n6240), .ZN(n6241) );
  NAND2_X1 U8047 ( .A1(n6241), .A2(n6608), .ZN(n9364) );
  NOR2_X1 U8048 ( .A1(n6697), .A2(n9364), .ZN(n6750) );
  NAND2_X1 U8049 ( .A1(n9391), .A2(n8169), .ZN(n6654) );
  NAND2_X1 U8050 ( .A1(n6615), .A2(n6654), .ZN(n6536) );
  NAND2_X1 U8051 ( .A1(n6536), .A2(n6616), .ZN(n6686) );
  INV_X1 U8052 ( .A(n6686), .ZN(n6242) );
  XNOR2_X1 U8053 ( .A(n9356), .B(n9158), .ZN(n9349) );
  OR2_X1 U8054 ( .A1(n9356), .A2(n9053), .ZN(n6622) );
  XNOR2_X1 U8055 ( .A(n9463), .B(n9157), .ZN(n9339) );
  INV_X1 U8056 ( .A(n9339), .ZN(n9334) );
  NAND2_X1 U8057 ( .A1(n9463), .A2(n9107), .ZN(n6679) );
  XNOR2_X1 U8058 ( .A(n9326), .B(n9156), .ZN(n9321) );
  NAND2_X1 U8059 ( .A1(n9322), .A2(n9321), .ZN(n9320) );
  OR2_X1 U8060 ( .A1(n9326), .A2(n6625), .ZN(n6681) );
  NAND2_X1 U8061 ( .A1(n9320), .A2(n6681), .ZN(n9304) );
  NAND2_X1 U8062 ( .A1(n9454), .A2(n6243), .ZN(n6631) );
  NAND2_X1 U8063 ( .A1(n9283), .A2(n6631), .ZN(n9302) );
  INV_X1 U8064 ( .A(n9302), .ZN(n9305) );
  NAND2_X2 U8065 ( .A1(n9304), .A2(n9305), .ZN(n9303) );
  OR2_X1 U8066 ( .A1(n9293), .A2(n6787), .ZN(n6636) );
  NAND2_X1 U8067 ( .A1(n9293), .A2(n6787), .ZN(n6634) );
  NAND2_X1 U8068 ( .A1(n6636), .A2(n6634), .ZN(n9284) );
  NOR2_X1 U8069 ( .A1(n9284), .A2(n6632), .ZN(n6244) );
  INV_X1 U8070 ( .A(n6668), .ZN(n9275) );
  INV_X1 U8071 ( .A(n9257), .ZN(n9253) );
  NAND2_X1 U8072 ( .A1(n9252), .A2(n9253), .ZN(n9251) );
  NAND2_X1 U8073 ( .A1(n9251), .A2(n6642), .ZN(n6246) );
  XNOR2_X1 U8074 ( .A(n6246), .B(n6245), .ZN(n6255) );
  NAND2_X1 U8075 ( .A1(n6219), .A2(n6220), .ZN(n6247) );
  NAND2_X1 U8076 ( .A1(n6655), .A2(n6742), .ZN(n6771) );
  NAND2_X1 U8077 ( .A1(n6247), .A2(n6771), .ZN(n9868) );
  AND2_X1 U8078 ( .A1(n7182), .A2(n6911), .ZN(n9131) );
  INV_X1 U8079 ( .A(n9131), .ZN(n9117) );
  INV_X1 U8080 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U8081 ( .A1(n6248), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U8082 ( .A1(n6249), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6250) );
  OAI211_X1 U8083 ( .C1(n6197), .C2(n6252), .A(n6251), .B(n6250), .ZN(n9151)
         );
  INV_X1 U8084 ( .A(n9151), .ZN(n6671) );
  OAI22_X1 U8085 ( .A1(n7251), .A2(n9117), .B1(n6671), .B2(n6253), .ZN(n6254)
         );
  INV_X1 U8086 ( .A(n6256), .ZN(n9260) );
  OAI211_X1 U8087 ( .C1(n8178), .C2(n9260), .A(n9901), .B(n6504), .ZN(n8175)
         );
  NOR2_X1 U8088 ( .A1(n8178), .A2(n9667), .ZN(n6257) );
  AND2_X1 U8089 ( .A1(n6655), .A2(n6745), .ZN(n6263) );
  NAND2_X1 U8090 ( .A1(n6219), .A2(n6263), .ZN(n7353) );
  NAND2_X4 U8091 ( .A1(n6259), .A2(n4292), .ZN(n6827) );
  NAND2_X1 U8092 ( .A1(n6260), .A2(n7643), .ZN(n6261) );
  NAND2_X1 U8093 ( .A1(n6261), .A2(n6771), .ZN(n6262) );
  NAND2_X4 U8094 ( .A1(n6262), .A2(n6847), .ZN(n6794) );
  AOI22_X1 U8095 ( .A1(n9454), .A2(n4277), .B1(n6825), .B2(n9155), .ZN(n6264)
         );
  XNOR2_X1 U8096 ( .A(n6264), .B(n6794), .ZN(n6791) );
  INV_X2 U8097 ( .A(n6827), .ZN(n6451) );
  NAND2_X1 U8098 ( .A1(n9155), .A2(n6451), .ZN(n6265) );
  NAND2_X1 U8099 ( .A1(n6266), .A2(n6265), .ZN(n6789) );
  XNOR2_X1 U8100 ( .A(n6791), .B(n6789), .ZN(n6462) );
  INV_X1 U8101 ( .A(n6288), .ZN(n6276) );
  INV_X2 U8102 ( .A(n6276), .ZN(n6825) );
  NAND2_X1 U8103 ( .A1(n4277), .A2(n4278), .ZN(n6270) );
  NAND2_X1 U8104 ( .A1(n6268), .A2(n6288), .ZN(n6269) );
  NAND2_X1 U8105 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  XNOR2_X1 U8106 ( .A(n6282), .B(n6281), .ZN(n7142) );
  NAND2_X1 U8107 ( .A1(n6286), .A2(n7135), .ZN(n6273) );
  NAND2_X1 U8108 ( .A1(n6275), .A2(n6288), .ZN(n6272) );
  NAND2_X1 U8109 ( .A1(n6273), .A2(n6272), .ZN(n6279) );
  INV_X1 U8110 ( .A(n6279), .ZN(n6274) );
  INV_X1 U8111 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U8112 ( .A1(n6275), .A2(n6451), .ZN(n6278) );
  OR2_X1 U8113 ( .A1(n9902), .A2(n6276), .ZN(n6277) );
  OAI211_X1 U8114 ( .C1(n5599), .C2(n6847), .A(n6278), .B(n6277), .ZN(n7090)
         );
  NAND2_X1 U8115 ( .A1(n7091), .A2(n7090), .ZN(n7089) );
  OR2_X1 U8116 ( .A1(n6279), .A2(n6794), .ZN(n6280) );
  AND2_X1 U8117 ( .A1(n7089), .A2(n6280), .ZN(n7143) );
  NAND2_X1 U8118 ( .A1(n7142), .A2(n7143), .ZN(n6285) );
  INV_X1 U8119 ( .A(n6281), .ZN(n6283) );
  NAND2_X1 U8120 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  NAND2_X1 U8121 ( .A1(n6285), .A2(n6284), .ZN(n7211) );
  NAND2_X1 U8122 ( .A1(n9176), .A2(n6288), .ZN(n6287) );
  INV_X1 U8123 ( .A(n6288), .ZN(n6796) );
  OR2_X1 U8124 ( .A1(n9924), .A2(n6796), .ZN(n6290) );
  NAND2_X1 U8125 ( .A1(n9176), .A2(n6451), .ZN(n6289) );
  NAND2_X1 U8126 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  XNOR2_X1 U8127 ( .A(n6293), .B(n6291), .ZN(n7212) );
  NAND2_X1 U8128 ( .A1(n7211), .A2(n7212), .ZN(n6295) );
  INV_X1 U8129 ( .A(n6291), .ZN(n6292) );
  NAND2_X1 U8130 ( .A1(n6293), .A2(n6292), .ZN(n6294) );
  NAND2_X1 U8131 ( .A1(n6295), .A2(n6294), .ZN(n7280) );
  NAND2_X1 U8132 ( .A1(n9870), .A2(n6286), .ZN(n6296) );
  XNOR2_X1 U8133 ( .A(n6298), .B(n6823), .ZN(n6302) );
  NAND2_X1 U8134 ( .A1(n9870), .A2(n6288), .ZN(n6299) );
  OAI21_X1 U8135 ( .B1(n6297), .B2(n6827), .A(n6299), .ZN(n6300) );
  XNOR2_X1 U8136 ( .A(n6302), .B(n6300), .ZN(n7281) );
  NAND2_X1 U8137 ( .A1(n7280), .A2(n7281), .ZN(n6304) );
  INV_X1 U8138 ( .A(n6300), .ZN(n6301) );
  NAND2_X1 U8139 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  NAND2_X1 U8140 ( .A1(n9174), .A2(n6288), .ZN(n6305) );
  OAI21_X1 U8141 ( .B1(n7485), .B2(n6793), .A(n6305), .ZN(n6306) );
  XNOR2_X1 U8142 ( .A(n6306), .B(n6794), .ZN(n6310) );
  OR2_X1 U8143 ( .A1(n7485), .A2(n6796), .ZN(n6308) );
  NAND2_X1 U8144 ( .A1(n9174), .A2(n6451), .ZN(n6307) );
  NAND2_X1 U8145 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  NAND2_X1 U8146 ( .A1(n6310), .A2(n6309), .ZN(n6317) );
  OR2_X1 U8147 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  NAND2_X1 U8148 ( .A1(n6317), .A2(n6311), .ZN(n7489) );
  NAND2_X1 U8149 ( .A1(n9859), .A2(n6286), .ZN(n6313) );
  OAI21_X1 U8150 ( .B1(n7361), .B2(n6796), .A(n6313), .ZN(n6314) );
  XNOR2_X1 U8151 ( .A(n6314), .B(n6823), .ZN(n6318) );
  AND2_X1 U8152 ( .A1(n6317), .A2(n6318), .ZN(n6315) );
  NAND2_X1 U8153 ( .A1(n9859), .A2(n6288), .ZN(n6316) );
  OAI21_X1 U8154 ( .B1(n7361), .B2(n6827), .A(n6316), .ZN(n7463) );
  INV_X1 U8155 ( .A(n6318), .ZN(n6319) );
  NAND2_X1 U8156 ( .A1(n9172), .A2(n6288), .ZN(n6321) );
  OAI21_X1 U8157 ( .B1(n9953), .B2(n6793), .A(n6321), .ZN(n6322) );
  XNOR2_X1 U8158 ( .A(n6322), .B(n6794), .ZN(n6326) );
  OR2_X1 U8159 ( .A1(n9953), .A2(n6796), .ZN(n6324) );
  NAND2_X1 U8160 ( .A1(n9172), .A2(n6451), .ZN(n6323) );
  NAND2_X1 U8161 ( .A1(n6324), .A2(n6323), .ZN(n6327) );
  XNOR2_X1 U8162 ( .A(n6326), .B(n6327), .ZN(n7503) );
  INV_X1 U8163 ( .A(n6326), .ZN(n6329) );
  INV_X1 U8164 ( .A(n6327), .ZN(n6328) );
  NAND2_X1 U8165 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  NAND2_X1 U8166 ( .A1(n7501), .A2(n6330), .ZN(n7583) );
  NAND2_X1 U8167 ( .A1(n9171), .A2(n6825), .ZN(n6331) );
  OAI21_X1 U8168 ( .B1(n9959), .B2(n6793), .A(n6331), .ZN(n6332) );
  XNOR2_X1 U8169 ( .A(n6332), .B(n6823), .ZN(n7585) );
  OR2_X1 U8170 ( .A1(n9959), .A2(n6796), .ZN(n6334) );
  NAND2_X1 U8171 ( .A1(n9171), .A2(n6451), .ZN(n6333) );
  AND2_X1 U8172 ( .A1(n6334), .A2(n6333), .ZN(n6336) );
  AND2_X1 U8173 ( .A1(n7585), .A2(n6336), .ZN(n6335) );
  INV_X1 U8174 ( .A(n7585), .ZN(n6337) );
  INV_X1 U8175 ( .A(n6336), .ZN(n7584) );
  NAND2_X1 U8176 ( .A1(n6337), .A2(n7584), .ZN(n6338) );
  NAND2_X1 U8177 ( .A1(n9967), .A2(n6286), .ZN(n6340) );
  NAND2_X1 U8178 ( .A1(n9170), .A2(n6288), .ZN(n6339) );
  NAND2_X1 U8179 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  XNOR2_X1 U8180 ( .A(n6341), .B(n6823), .ZN(n7796) );
  NAND2_X1 U8181 ( .A1(n9967), .A2(n6825), .ZN(n6343) );
  NAND2_X1 U8182 ( .A1(n9170), .A2(n6451), .ZN(n6342) );
  NAND2_X1 U8183 ( .A1(n9976), .A2(n6286), .ZN(n6346) );
  INV_X1 U8184 ( .A(n7680), .ZN(n9169) );
  NAND2_X1 U8185 ( .A1(n9169), .A2(n6825), .ZN(n6345) );
  NAND2_X1 U8186 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  XNOR2_X1 U8187 ( .A(n6347), .B(n6823), .ZN(n7858) );
  NOR2_X1 U8188 ( .A1(n7680), .A2(n6827), .ZN(n6348) );
  AOI21_X1 U8189 ( .B1(n9976), .B2(n6825), .A(n6348), .ZN(n6350) );
  AOI22_X1 U8190 ( .A1(n7858), .A2(n6350), .B1(n7800), .B2(n7796), .ZN(n6349)
         );
  INV_X1 U8191 ( .A(n7858), .ZN(n6351) );
  INV_X1 U8192 ( .A(n6350), .ZN(n7857) );
  INV_X1 U8193 ( .A(n6357), .ZN(n6354) );
  OAI22_X1 U8194 ( .A1(n5674), .A2(n6793), .B1(n7960), .B2(n6796), .ZN(n6353)
         );
  XOR2_X1 U8195 ( .A(n6794), .B(n6353), .Z(n6355) );
  INV_X1 U8196 ( .A(n6355), .ZN(n6356) );
  OAI22_X1 U8197 ( .A1(n5674), .A2(n6796), .B1(n7960), .B2(n6827), .ZN(n9748)
         );
  NAND2_X1 U8198 ( .A1(n9811), .A2(n6286), .ZN(n6360) );
  NAND2_X1 U8199 ( .A1(n9167), .A2(n6825), .ZN(n6359) );
  NAND2_X1 U8200 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  XNOR2_X1 U8201 ( .A(n6361), .B(n6823), .ZN(n6363) );
  NOR2_X1 U8202 ( .A1(n7726), .A2(n6827), .ZN(n6362) );
  AOI21_X1 U8203 ( .B1(n9811), .B2(n6825), .A(n6362), .ZN(n6364) );
  NAND2_X1 U8204 ( .A1(n6363), .A2(n6364), .ZN(n8030) );
  INV_X1 U8205 ( .A(n6363), .ZN(n6366) );
  INV_X1 U8206 ( .A(n6364), .ZN(n6365) );
  NAND2_X1 U8207 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  NAND2_X1 U8208 ( .A1(n7768), .A2(n6286), .ZN(n6369) );
  NAND2_X1 U8209 ( .A1(n9166), .A2(n6825), .ZN(n6368) );
  NAND2_X1 U8210 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  XNOR2_X1 U8211 ( .A(n6370), .B(n6823), .ZN(n6372) );
  NOR2_X1 U8212 ( .A1(n7961), .A2(n6827), .ZN(n6371) );
  AOI21_X1 U8213 ( .B1(n7768), .B2(n6825), .A(n6371), .ZN(n6373) );
  NAND2_X1 U8214 ( .A1(n6372), .A2(n6373), .ZN(n6377) );
  INV_X1 U8215 ( .A(n6372), .ZN(n6375) );
  INV_X1 U8216 ( .A(n6373), .ZN(n6374) );
  NAND2_X1 U8217 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  NAND2_X1 U8218 ( .A1(n6377), .A2(n6376), .ZN(n8029) );
  INV_X1 U8219 ( .A(n6377), .ZN(n6378) );
  AOI22_X1 U8220 ( .A1(n8089), .A2(n6288), .B1(n6451), .B2(n9165), .ZN(n6383)
         );
  NAND2_X1 U8221 ( .A1(n8089), .A2(n6286), .ZN(n6380) );
  NAND2_X1 U8222 ( .A1(n9165), .A2(n6825), .ZN(n6379) );
  NAND2_X1 U8223 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  XNOR2_X1 U8224 ( .A(n6381), .B(n6794), .ZN(n6382) );
  XOR2_X1 U8225 ( .A(n6383), .B(n6382), .Z(n8083) );
  INV_X1 U8226 ( .A(n6382), .ZN(n6384) );
  AOI22_X1 U8227 ( .A1(n9033), .A2(n6286), .B1(n6825), .B2(n9164), .ZN(n6385)
         );
  AOI22_X1 U8228 ( .A1(n9033), .A2(n6825), .B1(n6451), .B2(n9164), .ZN(n9027)
         );
  OAI22_X1 U8229 ( .A1(n8102), .A2(n6793), .B1(n8121), .B2(n6796), .ZN(n6386)
         );
  XNOR2_X1 U8230 ( .A(n6386), .B(n6794), .ZN(n6392) );
  NOR2_X1 U8231 ( .A1(n6393), .A2(n6392), .ZN(n6395) );
  INV_X1 U8232 ( .A(n6395), .ZN(n9061) );
  OAI22_X1 U8233 ( .A1(n9082), .A2(n6796), .B1(n9118), .B2(n6827), .ZN(n6407)
         );
  NAND2_X1 U8234 ( .A1(n9624), .A2(n6286), .ZN(n6388) );
  NAND2_X1 U8235 ( .A1(n9163), .A2(n6825), .ZN(n6387) );
  NAND2_X1 U8236 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  XNOR2_X1 U8237 ( .A(n6389), .B(n6794), .ZN(n6406) );
  XOR2_X1 U8238 ( .A(n6407), .B(n6406), .Z(n9075) );
  INV_X1 U8239 ( .A(n9075), .ZN(n6391) );
  OAI22_X1 U8240 ( .A1(n9668), .A2(n6793), .B1(n8146), .B2(n6796), .ZN(n6390)
         );
  XNOR2_X1 U8241 ( .A(n6390), .B(n6794), .ZN(n6400) );
  OAI22_X1 U8242 ( .A1(n9668), .A2(n6796), .B1(n8146), .B2(n6827), .ZN(n6399)
         );
  NOR2_X1 U8243 ( .A1(n6400), .A2(n6399), .ZN(n6398) );
  INV_X1 U8244 ( .A(n6398), .ZN(n9071) );
  AOI22_X1 U8245 ( .A1(n9142), .A2(n6825), .B1(n6451), .B2(n6096), .ZN(n9140)
         );
  NAND2_X1 U8246 ( .A1(n6396), .A2(n9060), .ZN(n6404) );
  INV_X1 U8247 ( .A(n6397), .ZN(n6402) );
  AOI21_X1 U8248 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n9063) );
  AND2_X1 U8249 ( .A1(n9063), .A2(n9075), .ZN(n6401) );
  OAI22_X1 U8250 ( .A1(n9662), .A2(n6793), .B1(n8168), .B2(n6796), .ZN(n6405)
         );
  XOR2_X1 U8251 ( .A(n6794), .B(n6405), .Z(n6411) );
  INV_X1 U8252 ( .A(n6411), .ZN(n6408) );
  OR2_X1 U8253 ( .A1(n6407), .A2(n6406), .ZN(n6410) );
  AND2_X1 U8254 ( .A1(n6408), .A2(n6410), .ZN(n6409) );
  AOI22_X1 U8255 ( .A1(n9426), .A2(n6825), .B1(n6451), .B2(n9162), .ZN(n9115)
         );
  NAND2_X1 U8256 ( .A1(n9483), .A2(n6286), .ZN(n6413) );
  NAND2_X1 U8257 ( .A1(n9161), .A2(n6825), .ZN(n6412) );
  NAND2_X1 U8258 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  XNOR2_X1 U8259 ( .A(n6414), .B(n6794), .ZN(n6420) );
  INV_X1 U8260 ( .A(n6420), .ZN(n6418) );
  NAND2_X1 U8261 ( .A1(n9483), .A2(n6825), .ZN(n6416) );
  NAND2_X1 U8262 ( .A1(n9161), .A2(n6451), .ZN(n6415) );
  NAND2_X1 U8263 ( .A1(n6416), .A2(n6415), .ZN(n6419) );
  INV_X1 U8264 ( .A(n6419), .ZN(n6417) );
  OAI22_X1 U8265 ( .A1(n9657), .A2(n6796), .B1(n8169), .B2(n6827), .ZN(n6424)
         );
  NAND2_X1 U8266 ( .A1(n9391), .A2(n6286), .ZN(n6422) );
  NAND2_X1 U8267 ( .A1(n9160), .A2(n6825), .ZN(n6421) );
  NAND2_X1 U8268 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  XNOR2_X1 U8269 ( .A(n6423), .B(n6794), .ZN(n6425) );
  XOR2_X1 U8270 ( .A(n6424), .B(n6425), .Z(n9096) );
  NAND2_X1 U8271 ( .A1(n9094), .A2(n9096), .ZN(n9095) );
  NAND2_X1 U8272 ( .A1(n9375), .A2(n4277), .ZN(n6428) );
  NAND2_X1 U8273 ( .A1(n9159), .A2(n6825), .ZN(n6427) );
  NAND2_X1 U8274 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  XNOR2_X1 U8275 ( .A(n6429), .B(n6794), .ZN(n6431) );
  XOR2_X1 U8276 ( .A(n6430), .B(n6431), .Z(n9052) );
  NAND2_X1 U8277 ( .A1(n9356), .A2(n6825), .ZN(n6433) );
  OR2_X1 U8278 ( .A1(n9053), .A2(n6827), .ZN(n6432) );
  NAND2_X1 U8279 ( .A1(n9356), .A2(n4277), .ZN(n6435) );
  OR2_X1 U8280 ( .A1(n9053), .A2(n6796), .ZN(n6434) );
  NAND2_X1 U8281 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  XNOR2_X1 U8282 ( .A(n6436), .B(n6794), .ZN(n6442) );
  NAND2_X1 U8283 ( .A1(n9463), .A2(n4277), .ZN(n6438) );
  NAND2_X1 U8284 ( .A1(n9157), .A2(n6825), .ZN(n6437) );
  NAND2_X1 U8285 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  XNOR2_X1 U8286 ( .A(n6439), .B(n6823), .ZN(n9041) );
  NOR2_X1 U8287 ( .A1(n9107), .A2(n6827), .ZN(n6440) );
  NOR2_X1 U8288 ( .A1(n9041), .A2(n9040), .ZN(n9039) );
  AOI21_X1 U8289 ( .B1(n9104), .B2(n6442), .A(n9039), .ZN(n6441) );
  INV_X1 U8290 ( .A(n9104), .ZN(n6443) );
  AOI21_X1 U8291 ( .B1(n9037), .B2(n6443), .A(n9040), .ZN(n6446) );
  INV_X1 U8292 ( .A(n9041), .ZN(n6445) );
  NAND3_X1 U8293 ( .A1(n9040), .A2(n6443), .A3(n9037), .ZN(n6444) );
  NAND2_X1 U8294 ( .A1(n9326), .A2(n6286), .ZN(n6449) );
  NAND2_X1 U8295 ( .A1(n9156), .A2(n6825), .ZN(n6448) );
  NAND2_X1 U8296 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  XNOR2_X1 U8297 ( .A(n6450), .B(n6794), .ZN(n6455) );
  NAND2_X1 U8298 ( .A1(n9326), .A2(n6825), .ZN(n6453) );
  NAND2_X1 U8299 ( .A1(n9156), .A2(n6451), .ZN(n6452) );
  NAND2_X1 U8300 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NOR2_X1 U8301 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  AOI21_X1 U8302 ( .B1(n6455), .B2(n6454), .A(n6456), .ZN(n9084) );
  NAND2_X1 U8303 ( .A1(n6460), .A2(n9084), .ZN(n9083) );
  INV_X1 U8304 ( .A(n6456), .ZN(n6457) );
  NAND2_X1 U8305 ( .A1(n9083), .A2(n6457), .ZN(n6461) );
  AND2_X1 U8306 ( .A1(n9084), .A2(n6462), .ZN(n6459) );
  INV_X1 U8307 ( .A(n6462), .ZN(n6458) );
  OAI21_X1 U8308 ( .B1(n6462), .B2(n6461), .A(n9125), .ZN(n6466) );
  NOR2_X1 U8309 ( .A1(n6464), .A2(n6463), .ZN(n7356) );
  NAND2_X1 U8310 ( .A1(n7356), .A2(n6524), .ZN(n6477) );
  INV_X1 U8311 ( .A(n6477), .ZN(n6469) );
  AND3_X1 U8312 ( .A1(n6896), .A2(n9991), .A3(n6470), .ZN(n6465) );
  AND2_X1 U8313 ( .A1(n6469), .A2(n6465), .ZN(n9148) );
  NAND2_X1 U8314 ( .A1(n6466), .A2(n9148), .ZN(n6484) );
  NAND2_X1 U8315 ( .A1(n7136), .A2(n6742), .ZN(n9880) );
  INV_X1 U8316 ( .A(n9880), .ZN(n7364) );
  NAND3_X1 U8317 ( .A1(n6469), .A2(n6896), .A3(n7364), .ZN(n6468) );
  AND2_X1 U8318 ( .A1(n6468), .A2(n9878), .ZN(n9749) );
  OAI22_X1 U8319 ( .A1(n6787), .A2(n9129), .B1(n6625), .B2(n9117), .ZN(n9306)
         );
  NOR2_X1 U8320 ( .A1(n6913), .A2(n6768), .ZN(n6780) );
  NAND2_X1 U8321 ( .A1(n6469), .A2(n6780), .ZN(n9090) );
  INV_X1 U8322 ( .A(n9090), .ZN(n9753) );
  AOI22_X1 U8323 ( .A1(n9306), .A2(n9753), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n6481) );
  NAND2_X1 U8324 ( .A1(n6477), .A2(n9991), .ZN(n6471) );
  NAND2_X1 U8325 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  NAND2_X1 U8326 ( .A1(n6472), .A2(n6768), .ZN(n6474) );
  AND2_X1 U8327 ( .A1(n6847), .A2(n6910), .ZN(n6473) );
  NAND2_X1 U8328 ( .A1(n6474), .A2(n6473), .ZN(n6479) );
  NOR2_X1 U8329 ( .A1(n9880), .A2(P1_U3086), .ZN(n6475) );
  OR2_X1 U8330 ( .A1(n6780), .A2(n6475), .ZN(n6476) );
  AND2_X1 U8331 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  AOI21_X1 U8332 ( .B1(n6479), .B2(P1_STATE_REG_SCAN_IN), .A(n6478), .ZN(n9135) );
  INV_X1 U8333 ( .A(n9135), .ZN(n9097) );
  NAND2_X1 U8334 ( .A1(n9097), .A2(n9312), .ZN(n6480) );
  OAI211_X1 U8335 ( .C1(n9315), .C2(n9749), .A(n6481), .B(n6480), .ZN(n6482)
         );
  NAND2_X1 U8336 ( .A1(n6484), .A2(n6483), .ZN(P1_U3225) );
  NOR2_X1 U8337 ( .A1(n8530), .A2(n8565), .ZN(n6485) );
  NAND2_X1 U8338 ( .A1(n8153), .A2(n8325), .ZN(n6488) );
  NAND2_X1 U8339 ( .A1(n4926), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8340 ( .A1(n8375), .A2(n8378), .ZN(n8376) );
  XOR2_X1 U8341 ( .A(n8365), .B(n8331), .Z(n8199) );
  NOR2_X1 U8342 ( .A1(n8530), .A2(n8529), .ZN(n6489) );
  AOI21_X1 U8343 ( .B1(n6490), .B2(n8330), .A(n6489), .ZN(n6491) );
  XNOR2_X1 U8344 ( .A(n6491), .B(n8331), .ZN(n6500) );
  INV_X1 U8345 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8346 ( .A1(n4959), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8347 ( .A1(n8316), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6492) );
  OAI211_X1 U8348 ( .C1(n6494), .C2(n4960), .A(n6493), .B(n6492), .ZN(n6495)
         );
  INV_X1 U8349 ( .A(n6495), .ZN(n6496) );
  AND2_X1 U8350 ( .A1(n8324), .A2(n6496), .ZN(n8329) );
  INV_X1 U8351 ( .A(n8867), .ZN(n8932) );
  NAND2_X1 U8352 ( .A1(n6497), .A2(P2_B_REG_SCAN_IN), .ZN(n6498) );
  NAND2_X1 U8353 ( .A1(n8932), .A2(n6498), .ZN(n8700) );
  OAI22_X1 U8354 ( .A1(n8529), .A2(n8865), .B1(n8329), .B2(n8700), .ZN(n6499)
         );
  AOI21_X2 U8355 ( .B1(n6500), .B2(n8928), .A(n6499), .ZN(n8203) );
  OAI21_X1 U8356 ( .B1(n8940), .B2(n8199), .A(n8203), .ZN(n6532) );
  NAND2_X1 U8357 ( .A1(n8944), .A2(n6501), .ZN(n6502) );
  OAI21_X1 U8358 ( .B1(n6532), .B2(n8944), .A(n6502), .ZN(n6503) );
  INV_X1 U8359 ( .A(n8375), .ZN(n6533) );
  OR2_X1 U8360 ( .A1(n8944), .A2(n8939), .ZN(n8908) );
  NAND2_X1 U8361 ( .A1(n6503), .A2(n4773), .ZN(P2_U3488) );
  INV_X1 U8362 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6509) );
  INV_X1 U8363 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6508) );
  MUX2_X1 U8364 ( .A(n6509), .B(n6508), .S(n6853), .Z(n6510) );
  XNOR2_X1 U8365 ( .A(n6510), .B(SI_31_), .ZN(n6511) );
  XNOR2_X1 U8366 ( .A(n6512), .B(n6511), .ZN(n9016) );
  XNOR2_X1 U8367 ( .A(n6516), .B(n8188), .ZN(n6517) );
  OR2_X1 U8368 ( .A1(n6526), .A2(n9998), .ZN(n6523) );
  INV_X1 U8369 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U8370 ( .A1(n6523), .A2(n6522), .ZN(P1_U3521) );
  INV_X1 U8371 ( .A(n6524), .ZN(n7357) );
  INV_X2 U8372 ( .A(n10013), .ZN(n10015) );
  OR2_X1 U8373 ( .A1(n6526), .A2(n10013), .ZN(n6531) );
  NAND2_X1 U8374 ( .A1(n10015), .A2(n9977), .ZN(n9633) );
  NOR2_X1 U8375 ( .A1(n10015), .A2(n6527), .ZN(n6528) );
  NAND2_X1 U8376 ( .A1(n6531), .A2(n6530), .ZN(P1_U3553) );
  OAI21_X1 U8377 ( .B1(n6532), .B2(n10060), .A(n4762), .ZN(n6534) );
  OR2_X1 U8378 ( .A1(n10060), .A2(n8939), .ZN(n8989) );
  NAND2_X1 U8379 ( .A1(n6534), .A2(n4765), .ZN(P2_U3456) );
  OAI21_X1 U8380 ( .B1(n6672), .B2(n6649), .A(n9151), .ZN(n6650) );
  NAND2_X1 U8381 ( .A1(n9356), .A2(n9053), .ZN(n6535) );
  NAND2_X1 U8382 ( .A1(n6679), .A2(n6535), .ZN(n6685) );
  MUX2_X1 U8383 ( .A(n6536), .B(n6697), .S(n6649), .Z(n6537) );
  INV_X1 U8384 ( .A(n6537), .ZN(n6620) );
  INV_X1 U8385 ( .A(n6700), .ZN(n6540) );
  OAI211_X1 U8386 ( .C1(n6538), .C2(n6540), .A(n9851), .B(n6539), .ZN(n6541)
         );
  NAND3_X1 U8387 ( .A1(n6541), .A2(n6704), .A3(n4792), .ZN(n6543) );
  NAND3_X1 U8388 ( .A1(n6543), .A2(n6546), .A3(n6542), .ZN(n6544) );
  NAND2_X1 U8389 ( .A1(n6544), .A2(n6545), .ZN(n6548) );
  NAND2_X1 U8390 ( .A1(n7470), .A2(n6545), .ZN(n6547) );
  NAND2_X1 U8391 ( .A1(n6547), .A2(n6546), .ZN(n9839) );
  MUX2_X1 U8392 ( .A(n6548), .B(n9839), .S(n6649), .Z(n6549) );
  NAND2_X1 U8393 ( .A1(n6549), .A2(n7557), .ZN(n6555) );
  NAND2_X1 U8394 ( .A1(n9818), .A2(n6550), .ZN(n6552) );
  MUX2_X1 U8395 ( .A(n6552), .B(n6551), .S(n6649), .Z(n6553) );
  INV_X1 U8396 ( .A(n6553), .ZN(n6554) );
  NAND2_X1 U8397 ( .A1(n6555), .A2(n6554), .ZN(n6561) );
  NAND2_X1 U8398 ( .A1(n6563), .A2(n6556), .ZN(n6558) );
  MUX2_X1 U8399 ( .A(n6558), .B(n6557), .S(n6649), .Z(n6559) );
  INV_X1 U8400 ( .A(n6559), .ZN(n6560) );
  NAND2_X1 U8401 ( .A1(n6561), .A2(n6560), .ZN(n6570) );
  INV_X1 U8402 ( .A(n6708), .ZN(n6562) );
  AOI21_X1 U8403 ( .B1(n6570), .B2(n6563), .A(n6562), .ZN(n6565) );
  OR2_X1 U8404 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  INV_X1 U8405 ( .A(n6715), .ZN(n7777) );
  AOI21_X1 U8406 ( .B1(n6566), .B2(n6713), .A(n7777), .ZN(n6568) );
  NAND4_X1 U8407 ( .A1(n6722), .A2(n6718), .A3(n7991), .A4(n6649), .ZN(n6567)
         );
  NAND2_X1 U8408 ( .A1(n6570), .A2(n6569), .ZN(n6571) );
  NAND2_X1 U8409 ( .A1(n6571), .A2(n9803), .ZN(n6572) );
  NAND3_X1 U8410 ( .A1(n6572), .A2(n6708), .A3(n7722), .ZN(n6574) );
  NAND3_X1 U8411 ( .A1(n6574), .A2(n6715), .A3(n6573), .ZN(n6576) );
  NAND2_X1 U8412 ( .A1(n6576), .A2(n6575), .ZN(n6578) );
  NAND2_X1 U8413 ( .A1(n9033), .A2(n7997), .ZN(n6577) );
  AND2_X1 U8414 ( .A1(n6589), .A2(n6577), .ZN(n6721) );
  INV_X1 U8415 ( .A(n6649), .ZN(n6641) );
  NAND4_X1 U8416 ( .A1(n6578), .A2(n6721), .A3(n6641), .A4(n6716), .ZN(n6592)
         );
  NAND2_X1 U8417 ( .A1(n9165), .A2(n6641), .ZN(n6579) );
  OAI22_X1 U8418 ( .A1(n7991), .A2(n6649), .B1(n8089), .B2(n6579), .ZN(n6580)
         );
  NAND2_X1 U8419 ( .A1(n6721), .A2(n6580), .ZN(n6588) );
  NOR2_X1 U8420 ( .A1(n9165), .A2(n6641), .ZN(n6581) );
  NAND2_X1 U8421 ( .A1(n8089), .A2(n6581), .ZN(n6582) );
  OAI21_X1 U8422 ( .B1(n6641), .B2(n9164), .A(n6582), .ZN(n6584) );
  INV_X1 U8423 ( .A(n6582), .ZN(n6583) );
  AOI22_X1 U8424 ( .A1(n6584), .A2(n9033), .B1(n6583), .B2(n7997), .ZN(n6585)
         );
  NAND2_X1 U8425 ( .A1(n6722), .A2(n6585), .ZN(n6586) );
  OAI21_X1 U8426 ( .B1(n6722), .B2(n6641), .A(n6586), .ZN(n6587) );
  OAI211_X1 U8427 ( .C1(n6641), .C2(n6589), .A(n6588), .B(n6587), .ZN(n6590)
         );
  NOR2_X1 U8428 ( .A1(n6590), .A2(n8117), .ZN(n6591) );
  NAND3_X1 U8429 ( .A1(n6593), .A2(n6592), .A3(n6591), .ZN(n6597) );
  AOI21_X1 U8430 ( .B1(n6604), .B2(n6724), .A(n6649), .ZN(n6595) );
  NOR2_X1 U8431 ( .A1(n6595), .A2(n6594), .ZN(n6596) );
  AND2_X1 U8432 ( .A1(n6606), .A2(n6598), .ZN(n6728) );
  NAND2_X1 U8433 ( .A1(n6610), .A2(n6728), .ZN(n6599) );
  NAND3_X1 U8434 ( .A1(n6599), .A2(n9404), .A3(n6729), .ZN(n6600) );
  AND2_X1 U8435 ( .A1(n6654), .A2(n6729), .ZN(n6601) );
  NAND2_X1 U8436 ( .A1(n9366), .A2(n6608), .ZN(n6612) );
  NAND2_X1 U8437 ( .A1(n9404), .A2(n6604), .ZN(n6726) );
  OR2_X1 U8438 ( .A1(n6726), .A2(n6605), .ZN(n6607) );
  AND3_X1 U8439 ( .A1(n6608), .A2(n6607), .A3(n6606), .ZN(n6698) );
  INV_X1 U8440 ( .A(n6726), .ZN(n6609) );
  AOI21_X1 U8441 ( .B1(n6610), .B2(n6609), .A(n6641), .ZN(n6611) );
  AOI22_X1 U8442 ( .A1(n6612), .A2(n6641), .B1(n6698), .B2(n6611), .ZN(n6613)
         );
  NAND2_X1 U8443 ( .A1(n6614), .A2(n6613), .ZN(n6619) );
  MUX2_X1 U8444 ( .A(n6616), .B(n6615), .S(n6649), .Z(n6617) );
  INV_X1 U8445 ( .A(n6617), .ZN(n6618) );
  OR2_X1 U8446 ( .A1(n9463), .A2(n9107), .ZN(n6623) );
  AND2_X1 U8447 ( .A1(n6623), .A2(n6622), .ZN(n6678) );
  NAND2_X1 U8448 ( .A1(n6624), .A2(n9321), .ZN(n6627) );
  NAND2_X1 U8449 ( .A1(n9326), .A2(n6625), .ZN(n6687) );
  MUX2_X1 U8450 ( .A(n6687), .B(n6681), .S(n6649), .Z(n6626) );
  NAND2_X1 U8451 ( .A1(n6633), .A2(n9283), .ZN(n6628) );
  AND2_X1 U8452 ( .A1(n6634), .A2(n6631), .ZN(n6677) );
  NAND2_X1 U8453 ( .A1(n6637), .A2(n6636), .ZN(n6696) );
  AOI21_X1 U8454 ( .B1(n6628), .B2(n6677), .A(n6696), .ZN(n6629) );
  NAND2_X1 U8455 ( .A1(n6642), .A2(n6635), .ZN(n6694) );
  OAI21_X1 U8456 ( .B1(n6629), .B2(n6694), .A(n6675), .ZN(n6630) );
  NAND2_X1 U8457 ( .A1(n6630), .A2(n6641), .ZN(n6646) );
  NAND2_X1 U8458 ( .A1(n6675), .A2(n6637), .ZN(n6638) );
  NAND2_X1 U8459 ( .A1(n6640), .A2(n6639), .ZN(n6645) );
  NOR2_X1 U8460 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  MUX2_X1 U8461 ( .A(n6737), .B(n6676), .S(n6649), .Z(n6647) );
  AND2_X1 U8462 ( .A1(n6915), .A2(n9151), .ZN(n6648) );
  AOI21_X1 U8463 ( .B1(n6672), .B2(n6649), .A(n6648), .ZN(n6651) );
  NAND2_X1 U8464 ( .A1(n6652), .A2(n6760), .ZN(n6653) );
  NAND2_X1 U8465 ( .A1(n6653), .A2(n6770), .ZN(n6774) );
  OAI21_X1 U8466 ( .B1(n6774), .B2(n7772), .A(n6655), .ZN(n6674) );
  OR2_X1 U8467 ( .A1(n6672), .A2(n6671), .ZN(n6755) );
  INV_X1 U8468 ( .A(n9321), .ZN(n9319) );
  NAND2_X1 U8469 ( .A1(n9366), .A2(n6654), .ZN(n9365) );
  INV_X1 U8470 ( .A(n8117), .ZN(n8119) );
  XOR2_X1 U8471 ( .A(n9811), .B(n9167), .Z(n9804) );
  NOR3_X1 U8472 ( .A1(n7359), .A2(n6655), .A3(n9881), .ZN(n6656) );
  AND2_X1 U8473 ( .A1(n6275), .A2(n9902), .ZN(n6702) );
  NOR2_X1 U8474 ( .A1(n9893), .A2(n6702), .ZN(n7380) );
  NAND4_X1 U8475 ( .A1(n7348), .A2(n6656), .A3(n7380), .A4(n9892), .ZN(n6657)
         );
  NOR4_X1 U8476 ( .A1(n6659), .A2(n6658), .A3(n9861), .A4(n6657), .ZN(n6660)
         );
  NAND4_X1 U8477 ( .A1(n7730), .A2(n7683), .A3(n6661), .A4(n6660), .ZN(n6662)
         );
  NOR4_X1 U8478 ( .A1(n8001), .A2(n9804), .A3(n7786), .A4(n6662), .ZN(n6664)
         );
  NAND4_X1 U8479 ( .A1(n8145), .A2(n8119), .A3(n6664), .A4(n6663), .ZN(n6665)
         );
  NOR4_X1 U8480 ( .A1(n9365), .A2(n9405), .A3(n9421), .A4(n6665), .ZN(n6666)
         );
  NAND4_X1 U8481 ( .A1(n9339), .A2(n9367), .A3(n6666), .A4(n9349), .ZN(n6667)
         );
  OR4_X1 U8482 ( .A1(n6668), .A2(n9319), .A3(n9302), .A4(n6667), .ZN(n6670) );
  NOR4_X1 U8483 ( .A1(n6670), .A2(n6669), .A3(n9257), .A4(n9284), .ZN(n6673)
         );
  NAND2_X1 U8484 ( .A1(n6672), .A2(n6671), .ZN(n6738) );
  NAND4_X1 U8485 ( .A1(n6740), .A2(n6673), .A3(n6738), .A4(n6770), .ZN(n6763)
         );
  NAND2_X1 U8486 ( .A1(n6674), .A2(n6763), .ZN(n6746) );
  NAND2_X1 U8487 ( .A1(n6676), .A2(n6675), .ZN(n6752) );
  INV_X1 U8488 ( .A(n6677), .ZN(n6691) );
  INV_X1 U8489 ( .A(n6678), .ZN(n6680) );
  NAND2_X1 U8490 ( .A1(n6680), .A2(n6679), .ZN(n6682) );
  NAND2_X1 U8491 ( .A1(n6682), .A2(n6681), .ZN(n6683) );
  NAND2_X1 U8492 ( .A1(n6683), .A2(n6687), .ZN(n6684) );
  NAND2_X1 U8493 ( .A1(n9283), .A2(n6684), .ZN(n6695) );
  INV_X1 U8494 ( .A(n6685), .ZN(n6688) );
  AND3_X1 U8495 ( .A1(n6688), .A2(n6687), .A3(n6686), .ZN(n6689) );
  NOR2_X1 U8496 ( .A1(n6695), .A2(n6689), .ZN(n6690) );
  NOR2_X1 U8497 ( .A1(n6691), .A2(n6690), .ZN(n6692) );
  NOR2_X1 U8498 ( .A1(n6692), .A2(n6696), .ZN(n6693) );
  OR2_X1 U8499 ( .A1(n6694), .A2(n6693), .ZN(n6748) );
  OR2_X1 U8500 ( .A1(n6696), .A2(n6695), .ZN(n6749) );
  INV_X1 U8501 ( .A(n6697), .ZN(n6733) );
  INV_X1 U8502 ( .A(n6698), .ZN(n6731) );
  AND3_X1 U8503 ( .A1(n6700), .A2(n4792), .A3(n6699), .ZN(n6706) );
  AOI21_X1 U8504 ( .B1(n6701), .B2(n6268), .A(n7643), .ZN(n6705) );
  INV_X1 U8505 ( .A(n6702), .ZN(n6703) );
  AND4_X1 U8506 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n6709)
         );
  OAI211_X1 U8507 ( .C1(n6710), .C2(n6709), .A(n6708), .B(n6707), .ZN(n6712)
         );
  NAND2_X1 U8508 ( .A1(n6712), .A2(n6711), .ZN(n6714) );
  NAND2_X1 U8509 ( .A1(n6714), .A2(n6713), .ZN(n6717) );
  NAND3_X1 U8510 ( .A1(n6717), .A2(n6716), .A3(n6715), .ZN(n6719) );
  NAND3_X1 U8511 ( .A1(n6719), .A2(n6718), .A3(n7991), .ZN(n6720) );
  NAND2_X1 U8512 ( .A1(n6721), .A2(n6720), .ZN(n6723) );
  NAND2_X1 U8513 ( .A1(n6723), .A2(n6722), .ZN(n6725) );
  NAND2_X1 U8514 ( .A1(n6725), .A2(n6724), .ZN(n6727) );
  AOI21_X1 U8515 ( .B1(n6728), .B2(n6727), .A(n6726), .ZN(n6730) );
  OAI21_X1 U8516 ( .B1(n6731), .B2(n6730), .A(n6729), .ZN(n6732) );
  NAND2_X1 U8517 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  NOR2_X1 U8518 ( .A1(n6749), .A2(n6734), .ZN(n6735) );
  NOR2_X1 U8519 ( .A1(n6748), .A2(n6735), .ZN(n6736) );
  NOR2_X1 U8520 ( .A1(n6752), .A2(n6736), .ZN(n6739) );
  NAND2_X1 U8521 ( .A1(n6738), .A2(n6737), .ZN(n6757) );
  NAND2_X1 U8522 ( .A1(n6740), .A2(n4784), .ZN(n6741) );
  NAND2_X1 U8523 ( .A1(n6741), .A2(n6770), .ZN(n6767) );
  OAI21_X1 U8524 ( .B1(n6767), .B2(n6742), .A(n6760), .ZN(n6743) );
  INV_X1 U8525 ( .A(n6743), .ZN(n6744) );
  OAI21_X1 U8526 ( .B1(n6746), .B2(n6745), .A(n6744), .ZN(n6747) );
  NAND2_X1 U8527 ( .A1(n6747), .A2(n6219), .ZN(n6766) );
  INV_X1 U8528 ( .A(n6748), .ZN(n6754) );
  INV_X1 U8529 ( .A(n6749), .ZN(n6751) );
  NAND2_X1 U8530 ( .A1(n6751), .A2(n6750), .ZN(n6753) );
  AOI21_X1 U8531 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(n6758) );
  INV_X1 U8532 ( .A(n6915), .ZN(n6756) );
  OAI22_X1 U8533 ( .A1(n6758), .A2(n6757), .B1(n6756), .B2(n6755), .ZN(n6759)
         );
  OAI211_X1 U8534 ( .C1(n5759), .C2(n6915), .A(n6759), .B(n6770), .ZN(n6761)
         );
  NAND3_X1 U8535 ( .A1(n6761), .A2(n6911), .A3(n6760), .ZN(n6762) );
  AOI21_X1 U8536 ( .B1(n6763), .B2(n6762), .A(n6745), .ZN(n6764) );
  NAND2_X1 U8537 ( .A1(n6764), .A2(n8189), .ZN(n6765) );
  NAND2_X1 U8538 ( .A1(n6766), .A2(n6765), .ZN(n6779) );
  INV_X1 U8539 ( .A(n6767), .ZN(n6769) );
  INV_X1 U8540 ( .A(n6770), .ZN(n6772) );
  AOI211_X1 U8541 ( .C1(n6772), .C2(n6219), .A(n6220), .B(n6771), .ZN(n6773)
         );
  NAND2_X1 U8542 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  NAND2_X1 U8543 ( .A1(n4775), .A2(n6775), .ZN(n6778) );
  INV_X1 U8544 ( .A(n6910), .ZN(n6776) );
  NAND2_X1 U8545 ( .A1(n6776), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7760) );
  INV_X1 U8546 ( .A(n7760), .ZN(n6777) );
  OAI21_X1 U8547 ( .B1(n6779), .B2(n6778), .A(n6777), .ZN(n6783) );
  INV_X1 U8548 ( .A(n5779), .ZN(n9761) );
  NAND3_X1 U8549 ( .A1(n9131), .A2(n6780), .A3(n9761), .ZN(n6781) );
  OAI211_X1 U8550 ( .C1(n6220), .C2(n7760), .A(n6781), .B(P1_B_REG_SCAN_IN), 
        .ZN(n6782) );
  NAND2_X1 U8551 ( .A1(n6783), .A2(n6782), .ZN(P1_U3242) );
  NAND2_X1 U8552 ( .A1(n9293), .A2(n6286), .ZN(n6785) );
  INV_X1 U8553 ( .A(n6787), .ZN(n9154) );
  NAND2_X1 U8554 ( .A1(n9154), .A2(n6825), .ZN(n6784) );
  NAND2_X1 U8555 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  XNOR2_X1 U8556 ( .A(n6786), .B(n6794), .ZN(n6801) );
  NOR2_X1 U8557 ( .A1(n6787), .A2(n6827), .ZN(n6788) );
  AOI21_X1 U8558 ( .B1(n9293), .B2(n6825), .A(n6788), .ZN(n6799) );
  XNOR2_X1 U8559 ( .A(n6801), .B(n6799), .ZN(n9127) );
  INV_X1 U8560 ( .A(n6789), .ZN(n6790) );
  NAND2_X1 U8561 ( .A1(n6791), .A2(n6790), .ZN(n9124) );
  OAI22_X1 U8562 ( .A1(n9272), .A2(n6793), .B1(n9130), .B2(n6796), .ZN(n6795)
         );
  XNOR2_X1 U8563 ( .A(n6795), .B(n6794), .ZN(n6798) );
  OAI22_X1 U8564 ( .A1(n9272), .A2(n6796), .B1(n9130), .B2(n6827), .ZN(n6797)
         );
  NOR2_X1 U8565 ( .A1(n6798), .A2(n6797), .ZN(n6833) );
  AOI21_X1 U8566 ( .B1(n6798), .B2(n6797), .A(n6833), .ZN(n6805) );
  INV_X1 U8567 ( .A(n6805), .ZN(n6803) );
  INV_X1 U8568 ( .A(n6799), .ZN(n6800) );
  NAND2_X1 U8569 ( .A1(n6801), .A2(n6800), .ZN(n6806) );
  INV_X1 U8570 ( .A(n6806), .ZN(n6802) );
  NOR2_X1 U8571 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  AOI21_X1 U8572 ( .B1(n9126), .B2(n6806), .A(n6805), .ZN(n6807) );
  OAI21_X1 U8573 ( .B1(n6842), .B2(n6807), .A(n9148), .ZN(n6815) );
  OR2_X1 U8574 ( .A1(n7251), .A2(n9129), .ZN(n6809) );
  NAND2_X1 U8575 ( .A1(n9154), .A2(n9131), .ZN(n6808) );
  AND2_X1 U8576 ( .A1(n6809), .A2(n6808), .ZN(n9276) );
  OAI22_X1 U8577 ( .A1(n9276), .A2(n9090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6810), .ZN(n6811) );
  AOI21_X1 U8578 ( .B1(n9270), .B2(n9097), .A(n6811), .ZN(n6812) );
  NAND2_X1 U8579 ( .A1(n6815), .A2(n6814), .ZN(P1_U3214) );
  NAND2_X1 U8580 ( .A1(n6816), .A2(n10015), .ZN(n6820) );
  NAND2_X1 U8581 ( .A1(n10013), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6817) );
  INV_X1 U8582 ( .A(n6818), .ZN(n6819) );
  NAND2_X1 U8583 ( .A1(n6820), .A2(n6819), .ZN(P1_U3551) );
  INV_X1 U8584 ( .A(n6842), .ZN(n6832) );
  INV_X1 U8585 ( .A(n6833), .ZN(n6831) );
  NAND2_X1 U8586 ( .A1(n9261), .A2(n4277), .ZN(n6822) );
  OR2_X1 U8587 ( .A1(n7251), .A2(n6796), .ZN(n6821) );
  NAND2_X1 U8588 ( .A1(n6822), .A2(n6821), .ZN(n6824) );
  XNOR2_X1 U8589 ( .A(n6824), .B(n6823), .ZN(n6829) );
  NAND2_X1 U8590 ( .A1(n9261), .A2(n6825), .ZN(n6826) );
  OAI21_X1 U8591 ( .B1(n7251), .B2(n6827), .A(n6826), .ZN(n6828) );
  XNOR2_X1 U8592 ( .A(n6829), .B(n6828), .ZN(n6834) );
  INV_X1 U8593 ( .A(n6834), .ZN(n6830) );
  NAND2_X1 U8594 ( .A1(n6832), .A2(n4772), .ZN(n6844) );
  AND2_X1 U8595 ( .A1(n6834), .A2(n9148), .ZN(n6841) );
  NAND3_X1 U8596 ( .A1(n6834), .A2(n9148), .A3(n6833), .ZN(n6839) );
  INV_X1 U8597 ( .A(n9749), .ZN(n9141) );
  INV_X1 U8598 ( .A(n9130), .ZN(n9153) );
  INV_X1 U8599 ( .A(n6835), .ZN(n9152) );
  INV_X1 U8600 ( .A(n9129), .ZN(n9086) );
  AOI22_X1 U8601 ( .A1(n9153), .A2(n9131), .B1(n9152), .B2(n9086), .ZN(n9254)
         );
  AOI22_X1 U8602 ( .A1(n9262), .A2(n9097), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6836) );
  OAI21_X1 U8603 ( .B1(n9254), .B2(n9090), .A(n6836), .ZN(n6837) );
  AOI21_X1 U8604 ( .B1(n9261), .B2(n9141), .A(n6837), .ZN(n6838) );
  NAND2_X1 U8605 ( .A1(n6844), .A2(n6843), .ZN(P1_U3220) );
  INV_X1 U8606 ( .A(n6845), .ZN(n6846) );
  INV_X1 U8607 ( .A(n9177), .ZN(P1_U3973) );
  XNOR2_X1 U8608 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U8609 ( .A(n6849), .B(n5599), .S(P1_STATE_REG_SCAN_IN), .Z(n6850) );
  INV_X1 U8610 ( .A(n6850), .ZN(P1_U3355) );
  OR2_X1 U8611 ( .A1(n6853), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8194) );
  OAI222_X1 U8612 ( .A1(n8194), .A2(n6851), .B1(n9675), .B2(n6858), .C1(
        P1_U3086), .C2(n6979), .ZN(P1_U3352) );
  OAI222_X1 U8613 ( .A1(n8194), .A2(n6852), .B1(n9675), .B2(n6856), .C1(
        P1_U3086), .C2(n9797), .ZN(P1_U3351) );
  AND2_X1 U8614 ( .A1(n6853), .A2(P2_U3151), .ZN(n8093) );
  INV_X2 U8615 ( .A(n8093), .ZN(n9021) );
  OR2_X1 U8616 ( .A1(n6853), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9024) );
  CLKBUF_X1 U8617 ( .A(n9024), .Z(n8056) );
  OAI222_X1 U8618 ( .A1(n9021), .A2(n6854), .B1(n8056), .B2(n6869), .C1(n7028), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  OAI222_X1 U8619 ( .A1(n7068), .A2(P2_U3151), .B1(n8056), .B2(n6856), .C1(
        n6855), .C2(n9021), .ZN(P2_U3291) );
  OAI222_X1 U8620 ( .A1(P2_U3151), .A2(n7118), .B1(n8056), .B2(n6873), .C1(
        n4843), .C2(n9021), .ZN(P2_U3290) );
  OAI222_X1 U8621 ( .A1(n7045), .A2(P2_U3151), .B1(n9024), .B2(n6867), .C1(
        n6857), .C2(n9021), .ZN(P2_U3293) );
  OAI222_X1 U8622 ( .A1(n6859), .A2(P2_U3151), .B1(n8056), .B2(n6858), .C1(
        n4407), .C2(n9021), .ZN(P2_U3292) );
  NAND2_X1 U8623 ( .A1(n6861), .A2(n6860), .ZN(n6883) );
  NOR2_X1 U8624 ( .A1(n6863), .A2(n6862), .ZN(n6865) );
  AOI22_X1 U8625 ( .A1(n6883), .A2(n6864), .B1(n6865), .B2(n7970), .ZN(
        P2_U3377) );
  AOI22_X1 U8626 ( .A1(n6883), .A2(n6866), .B1(n6865), .B2(n7933), .ZN(
        P2_U3376) );
  OAI222_X1 U8627 ( .A1(n8194), .A2(n6868), .B1(n9675), .B2(n6867), .C1(
        P1_U3086), .C2(n7193), .ZN(P1_U3353) );
  INV_X1 U8628 ( .A(n8194), .ZN(n9673) );
  INV_X1 U8629 ( .A(n9673), .ZN(n8195) );
  OAI222_X1 U8630 ( .A1(n8195), .A2(n6870), .B1(n9675), .B2(n6869), .C1(
        P1_U3086), .C2(n6930), .ZN(P1_U3354) );
  OAI222_X1 U8631 ( .A1(n9675), .A2(n6873), .B1(n6872), .B2(P1_U3086), .C1(
        n6871), .C2(n8195), .ZN(P1_U3350) );
  INV_X1 U8632 ( .A(n6874), .ZN(n6877) );
  OAI222_X1 U8633 ( .A1(n8194), .A2(n6875), .B1(n9675), .B2(n6877), .C1(
        P1_U3086), .C2(n7005), .ZN(P1_U3349) );
  OAI222_X1 U8634 ( .A1(n6878), .A2(P2_U3151), .B1(n8056), .B2(n6877), .C1(
        n6876), .C2(n9021), .ZN(P2_U3289) );
  INV_X1 U8635 ( .A(n6879), .ZN(n6882) );
  INV_X1 U8636 ( .A(n7099), .ZN(n7012) );
  OAI222_X1 U8637 ( .A1(n8194), .A2(n6880), .B1(n9675), .B2(n6882), .C1(
        P1_U3086), .C2(n7012), .ZN(P1_U3348) );
  OAI222_X1 U8638 ( .A1(n7392), .A2(P2_U3151), .B1(n8056), .B2(n6882), .C1(
        n6881), .C2(n9021), .ZN(P2_U3288) );
  INV_X1 U8639 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6884) );
  NOR2_X1 U8640 ( .A1(n6943), .A2(n6884), .ZN(P2_U3257) );
  INV_X1 U8641 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6885) );
  NOR2_X1 U8642 ( .A1(n6943), .A2(n6885), .ZN(P2_U3246) );
  INV_X1 U8643 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6886) );
  NOR2_X1 U8644 ( .A1(n6943), .A2(n6886), .ZN(P2_U3247) );
  INV_X1 U8645 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6887) );
  NOR2_X1 U8646 ( .A1(n6943), .A2(n6887), .ZN(P2_U3255) );
  INV_X1 U8647 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6888) );
  NOR2_X1 U8648 ( .A1(n6943), .A2(n6888), .ZN(P2_U3256) );
  INV_X1 U8649 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6889) );
  NOR2_X1 U8650 ( .A1(n6943), .A2(n6889), .ZN(P2_U3254) );
  INV_X1 U8651 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6890) );
  NOR2_X1 U8652 ( .A1(n6943), .A2(n6890), .ZN(P2_U3252) );
  INV_X1 U8653 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6891) );
  NOR2_X1 U8654 ( .A1(n6943), .A2(n6891), .ZN(P2_U3253) );
  INV_X1 U8655 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6892) );
  NOR2_X1 U8656 ( .A1(n6943), .A2(n6892), .ZN(P2_U3249) );
  INV_X1 U8657 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6893) );
  NOR2_X1 U8658 ( .A1(n6943), .A2(n6893), .ZN(P2_U3248) );
  INV_X1 U8659 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6894) );
  NOR2_X1 U8660 ( .A1(n6943), .A2(n6894), .ZN(P2_U3250) );
  INV_X1 U8661 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6895) );
  NOR2_X1 U8662 ( .A1(n6943), .A2(n6895), .ZN(P2_U3251) );
  AND2_X1 U8663 ( .A1(n6897), .A2(n6896), .ZN(n9915) );
  INV_X1 U8664 ( .A(n9915), .ZN(n9916) );
  NAND2_X1 U8665 ( .A1(n9916), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6898) );
  OAI21_X1 U8666 ( .B1(n9916), .B2(n6899), .A(n6898), .ZN(P1_U3439) );
  INV_X1 U8667 ( .A(n6900), .ZN(n6903) );
  OAI222_X1 U8668 ( .A1(n8194), .A2(n6901), .B1(n9675), .B2(n6903), .C1(
        P1_U3086), .C2(n4480), .ZN(P1_U3347) );
  OAI222_X1 U8669 ( .A1(n8587), .A2(P2_U3151), .B1(n8056), .B2(n6903), .C1(
        n6902), .C2(n9021), .ZN(P2_U3287) );
  INV_X1 U8670 ( .A(P2_U3893), .ZN(n8687) );
  NAND2_X1 U8671 ( .A1(n8687), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n6904) );
  OAI21_X1 U8672 ( .B1(n8866), .B2(n8687), .A(n6904), .ZN(P2_U3505) );
  INV_X1 U8673 ( .A(n6905), .ZN(n6908) );
  INV_X1 U8674 ( .A(n7291), .ZN(n7162) );
  OAI222_X1 U8675 ( .A1(n9675), .A2(n6908), .B1(n7162), .B2(P1_U3086), .C1(
        n6906), .C2(n8194), .ZN(P1_U3346) );
  OAI222_X1 U8676 ( .A1(P2_U3151), .A2(n6909), .B1(n8056), .B2(n6908), .C1(
        n6907), .C2(n9021), .ZN(P2_U3286) );
  NAND2_X1 U8677 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  NAND2_X1 U8678 ( .A1(n5621), .A2(n6912), .ZN(n6923) );
  AND2_X1 U8679 ( .A1(n6913), .A2(n7760), .ZN(n6922) );
  INV_X1 U8680 ( .A(n6922), .ZN(n6914) );
  AND2_X1 U8681 ( .A1(n6923), .A2(n6914), .ZN(n9794) );
  NOR2_X1 U8682 ( .A1(n9794), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8683 ( .A1(n6915), .A2(P1_U3973), .ZN(n6916) );
  OAI21_X1 U8684 ( .B1(n6509), .B2(P1_U3973), .A(n6916), .ZN(P1_U3585) );
  NAND2_X1 U8685 ( .A1(n9177), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6917) );
  OAI21_X1 U8686 ( .B1(n8146), .B2(n9177), .A(n6917), .ZN(P1_U3570) );
  INV_X1 U8687 ( .A(n6918), .ZN(n6921) );
  INV_X1 U8688 ( .A(n7429), .ZN(n7434) );
  INV_X1 U8689 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6919) );
  OAI222_X1 U8690 ( .A1(n9675), .A2(n6921), .B1(n7434), .B2(P1_U3086), .C1(
        n6919), .C2(n8195), .ZN(P1_U3345) );
  OAI222_X1 U8691 ( .A1(P2_U3151), .A2(n7742), .B1(n8056), .B2(n6921), .C1(
        n6920), .C2(n9021), .ZN(P2_U3285) );
  OR2_X1 U8692 ( .A1(n6923), .A2(n6922), .ZN(n9770) );
  OR2_X1 U8693 ( .A1(n9770), .A2(n7182), .ZN(n9798) );
  INV_X1 U8694 ( .A(n9798), .ZN(n9776) );
  OR2_X1 U8695 ( .A1(n9770), .A2(n9761), .ZN(n9242) );
  INV_X1 U8696 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10005) );
  MUX2_X1 U8697 ( .A(n10005), .B(P1_REG1_REG_4__SCAN_IN), .S(n9797), .Z(n9791)
         );
  MUX2_X1 U8698 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6924), .S(n6934), .Z(n6974)
         );
  INV_X1 U8699 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U8700 ( .A1(n6932), .A2(P1_REG1_REG_2__SCAN_IN), .B1(n10002), .B2(
        n7193), .ZN(n7185) );
  MUX2_X1 U8701 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6925), .S(n9775), .Z(n9779)
         );
  NAND3_X1 U8702 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n9779), .ZN(n9778) );
  OAI21_X1 U8703 ( .B1(n6925), .B2(n6930), .A(n9778), .ZN(n7184) );
  NAND2_X1 U8704 ( .A1(n7185), .A2(n7184), .ZN(n6926) );
  OAI21_X1 U8705 ( .B1(n10002), .B2(n7193), .A(n6926), .ZN(n6975) );
  NAND2_X1 U8706 ( .A1(n6974), .A2(n6975), .ZN(n6973) );
  OAI21_X1 U8707 ( .B1(n6979), .B2(n6924), .A(n6973), .ZN(n9790) );
  NAND2_X1 U8708 ( .A1(n9791), .A2(n9790), .ZN(n9788) );
  OAI21_X1 U8709 ( .B1(n10005), .B2(n9797), .A(n9788), .ZN(n6988) );
  MUX2_X1 U8710 ( .A(n6013), .B(P1_REG1_REG_5__SCAN_IN), .S(n6986), .Z(n6987)
         );
  XOR2_X1 U8711 ( .A(n6988), .B(n6987), .Z(n6929) );
  INV_X1 U8712 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9575) );
  NOR2_X1 U8713 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9575), .ZN(n6927) );
  AOI21_X1 U8714 ( .B1(n9794), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6927), .ZN(
        n6928) );
  OAI21_X1 U8715 ( .B1(n9242), .B2(n6929), .A(n6928), .ZN(n6941) );
  INV_X1 U8716 ( .A(n9797), .ZN(n6935) );
  INV_X1 U8717 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U8718 ( .A1(n9775), .A2(n6931), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n6930), .ZN(n9772) );
  NAND2_X1 U8719 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9773) );
  NOR2_X1 U8720 ( .A1(n9772), .A2(n9773), .ZN(n9771) );
  AOI21_X1 U8721 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9775), .A(n9771), .ZN(
        n7187) );
  INV_X1 U8722 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U8723 ( .A1(n6932), .A2(n9889), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n7193), .ZN(n7188) );
  NOR2_X1 U8724 ( .A1(n7187), .A2(n7188), .ZN(n7186) );
  NAND2_X1 U8725 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6934), .ZN(n6933) );
  OAI21_X1 U8726 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6934), .A(n6933), .ZN(
        n6971) );
  NOR2_X1 U8727 ( .A1(n6972), .A2(n6971), .ZN(n6970) );
  INV_X1 U8728 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7363) );
  MUX2_X1 U8729 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7363), .S(n9797), .Z(n9786)
         );
  NOR2_X1 U8730 ( .A1(n9787), .A2(n9786), .ZN(n9785) );
  AOI21_X1 U8731 ( .B1(n6935), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9785), .ZN(
        n6939) );
  NAND2_X1 U8732 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6986), .ZN(n6936) );
  OAI21_X1 U8733 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6986), .A(n6936), .ZN(
        n6938) );
  NOR2_X1 U8734 ( .A1(n6939), .A2(n6938), .ZN(n6982) );
  OR2_X1 U8735 ( .A1(n5778), .A2(n5779), .ZN(n6937) );
  OR2_X1 U8736 ( .A1(n9770), .A2(n6937), .ZN(n9784) );
  AOI211_X1 U8737 ( .C1(n6939), .C2(n6938), .A(n6982), .B(n9784), .ZN(n6940)
         );
  AOI211_X1 U8738 ( .C1(n9776), .C2(n6986), .A(n6941), .B(n6940), .ZN(n6942)
         );
  INV_X1 U8739 ( .A(n6942), .ZN(P1_U3248) );
  INV_X1 U8740 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6944) );
  NOR2_X1 U8741 ( .A1(n6943), .A2(n6944), .ZN(P2_U3242) );
  INV_X1 U8742 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6945) );
  NOR2_X1 U8743 ( .A1(n6943), .A2(n6945), .ZN(P2_U3238) );
  INV_X1 U8744 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6946) );
  NOR2_X1 U8745 ( .A1(n6943), .A2(n6946), .ZN(P2_U3244) );
  INV_X1 U8746 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6947) );
  NOR2_X1 U8747 ( .A1(n6943), .A2(n6947), .ZN(P2_U3241) );
  INV_X1 U8748 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6948) );
  NOR2_X1 U8749 ( .A1(n6943), .A2(n6948), .ZN(P2_U3258) );
  INV_X1 U8750 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6949) );
  NOR2_X1 U8751 ( .A1(n6943), .A2(n6949), .ZN(P2_U3239) );
  INV_X1 U8752 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6950) );
  NOR2_X1 U8753 ( .A1(n6943), .A2(n6950), .ZN(P2_U3245) );
  INV_X1 U8754 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6951) );
  NOR2_X1 U8755 ( .A1(n6943), .A2(n6951), .ZN(P2_U3263) );
  INV_X1 U8756 ( .A(n8689), .ZN(n8665) );
  OAI21_X1 U8757 ( .B1(n8665), .B2(n6954), .A(n6953), .ZN(n6955) );
  OAI21_X1 U8758 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6956), .A(n6955), .ZN(n6957) );
  AOI21_X1 U8759 ( .B1(n7394), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6957), .ZN(
        n6958) );
  OAI21_X1 U8760 ( .B1(n6959), .B2(n8686), .A(n6958), .ZN(P2_U3182) );
  INV_X1 U8761 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6960) );
  NOR2_X1 U8762 ( .A1(n6943), .A2(n6960), .ZN(P2_U3261) );
  INV_X1 U8763 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6961) );
  NOR2_X1 U8764 ( .A1(n6943), .A2(n6961), .ZN(P2_U3260) );
  INV_X1 U8765 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6962) );
  NOR2_X1 U8766 ( .A1(n6943), .A2(n6962), .ZN(P2_U3243) );
  INV_X1 U8767 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6963) );
  NOR2_X1 U8768 ( .A1(n6943), .A2(n6963), .ZN(P2_U3234) );
  INV_X1 U8769 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6964) );
  NOR2_X1 U8770 ( .A1(n6943), .A2(n6964), .ZN(P2_U3262) );
  INV_X1 U8771 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6965) );
  NOR2_X1 U8772 ( .A1(n6943), .A2(n6965), .ZN(P2_U3240) );
  INV_X1 U8773 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6966) );
  NOR2_X1 U8774 ( .A1(n6943), .A2(n6966), .ZN(P2_U3237) );
  INV_X1 U8775 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6967) );
  NOR2_X1 U8776 ( .A1(n6943), .A2(n6967), .ZN(P2_U3259) );
  INV_X1 U8777 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6968) );
  NOR2_X1 U8778 ( .A1(n6943), .A2(n6968), .ZN(P2_U3236) );
  INV_X1 U8779 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6969) );
  NOR2_X1 U8780 ( .A1(n6943), .A2(n6969), .ZN(P2_U3235) );
  AOI211_X1 U8781 ( .C1(n6972), .C2(n6971), .A(n6970), .B(n9784), .ZN(n6981)
         );
  INV_X1 U8782 ( .A(n9242), .ZN(n9789) );
  OAI211_X1 U8783 ( .C1(n6975), .C2(n6974), .A(n9789), .B(n6973), .ZN(n6978)
         );
  AND2_X1 U8784 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6976) );
  AOI21_X1 U8785 ( .B1(n9794), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6976), .ZN(
        n6977) );
  OAI211_X1 U8786 ( .C1(n9798), .C2(n6979), .A(n6978), .B(n6977), .ZN(n6980)
         );
  OR2_X1 U8787 ( .A1(n6981), .A2(n6980), .ZN(P1_U3246) );
  INV_X1 U8788 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U8789 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n7005), .B1(n7001), .B2(
        n6983), .ZN(n6984) );
  NOR2_X1 U8790 ( .A1(n6985), .A2(n6984), .ZN(n7000) );
  AOI211_X1 U8791 ( .C1(n6985), .C2(n6984), .A(n7000), .B(n9784), .ZN(n6999)
         );
  NAND2_X1 U8792 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6986), .ZN(n6991) );
  INV_X1 U8793 ( .A(n6987), .ZN(n6989) );
  NAND2_X1 U8794 ( .A1(n6989), .A2(n6988), .ZN(n6990) );
  NAND2_X1 U8795 ( .A1(n6991), .A2(n6990), .ZN(n6994) );
  INV_X1 U8796 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6992) );
  MUX2_X1 U8797 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6992), .S(n7001), .Z(n6993)
         );
  NAND2_X1 U8798 ( .A1(n6993), .A2(n6994), .ZN(n7004) );
  OAI211_X1 U8799 ( .C1(n6994), .C2(n6993), .A(n9789), .B(n7004), .ZN(n6997)
         );
  AND2_X1 U8800 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6995) );
  AOI21_X1 U8801 ( .B1(n9794), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6995), .ZN(
        n6996) );
  OAI211_X1 U8802 ( .C1(n9798), .C2(n7005), .A(n6997), .B(n6996), .ZN(n6998)
         );
  OR2_X1 U8803 ( .A1(n6999), .A2(n6998), .ZN(P1_U3249) );
  AOI21_X1 U8804 ( .B1(n7001), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7000), .ZN(
        n7003) );
  INV_X1 U8805 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9524) );
  AOI22_X1 U8806 ( .A1(n7099), .A2(n9524), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n7012), .ZN(n7002) );
  NOR2_X1 U8807 ( .A1(n7003), .A2(n7002), .ZN(n7095) );
  AOI211_X1 U8808 ( .C1(n7003), .C2(n7002), .A(n7095), .B(n9784), .ZN(n7014)
         );
  OAI21_X1 U8809 ( .B1(n7005), .B2(n6992), .A(n7004), .ZN(n7008) );
  INV_X1 U8810 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7006) );
  MUX2_X1 U8811 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7006), .S(n7099), .Z(n7007)
         );
  NAND2_X1 U8812 ( .A1(n7007), .A2(n7008), .ZN(n7100) );
  OAI211_X1 U8813 ( .C1(n7008), .C2(n7007), .A(n9789), .B(n7100), .ZN(n7011)
         );
  AND2_X1 U8814 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7009) );
  AOI21_X1 U8815 ( .B1(n9794), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7009), .ZN(
        n7010) );
  OAI211_X1 U8816 ( .C1(n9798), .C2(n7012), .A(n7011), .B(n7010), .ZN(n7013)
         );
  OR2_X1 U8817 ( .A1(n7014), .A2(n7013), .ZN(P1_U3250) );
  OAI211_X1 U8818 ( .C1(n7017), .C2(n7016), .A(n8665), .B(n7015), .ZN(n7018)
         );
  OAI21_X1 U8819 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n4920), .A(n7018), .ZN(n7026) );
  INV_X1 U8820 ( .A(n8697), .ZN(n8675) );
  INV_X1 U8821 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7209) );
  AOI21_X1 U8822 ( .B1(n7209), .B2(n4349), .A(n7019), .ZN(n7024) );
  INV_X1 U8823 ( .A(n7020), .ZN(n7021) );
  AOI21_X1 U8824 ( .B1(n7262), .B2(n7022), .A(n7021), .ZN(n7023) );
  OAI22_X1 U8825 ( .A1(n8675), .A2(n7024), .B1(n7023), .B2(n8698), .ZN(n7025)
         );
  AOI211_X1 U8826 ( .C1(n7394), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7026), .B(
        n7025), .ZN(n7027) );
  OAI21_X1 U8827 ( .B1(n7028), .B2(n8686), .A(n7027), .ZN(P2_U3183) );
  INV_X1 U8828 ( .A(n8698), .ZN(n8601) );
  OAI21_X1 U8829 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(n7039) );
  INV_X1 U8830 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7032) );
  NOR2_X1 U8831 ( .A1(n8695), .A2(n7032), .ZN(n7038) );
  AOI21_X1 U8832 ( .B1(n7035), .B2(n7034), .A(n7033), .ZN(n7036) );
  OAI22_X1 U8833 ( .A1(n8675), .A2(n7036), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7331), .ZN(n7037) );
  AOI211_X1 U8834 ( .C1(n8601), .C2(n7039), .A(n7038), .B(n7037), .ZN(n7044)
         );
  OAI211_X1 U8835 ( .C1(n7042), .C2(n7041), .A(n7040), .B(n8665), .ZN(n7043)
         );
  OAI211_X1 U8836 ( .C1(n8686), .C2(n7045), .A(n7044), .B(n7043), .ZN(P2_U3184) );
  INV_X1 U8837 ( .A(n7046), .ZN(n7049) );
  INV_X1 U8838 ( .A(n7603), .ZN(n7595) );
  OAI222_X1 U8839 ( .A1(n8194), .A2(n7047), .B1(n9675), .B2(n7049), .C1(
        P1_U3086), .C2(n7595), .ZN(P1_U3344) );
  OAI222_X1 U8840 ( .A1(n7050), .A2(P2_U3151), .B1(n8056), .B2(n7049), .C1(
        n7048), .C2(n9021), .ZN(P2_U3284) );
  INV_X1 U8841 ( .A(n7051), .ZN(n7053) );
  NAND3_X1 U8842 ( .A1(n7072), .A2(n7053), .A3(n7052), .ZN(n7054) );
  AOI21_X1 U8843 ( .B1(n7055), .B2(n7054), .A(n8698), .ZN(n7062) );
  AND3_X1 U8844 ( .A1(n7078), .A2(n7057), .A3(n7056), .ZN(n7058) );
  OAI21_X1 U8845 ( .B1(n7059), .B2(n7058), .A(n8697), .ZN(n7060) );
  NAND2_X1 U8846 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U8847 ( .A1(n7060), .A2(n7311), .ZN(n7061) );
  AOI211_X1 U8848 ( .C1(n7394), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7062), .B(
        n7061), .ZN(n7067) );
  OAI211_X1 U8849 ( .C1(n7065), .C2(n7064), .A(n7063), .B(n8665), .ZN(n7066)
         );
  OAI211_X1 U8850 ( .C1(n8686), .C2(n7068), .A(n7067), .B(n7066), .ZN(P2_U3186) );
  AOI21_X1 U8851 ( .B1(n7071), .B2(n7070), .A(n7069), .ZN(n7086) );
  INV_X1 U8852 ( .A(n8686), .ZN(n8674) );
  INV_X1 U8853 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7076) );
  INV_X1 U8854 ( .A(n7072), .ZN(n7073) );
  AOI21_X1 U8855 ( .B1(n5530), .B2(n7074), .A(n7073), .ZN(n7075) );
  OAI22_X1 U8856 ( .A1(n8695), .A2(n7076), .B1(n8698), .B2(n7075), .ZN(n7083)
         );
  INV_X1 U8857 ( .A(n7077), .ZN(n7080) );
  INV_X1 U8858 ( .A(n7078), .ZN(n7079) );
  AOI21_X1 U8859 ( .B1(n5529), .B2(n7080), .A(n7079), .ZN(n7081) );
  NAND2_X1 U8860 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7336) );
  OAI21_X1 U8861 ( .B1(n7081), .B2(n8675), .A(n7336), .ZN(n7082) );
  AOI211_X1 U8862 ( .C1(n7084), .C2(n8674), .A(n7083), .B(n7082), .ZN(n7085)
         );
  OAI21_X1 U8863 ( .B1(n7086), .B2(n8689), .A(n7085), .ZN(P2_U3185) );
  INV_X1 U8864 ( .A(n7087), .ZN(n7111) );
  AOI22_X1 U8865 ( .A1(n7620), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9673), .ZN(n7088) );
  OAI21_X1 U8866 ( .B1(n7111), .B2(n9675), .A(n7088), .ZN(P1_U3343) );
  OAI21_X1 U8867 ( .B1(n7091), .B2(n7090), .A(n7089), .ZN(n7179) );
  INV_X1 U8868 ( .A(n9148), .ZN(n9755) );
  NAND2_X1 U8869 ( .A1(n9135), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7214) );
  NAND2_X1 U8870 ( .A1(n7214), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7094) );
  NOR2_X1 U8871 ( .A1(n7092), .A2(n9129), .ZN(n7377) );
  AOI22_X1 U8872 ( .A1(n7135), .A2(n9141), .B1(n7377), .B2(n9753), .ZN(n7093)
         );
  OAI211_X1 U8873 ( .C1(n7179), .C2(n9755), .A(n7094), .B(n7093), .ZN(P1_U3232) );
  NAND2_X1 U8874 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7158), .ZN(n7096) );
  OAI21_X1 U8875 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7158), .A(n7096), .ZN(
        n7097) );
  AOI211_X1 U8876 ( .C1(n7098), .C2(n7097), .A(n7157), .B(n9784), .ZN(n7109)
         );
  NAND2_X1 U8877 ( .A1(n7099), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7101) );
  NAND2_X1 U8878 ( .A1(n7101), .A2(n7100), .ZN(n7104) );
  MUX2_X1 U8879 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7102), .S(n7158), .Z(n7103)
         );
  NAND2_X1 U8880 ( .A1(n7103), .A2(n7104), .ZN(n7153) );
  OAI211_X1 U8881 ( .C1(n7104), .C2(n7103), .A(n9789), .B(n7153), .ZN(n7107)
         );
  INV_X1 U8882 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7105) );
  NOR2_X1 U8883 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7105), .ZN(n7801) );
  AOI21_X1 U8884 ( .B1(n9794), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7801), .ZN(
        n7106) );
  OAI211_X1 U8885 ( .C1(n9798), .C2(n4480), .A(n7107), .B(n7106), .ZN(n7108)
         );
  OR2_X1 U8886 ( .A1(n7109), .A2(n7108), .ZN(P1_U3251) );
  OAI222_X1 U8887 ( .A1(P2_U3151), .A2(n7112), .B1(n8056), .B2(n7111), .C1(
        n7110), .C2(n9021), .ZN(P2_U3283) );
  NAND2_X1 U8888 ( .A1(n7113), .A2(n7114), .ZN(n8395) );
  NAND2_X1 U8889 ( .A1(n8391), .A2(n8395), .ZN(n8335) );
  INV_X1 U8890 ( .A(n8335), .ZN(n7254) );
  INV_X1 U8891 ( .A(n8305), .ZN(n8067) );
  NAND2_X1 U8892 ( .A1(n8067), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7172) );
  NAND2_X1 U8893 ( .A1(n7172), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7116) );
  AOI22_X1 U8894 ( .A1(n8310), .A2(n7257), .B1(n8304), .B2(n8582), .ZN(n7115)
         );
  OAI211_X1 U8895 ( .C1(n7254), .C2(n8312), .A(n7116), .B(n7115), .ZN(P2_U3172) );
  AOI21_X1 U8896 ( .B1(n4986), .B2(n7117), .A(n7230), .ZN(n7119) );
  OAI22_X1 U8897 ( .A1(n7119), .A2(n8675), .B1(n7118), .B2(n8686), .ZN(n7128)
         );
  NAND2_X1 U8898 ( .A1(n7120), .A2(n7452), .ZN(n7121) );
  AOI21_X1 U8899 ( .B1(n7122), .B2(n7121), .A(n8698), .ZN(n7127) );
  INV_X1 U8900 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7125) );
  NOR2_X1 U8901 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7123), .ZN(n7414) );
  INV_X1 U8902 ( .A(n7414), .ZN(n7124) );
  OAI21_X1 U8903 ( .B1(n8695), .B2(n7125), .A(n7124), .ZN(n7126) );
  NOR3_X1 U8904 ( .A1(n7128), .A2(n7127), .A3(n7126), .ZN(n7133) );
  OAI211_X1 U8905 ( .C1(n7131), .C2(n7130), .A(n7129), .B(n8665), .ZN(n7132)
         );
  NAND2_X1 U8906 ( .A1(n7133), .A2(n7132), .ZN(P2_U3187) );
  INV_X1 U8907 ( .A(n9868), .ZN(n9895) );
  AOI21_X1 U8908 ( .B1(n9941), .B2(n9895), .A(n7380), .ZN(n7134) );
  AOI211_X1 U8909 ( .C1(n7136), .C2(n7135), .A(n7377), .B(n7134), .ZN(n7175)
         );
  NAND2_X1 U8910 ( .A1(n10013), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7137) );
  OAI21_X1 U8911 ( .B1(n7175), .B2(n10013), .A(n7137), .ZN(P1_U3522) );
  INV_X1 U8912 ( .A(n7138), .ZN(n7140) );
  INV_X1 U8913 ( .A(n7707), .ZN(n7714) );
  OAI222_X1 U8914 ( .A1(n8194), .A2(n7139), .B1(n9675), .B2(n7140), .C1(
        P1_U3086), .C2(n7714), .ZN(P1_U3342) );
  OAI222_X1 U8915 ( .A1(n7141), .A2(P2_U3151), .B1(n8056), .B2(n7140), .C1(
        n9523), .C2(n9021), .ZN(P2_U3282) );
  XOR2_X1 U8916 ( .A(n7143), .B(n7142), .Z(n7146) );
  AOI22_X1 U8917 ( .A1(n9131), .A2(n6275), .B1(n9176), .B2(n9086), .ZN(n9894)
         );
  OAI22_X1 U8918 ( .A1(n9894), .A2(n9090), .B1(n9749), .B2(n6701), .ZN(n7144)
         );
  AOI21_X1 U8919 ( .B1(n7214), .B2(P1_REG3_REG_1__SCAN_IN), .A(n7144), .ZN(
        n7145) );
  OAI21_X1 U8920 ( .B1(n7146), .B2(n9755), .A(n7145), .ZN(P1_U3222) );
  XOR2_X1 U8921 ( .A(n7148), .B(n7147), .Z(n7152) );
  INV_X1 U8922 ( .A(n8310), .ZN(n8299) );
  INV_X1 U8923 ( .A(n8308), .ZN(n8293) );
  AOI22_X1 U8924 ( .A1(n8293), .A2(n8582), .B1(n8304), .B2(n8580), .ZN(n7149)
         );
  OAI21_X1 U8925 ( .B1(n8299), .B2(n8402), .A(n7149), .ZN(n7150) );
  AOI21_X1 U8926 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7172), .A(n7150), .ZN(
        n7151) );
  OAI21_X1 U8927 ( .B1(n7152), .B2(n8312), .A(n7151), .ZN(P2_U3177) );
  AOI22_X1 U8928 ( .A1(n7291), .A2(n6041), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n7162), .ZN(n7156) );
  NAND2_X1 U8929 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7158), .ZN(n7154) );
  NAND2_X1 U8930 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  NOR2_X1 U8931 ( .A1(n7156), .A2(n7155), .ZN(n7292) );
  AOI21_X1 U8932 ( .B1(n7156), .B2(n7155), .A(n7292), .ZN(n7166) );
  AOI22_X1 U8933 ( .A1(n7291), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6042), .B2(
        n7162), .ZN(n7160) );
  OAI21_X1 U8934 ( .B1(n7160), .B2(n7159), .A(n7288), .ZN(n7161) );
  INV_X1 U8935 ( .A(n9784), .ZN(n9214) );
  NAND2_X1 U8936 ( .A1(n7161), .A2(n9214), .ZN(n7165) );
  AND2_X1 U8937 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7861) );
  NOR2_X1 U8938 ( .A1(n9798), .A2(n7162), .ZN(n7163) );
  AOI211_X1 U8939 ( .C1(n9794), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7861), .B(
        n7163), .ZN(n7164) );
  OAI211_X1 U8940 ( .C1(n7166), .C2(n9242), .A(n7165), .B(n7164), .ZN(P1_U3252) );
  XOR2_X1 U8941 ( .A(n7168), .B(n7167), .Z(n7174) );
  AOI22_X1 U8942 ( .A1(n8293), .A2(n7113), .B1(n8304), .B2(n8581), .ZN(n7169)
         );
  OAI21_X1 U8943 ( .B1(n8299), .B2(n7170), .A(n7169), .ZN(n7171) );
  AOI21_X1 U8944 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7172), .A(n7171), .ZN(
        n7173) );
  OAI21_X1 U8945 ( .B1(n7174), .B2(n8312), .A(n7173), .ZN(P2_U3162) );
  INV_X1 U8946 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7177) );
  OR2_X1 U8947 ( .A1(n7175), .A2(n9998), .ZN(n7176) );
  OAI21_X1 U8948 ( .B1(n10000), .B2(n7177), .A(n7176), .ZN(P1_U3453) );
  INV_X1 U8949 ( .A(n9773), .ZN(n7178) );
  MUX2_X1 U8950 ( .A(n7179), .B(n7178), .S(n9761), .Z(n7183) );
  NOR2_X1 U8951 ( .A1(n5779), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7180) );
  OR2_X1 U8952 ( .A1(n7180), .A2(n5778), .ZN(n9762) );
  NAND2_X1 U8953 ( .A1(n9762), .A2(n5599), .ZN(n9766) );
  NAND2_X1 U8954 ( .A1(n9766), .A2(P1_U3973), .ZN(n7181) );
  AOI21_X1 U8955 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(n9801) );
  XOR2_X1 U8956 ( .A(n7185), .B(n7184), .Z(n7190) );
  AOI211_X1 U8957 ( .C1(n7188), .C2(n7187), .A(n7186), .B(n9784), .ZN(n7189)
         );
  AOI21_X1 U8958 ( .B1(n9789), .B2(n7190), .A(n7189), .ZN(n7192) );
  AOI22_X1 U8959 ( .A1(n9794), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7191) );
  OAI211_X1 U8960 ( .C1(n7193), .C2(n9798), .A(n7192), .B(n7191), .ZN(n7194)
         );
  OR2_X1 U8961 ( .A1(n9801), .A2(n7194), .ZN(P1_U3245) );
  INV_X1 U8962 ( .A(n7195), .ZN(n7198) );
  OAI222_X1 U8963 ( .A1(n7197), .A2(P2_U3151), .B1(n8056), .B2(n7198), .C1(
        n7196), .C2(n9021), .ZN(P2_U3281) );
  INV_X1 U8964 ( .A(n7980), .ZN(n7983) );
  OAI222_X1 U8965 ( .A1(n8195), .A2(n7199), .B1(n9675), .B2(n7198), .C1(
        P1_U3086), .C2(n7983), .ZN(P1_U3341) );
  XNOR2_X1 U8966 ( .A(n7200), .B(n7201), .ZN(n7202) );
  NAND2_X1 U8967 ( .A1(n7202), .A2(n8928), .ZN(n7204) );
  INV_X1 U8968 ( .A(n8865), .ZN(n8934) );
  AOI22_X1 U8969 ( .A1(n8934), .A2(n7113), .B1(n8581), .B2(n8932), .ZN(n7203)
         );
  AND2_X1 U8970 ( .A1(n7204), .A2(n7203), .ZN(n7263) );
  NAND2_X1 U8971 ( .A1(n7200), .A2(n8391), .ZN(n7205) );
  NAND2_X1 U8972 ( .A1(n7206), .A2(n7205), .ZN(n7261) );
  INV_X1 U8973 ( .A(n7950), .ZN(n7278) );
  AOI22_X1 U8974 ( .A1(n7261), .A2(n7278), .B1(n8915), .B2(n7264), .ZN(n7208)
         );
  INV_X1 U8975 ( .A(n7848), .ZN(n7275) );
  NAND2_X1 U8976 ( .A1(n7261), .A2(n7275), .ZN(n7207) );
  AND3_X1 U8977 ( .A1(n7263), .A2(n7208), .A3(n7207), .ZN(n10037) );
  MUX2_X1 U8978 ( .A(n7209), .B(n10037), .S(n8942), .Z(n7210) );
  INV_X1 U8979 ( .A(n7210), .ZN(P2_U3460) );
  XOR2_X1 U8980 ( .A(n7211), .B(n7212), .Z(n7216) );
  AOI22_X1 U8981 ( .A1(n9175), .A2(n9086), .B1(n9131), .B2(n6268), .ZN(n9883)
         );
  OAI22_X1 U8982 ( .A1(n9883), .A2(n9090), .B1(n9924), .B2(n9749), .ZN(n7213)
         );
  AOI21_X1 U8983 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7214), .A(n7213), .ZN(
        n7215) );
  OAI21_X1 U8984 ( .B1(n7216), .B2(n9755), .A(n7215), .ZN(P1_U3237) );
  AOI21_X1 U8985 ( .B1(n7219), .B2(n7218), .A(n7217), .ZN(n7237) );
  INV_X1 U8986 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U8987 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7571) );
  OAI21_X1 U8988 ( .B1(n8695), .B2(n7220), .A(n7571), .ZN(n7227) );
  OR3_X1 U8989 ( .A1(n7223), .A2(n7222), .A3(n7221), .ZN(n7224) );
  AOI21_X1 U8990 ( .B1(n7225), .B2(n7224), .A(n8698), .ZN(n7226) );
  AOI211_X1 U8991 ( .C1(n8674), .C2(n7228), .A(n7227), .B(n7226), .ZN(n7236)
         );
  INV_X1 U8992 ( .A(n7229), .ZN(n7234) );
  NOR3_X1 U8993 ( .A1(n7232), .A2(n7231), .A3(n7230), .ZN(n7233) );
  OAI21_X1 U8994 ( .B1(n7234), .B2(n7233), .A(n8697), .ZN(n7235) );
  OAI211_X1 U8995 ( .C1(n7237), .C2(n8689), .A(n7236), .B(n7235), .ZN(P2_U3188) );
  INV_X1 U8996 ( .A(n7238), .ZN(n7244) );
  OR2_X1 U8997 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  NAND4_X1 U8998 ( .A1(n7244), .A2(n7243), .A3(n7242), .A4(n7241), .ZN(n7245)
         );
  OR2_X1 U8999 ( .A1(n7245), .A2(n9738), .ZN(n10020) );
  INV_X1 U9000 ( .A(n10017), .ZN(n10028) );
  AOI22_X1 U9001 ( .A1(n10026), .A2(n7257), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10028), .ZN(n7249) );
  NOR2_X1 U9002 ( .A1(n7254), .A2(n7246), .ZN(n7247) );
  NOR2_X1 U9003 ( .A1(n7272), .A2(n8867), .ZN(n7256) );
  OAI21_X1 U9004 ( .B1(n7247), .B2(n7256), .A(n4275), .ZN(n7248) );
  OAI211_X1 U9005 ( .C1(n4933), .C2(n4275), .A(n7249), .B(n7248), .ZN(P2_U3233) );
  NAND2_X1 U9006 ( .A1(n9177), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7250) );
  OAI21_X1 U9007 ( .B1(n7251), .B2(n9177), .A(n7250), .ZN(P1_U3582) );
  INV_X1 U9008 ( .A(n7252), .ZN(n7260) );
  INV_X1 U9009 ( .A(n9182), .ZN(n9187) );
  INV_X1 U9010 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7253) );
  OAI222_X1 U9011 ( .A1(n9675), .A2(n7260), .B1(n9187), .B2(P1_U3086), .C1(
        n7253), .C2(n8195), .ZN(P1_U3340) );
  AOI21_X1 U9012 ( .B1(n8940), .B2(n8862), .A(n7254), .ZN(n7255) );
  AOI211_X1 U9013 ( .C1(n8915), .C2(n7257), .A(n7256), .B(n7255), .ZN(n10035)
         );
  OR2_X1 U9014 ( .A1(n10035), .A2(n8944), .ZN(n7258) );
  OAI21_X1 U9015 ( .B1(n8942), .B2(n5477), .A(n7258), .ZN(P2_U3459) );
  INV_X1 U9016 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7259) );
  OAI222_X1 U9017 ( .A1(P2_U3151), .A2(n5505), .B1(n8056), .B2(n7260), .C1(
        n7259), .C2(n9021), .ZN(P2_U3280) );
  INV_X1 U9018 ( .A(n7261), .ZN(n7267) );
  OR2_X1 U9019 ( .A1(n5819), .A2(n8390), .ZN(n7326) );
  NAND2_X1 U9020 ( .A1(n7848), .A2(n7326), .ZN(n9735) );
  NAND2_X1 U9021 ( .A1(n4275), .A2(n9735), .ZN(n10025) );
  MUX2_X1 U9022 ( .A(n7263), .B(n7262), .S(n10034), .Z(n7266) );
  AOI22_X1 U9023 ( .A1(n10026), .A2(n7264), .B1(n10028), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7265) );
  OAI211_X1 U9024 ( .C1(n7267), .C2(n10025), .A(n7266), .B(n7265), .ZN(
        P2_U3232) );
  XNOR2_X1 U9025 ( .A(n7268), .B(n8399), .ZN(n7327) );
  AND2_X1 U9026 ( .A1(n7269), .A2(n8915), .ZN(n7328) );
  XNOR2_X1 U9027 ( .A(n7270), .B(n8399), .ZN(n7274) );
  OAI22_X1 U9028 ( .A1(n7272), .A2(n8865), .B1(n7271), .B2(n8867), .ZN(n7273)
         );
  AOI21_X1 U9029 ( .B1(n7274), .B2(n8928), .A(n7273), .ZN(n7277) );
  NAND2_X1 U9030 ( .A1(n7327), .A2(n7275), .ZN(n7276) );
  NAND2_X1 U9031 ( .A1(n7277), .A2(n7276), .ZN(n7333) );
  AOI211_X1 U9032 ( .C1(n7278), .C2(n7327), .A(n7328), .B(n7333), .ZN(n10038)
         );
  NAND2_X1 U9033 ( .A1(n8944), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7279) );
  OAI21_X1 U9034 ( .B1(n10038), .B2(n8944), .A(n7279), .ZN(P2_U3461) );
  XOR2_X1 U9035 ( .A(n7281), .B(n7280), .Z(n7286) );
  OAI22_X1 U9036 ( .A1(n7283), .A2(n9129), .B1(n7282), .B2(n9117), .ZN(n9867)
         );
  AOI22_X1 U9037 ( .A1(n9867), .A2(n9753), .B1(n9141), .B2(n9870), .ZN(n7285)
         );
  MUX2_X1 U9038 ( .A(n9135), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7284) );
  OAI211_X1 U9039 ( .C1(n7286), .C2(n9755), .A(n7285), .B(n7284), .ZN(P1_U3218) );
  NAND2_X1 U9040 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7429), .ZN(n7287) );
  OAI21_X1 U9041 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7429), .A(n7287), .ZN(
        n7290) );
  OAI21_X1 U9042 ( .B1(n7291), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7288), .ZN(
        n7289) );
  NOR2_X1 U9043 ( .A1(n7290), .A2(n7289), .ZN(n7428) );
  AOI211_X1 U9044 ( .C1(n7290), .C2(n7289), .A(n7428), .B(n9784), .ZN(n7300)
         );
  NOR2_X1 U9045 ( .A1(n7291), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7293) );
  NOR2_X1 U9046 ( .A1(n7293), .A2(n7292), .ZN(n7296) );
  MUX2_X1 U9047 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7294), .S(n7429), .Z(n7295)
         );
  NAND2_X1 U9048 ( .A1(n7295), .A2(n7296), .ZN(n7433) );
  OAI211_X1 U9049 ( .C1(n7296), .C2(n7295), .A(n7433), .B(n9789), .ZN(n7298)
         );
  NOR2_X1 U9050 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6047), .ZN(n9751) );
  AOI21_X1 U9051 ( .B1(n9794), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9751), .ZN(
        n7297) );
  OAI211_X1 U9052 ( .C1(n9798), .C2(n7434), .A(n7298), .B(n7297), .ZN(n7299)
         );
  OR2_X1 U9053 ( .A1(n7300), .A2(n7299), .ZN(P1_U3253) );
  INV_X1 U9054 ( .A(n7301), .ZN(n7304) );
  OAI222_X1 U9055 ( .A1(n7303), .A2(P2_U3151), .B1(n8056), .B2(n7304), .C1(
        n7302), .C2(n9021), .ZN(P2_U3279) );
  INV_X1 U9056 ( .A(n9196), .ZN(n9204) );
  OAI222_X1 U9057 ( .A1(n8195), .A2(n7305), .B1(n9675), .B2(n7304), .C1(
        P1_U3086), .C2(n9204), .ZN(P1_U3339) );
  INV_X1 U9058 ( .A(n7306), .ZN(n7307) );
  AOI21_X1 U9059 ( .B1(n7309), .B2(n7308), .A(n7307), .ZN(n7317) );
  INV_X1 U9060 ( .A(n7310), .ZN(n10029) );
  INV_X1 U9061 ( .A(n7311), .ZN(n7312) );
  AOI21_X1 U9062 ( .B1(n8293), .B2(n8580), .A(n7312), .ZN(n7314) );
  NAND2_X1 U9063 ( .A1(n8310), .A2(n10027), .ZN(n7313) );
  OAI211_X1 U9064 ( .C1(n7549), .C2(n8295), .A(n7314), .B(n7313), .ZN(n7315)
         );
  AOI21_X1 U9065 ( .B1(n10029), .B2(n8305), .A(n7315), .ZN(n7316) );
  OAI21_X1 U9066 ( .B1(n7317), .B2(n8312), .A(n7316), .ZN(P2_U3170) );
  OAI21_X1 U9067 ( .B1(n7319), .B2(n8337), .A(n7318), .ZN(n7374) );
  NOR2_X1 U9068 ( .A1(n7320), .A2(n8939), .ZN(n7324) );
  XNOR2_X1 U9069 ( .A(n7321), .B(n8337), .ZN(n7322) );
  OAI222_X1 U9070 ( .A1(n8867), .A2(n8410), .B1(n8865), .B2(n7323), .C1(n8862), 
        .C2(n7322), .ZN(n7369) );
  AOI211_X1 U9071 ( .C1(n8905), .C2(n7374), .A(n7324), .B(n7369), .ZN(n10039)
         );
  OR2_X1 U9072 ( .A1(n10039), .A2(n8944), .ZN(n7325) );
  OAI21_X1 U9073 ( .B1(n8942), .B2(n5529), .A(n7325), .ZN(P2_U3462) );
  INV_X1 U9074 ( .A(n7326), .ZN(n7533) );
  NAND2_X1 U9075 ( .A1(n7327), .A2(n7533), .ZN(n7330) );
  NAND2_X1 U9076 ( .A1(n7328), .A2(n5819), .ZN(n7329) );
  OAI211_X1 U9077 ( .C1(n10017), .C2(n7331), .A(n7330), .B(n7329), .ZN(n7332)
         );
  NOR2_X1 U9078 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  MUX2_X1 U9079 ( .A(n9594), .B(n7334), .S(n4275), .Z(n7335) );
  INV_X1 U9080 ( .A(n7335), .ZN(P2_U3231) );
  INV_X1 U9081 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7370) );
  INV_X1 U9082 ( .A(n7336), .ZN(n7337) );
  AOI21_X1 U9083 ( .B1(n8293), .B2(n8581), .A(n7337), .ZN(n7339) );
  NAND2_X1 U9084 ( .A1(n8310), .A2(n7371), .ZN(n7338) );
  OAI211_X1 U9085 ( .C1(n8410), .C2(n8295), .A(n7339), .B(n7338), .ZN(n7345)
         );
  INV_X1 U9086 ( .A(n7340), .ZN(n7341) );
  AOI211_X1 U9087 ( .C1(n7343), .C2(n7342), .A(n8312), .B(n7341), .ZN(n7344)
         );
  AOI211_X1 U9088 ( .C1(n7370), .C2(n8305), .A(n7345), .B(n7344), .ZN(n7346)
         );
  INV_X1 U9089 ( .A(n7346), .ZN(P2_U3158) );
  NAND2_X1 U9090 ( .A1(n7347), .A2(n6007), .ZN(n7350) );
  NAND2_X1 U9091 ( .A1(n7350), .A2(n7349), .ZN(n7351) );
  XOR2_X1 U9092 ( .A(n7359), .B(n7351), .Z(n9940) );
  INV_X1 U9093 ( .A(n7352), .ZN(n9973) );
  INV_X1 U9094 ( .A(n7353), .ZN(n9812) );
  INV_X1 U9095 ( .A(n7354), .ZN(n7355) );
  NAND3_X1 U9096 ( .A1(n7357), .A2(n7356), .A3(n7355), .ZN(n7358) );
  OAI21_X2 U9097 ( .B1(n9973), .B2(n9812), .A(n9836), .ZN(n9412) );
  XNOR2_X1 U9098 ( .A(n7360), .B(n7359), .ZN(n7362) );
  OAI22_X1 U9099 ( .A1(n7361), .A2(n9129), .B1(n6297), .B2(n9117), .ZN(n7483)
         );
  AOI21_X1 U9100 ( .B1(n7362), .B2(n9868), .A(n7483), .ZN(n9938) );
  INV_X2 U9101 ( .A(n9836), .ZN(n9898) );
  MUX2_X1 U9102 ( .A(n9938), .B(n7363), .S(n9898), .Z(n7368) );
  AOI211_X1 U9103 ( .C1(n9937), .C2(n9872), .A(n9425), .B(n9863), .ZN(n9936)
         );
  NAND2_X1 U9104 ( .A1(n9836), .A2(n8189), .ZN(n9831) );
  INV_X2 U9105 ( .A(n9831), .ZN(n9905) );
  NAND2_X1 U9106 ( .A1(n9836), .A2(n7364), .ZN(n9427) );
  INV_X1 U9107 ( .A(n7492), .ZN(n7365) );
  OAI22_X1 U9108 ( .A1(n9427), .A2(n7485), .B1(n7365), .B2(n9878), .ZN(n7366)
         );
  AOI21_X1 U9109 ( .B1(n9936), .B2(n9905), .A(n7366), .ZN(n7367) );
  OAI211_X1 U9110 ( .C1(n9940), .C2(n9412), .A(n7368), .B(n7367), .ZN(P1_U3289) );
  INV_X1 U9111 ( .A(n7369), .ZN(n7376) );
  INV_X1 U9112 ( .A(n10025), .ZN(n10030) );
  AOI22_X1 U9113 ( .A1(n10026), .A2(n7371), .B1(n10028), .B2(n7370), .ZN(n7372) );
  OAI21_X1 U9114 ( .B1(n5530), .B2(n4275), .A(n7372), .ZN(n7373) );
  AOI21_X1 U9115 ( .B1(n7374), .B2(n10030), .A(n7373), .ZN(n7375) );
  OAI21_X1 U9116 ( .B1(n7376), .B2(n10034), .A(n7375), .ZN(P2_U3230) );
  INV_X1 U9117 ( .A(n9427), .ZN(n9906) );
  AOI21_X1 U9118 ( .B1(n9905), .B2(n9901), .A(n9906), .ZN(n7386) );
  INV_X1 U9119 ( .A(n7377), .ZN(n7378) );
  OAI21_X1 U9120 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7384) );
  INV_X1 U9121 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7382) );
  INV_X1 U9122 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7381) );
  OAI22_X1 U9123 ( .A1(n9836), .A2(n7382), .B1(n7381), .B2(n9878), .ZN(n7383)
         );
  AOI21_X1 U9124 ( .B1(n7384), .B2(n9836), .A(n7383), .ZN(n7385) );
  OAI21_X1 U9125 ( .B1(n7386), .B2(n9902), .A(n7385), .ZN(P1_U3293) );
  XNOR2_X1 U9126 ( .A(n7388), .B(n7387), .ZN(n7401) );
  INV_X1 U9127 ( .A(n7389), .ZN(n8600) );
  AOI21_X1 U9128 ( .B1(n7536), .B2(n7390), .A(n8600), .ZN(n7396) );
  INV_X1 U9129 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7391) );
  NOR2_X1 U9130 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7391), .ZN(n7514) );
  NOR2_X1 U9131 ( .A1(n8686), .A2(n7392), .ZN(n7393) );
  AOI211_X1 U9132 ( .C1(n7394), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7514), .B(
        n7393), .ZN(n7395) );
  OAI21_X1 U9133 ( .B1(n7396), .B2(n8698), .A(n7395), .ZN(n7400) );
  NAND2_X1 U9134 ( .A1(n7397), .A2(n4913), .ZN(n7398) );
  AOI21_X1 U9135 ( .B1(n8594), .B2(n7398), .A(n8675), .ZN(n7399) );
  AOI211_X1 U9136 ( .C1(n8665), .C2(n7401), .A(n7400), .B(n7399), .ZN(n7402)
         );
  INV_X1 U9137 ( .A(n7402), .ZN(P2_U3189) );
  INV_X1 U9138 ( .A(n7403), .ZN(n7406) );
  OAI222_X1 U9139 ( .A1(n7405), .A2(P2_U3151), .B1(n8056), .B2(n7406), .C1(
        n7404), .C2(n9021), .ZN(P2_U3278) );
  INV_X1 U9140 ( .A(n9222), .ZN(n9211) );
  OAI222_X1 U9141 ( .A1(n8195), .A2(n7407), .B1(n9675), .B2(n7406), .C1(
        P1_U3086), .C2(n9211), .ZN(P1_U3338) );
  NAND2_X1 U9142 ( .A1(n8687), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7408) );
  OAI21_X1 U9143 ( .B1(n8744), .B2(n8687), .A(n7408), .ZN(P2_U3516) );
  INV_X1 U9144 ( .A(n7409), .ZN(n7444) );
  AOI22_X1 U9145 ( .A1(n9235), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9673), .ZN(n7410) );
  OAI21_X1 U9146 ( .B1(n7444), .B2(n9675), .A(n7410), .ZN(P1_U3337) );
  XOR2_X1 U9147 ( .A(n7412), .B(n7411), .Z(n7420) );
  INV_X1 U9148 ( .A(n7413), .ZN(n7453) );
  AOI21_X1 U9149 ( .B1(n8293), .B2(n8579), .A(n7414), .ZN(n7416) );
  NAND2_X1 U9150 ( .A1(n8310), .A2(n7454), .ZN(n7415) );
  OAI211_X1 U9151 ( .C1(n7417), .C2(n8295), .A(n7416), .B(n7415), .ZN(n7418)
         );
  AOI21_X1 U9152 ( .B1(n7453), .B2(n8305), .A(n7418), .ZN(n7419) );
  OAI21_X1 U9153 ( .B1(n7420), .B2(n8312), .A(n7419), .ZN(P2_U3167) );
  XNOR2_X1 U9154 ( .A(n7421), .B(n8339), .ZN(n10031) );
  XNOR2_X1 U9155 ( .A(n7422), .B(n8339), .ZN(n7423) );
  AOI222_X1 U9156 ( .A1(n8928), .A2(n7423), .B1(n8578), .B2(n8932), .C1(n8580), 
        .C2(n8934), .ZN(n10033) );
  OAI21_X1 U9157 ( .B1(n7424), .B2(n8939), .A(n10033), .ZN(n7425) );
  AOI21_X1 U9158 ( .B1(n8905), .B2(n10031), .A(n7425), .ZN(n10041) );
  INV_X1 U9159 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7426) );
  OR2_X1 U9160 ( .A1(n8942), .A2(n7426), .ZN(n7427) );
  OAI21_X1 U9161 ( .B1(n10041), .B2(n8944), .A(n7427), .ZN(P2_U3463) );
  NAND2_X1 U9162 ( .A1(n7603), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7430) );
  OAI21_X1 U9163 ( .B1(n7603), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7430), .ZN(
        n7431) );
  AOI211_X1 U9164 ( .C1(n7432), .C2(n7431), .A(n7602), .B(n9784), .ZN(n7443)
         );
  OAI21_X1 U9165 ( .B1(n7434), .B2(n7294), .A(n7433), .ZN(n7437) );
  MUX2_X1 U9166 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7435), .S(n7603), .Z(n7436)
         );
  NAND2_X1 U9167 ( .A1(n7436), .A2(n7437), .ZN(n7594) );
  OAI211_X1 U9168 ( .C1(n7437), .C2(n7436), .A(n9789), .B(n7594), .ZN(n7441)
         );
  NOR2_X1 U9169 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7438), .ZN(n7439) );
  AOI21_X1 U9170 ( .B1(n9794), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7439), .ZN(
        n7440) );
  OAI211_X1 U9171 ( .C1(n9798), .C2(n7595), .A(n7441), .B(n7440), .ZN(n7442)
         );
  OR2_X1 U9172 ( .A1(n7443), .A2(n7442), .ZN(P1_U3254) );
  INV_X1 U9173 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7445) );
  OAI222_X1 U9174 ( .A1(n9021), .A2(n7445), .B1(n8056), .B2(n7444), .C1(
        P2_U3151), .C2(n8691), .ZN(P2_U3277) );
  INV_X1 U9175 ( .A(n7447), .ZN(n7449) );
  OR2_X1 U9176 ( .A1(n7449), .A2(n7448), .ZN(n8336) );
  XNOR2_X1 U9177 ( .A(n7446), .B(n8336), .ZN(n7497) );
  INV_X1 U9178 ( .A(n7497), .ZN(n7457) );
  XOR2_X1 U9179 ( .A(n8336), .B(n7450), .Z(n7451) );
  AOI222_X1 U9180 ( .A1(n8928), .A2(n7451), .B1(n8577), .B2(n8932), .C1(n8579), 
        .C2(n8934), .ZN(n7494) );
  MUX2_X1 U9181 ( .A(n7452), .B(n7494), .S(n4275), .Z(n7456) );
  AOI22_X1 U9182 ( .A1(n10026), .A2(n7454), .B1(n10028), .B2(n7453), .ZN(n7455) );
  OAI211_X1 U9183 ( .C1(n7457), .C2(n10025), .A(n7456), .B(n7455), .ZN(
        P2_U3228) );
  INV_X1 U9184 ( .A(n7458), .ZN(n7465) );
  INV_X1 U9185 ( .A(n7460), .ZN(n7462) );
  NAND2_X1 U9186 ( .A1(n7462), .A2(n7461), .ZN(n7464) );
  AOI22_X1 U9187 ( .A1(n7465), .A2(n7459), .B1(n7464), .B2(n7463), .ZN(n7469)
         );
  AOI22_X1 U9188 ( .A1(n9131), .A2(n9174), .B1(n9172), .B2(n9086), .ZN(n9854)
         );
  OAI22_X1 U9189 ( .A1(n9854), .A2(n9090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9575), .ZN(n7467) );
  NOR2_X1 U9190 ( .A1(n9760), .A2(n9857), .ZN(n7466) );
  AOI211_X1 U9191 ( .C1(n9859), .C2(n9141), .A(n7467), .B(n7466), .ZN(n7468)
         );
  OAI21_X1 U9192 ( .B1(n7469), .B2(n9755), .A(n7468), .ZN(P1_U3227) );
  XNOR2_X1 U9193 ( .A(n7470), .B(n7474), .ZN(n7471) );
  NAND2_X1 U9194 ( .A1(n7471), .A2(n9868), .ZN(n7472) );
  AOI22_X1 U9195 ( .A1(n9173), .A2(n9131), .B1(n9086), .B2(n9171), .ZN(n7505)
         );
  NAND2_X1 U9196 ( .A1(n7472), .A2(n7505), .ZN(n9956) );
  INV_X1 U9197 ( .A(n9956), .ZN(n7482) );
  XNOR2_X1 U9198 ( .A(n7473), .B(n7474), .ZN(n9951) );
  INV_X1 U9199 ( .A(n9412), .ZN(n9874) );
  AOI21_X1 U9200 ( .B1(n9862), .B2(n7477), .A(n9425), .ZN(n7476) );
  NAND2_X1 U9201 ( .A1(n7476), .A2(n7475), .ZN(n9952) );
  INV_X1 U9202 ( .A(n9878), .ZN(n9899) );
  AOI22_X1 U9203 ( .A1(n9898), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7508), .B2(
        n9899), .ZN(n7479) );
  NAND2_X1 U9204 ( .A1(n9906), .A2(n7477), .ZN(n7478) );
  OAI211_X1 U9205 ( .C1(n9952), .C2(n9831), .A(n7479), .B(n7478), .ZN(n7480)
         );
  AOI21_X1 U9206 ( .B1(n9951), .B2(n9874), .A(n7480), .ZN(n7481) );
  OAI21_X1 U9207 ( .B1(n7482), .B2(n9898), .A(n7481), .ZN(P1_U3287) );
  NAND2_X1 U9208 ( .A1(n7483), .A2(n9753), .ZN(n7484) );
  NAND2_X1 U9209 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9792) );
  OAI211_X1 U9210 ( .C1(n7485), .C2(n9749), .A(n7484), .B(n9792), .ZN(n7491)
         );
  INV_X1 U9211 ( .A(n7487), .ZN(n7488) );
  AOI211_X1 U9212 ( .C1(n7489), .C2(n7486), .A(n9755), .B(n7488), .ZN(n7490)
         );
  AOI211_X1 U9213 ( .C1(n7492), .C2(n9097), .A(n7491), .B(n7490), .ZN(n7493)
         );
  INV_X1 U9214 ( .A(n7493), .ZN(P1_U3230) );
  OAI21_X1 U9215 ( .B1(n7495), .B2(n8939), .A(n7494), .ZN(n7496) );
  AOI21_X1 U9216 ( .B1(n8905), .B2(n7497), .A(n7496), .ZN(n10043) );
  OR2_X1 U9217 ( .A1(n8942), .A2(n4986), .ZN(n7498) );
  OAI21_X1 U9218 ( .B1(n10043), .B2(n8944), .A(n7498), .ZN(P2_U3464) );
  INV_X1 U9219 ( .A(n7499), .ZN(n8190) );
  OAI222_X1 U9220 ( .A1(P2_U3151), .A2(n8373), .B1(n8056), .B2(n8190), .C1(
        n7500), .C2(n9021), .ZN(P2_U3276) );
  INV_X1 U9221 ( .A(n7501), .ZN(n7502) );
  AOI21_X1 U9222 ( .B1(n7503), .B2(n7458), .A(n7502), .ZN(n7510) );
  NOR2_X1 U9223 ( .A1(n9749), .A2(n9953), .ZN(n7507) );
  INV_X1 U9224 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7504) );
  OAI22_X1 U9225 ( .A1(n7505), .A2(n9090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7504), .ZN(n7506) );
  AOI211_X1 U9226 ( .C1(n7508), .C2(n9097), .A(n7507), .B(n7506), .ZN(n7509)
         );
  OAI21_X1 U9227 ( .B1(n7510), .B2(n9755), .A(n7509), .ZN(P1_U3239) );
  OAI21_X1 U9228 ( .B1(n7512), .B2(n4346), .A(n7511), .ZN(n7520) );
  NOR2_X1 U9229 ( .A1(n8299), .A2(n7530), .ZN(n7519) );
  INV_X1 U9230 ( .A(n7535), .ZN(n7513) );
  NAND2_X1 U9231 ( .A1(n8305), .A2(n7513), .ZN(n7516) );
  AOI21_X1 U9232 ( .B1(n8293), .B2(n8577), .A(n7514), .ZN(n7515) );
  OAI211_X1 U9233 ( .C1(n7517), .C2(n8295), .A(n7516), .B(n7515), .ZN(n7518)
         );
  AOI211_X1 U9234 ( .C1(n7520), .C2(n5916), .A(n7519), .B(n7518), .ZN(n7521)
         );
  INV_X1 U9235 ( .A(n7521), .ZN(P2_U3153) );
  INV_X1 U9236 ( .A(n7522), .ZN(n7543) );
  OAI222_X1 U9237 ( .A1(n9675), .A2(n7543), .B1(n6745), .B2(P1_U3086), .C1(
        n7523), .C2(n8195), .ZN(P1_U3335) );
  OAI21_X1 U9238 ( .B1(n7525), .B2(n4279), .A(n7524), .ZN(n7541) );
  XNOR2_X1 U9239 ( .A(n7526), .B(n4279), .ZN(n7527) );
  NAND2_X1 U9240 ( .A1(n7527), .A2(n8928), .ZN(n7529) );
  AOI22_X1 U9241 ( .A1(n8934), .A2(n8577), .B1(n8575), .B2(n8932), .ZN(n7528)
         );
  OAI211_X1 U9242 ( .C1(n7848), .C2(n7541), .A(n7529), .B(n7528), .ZN(n7534)
         );
  OAI22_X1 U9243 ( .A1(n7541), .A2(n7950), .B1(n7530), .B2(n8939), .ZN(n7531)
         );
  NOR2_X1 U9244 ( .A1(n7534), .A2(n7531), .ZN(n10047) );
  OR2_X1 U9245 ( .A1(n8942), .A2(n4913), .ZN(n7532) );
  OAI21_X1 U9246 ( .B1(n10047), .B2(n8944), .A(n7532), .ZN(P2_U3466) );
  NAND2_X1 U9247 ( .A1(n4275), .A2(n7533), .ZN(n7853) );
  NAND2_X1 U9248 ( .A1(n7534), .A2(n4275), .ZN(n7540) );
  OAI22_X1 U9249 ( .A1(n4275), .A2(n7536), .B1(n7535), .B2(n10017), .ZN(n7537)
         );
  AOI21_X1 U9250 ( .B1(n10026), .B2(n7538), .A(n7537), .ZN(n7539) );
  OAI211_X1 U9251 ( .C1(n7541), .C2(n7853), .A(n7540), .B(n7539), .ZN(P2_U3226) );
  OAI222_X1 U9252 ( .A1(n7544), .A2(P2_U3151), .B1(n8056), .B2(n7543), .C1(
        n7542), .C2(n9021), .ZN(P2_U3275) );
  NAND2_X1 U9253 ( .A1(n7545), .A2(n8432), .ZN(n7546) );
  AND2_X1 U9254 ( .A1(n8438), .A2(n8436), .ZN(n8340) );
  XNOR2_X1 U9255 ( .A(n7546), .B(n8340), .ZN(n10024) );
  NOR2_X1 U9256 ( .A1(n10024), .A2(n8940), .ZN(n7550) );
  XOR2_X1 U9257 ( .A(n7547), .B(n8340), .Z(n7548) );
  OAI222_X1 U9258 ( .A1(n8867), .A2(n7637), .B1(n8865), .B2(n7549), .C1(n7548), 
        .C2(n8862), .ZN(n10016) );
  AOI211_X1 U9259 ( .C1(n8915), .C2(n7581), .A(n7550), .B(n10016), .ZN(n10045)
         );
  OR2_X1 U9260 ( .A1(n10045), .A2(n8944), .ZN(n7551) );
  OAI21_X1 U9261 ( .B1(n8942), .B2(n7552), .A(n7551), .ZN(P2_U3465) );
  NAND2_X1 U9262 ( .A1(n8687), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7553) );
  OAI21_X1 U9263 ( .B1(n8329), .B2(n8687), .A(n7553), .ZN(P2_U3521) );
  XOR2_X1 U9264 ( .A(n7554), .B(n7558), .Z(n9970) );
  INV_X1 U9265 ( .A(n7555), .ZN(n7556) );
  AOI21_X1 U9266 ( .B1(n9839), .B2(n7557), .A(n7556), .ZN(n7559) );
  NAND2_X1 U9267 ( .A1(n7559), .A2(n7558), .ZN(n9819) );
  OAI211_X1 U9268 ( .C1(n7559), .C2(n7558), .A(n9819), .B(n9868), .ZN(n7562)
         );
  NAND2_X1 U9269 ( .A1(n9171), .A2(n9131), .ZN(n7560) );
  OAI21_X1 U9270 ( .B1(n7680), .B2(n9129), .A(n7560), .ZN(n7802) );
  INV_X1 U9271 ( .A(n7802), .ZN(n7561) );
  NAND2_X1 U9272 ( .A1(n7562), .A2(n7561), .ZN(n9965) );
  OAI21_X1 U9273 ( .B1(n9846), .B2(n6039), .A(n9901), .ZN(n7564) );
  NOR2_X1 U9274 ( .A1(n7564), .A2(n7563), .ZN(n9966) );
  NAND2_X1 U9275 ( .A1(n9966), .A2(n9905), .ZN(n7567) );
  OAI22_X1 U9276 ( .A1(n9836), .A2(n4479), .B1(n7804), .B2(n9878), .ZN(n7565)
         );
  AOI21_X1 U9277 ( .B1(n9906), .B2(n9967), .A(n7565), .ZN(n7566) );
  NAND2_X1 U9278 ( .A1(n7567), .A2(n7566), .ZN(n7568) );
  AOI21_X1 U9279 ( .B1(n9965), .B2(n9836), .A(n7568), .ZN(n7569) );
  OAI21_X1 U9280 ( .B1(n9970), .B2(n9412), .A(n7569), .ZN(P1_U3285) );
  INV_X1 U9281 ( .A(n10018), .ZN(n7570) );
  NAND2_X1 U9282 ( .A1(n8305), .A2(n7570), .ZN(n7574) );
  INV_X1 U9283 ( .A(n7571), .ZN(n7572) );
  AOI21_X1 U9284 ( .B1(n8293), .B2(n8578), .A(n7572), .ZN(n7573) );
  OAI211_X1 U9285 ( .C1(n7637), .C2(n8295), .A(n7574), .B(n7573), .ZN(n7580)
         );
  INV_X1 U9286 ( .A(n7576), .ZN(n7577) );
  AOI211_X1 U9287 ( .C1(n7578), .C2(n7575), .A(n8312), .B(n7577), .ZN(n7579)
         );
  AOI211_X1 U9288 ( .C1(n7581), .C2(n8310), .A(n7580), .B(n7579), .ZN(n7582)
         );
  INV_X1 U9289 ( .A(n7582), .ZN(P2_U3179) );
  XNOR2_X1 U9290 ( .A(n7585), .B(n7584), .ZN(n7586) );
  XNOR2_X1 U9291 ( .A(n7583), .B(n7586), .ZN(n7592) );
  NAND2_X1 U9292 ( .A1(n9172), .A2(n9131), .ZN(n7587) );
  OAI21_X1 U9293 ( .B1(n7588), .B2(n9129), .A(n7587), .ZN(n9842) );
  AOI22_X1 U9294 ( .A1(n9842), .A2(n9753), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7590) );
  OR2_X1 U9295 ( .A1(n9749), .A2(n9959), .ZN(n7589) );
  OAI211_X1 U9296 ( .C1(n9135), .C2(n9843), .A(n7590), .B(n7589), .ZN(n7591)
         );
  AOI21_X1 U9297 ( .B1(n7592), .B2(n9148), .A(n7591), .ZN(n7593) );
  INV_X1 U9298 ( .A(n7593), .ZN(P1_U3213) );
  OAI21_X1 U9299 ( .B1(n7595), .B2(n7435), .A(n7594), .ZN(n7599) );
  NOR2_X1 U9300 ( .A1(n7620), .A2(n7596), .ZN(n7597) );
  AOI21_X1 U9301 ( .B1(n7596), .B2(n7620), .A(n7597), .ZN(n7598) );
  NOR2_X1 U9302 ( .A1(n7599), .A2(n7598), .ZN(n7621) );
  AOI21_X1 U9303 ( .B1(n7599), .B2(n7598), .A(n7621), .ZN(n7601) );
  AND2_X1 U9304 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8034) );
  AOI21_X1 U9305 ( .B1(n9794), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8034), .ZN(
        n7600) );
  OAI21_X1 U9306 ( .B1(n9242), .B2(n7601), .A(n7600), .ZN(n7608) );
  NOR2_X1 U9307 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7620), .ZN(n7604) );
  AOI21_X1 U9308 ( .B1(n7620), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7604), .ZN(
        n7605) );
  AOI221_X1 U9309 ( .B1(n7606), .B2(n7617), .C1(n7605), .C2(n7617), .A(n9784), 
        .ZN(n7607) );
  AOI211_X1 U9310 ( .C1(n9776), .C2(n7620), .A(n7608), .B(n7607), .ZN(n7609)
         );
  INV_X1 U9311 ( .A(n7609), .ZN(P1_U3255) );
  XOR2_X1 U9312 ( .A(n7611), .B(n7610), .Z(n7616) );
  NAND2_X1 U9313 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n8588) );
  OAI21_X1 U9314 ( .B1(n8308), .B2(n7637), .A(n8588), .ZN(n7612) );
  AOI21_X1 U9315 ( .B1(n8304), .B2(n8574), .A(n7612), .ZN(n7613) );
  OAI21_X1 U9316 ( .B1(n8067), .B2(n4787), .A(n7613), .ZN(n7614) );
  AOI21_X1 U9317 ( .B1(n7646), .B2(n8310), .A(n7614), .ZN(n7615) );
  OAI21_X1 U9318 ( .B1(n7616), .B2(n8312), .A(n7615), .ZN(P2_U3161) );
  AOI22_X1 U9319 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7714), .B1(n7707), .B2(
        n6072), .ZN(n7619) );
  OAI21_X1 U9320 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7620), .A(n7617), .ZN(
        n7618) );
  NOR2_X1 U9321 ( .A1(n7619), .A2(n7618), .ZN(n7706) );
  AOI211_X1 U9322 ( .C1(n7619), .C2(n7618), .A(n7706), .B(n9784), .ZN(n7633)
         );
  OR2_X1 U9323 ( .A1(n7620), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7623) );
  INV_X1 U9324 ( .A(n7621), .ZN(n7622) );
  AND2_X1 U9325 ( .A1(n7623), .A2(n7622), .ZN(n7627) );
  OR2_X1 U9326 ( .A1(n7707), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9327 ( .A1(n7707), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7624) );
  AND2_X1 U9328 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U9329 ( .A1(n7626), .A2(n7627), .ZN(n7713) );
  OAI211_X1 U9330 ( .C1(n7627), .C2(n7626), .A(n9789), .B(n7713), .ZN(n7631)
         );
  NOR2_X1 U9331 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7628), .ZN(n7629) );
  AOI21_X1 U9332 ( .B1(n9794), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7629), .ZN(
        n7630) );
  OAI211_X1 U9333 ( .C1(n9798), .C2(n7714), .A(n7631), .B(n7630), .ZN(n7632)
         );
  OR2_X1 U9334 ( .A1(n7633), .A2(n7632), .ZN(P1_U3256) );
  INV_X1 U9335 ( .A(n8420), .ZN(n7634) );
  OR2_X1 U9336 ( .A1(n7634), .A2(n8422), .ZN(n8343) );
  XNOR2_X1 U9337 ( .A(n7635), .B(n8343), .ZN(n7636) );
  OAI222_X1 U9338 ( .A1(n8867), .A2(n7825), .B1(n8865), .B2(n7637), .C1(n8862), 
        .C2(n7636), .ZN(n7644) );
  NAND2_X1 U9339 ( .A1(n7524), .A2(n7638), .ZN(n7639) );
  XOR2_X1 U9340 ( .A(n8343), .B(n7639), .Z(n7649) );
  OAI22_X1 U9341 ( .A1(n7649), .A2(n8940), .B1(n7640), .B2(n8939), .ZN(n7641)
         );
  NOR2_X1 U9342 ( .A1(n7644), .A2(n7641), .ZN(n10049) );
  OR2_X1 U9343 ( .A1(n8942), .A2(n5490), .ZN(n7642) );
  OAI21_X1 U9344 ( .B1(n10049), .B2(n8944), .A(n7642), .ZN(P2_U3467) );
  INV_X1 U9345 ( .A(n5725), .ZN(n7651) );
  OAI222_X1 U9346 ( .A1(n9675), .A2(n7651), .B1(P1_U3086), .B2(n7643), .C1(
        n9514), .C2(n8194), .ZN(P1_U3334) );
  NAND2_X1 U9347 ( .A1(n7644), .A2(n4275), .ZN(n7648) );
  OAI22_X1 U9348 ( .A1(n4275), .A2(n4888), .B1(n4787), .B2(n10017), .ZN(n7645)
         );
  AOI21_X1 U9349 ( .B1(n10026), .B2(n7646), .A(n7645), .ZN(n7647) );
  OAI211_X1 U9350 ( .C1(n7649), .C2(n10025), .A(n7648), .B(n7647), .ZN(
        P2_U3225) );
  INV_X1 U9351 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7650) );
  OAI222_X1 U9352 ( .A1(n8390), .A2(P2_U3151), .B1(n8056), .B2(n7651), .C1(
        n7650), .C2(n9021), .ZN(P2_U3274) );
  AOI21_X1 U9353 ( .B1(n7652), .B2(n7653), .A(n8312), .ZN(n7655) );
  NAND2_X1 U9354 ( .A1(n7655), .A2(n7654), .ZN(n7660) );
  INV_X1 U9355 ( .A(n7700), .ZN(n7658) );
  NOR2_X1 U9356 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5020), .ZN(n7663) );
  AOI21_X1 U9357 ( .B1(n8293), .B2(n8575), .A(n7663), .ZN(n7656) );
  OAI21_X1 U9358 ( .B1(n7936), .B2(n8295), .A(n7656), .ZN(n7657) );
  AOI21_X1 U9359 ( .B1(n7658), .B2(n8305), .A(n7657), .ZN(n7659) );
  OAI211_X1 U9360 ( .C1(n7696), .C2(n8299), .A(n7660), .B(n7659), .ZN(P2_U3171) );
  AOI21_X1 U9361 ( .B1(n7662), .B2(n5018), .A(n7661), .ZN(n7677) );
  INV_X1 U9362 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9694) );
  INV_X1 U9363 ( .A(n7663), .ZN(n7669) );
  OAI21_X1 U9364 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7667) );
  NAND2_X1 U9365 ( .A1(n8665), .A2(n7667), .ZN(n7668) );
  OAI211_X1 U9366 ( .C1(n8695), .C2(n9694), .A(n7669), .B(n7668), .ZN(n7674)
         );
  AOI21_X1 U9367 ( .B1(n5019), .B2(n7671), .A(n7670), .ZN(n7672) );
  NOR2_X1 U9368 ( .A1(n7672), .A2(n8698), .ZN(n7673) );
  AOI211_X1 U9369 ( .C1(n8674), .C2(n7675), .A(n7674), .B(n7673), .ZN(n7676)
         );
  OAI21_X1 U9370 ( .B1(n7677), .B2(n8675), .A(n7676), .ZN(P2_U3191) );
  OAI21_X1 U9371 ( .B1(n7683), .B2(n7679), .A(n7678), .ZN(n7681) );
  OAI22_X1 U9372 ( .A1(n7726), .A2(n9129), .B1(n7680), .B2(n9117), .ZN(n9752)
         );
  AOI21_X1 U9373 ( .B1(n7681), .B2(n9868), .A(n9752), .ZN(n9985) );
  XNOR2_X1 U9374 ( .A(n7682), .B(n7683), .ZN(n9988) );
  NAND2_X1 U9375 ( .A1(n9988), .A2(n9874), .ZN(n7689) );
  OAI22_X1 U9376 ( .A1(n9836), .A2(n7684), .B1(n9759), .B2(n9878), .ZN(n7686)
         );
  OAI211_X1 U9377 ( .C1(n5675), .C2(n5674), .A(n9901), .B(n9813), .ZN(n9984)
         );
  NOR2_X1 U9378 ( .A1(n9984), .A2(n9831), .ZN(n7685) );
  AOI211_X1 U9379 ( .C1(n9906), .C2(n7687), .A(n7686), .B(n7685), .ZN(n7688)
         );
  OAI211_X1 U9380 ( .C1(n9898), .C2(n9985), .A(n7689), .B(n7688), .ZN(P1_U3283) );
  OAI21_X1 U9381 ( .B1(n7691), .B2(n8345), .A(n7690), .ZN(n7705) );
  XNOR2_X1 U9382 ( .A(n7692), .B(n8345), .ZN(n7693) );
  NAND2_X1 U9383 ( .A1(n7693), .A2(n8928), .ZN(n7695) );
  AOI22_X1 U9384 ( .A1(n8934), .A2(n8575), .B1(n8573), .B2(n8932), .ZN(n7694)
         );
  OAI211_X1 U9385 ( .C1(n7848), .C2(n7705), .A(n7695), .B(n7694), .ZN(n7699)
         );
  OAI22_X1 U9386 ( .A1(n7705), .A2(n7950), .B1(n7696), .B2(n8939), .ZN(n7697)
         );
  NOR2_X1 U9387 ( .A1(n7699), .A2(n7697), .ZN(n10051) );
  OR2_X1 U9388 ( .A1(n8942), .A2(n5018), .ZN(n7698) );
  OAI21_X1 U9389 ( .B1(n10051), .B2(n8944), .A(n7698), .ZN(P2_U3468) );
  NAND2_X1 U9390 ( .A1(n7699), .A2(n4275), .ZN(n7704) );
  OAI22_X1 U9391 ( .A1(n4275), .A2(n5019), .B1(n7700), .B2(n10017), .ZN(n7701)
         );
  AOI21_X1 U9392 ( .B1(n7702), .B2(n10026), .A(n7701), .ZN(n7703) );
  OAI211_X1 U9393 ( .C1(n7705), .C2(n7853), .A(n7704), .B(n7703), .ZN(P2_U3224) );
  NAND2_X1 U9394 ( .A1(n7980), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7708) );
  OAI21_X1 U9395 ( .B1(n7980), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7708), .ZN(
        n7709) );
  AOI211_X1 U9396 ( .C1(n7710), .C2(n7709), .A(n7979), .B(n9784), .ZN(n7721)
         );
  NOR2_X1 U9397 ( .A1(n7983), .A2(n7711), .ZN(n7712) );
  AOI21_X1 U9398 ( .B1(n7711), .B2(n7983), .A(n7712), .ZN(n7716) );
  OAI21_X1 U9399 ( .B1(n7714), .B2(n6071), .A(n7713), .ZN(n7715) );
  NAND2_X1 U9400 ( .A1(n7716), .A2(n7715), .ZN(n7982) );
  OAI211_X1 U9401 ( .C1(n7716), .C2(n7715), .A(n9789), .B(n7982), .ZN(n7719)
         );
  AND2_X1 U9402 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7717) );
  AOI21_X1 U9403 ( .B1(n9794), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7717), .ZN(
        n7718) );
  OAI211_X1 U9404 ( .C1(n9798), .C2(n7983), .A(n7719), .B(n7718), .ZN(n7720)
         );
  OR2_X1 U9405 ( .A1(n7721), .A2(n7720), .ZN(P1_U3257) );
  NAND2_X1 U9406 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  XNOR2_X1 U9407 ( .A(n7724), .B(n4440), .ZN(n7725) );
  NAND2_X1 U9408 ( .A1(n7725), .A2(n9868), .ZN(n7728) );
  OAI22_X1 U9409 ( .A1(n7726), .A2(n9117), .B1(n7897), .B2(n9129), .ZN(n8035)
         );
  INV_X1 U9410 ( .A(n8035), .ZN(n7727) );
  NAND2_X1 U9411 ( .A1(n7728), .A2(n7727), .ZN(n7764) );
  INV_X1 U9412 ( .A(n7764), .ZN(n7737) );
  XNOR2_X1 U9413 ( .A(n7729), .B(n7730), .ZN(n7766) );
  NAND2_X1 U9414 ( .A1(n7766), .A2(n9874), .ZN(n7736) );
  AOI211_X1 U9415 ( .C1(n7768), .C2(n4343), .A(n9425), .B(n7731), .ZN(n7765)
         );
  NOR2_X1 U9416 ( .A1(n8038), .A2(n9427), .ZN(n7734) );
  OAI22_X1 U9417 ( .A1(n9836), .A2(n7732), .B1(n8032), .B2(n9878), .ZN(n7733)
         );
  AOI211_X1 U9418 ( .C1(n7765), .C2(n9905), .A(n7734), .B(n7733), .ZN(n7735)
         );
  OAI211_X1 U9419 ( .C1(n9898), .C2(n7737), .A(n7736), .B(n7735), .ZN(P1_U3281) );
  INV_X1 U9420 ( .A(n7738), .ZN(n7739) );
  AOI21_X1 U9421 ( .B1(n7741), .B2(n7740), .A(n7739), .ZN(n7757) );
  INV_X1 U9422 ( .A(n7742), .ZN(n7755) );
  INV_X1 U9423 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9698) );
  OAI21_X1 U9424 ( .B1(n7745), .B2(n7744), .A(n7743), .ZN(n7747) );
  INV_X1 U9425 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7746) );
  NOR2_X1 U9426 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7746), .ZN(n7827) );
  AOI21_X1 U9427 ( .B1(n7747), .B2(n8665), .A(n7827), .ZN(n7748) );
  OAI21_X1 U9428 ( .B1(n9698), .B2(n8695), .A(n7748), .ZN(n7754) );
  NAND2_X1 U9429 ( .A1(n7750), .A2(n7749), .ZN(n7751) );
  AOI21_X1 U9430 ( .B1(n7752), .B2(n7751), .A(n8675), .ZN(n7753) );
  AOI211_X1 U9431 ( .C1(n8674), .C2(n7755), .A(n7754), .B(n7753), .ZN(n7756)
         );
  OAI21_X1 U9432 ( .B1(n7757), .B2(n8698), .A(n7756), .ZN(P2_U3192) );
  INV_X1 U9433 ( .A(n7758), .ZN(n7763) );
  NAND2_X1 U9434 ( .A1(n9673), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7759) );
  OAI211_X1 U9435 ( .C1(n7763), .C2(n9675), .A(n7760), .B(n7759), .ZN(P1_U3332) );
  NAND2_X1 U9436 ( .A1(n7761), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8561) );
  NAND2_X1 U9437 ( .A1(n8093), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7762) );
  OAI211_X1 U9438 ( .C1(n7763), .C2(n9024), .A(n8561), .B(n7762), .ZN(P2_U3272) );
  INV_X1 U9439 ( .A(n9941), .ZN(n9987) );
  AOI211_X1 U9440 ( .C1(n7766), .C2(n9987), .A(n7765), .B(n7764), .ZN(n7770)
         );
  AOI22_X1 U9441 ( .A1(n7768), .A2(n6529), .B1(n10013), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7767) );
  OAI21_X1 U9442 ( .B1(n7770), .B2(n10013), .A(n7767), .ZN(P1_U3534) );
  AOI22_X1 U9443 ( .A1(n7768), .A2(n5816), .B1(n9998), .B2(
        P1_REG0_REG_12__SCAN_IN), .ZN(n7769) );
  OAI21_X1 U9444 ( .B1(n7770), .B2(n9998), .A(n7769), .ZN(P1_U3489) );
  INV_X1 U9445 ( .A(n7771), .ZN(n7774) );
  OAI222_X1 U9446 ( .A1(n8195), .A2(n9604), .B1(n9675), .B2(n7774), .C1(n7772), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  OAI222_X1 U9447 ( .A1(P2_U3151), .A2(n7775), .B1(n8056), .B2(n7774), .C1(
        n7773), .C2(n9021), .ZN(P2_U3273) );
  OAI21_X1 U9448 ( .B1(n7778), .B2(n7777), .A(n7776), .ZN(n7782) );
  INV_X1 U9449 ( .A(n7779), .ZN(n7780) );
  NAND2_X1 U9450 ( .A1(n7776), .A2(n7780), .ZN(n7781) );
  NAND3_X1 U9451 ( .A1(n7782), .A2(n7781), .A3(n9868), .ZN(n7784) );
  OAI22_X1 U9452 ( .A1(n7997), .A2(n9129), .B1(n7961), .B2(n9117), .ZN(n8085)
         );
  INV_X1 U9453 ( .A(n8085), .ZN(n7783) );
  NAND2_X1 U9454 ( .A1(n7784), .A2(n7783), .ZN(n7923) );
  INV_X1 U9455 ( .A(n7923), .ZN(n7794) );
  OAI21_X1 U9456 ( .B1(n7787), .B2(n7786), .A(n7785), .ZN(n7925) );
  NAND2_X1 U9457 ( .A1(n7925), .A2(n9874), .ZN(n7793) );
  INV_X1 U9458 ( .A(n7731), .ZN(n7789) );
  INV_X1 U9459 ( .A(n7903), .ZN(n7788) );
  AOI211_X1 U9460 ( .C1(n8089), .C2(n7789), .A(n9425), .B(n7788), .ZN(n7924)
         );
  NOR2_X1 U9461 ( .A1(n7930), .A2(n9427), .ZN(n7791) );
  OAI22_X1 U9462 ( .A1(n9836), .A2(n6072), .B1(n8087), .B2(n9878), .ZN(n7790)
         );
  AOI211_X1 U9463 ( .C1(n7924), .C2(n9905), .A(n7791), .B(n7790), .ZN(n7792)
         );
  OAI211_X1 U9464 ( .C1(n9898), .C2(n7794), .A(n7793), .B(n7792), .ZN(P1_U3280) );
  INV_X1 U9465 ( .A(n7796), .ZN(n7798) );
  INV_X1 U9466 ( .A(n7795), .ZN(n7797) );
  AND2_X1 U9467 ( .A1(n7795), .A2(n7796), .ZN(n7854) );
  AOI21_X1 U9468 ( .B1(n7798), .B2(n7797), .A(n7854), .ZN(n7799) );
  NAND2_X1 U9469 ( .A1(n7799), .A2(n7800), .ZN(n7856) );
  OAI21_X1 U9470 ( .B1(n7800), .B2(n7799), .A(n7856), .ZN(n7807) );
  NOR2_X1 U9471 ( .A1(n6039), .A2(n9749), .ZN(n7806) );
  AOI21_X1 U9472 ( .B1(n7802), .B2(n9753), .A(n7801), .ZN(n7803) );
  OAI21_X1 U9473 ( .B1(n9760), .B2(n7804), .A(n7803), .ZN(n7805) );
  AOI211_X1 U9474 ( .C1(n7807), .C2(n9148), .A(n7806), .B(n7805), .ZN(n7808)
         );
  INV_X1 U9475 ( .A(n7808), .ZN(P1_U3221) );
  AOI21_X1 U9476 ( .B1(n7810), .B2(n5048), .A(n7809), .ZN(n7824) );
  INV_X1 U9477 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9702) );
  AND2_X1 U9478 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7873) );
  INV_X1 U9479 ( .A(n7873), .ZN(n7816) );
  OAI21_X1 U9480 ( .B1(n7813), .B2(n7812), .A(n7811), .ZN(n7814) );
  NAND2_X1 U9481 ( .A1(n8665), .A2(n7814), .ZN(n7815) );
  OAI211_X1 U9482 ( .C1(n8695), .C2(n9702), .A(n7816), .B(n7815), .ZN(n7821)
         );
  AOI21_X1 U9483 ( .B1(n5049), .B2(n7818), .A(n7817), .ZN(n7819) );
  NOR2_X1 U9484 ( .A1(n7819), .A2(n8698), .ZN(n7820) );
  AOI211_X1 U9485 ( .C1(n8674), .C2(n7822), .A(n7821), .B(n7820), .ZN(n7823)
         );
  OAI21_X1 U9486 ( .B1(n7824), .B2(n8675), .A(n7823), .ZN(P2_U3193) );
  XNOR2_X1 U9487 ( .A(n7867), .B(n8573), .ZN(n7869) );
  XOR2_X1 U9488 ( .A(n7868), .B(n7869), .Z(n7831) );
  NOR2_X1 U9489 ( .A1(n8308), .A2(n7825), .ZN(n7826) );
  AOI211_X1 U9490 ( .C1(n8304), .C2(n8572), .A(n7827), .B(n7826), .ZN(n7828)
         );
  OAI21_X1 U9491 ( .B1(n7849), .B2(n8067), .A(n7828), .ZN(n7829) );
  AOI21_X1 U9492 ( .B1(n7954), .B2(n8310), .A(n7829), .ZN(n7830) );
  OAI21_X1 U9493 ( .B1(n7831), .B2(n8312), .A(n7830), .ZN(P2_U3157) );
  OAI211_X1 U9494 ( .C1(n7834), .C2(n7833), .A(n7832), .B(n5916), .ZN(n7839)
         );
  INV_X1 U9495 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7835) );
  OR2_X1 U9496 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7835), .ZN(n7885) );
  OAI21_X1 U9497 ( .B1(n8308), .B2(n8044), .A(n7885), .ZN(n7837) );
  NOR2_X1 U9498 ( .A1(n8067), .A2(n8049), .ZN(n7836) );
  AOI211_X1 U9499 ( .C1(n8304), .C2(n8933), .A(n7837), .B(n7836), .ZN(n7838)
         );
  OAI211_X1 U9500 ( .C1(n8449), .C2(n8299), .A(n7839), .B(n7838), .ZN(P2_U3164) );
  NAND2_X1 U9501 ( .A1(n7690), .A2(n8421), .ZN(n7843) );
  INV_X1 U9502 ( .A(n7840), .ZN(n7842) );
  NAND2_X1 U9503 ( .A1(n7842), .A2(n7841), .ZN(n8346) );
  XNOR2_X1 U9504 ( .A(n7843), .B(n8346), .ZN(n7951) );
  XNOR2_X1 U9505 ( .A(n7844), .B(n8346), .ZN(n7845) );
  NAND2_X1 U9506 ( .A1(n7845), .A2(n8928), .ZN(n7847) );
  AOI22_X1 U9507 ( .A1(n8934), .A2(n8574), .B1(n8572), .B2(n8932), .ZN(n7846)
         );
  OAI211_X1 U9508 ( .C1(n7848), .C2(n7951), .A(n7847), .B(n7846), .ZN(n7952)
         );
  NAND2_X1 U9509 ( .A1(n7952), .A2(n4275), .ZN(n7852) );
  OAI22_X1 U9510 ( .A1(n4275), .A2(n5458), .B1(n7849), .B2(n10017), .ZN(n7850)
         );
  AOI21_X1 U9511 ( .B1(n7954), .B2(n10026), .A(n7850), .ZN(n7851) );
  OAI211_X1 U9512 ( .C1(n7951), .C2(n7853), .A(n7852), .B(n7851), .ZN(P2_U3223) );
  INV_X1 U9513 ( .A(n7854), .ZN(n7855) );
  NAND2_X1 U9514 ( .A1(n7856), .A2(n7855), .ZN(n7860) );
  XNOR2_X1 U9515 ( .A(n7858), .B(n7857), .ZN(n7859) );
  XNOR2_X1 U9516 ( .A(n7860), .B(n7859), .ZN(n7865) );
  NAND2_X1 U9517 ( .A1(n9170), .A2(n9131), .ZN(n9824) );
  NAND2_X1 U9518 ( .A1(n9168), .A2(n9086), .ZN(n9832) );
  NAND2_X1 U9519 ( .A1(n9824), .A2(n9832), .ZN(n9975) );
  AOI21_X1 U9520 ( .B1(n9975), .B2(n9753), .A(n7861), .ZN(n7863) );
  NAND2_X1 U9521 ( .A1(n9976), .A2(n9141), .ZN(n7862) );
  OAI211_X1 U9522 ( .C1(n9135), .C2(n9823), .A(n7863), .B(n7862), .ZN(n7864)
         );
  AOI21_X1 U9523 ( .B1(n7865), .B2(n9148), .A(n7864), .ZN(n7866) );
  INV_X1 U9524 ( .A(n7866), .ZN(P1_U3231) );
  OAI22_X1 U9525 ( .A1(n7869), .A2(n7868), .B1(n8573), .B2(n7867), .ZN(n7870)
         );
  XOR2_X1 U9526 ( .A(n7871), .B(n7870), .Z(n7877) );
  NOR2_X1 U9527 ( .A1(n8308), .A2(n7936), .ZN(n7872) );
  AOI211_X1 U9528 ( .C1(n8304), .C2(n8571), .A(n7873), .B(n7872), .ZN(n7874)
         );
  OAI21_X1 U9529 ( .B1(n7944), .B2(n8067), .A(n7874), .ZN(n7875) );
  AOI21_X1 U9530 ( .B1(n7946), .B2(n8310), .A(n7875), .ZN(n7876) );
  OAI21_X1 U9531 ( .B1(n7877), .B2(n8312), .A(n7876), .ZN(P2_U3176) );
  AOI21_X1 U9532 ( .B1(n7879), .B2(n7878), .A(n4335), .ZN(n7894) );
  INV_X1 U9533 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9706) );
  OAI21_X1 U9534 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7883) );
  NAND2_X1 U9535 ( .A1(n8665), .A2(n7883), .ZN(n7884) );
  OAI211_X1 U9536 ( .C1(n8695), .C2(n9706), .A(n7885), .B(n7884), .ZN(n7891)
         );
  NAND2_X1 U9537 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  AOI21_X1 U9538 ( .B1(n7889), .B2(n7888), .A(n8675), .ZN(n7890) );
  AOI211_X1 U9539 ( .C1(n8674), .C2(n7892), .A(n7891), .B(n7890), .ZN(n7893)
         );
  OAI21_X1 U9540 ( .B1(n7894), .B2(n8698), .A(n7893), .ZN(P2_U3194) );
  INV_X1 U9541 ( .A(n7992), .ZN(n7895) );
  AOI211_X1 U9542 ( .C1(n7900), .C2(n7896), .A(n9895), .B(n7895), .ZN(n7898)
         );
  OAI22_X1 U9543 ( .A1(n8121), .A2(n9129), .B1(n7897), .B2(n9117), .ZN(n9029)
         );
  OR2_X1 U9544 ( .A1(n7898), .A2(n9029), .ZN(n7971) );
  INV_X1 U9545 ( .A(n7971), .ZN(n7909) );
  OAI21_X1 U9546 ( .B1(n7901), .B2(n7900), .A(n7899), .ZN(n7973) );
  NAND2_X1 U9547 ( .A1(n7973), .A2(n9874), .ZN(n7908) );
  INV_X1 U9548 ( .A(n8004), .ZN(n7902) );
  AOI211_X1 U9549 ( .C1(n9033), .C2(n7903), .A(n9425), .B(n7902), .ZN(n7972)
         );
  INV_X1 U9550 ( .A(n9033), .ZN(n7978) );
  NOR2_X1 U9551 ( .A1(n7978), .A2(n9427), .ZN(n7906) );
  OAI22_X1 U9552 ( .A1(n9836), .A2(n7904), .B1(n9031), .B2(n9878), .ZN(n7905)
         );
  AOI211_X1 U9553 ( .C1(n7972), .C2(n9905), .A(n7906), .B(n7905), .ZN(n7907)
         );
  OAI211_X1 U9554 ( .C1(n9898), .C2(n7909), .A(n7908), .B(n7907), .ZN(P1_U3279) );
  INV_X1 U9555 ( .A(n7910), .ZN(n7932) );
  INV_X1 U9556 ( .A(n7911), .ZN(n7913) );
  OAI222_X1 U9557 ( .A1(n9675), .A2(n7932), .B1(P1_U3086), .B2(n7913), .C1(
        n7912), .C2(n8194), .ZN(P1_U3331) );
  XNOR2_X1 U9558 ( .A(n7914), .B(n8933), .ZN(n7915) );
  XNOR2_X1 U9559 ( .A(n7916), .B(n7915), .ZN(n7922) );
  NOR2_X1 U9560 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5070), .ZN(n8013) );
  NOR2_X1 U9561 ( .A1(n8295), .A2(n8866), .ZN(n7917) );
  AOI211_X1 U9562 ( .C1(n8293), .C2(n8571), .A(n8013), .B(n7917), .ZN(n7918)
         );
  OAI21_X1 U9563 ( .B1(n8876), .B2(n8067), .A(n7918), .ZN(n7919) );
  AOI21_X1 U9564 ( .B1(n7920), .B2(n8310), .A(n7919), .ZN(n7921) );
  OAI21_X1 U9565 ( .B1(n7922), .B2(n8312), .A(n7921), .ZN(P2_U3174) );
  AOI211_X1 U9566 ( .C1(n7925), .C2(n9987), .A(n7924), .B(n7923), .ZN(n7927)
         );
  MUX2_X1 U9567 ( .A(n6071), .B(n7927), .S(n10015), .Z(n7926) );
  OAI21_X1 U9568 ( .B1(n7930), .B2(n9633), .A(n7926), .ZN(P1_U3535) );
  INV_X1 U9569 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7928) );
  MUX2_X1 U9570 ( .A(n7928), .B(n7927), .S(n10000), .Z(n7929) );
  OAI21_X1 U9571 ( .B1(n7930), .B2(n9667), .A(n7929), .ZN(P1_U3492) );
  OAI222_X1 U9572 ( .A1(n7933), .A2(P2_U3151), .B1(n9024), .B2(n7932), .C1(
        n7931), .C2(n9021), .ZN(P2_U3271) );
  XNOR2_X1 U9573 ( .A(n7934), .B(n8348), .ZN(n7935) );
  OAI222_X1 U9574 ( .A1(n8867), .A2(n8134), .B1(n8865), .B2(n7936), .C1(n7935), 
        .C2(n8862), .ZN(n7943) );
  NAND2_X1 U9575 ( .A1(n7938), .A2(n7937), .ZN(n7939) );
  XNOR2_X1 U9576 ( .A(n7939), .B(n8348), .ZN(n7949) );
  OAI22_X1 U9577 ( .A1(n7949), .A2(n8940), .B1(n7940), .B2(n8939), .ZN(n7941)
         );
  NOR2_X1 U9578 ( .A1(n7943), .A2(n7941), .ZN(n10055) );
  OR2_X1 U9579 ( .A1(n8942), .A2(n5048), .ZN(n7942) );
  OAI21_X1 U9580 ( .B1(n10055), .B2(n8944), .A(n7942), .ZN(P2_U3470) );
  NAND2_X1 U9581 ( .A1(n7943), .A2(n4275), .ZN(n7948) );
  OAI22_X1 U9582 ( .A1(n4275), .A2(n5049), .B1(n7944), .B2(n10017), .ZN(n7945)
         );
  AOI21_X1 U9583 ( .B1(n7946), .B2(n10026), .A(n7945), .ZN(n7947) );
  OAI211_X1 U9584 ( .C1(n7949), .C2(n10025), .A(n7948), .B(n7947), .ZN(
        P2_U3222) );
  NOR2_X1 U9585 ( .A1(n7951), .A2(n7950), .ZN(n7953) );
  AOI211_X1 U9586 ( .C1(n8915), .C2(n7954), .A(n7953), .B(n7952), .ZN(n10053)
         );
  OR2_X1 U9587 ( .A1(n10053), .A2(n8944), .ZN(n7955) );
  OAI21_X1 U9588 ( .B1(n8942), .B2(n5494), .A(n7955), .ZN(P2_U3469) );
  INV_X1 U9589 ( .A(n7956), .ZN(n7959) );
  NOR3_X1 U9590 ( .A1(n4331), .A2(n4362), .A3(n7957), .ZN(n7958) );
  OAI21_X1 U9591 ( .B1(n7959), .B2(n7958), .A(n9148), .ZN(n7965) );
  OAI22_X1 U9592 ( .A1(n7961), .A2(n9129), .B1(n7960), .B2(n9117), .ZN(n9807)
         );
  AOI22_X1 U9593 ( .A1(n9807), .A2(n9753), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7962) );
  OAI21_X1 U9594 ( .B1(n9135), .B2(n9809), .A(n7962), .ZN(n7963) );
  AOI21_X1 U9595 ( .B1(n9811), .B2(n9141), .A(n7963), .ZN(n7964) );
  NAND2_X1 U9596 ( .A1(n7965), .A2(n7964), .ZN(P1_U3236) );
  INV_X1 U9597 ( .A(n7966), .ZN(n7969) );
  OAI222_X1 U9598 ( .A1(n9675), .A2(n7969), .B1(P1_U3086), .B2(n7967), .C1(
        n9517), .C2(n8194), .ZN(P1_U3330) );
  OAI222_X1 U9599 ( .A1(n7970), .A2(P2_U3151), .B1(n9024), .B2(n7969), .C1(
        n7968), .C2(n9021), .ZN(P2_U3270) );
  AOI211_X1 U9600 ( .C1(n7973), .C2(n9987), .A(n7972), .B(n7971), .ZN(n7975)
         );
  MUX2_X1 U9601 ( .A(n7711), .B(n7975), .S(n10015), .Z(n7974) );
  OAI21_X1 U9602 ( .B1(n7978), .B2(n9633), .A(n7974), .ZN(P1_U3536) );
  INV_X1 U9603 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7976) );
  MUX2_X1 U9604 ( .A(n7976), .B(n7975), .S(n10000), .Z(n7977) );
  OAI21_X1 U9605 ( .B1(n7978), .B2(n9667), .A(n7977), .ZN(P1_U3495) );
  NOR2_X1 U9606 ( .A1(n8005), .A2(n7981), .ZN(n9189) );
  AOI211_X1 U9607 ( .C1(n8005), .C2(n7981), .A(n9189), .B(n9784), .ZN(n7990)
         );
  OAI21_X1 U9608 ( .B1(n7711), .B2(n7983), .A(n7982), .ZN(n9181) );
  XNOR2_X1 U9609 ( .A(n9187), .B(n9181), .ZN(n7984) );
  NAND2_X1 U9610 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7984), .ZN(n9183) );
  OAI211_X1 U9611 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7984), .A(n9789), .B(
        n9183), .ZN(n7988) );
  NOR2_X1 U9612 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7985), .ZN(n7986) );
  AOI21_X1 U9613 ( .B1(n9794), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7986), .ZN(
        n7987) );
  OAI211_X1 U9614 ( .C1(n9798), .C2(n9187), .A(n7988), .B(n7987), .ZN(n7989)
         );
  OR2_X1 U9615 ( .A1(n7990), .A2(n7989), .ZN(P1_U3258) );
  NAND2_X1 U9616 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  NAND2_X1 U9617 ( .A1(n7993), .A2(n8001), .ZN(n7995) );
  NAND2_X1 U9618 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  NAND2_X1 U9619 ( .A1(n7996), .A2(n9868), .ZN(n7999) );
  OAI22_X1 U9620 ( .A1(n8146), .A2(n9129), .B1(n7997), .B2(n9117), .ZN(n9143)
         );
  INV_X1 U9621 ( .A(n9143), .ZN(n7998) );
  NAND2_X1 U9622 ( .A1(n7999), .A2(n7998), .ZN(n8095) );
  INV_X1 U9623 ( .A(n8095), .ZN(n8010) );
  OAI21_X1 U9624 ( .B1(n8002), .B2(n8001), .A(n4469), .ZN(n8097) );
  NAND2_X1 U9625 ( .A1(n8097), .A2(n9874), .ZN(n8009) );
  INV_X1 U9626 ( .A(n8003), .ZN(n8126) );
  AOI211_X1 U9627 ( .C1(n9142), .C2(n8004), .A(n9425), .B(n8126), .ZN(n8096)
         );
  NOR2_X1 U9628 ( .A1(n8102), .A2(n9427), .ZN(n8007) );
  OAI22_X1 U9629 ( .A1(n9836), .A2(n8005), .B1(n9146), .B2(n9878), .ZN(n8006)
         );
  AOI211_X1 U9630 ( .C1(n8096), .C2(n9905), .A(n8007), .B(n8006), .ZN(n8008)
         );
  OAI211_X1 U9631 ( .C1(n9898), .C2(n8010), .A(n8009), .B(n8008), .ZN(P1_U3278) );
  AOI21_X1 U9632 ( .B1(n8012), .B2(n5068), .A(n8011), .ZN(n8027) );
  INV_X1 U9633 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9710) );
  INV_X1 U9634 ( .A(n8013), .ZN(n8019) );
  OAI21_X1 U9635 ( .B1(n8016), .B2(n8015), .A(n8014), .ZN(n8017) );
  NAND2_X1 U9636 ( .A1(n8665), .A2(n8017), .ZN(n8018) );
  OAI211_X1 U9637 ( .C1(n8695), .C2(n9710), .A(n8019), .B(n8018), .ZN(n8024)
         );
  AOI21_X1 U9638 ( .B1(n5069), .B2(n8021), .A(n8020), .ZN(n8022) );
  NOR2_X1 U9639 ( .A1(n8022), .A2(n8698), .ZN(n8023) );
  AOI211_X1 U9640 ( .C1(n8674), .C2(n8025), .A(n8024), .B(n8023), .ZN(n8026)
         );
  OAI21_X1 U9641 ( .B1(n8027), .B2(n8675), .A(n8026), .ZN(P2_U3195) );
  AND3_X1 U9642 ( .A1(n7956), .A2(n8030), .A3(n8029), .ZN(n8031) );
  OAI21_X1 U9643 ( .B1(n8028), .B2(n8031), .A(n9148), .ZN(n8037) );
  NOR2_X1 U9644 ( .A1(n9760), .A2(n8032), .ZN(n8033) );
  AOI211_X1 U9645 ( .C1(n9753), .C2(n8035), .A(n8034), .B(n8033), .ZN(n8036)
         );
  OAI211_X1 U9646 ( .C1(n8038), .C2(n9749), .A(n8037), .B(n8036), .ZN(P1_U3224) );
  INV_X1 U9647 ( .A(n8039), .ZN(n8057) );
  OAI222_X1 U9648 ( .A1(n9675), .A2(n8057), .B1(P1_U3086), .B2(n8041), .C1(
        n8040), .C2(n8194), .ZN(P1_U3329) );
  XNOR2_X1 U9649 ( .A(n8042), .B(n8458), .ZN(n8043) );
  OAI222_X1 U9650 ( .A1(n8867), .A2(n8064), .B1(n8865), .B2(n8044), .C1(n8043), 
        .C2(n8862), .ZN(n8051) );
  OAI21_X1 U9651 ( .B1(n8046), .B2(n8458), .A(n8045), .ZN(n8055) );
  OAI22_X1 U9652 ( .A1(n8055), .A2(n8940), .B1(n8449), .B2(n8939), .ZN(n8047)
         );
  NOR2_X1 U9653 ( .A1(n8051), .A2(n8047), .ZN(n10058) );
  OR2_X1 U9654 ( .A1(n8942), .A2(n4808), .ZN(n8048) );
  OAI21_X1 U9655 ( .B1(n10058), .B2(n8944), .A(n8048), .ZN(P2_U3471) );
  NOR2_X1 U9656 ( .A1(n10017), .A2(n8049), .ZN(n8050) );
  OAI21_X1 U9657 ( .B1(n8051), .B2(n8050), .A(n4275), .ZN(n8054) );
  AOI22_X1 U9658 ( .A1(n8052), .A2(n10026), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n10034), .ZN(n8053) );
  OAI211_X1 U9659 ( .C1(n8055), .C2(n10025), .A(n8054), .B(n8053), .ZN(
        P2_U3221) );
  OAI222_X1 U9660 ( .A1(n9021), .A2(n8059), .B1(P2_U3151), .B2(n8058), .C1(
        n8057), .C2(n8056), .ZN(P2_U3269) );
  INV_X1 U9661 ( .A(n8074), .ZN(n8060) );
  AOI21_X1 U9662 ( .B1(n8062), .B2(n8061), .A(n8060), .ZN(n8070) );
  INV_X1 U9663 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8063) );
  OR2_X1 U9664 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8063), .ZN(n8616) );
  OAI21_X1 U9665 ( .B1(n8308), .B2(n8064), .A(n8616), .ZN(n8065) );
  AOI21_X1 U9666 ( .B1(n8304), .B2(n5118), .A(n8065), .ZN(n8066) );
  OAI21_X1 U9667 ( .B1(n8067), .B2(n9743), .A(n8066), .ZN(n8068) );
  AOI21_X1 U9668 ( .B1(n8468), .B2(n8310), .A(n8068), .ZN(n8069) );
  OAI21_X1 U9669 ( .B1(n8070), .B2(n8312), .A(n8069), .ZN(P2_U3155) );
  INV_X1 U9670 ( .A(n8071), .ZN(n8163) );
  OAI222_X1 U9671 ( .A1(n8072), .A2(P2_U3151), .B1(n9024), .B2(n8163), .C1(
        n9576), .C2(n9021), .ZN(P2_U3268) );
  AND2_X1 U9672 ( .A1(n8074), .A2(n8073), .ZN(n8076) );
  OAI211_X1 U9673 ( .C1(n8076), .C2(n8075), .A(n5916), .B(n8108), .ZN(n8080)
         );
  AND2_X1 U9674 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8630) );
  AOI21_X1 U9675 ( .B1(n8304), .B2(n8837), .A(n8630), .ZN(n8077) );
  OAI21_X1 U9676 ( .B1(n8866), .B2(n8308), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9677 ( .B1(n8873), .B2(n8305), .A(n8078), .ZN(n8079) );
  OAI211_X1 U9678 ( .C1(n8081), .C2(n8299), .A(n8080), .B(n8079), .ZN(P2_U3181) );
  AOI21_X1 U9679 ( .B1(n8084), .B2(n8083), .A(n8082), .ZN(n8091) );
  AOI22_X1 U9680 ( .A1(n8085), .A2(n9753), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n8086) );
  OAI21_X1 U9681 ( .B1(n9760), .B2(n8087), .A(n8086), .ZN(n8088) );
  AOI21_X1 U9682 ( .B1(n8089), .B2(n9141), .A(n8088), .ZN(n8090) );
  OAI21_X1 U9683 ( .B1(n8091), .B2(n9755), .A(n8090), .ZN(P1_U3234) );
  INV_X1 U9684 ( .A(n5955), .ZN(n8152) );
  AOI21_X1 U9685 ( .B1(n8093), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8092), .ZN(
        n8094) );
  OAI21_X1 U9686 ( .B1(n8152), .B2(n9024), .A(n8094), .ZN(P2_U3267) );
  INV_X1 U9687 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8098) );
  AOI211_X1 U9688 ( .C1(n8097), .C2(n9987), .A(n8096), .B(n8095), .ZN(n8100)
         );
  MUX2_X1 U9689 ( .A(n8098), .B(n8100), .S(n10000), .Z(n8099) );
  OAI21_X1 U9690 ( .B1(n8102), .B2(n9667), .A(n8099), .ZN(P1_U3498) );
  MUX2_X1 U9691 ( .A(n6089), .B(n8100), .S(n10015), .Z(n8101) );
  OAI21_X1 U9692 ( .B1(n8102), .B2(n9633), .A(n8101), .ZN(P1_U3537) );
  INV_X1 U9693 ( .A(n8103), .ZN(n8252) );
  INV_X1 U9694 ( .A(n8104), .ZN(n8107) );
  INV_X1 U9695 ( .A(n8105), .ZN(n8106) );
  AOI21_X1 U9696 ( .B1(n8108), .B2(n8107), .A(n8106), .ZN(n8109) );
  OAI21_X1 U9697 ( .B1(n8252), .B2(n8109), .A(n5916), .ZN(n8114) );
  INV_X1 U9698 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8110) );
  NOR2_X1 U9699 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8110), .ZN(n8644) );
  AOI21_X1 U9700 ( .B1(n8293), .B2(n5118), .A(n8644), .ZN(n8111) );
  OAI21_X1 U9701 ( .B1(n8851), .B2(n8295), .A(n8111), .ZN(n8112) );
  AOI21_X1 U9702 ( .B1(n8856), .B2(n8305), .A(n8112), .ZN(n8113) );
  OAI211_X1 U9703 ( .C1(n8115), .C2(n8299), .A(n8114), .B(n8113), .ZN(P2_U3166) );
  OAI21_X1 U9704 ( .B1(n8118), .B2(n8117), .A(n8116), .ZN(n9630) );
  XNOR2_X1 U9705 ( .A(n8120), .B(n8119), .ZN(n8122) );
  OAI22_X1 U9706 ( .A1(n9118), .A2(n9129), .B1(n8121), .B2(n9117), .ZN(n9068)
         );
  AOI21_X1 U9707 ( .B1(n8122), .B2(n9868), .A(n9068), .ZN(n9629) );
  INV_X1 U9708 ( .A(n9629), .ZN(n8129) );
  INV_X1 U9709 ( .A(n9066), .ZN(n8123) );
  AOI22_X1 U9710 ( .A1(n9898), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8123), .B2(
        n9899), .ZN(n8124) );
  OAI21_X1 U9711 ( .B1(n9668), .B2(n9427), .A(n8124), .ZN(n8128) );
  INV_X1 U9712 ( .A(n8125), .ZN(n8141) );
  OAI211_X1 U9713 ( .C1(n9668), .C2(n8126), .A(n8141), .B(n9901), .ZN(n9628)
         );
  NOR2_X1 U9714 ( .A1(n9628), .A2(n9831), .ZN(n8127) );
  AOI211_X1 U9715 ( .C1(n9836), .C2(n8129), .A(n8128), .B(n8127), .ZN(n8130)
         );
  OAI21_X1 U9716 ( .B1(n9630), .B2(n9412), .A(n8130), .ZN(P1_U3277) );
  OR2_X1 U9717 ( .A1(n8131), .A2(n4325), .ZN(n8462) );
  XNOR2_X1 U9718 ( .A(n8132), .B(n8462), .ZN(n8133) );
  OAI222_X1 U9719 ( .A1(n8867), .A2(n8866), .B1(n8865), .B2(n8134), .C1(n8862), 
        .C2(n8133), .ZN(n8879) );
  XNOR2_X1 U9720 ( .A(n8135), .B(n8462), .ZN(n8882) );
  OAI22_X1 U9721 ( .A1(n8882), .A2(n8940), .B1(n8877), .B2(n8939), .ZN(n8136)
         );
  NOR2_X1 U9722 ( .A1(n8879), .A2(n8136), .ZN(n9745) );
  OR2_X1 U9723 ( .A1(n8942), .A2(n5068), .ZN(n8137) );
  OAI21_X1 U9724 ( .B1(n9745), .B2(n8944), .A(n8137), .ZN(P2_U3472) );
  XOR2_X1 U9725 ( .A(n8138), .B(n8145), .Z(n9627) );
  INV_X1 U9726 ( .A(n8139), .ZN(n8140) );
  AOI211_X1 U9727 ( .C1(n9624), .C2(n8141), .A(n9425), .B(n8140), .ZN(n9623)
         );
  INV_X1 U9728 ( .A(n9077), .ZN(n8142) );
  AOI22_X1 U9729 ( .A1(n9898), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8142), .B2(
        n9899), .ZN(n8143) );
  OAI21_X1 U9730 ( .B1(n9082), .B2(n9427), .A(n8143), .ZN(n8149) );
  XOR2_X1 U9731 ( .A(n8145), .B(n8144), .Z(n8147) );
  OAI22_X1 U9732 ( .A1(n8168), .A2(n9129), .B1(n8146), .B2(n9117), .ZN(n9079)
         );
  AOI21_X1 U9733 ( .B1(n8147), .B2(n9868), .A(n9079), .ZN(n9626) );
  NOR2_X1 U9734 ( .A1(n9626), .A2(n9898), .ZN(n8148) );
  AOI211_X1 U9735 ( .C1(n9623), .C2(n9905), .A(n8149), .B(n8148), .ZN(n8150)
         );
  OAI21_X1 U9736 ( .B1(n9627), .B2(n9412), .A(n8150), .ZN(P1_U3276) );
  OAI222_X1 U9737 ( .A1(n9675), .A2(n8152), .B1(P1_U3086), .B2(n5778), .C1(
        n8151), .C2(n8195), .ZN(P1_U3327) );
  INV_X1 U9738 ( .A(n8153), .ZN(n8196) );
  OAI222_X1 U9739 ( .A1(P2_U3151), .A2(n8155), .B1(n9024), .B2(n8196), .C1(
        n8154), .C2(n9021), .ZN(P2_U3266) );
  INV_X1 U9740 ( .A(n8227), .ZN(n8157) );
  OAI22_X1 U9741 ( .A1(n8157), .A2(n10017), .B1(n4275), .B2(n8156), .ZN(n8160)
         );
  NOR2_X1 U9742 ( .A1(n8158), .A2(n10025), .ZN(n8159) );
  AOI211_X1 U9743 ( .C1(n10026), .C2(n5967), .A(n8160), .B(n8159), .ZN(n8161)
         );
  OAI21_X1 U9744 ( .B1(n8162), .B2(n10034), .A(n8161), .ZN(P2_U3205) );
  OAI222_X1 U9745 ( .A1(n8194), .A2(n8164), .B1(n9675), .B2(n8163), .C1(
        P1_U3086), .C2(n5779), .ZN(P1_U3328) );
  NOR2_X1 U9746 ( .A1(n4337), .A2(n8166), .ZN(n8167) );
  XNOR2_X1 U9747 ( .A(n8165), .B(n8167), .ZN(n8173) );
  OAI22_X1 U9748 ( .A1(n8169), .A2(n9129), .B1(n8168), .B2(n9117), .ZN(n9407)
         );
  AOI22_X1 U9749 ( .A1(n9407), .A2(n9753), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n8170) );
  OAI21_X1 U9750 ( .B1(n9135), .B2(n9400), .A(n8170), .ZN(n8171) );
  AOI21_X1 U9751 ( .B1(n9483), .B2(n9141), .A(n8171), .ZN(n8172) );
  OAI21_X1 U9752 ( .B1(n8173), .B2(n9755), .A(n8172), .ZN(P1_U3219) );
  INV_X1 U9753 ( .A(n8174), .ZN(n8181) );
  NOR2_X1 U9754 ( .A1(n8175), .A2(n9831), .ZN(n8180) );
  AOI22_X1 U9755 ( .A1(n8176), .A2(n9899), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9898), .ZN(n8177) );
  OAI21_X1 U9756 ( .B1(n8178), .B2(n9427), .A(n8177), .ZN(n8179) );
  OAI21_X1 U9757 ( .B1(n8183), .B2(n9412), .A(n8182), .ZN(P1_U3356) );
  NAND2_X1 U9758 ( .A1(n8184), .A2(n9905), .ZN(n8187) );
  NOR2_X1 U9759 ( .A1(n9898), .A2(n8185), .ZN(n9248) );
  AOI21_X1 U9760 ( .B1(n9898), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9248), .ZN(
        n8186) );
  OAI211_X1 U9761 ( .C1(n8188), .C2(n9427), .A(n8187), .B(n8186), .ZN(P1_U3263) );
  OAI222_X1 U9762 ( .A1(n8195), .A2(n8191), .B1(n9675), .B2(n8190), .C1(
        P1_U3086), .C2(n8189), .ZN(P1_U3336) );
  INV_X1 U9763 ( .A(n8326), .ZN(n9023) );
  OAI222_X1 U9764 ( .A1(n8194), .A2(n8193), .B1(n9675), .B2(n9023), .C1(
        P1_U3086), .C2(n8192), .ZN(P1_U3325) );
  OAI222_X1 U9765 ( .A1(n9675), .A2(n8196), .B1(P1_U3086), .B2(n5775), .C1(
        n9607), .C2(n8195), .ZN(P1_U3326) );
  NAND2_X1 U9766 ( .A1(n8197), .A2(n10028), .ZN(n8702) );
  OAI21_X1 U9767 ( .B1(n4275), .B2(n8198), .A(n8702), .ZN(n8201) );
  NOR2_X1 U9768 ( .A1(n8199), .A2(n10025), .ZN(n8200) );
  OAI21_X1 U9769 ( .B1(n8203), .B2(n10034), .A(n8202), .ZN(P2_U3204) );
  INV_X1 U9770 ( .A(n8743), .ZN(n8780) );
  XNOR2_X1 U9771 ( .A(n8204), .B(n8780), .ZN(n8209) );
  AOI22_X1 U9772 ( .A1(n8792), .A2(n8293), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8206) );
  NAND2_X1 U9773 ( .A1(n8769), .A2(n8305), .ZN(n8205) );
  OAI211_X1 U9774 ( .C1(n8735), .C2(n8295), .A(n8206), .B(n8205), .ZN(n8207)
         );
  AOI21_X1 U9775 ( .B1(n8970), .B2(n8310), .A(n8207), .ZN(n8208) );
  OAI21_X1 U9776 ( .B1(n8209), .B2(n8312), .A(n8208), .ZN(P2_U3156) );
  INV_X1 U9777 ( .A(n8210), .ZN(n8212) );
  NAND2_X1 U9778 ( .A1(n8212), .A2(n8211), .ZN(n8213) );
  XNOR2_X1 U9779 ( .A(n8214), .B(n8213), .ZN(n8221) );
  NAND2_X1 U9780 ( .A1(n8293), .A2(n8838), .ZN(n8216) );
  OAI211_X1 U9781 ( .C1(n8568), .C2(n8295), .A(n8216), .B(n8215), .ZN(n8219)
         );
  NOR2_X1 U9782 ( .A1(n8217), .A2(n8299), .ZN(n8218) );
  AOI211_X1 U9783 ( .C1(n8812), .C2(n8305), .A(n8219), .B(n8218), .ZN(n8220)
         );
  OAI21_X1 U9784 ( .B1(n8221), .B2(n8312), .A(n8220), .ZN(P2_U3159) );
  INV_X1 U9785 ( .A(n8222), .ZN(n8223) );
  XOR2_X1 U9786 ( .A(n8225), .B(n8330), .Z(n8226) );
  NOR2_X1 U9787 ( .A1(n8378), .A2(n8295), .ZN(n8230) );
  AOI22_X1 U9788 ( .A1(n8227), .A2(n8305), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8228) );
  OAI21_X1 U9789 ( .B1(n8721), .B2(n8308), .A(n8228), .ZN(n8229) );
  AOI211_X1 U9790 ( .C1(n5967), .C2(n8310), .A(n8230), .B(n8229), .ZN(n8231)
         );
  XOR2_X1 U9791 ( .A(n8232), .B(n8233), .Z(n8240) );
  OAI22_X1 U9792 ( .A1(n8568), .A2(n8308), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8234), .ZN(n8237) );
  NOR2_X1 U9793 ( .A1(n8235), .A2(n8295), .ZN(n8236) );
  AOI211_X1 U9794 ( .C1(n8795), .C2(n8305), .A(n8237), .B(n8236), .ZN(n8239)
         );
  NAND2_X1 U9795 ( .A1(n8982), .A2(n8310), .ZN(n8238) );
  OAI211_X1 U9796 ( .C1(n8240), .C2(n8312), .A(n8239), .B(n8238), .ZN(P2_U3163) );
  XOR2_X1 U9797 ( .A(n8242), .B(n8241), .Z(n8248) );
  NAND2_X1 U9798 ( .A1(n8567), .A2(n8304), .ZN(n8244) );
  AOI22_X1 U9799 ( .A1(n8738), .A2(n8305), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8243) );
  OAI211_X1 U9800 ( .C1(n8735), .C2(n8308), .A(n8244), .B(n8243), .ZN(n8245)
         );
  AOI21_X1 U9801 ( .B1(n8246), .B2(n8310), .A(n8245), .ZN(n8247) );
  OAI21_X1 U9802 ( .B1(n8248), .B2(n8312), .A(n8247), .ZN(P2_U3165) );
  INV_X1 U9803 ( .A(n8249), .ZN(n8251) );
  NOR3_X1 U9804 ( .A1(n8252), .A2(n8251), .A3(n8250), .ZN(n8255) );
  INV_X1 U9805 ( .A(n8253), .ZN(n8254) );
  OAI21_X1 U9806 ( .B1(n8255), .B2(n8254), .A(n5916), .ZN(n8260) );
  NAND2_X1 U9807 ( .A1(n8293), .A2(n8837), .ZN(n8256) );
  NAND2_X1 U9808 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8667) );
  OAI211_X1 U9809 ( .C1(n8257), .C2(n8295), .A(n8256), .B(n8667), .ZN(n8258)
         );
  AOI21_X1 U9810 ( .B1(n8841), .B2(n8305), .A(n8258), .ZN(n8259) );
  OAI211_X1 U9811 ( .C1(n8261), .C2(n8299), .A(n8260), .B(n8259), .ZN(P2_U3168) );
  XOR2_X1 U9812 ( .A(n8263), .B(n8262), .Z(n8269) );
  AOI22_X1 U9813 ( .A1(n8780), .A2(n8293), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8265) );
  NAND2_X1 U9814 ( .A1(n8745), .A2(n8305), .ZN(n8264) );
  OAI211_X1 U9815 ( .C1(n8744), .C2(n8295), .A(n8265), .B(n8264), .ZN(n8266)
         );
  AOI21_X1 U9816 ( .B1(n8267), .B2(n8310), .A(n8266), .ZN(n8268) );
  OAI21_X1 U9817 ( .B1(n8269), .B2(n8312), .A(n8268), .ZN(P2_U3169) );
  XOR2_X1 U9818 ( .A(n8271), .B(n8270), .Z(n8277) );
  INV_X1 U9819 ( .A(n8801), .ZN(n8779) );
  AOI22_X1 U9820 ( .A1(n8779), .A2(n8304), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8273) );
  NAND2_X1 U9821 ( .A1(n8305), .A2(n8802), .ZN(n8272) );
  OAI211_X1 U9822 ( .C1(n8826), .C2(n8308), .A(n8273), .B(n8272), .ZN(n8274)
         );
  AOI21_X1 U9823 ( .B1(n8275), .B2(n8310), .A(n8274), .ZN(n8276) );
  OAI21_X1 U9824 ( .B1(n8277), .B2(n8312), .A(n8276), .ZN(P2_U3173) );
  NAND2_X1 U9825 ( .A1(n8279), .A2(n8278), .ZN(n8281) );
  AOI21_X1 U9826 ( .B1(n8281), .B2(n8280), .A(n8312), .ZN(n8283) );
  NAND2_X1 U9827 ( .A1(n8283), .A2(n8282), .ZN(n8287) );
  AOI22_X1 U9828 ( .A1(n8779), .A2(n8293), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8284) );
  OAI21_X1 U9829 ( .B1(n8743), .B2(n8295), .A(n8284), .ZN(n8285) );
  AOI21_X1 U9830 ( .B1(n8783), .B2(n8305), .A(n8285), .ZN(n8286) );
  OAI211_X1 U9831 ( .C1(n8288), .C2(n8299), .A(n8287), .B(n8286), .ZN(P2_U3175) );
  INV_X1 U9832 ( .A(n8914), .ZN(n8300) );
  OAI21_X1 U9833 ( .B1(n8291), .B2(n8290), .A(n8289), .ZN(n8292) );
  NAND2_X1 U9834 ( .A1(n8292), .A2(n5916), .ZN(n8298) );
  NAND2_X1 U9835 ( .A1(n8293), .A2(n8570), .ZN(n8294) );
  NAND2_X1 U9836 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8694) );
  OAI211_X1 U9837 ( .C1(n8826), .C2(n8295), .A(n8294), .B(n8694), .ZN(n8296)
         );
  AOI21_X1 U9838 ( .B1(n8827), .B2(n8305), .A(n8296), .ZN(n8297) );
  OAI211_X1 U9839 ( .C1(n8300), .C2(n8299), .A(n8298), .B(n8297), .ZN(P2_U3178) );
  XOR2_X1 U9840 ( .A(n8303), .B(n8301), .Z(n8313) );
  NAND2_X1 U9841 ( .A1(n8566), .A2(n8304), .ZN(n8307) );
  AOI22_X1 U9842 ( .A1(n8726), .A2(n8305), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8306) );
  OAI211_X1 U9843 ( .C1(n8744), .C2(n8308), .A(n8307), .B(n8306), .ZN(n8309)
         );
  AOI21_X1 U9844 ( .B1(n8954), .B2(n8310), .A(n8309), .ZN(n8311) );
  OAI21_X1 U9845 ( .B1(n8313), .B2(n8312), .A(n8311), .ZN(P2_U3180) );
  NAND2_X1 U9846 ( .A1(n9016), .A2(n8325), .ZN(n8315) );
  NAND2_X1 U9847 ( .A1(n4926), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8314) );
  INV_X1 U9848 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U9849 ( .A1(n8316), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8320) );
  INV_X1 U9850 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8317) );
  OR2_X1 U9851 ( .A1(n8318), .A2(n8317), .ZN(n8319) );
  OAI211_X1 U9852 ( .C1(n8321), .C2(n4960), .A(n8320), .B(n8319), .ZN(n8322)
         );
  INV_X1 U9853 ( .A(n8322), .ZN(n8323) );
  AND2_X1 U9854 ( .A1(n8324), .A2(n8323), .ZN(n8701) );
  NAND2_X1 U9855 ( .A1(n8945), .A2(n8701), .ZN(n8545) );
  INV_X1 U9856 ( .A(n8701), .ZN(n8563) );
  INV_X1 U9857 ( .A(n8548), .ZN(n8364) );
  NAND2_X1 U9858 ( .A1(n8326), .A2(n8325), .ZN(n8328) );
  NAND2_X1 U9859 ( .A1(n4926), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U9860 ( .A1(n8366), .A2(n8329), .ZN(n8539) );
  INV_X1 U9861 ( .A(n8331), .ZN(n8362) );
  INV_X1 U9862 ( .A(n8332), .ZN(n8519) );
  NAND2_X1 U9863 ( .A1(n8513), .A2(n8512), .ZN(n8751) );
  INV_X1 U9864 ( .A(n8334), .ZN(n8848) );
  INV_X1 U9865 ( .A(n8859), .ZN(n8863) );
  NOR2_X1 U9866 ( .A1(n7200), .A2(n8335), .ZN(n8338) );
  AND4_X1 U9867 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8399), .ZN(n8341)
         );
  NAND4_X1 U9868 ( .A1(n8341), .A2(n8340), .A3(n4279), .A4(n8339), .ZN(n8342)
         );
  NOR2_X1 U9869 ( .A1(n8343), .A2(n8342), .ZN(n8344) );
  NAND3_X1 U9870 ( .A1(n8346), .A2(n8345), .A3(n8344), .ZN(n8347) );
  NOR2_X1 U9871 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  NAND3_X1 U9872 ( .A1(n8462), .A2(n8349), .A3(n8458), .ZN(n8350) );
  NOR2_X1 U9873 ( .A1(n8350), .A2(n8930), .ZN(n8351) );
  NAND4_X1 U9874 ( .A1(n8848), .A2(n8863), .A3(n8351), .A4(n8387), .ZN(n8355)
         );
  INV_X1 U9875 ( .A(n8484), .ZN(n8354) );
  AND2_X1 U9876 ( .A1(n8487), .A2(n8352), .ZN(n8388) );
  INV_X1 U9877 ( .A(n8388), .ZN(n8353) );
  OR3_X1 U9878 ( .A1(n8355), .A2(n8354), .A3(n8353), .ZN(n8356) );
  NOR2_X1 U9879 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  NAND4_X1 U9880 ( .A1(n4290), .A2(n8789), .A3(n8803), .A4(n8358), .ZN(n8359)
         );
  OR2_X1 U9881 ( .A1(n8359), .A2(n8756), .ZN(n8360) );
  NOR2_X1 U9882 ( .A1(n8751), .A2(n8360), .ZN(n8361) );
  NAND4_X1 U9883 ( .A1(n8539), .A2(n5958), .A3(n8362), .A4(n4766), .ZN(n8363)
         );
  NOR4_X1 U9884 ( .A1(n4400), .A2(n8364), .A3(n8542), .A4(n8363), .ZN(n8372)
         );
  INV_X1 U9885 ( .A(n8366), .ZN(n8367) );
  NAND2_X1 U9886 ( .A1(n8543), .A2(n8563), .ZN(n8369) );
  XNOR2_X1 U9887 ( .A(n8374), .B(n8373), .ZN(n8555) );
  NAND2_X1 U9888 ( .A1(n8377), .A2(n8376), .ZN(n8380) );
  INV_X1 U9889 ( .A(n8378), .ZN(n8564) );
  NAND2_X1 U9890 ( .A1(n8380), .A2(n8379), .ZN(n8526) );
  INV_X1 U9891 ( .A(n8526), .ZN(n8527) );
  MUX2_X1 U9892 ( .A(n8529), .B(n8530), .S(n8540), .Z(n8534) );
  NAND2_X1 U9893 ( .A1(n8748), .A2(n8381), .ZN(n8382) );
  MUX2_X1 U9894 ( .A(n8383), .B(n8382), .S(n8540), .Z(n8384) );
  NOR2_X1 U9895 ( .A1(n8384), .A2(n4582), .ZN(n8511) );
  NAND2_X1 U9896 ( .A1(n8502), .A2(n8493), .ZN(n8386) );
  NAND2_X1 U9897 ( .A1(n8501), .A2(n8496), .ZN(n8385) );
  MUX2_X1 U9898 ( .A(n8386), .B(n8385), .S(n8540), .Z(n8505) );
  AND2_X1 U9899 ( .A1(n8484), .A2(n8387), .ZN(n8389) );
  MUX2_X1 U9900 ( .A(n8389), .B(n8388), .S(n8547), .Z(n8483) );
  NAND2_X1 U9901 ( .A1(n8391), .A2(n8390), .ZN(n8392) );
  NAND2_X1 U9902 ( .A1(n8392), .A2(n8395), .ZN(n8394) );
  NAND2_X1 U9903 ( .A1(n8396), .A2(n8540), .ZN(n8393) );
  AOI21_X1 U9904 ( .B1(n8394), .B2(n8400), .A(n8393), .ZN(n8398) );
  AOI21_X1 U9905 ( .B1(n8396), .B2(n8395), .A(n8540), .ZN(n8397) );
  OR2_X1 U9906 ( .A1(n8398), .A2(n8397), .ZN(n8409) );
  OAI21_X1 U9907 ( .B1(n8400), .B2(n8540), .A(n8399), .ZN(n8401) );
  INV_X1 U9908 ( .A(n8401), .ZN(n8408) );
  NAND2_X1 U9909 ( .A1(n8581), .A2(n8402), .ZN(n8403) );
  NAND2_X1 U9910 ( .A1(n8414), .A2(n8403), .ZN(n8406) );
  NAND2_X1 U9911 ( .A1(n8430), .A2(n8404), .ZN(n8405) );
  MUX2_X1 U9912 ( .A(n8406), .B(n8405), .S(n8540), .Z(n8407) );
  AOI21_X1 U9913 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(n8413) );
  NOR2_X1 U9914 ( .A1(n8410), .A2(n10027), .ZN(n8431) );
  INV_X1 U9915 ( .A(n8415), .ZN(n8411) );
  MUX2_X1 U9916 ( .A(n8431), .B(n8411), .S(n8547), .Z(n8412) );
  OR2_X1 U9917 ( .A1(n8413), .A2(n8412), .ZN(n8435) );
  INV_X1 U9918 ( .A(n8414), .ZN(n8416) );
  OAI211_X1 U9919 ( .C1(n8435), .C2(n8416), .A(n8415), .B(n4782), .ZN(n8418)
         );
  NAND2_X1 U9920 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  NAND3_X1 U9921 ( .A1(n8419), .A2(n4279), .A3(n8436), .ZN(n8428) );
  NAND2_X1 U9922 ( .A1(n8421), .A2(n8420), .ZN(n8423) );
  INV_X1 U9923 ( .A(n8422), .ZN(n8441) );
  NAND2_X1 U9924 ( .A1(n8446), .A2(n8441), .ZN(n8425) );
  MUX2_X1 U9925 ( .A(n8423), .B(n8425), .S(n8540), .Z(n8443) );
  OR2_X1 U9926 ( .A1(n8425), .A2(n8424), .ZN(n8426) );
  OAI211_X1 U9927 ( .C1(n8428), .C2(n8443), .A(n8427), .B(n8426), .ZN(n8429)
         );
  INV_X1 U9928 ( .A(n8430), .ZN(n8434) );
  INV_X1 U9929 ( .A(n8431), .ZN(n8433) );
  OAI211_X1 U9930 ( .C1(n8435), .C2(n8434), .A(n8433), .B(n8432), .ZN(n8437)
         );
  NAND3_X1 U9931 ( .A1(n8437), .A2(n8436), .A3(n4782), .ZN(n8439) );
  NAND3_X1 U9932 ( .A1(n8439), .A2(n4279), .A3(n8438), .ZN(n8442) );
  NAND3_X1 U9933 ( .A1(n8442), .A2(n8441), .A3(n8440), .ZN(n8445) );
  INV_X1 U9934 ( .A(n8443), .ZN(n8444) );
  NAND2_X1 U9935 ( .A1(n8445), .A2(n8444), .ZN(n8448) );
  OR2_X1 U9936 ( .A1(n8449), .A2(n8571), .ZN(n8460) );
  INV_X1 U9937 ( .A(n8450), .ZN(n8451) );
  NAND2_X1 U9938 ( .A1(n8452), .A2(n8451), .ZN(n8454) );
  NAND2_X1 U9939 ( .A1(n8454), .A2(n8453), .ZN(n8457) );
  INV_X1 U9940 ( .A(n8455), .ZN(n8456) );
  AOI21_X1 U9941 ( .B1(n8458), .B2(n8457), .A(n8456), .ZN(n8459) );
  MUX2_X1 U9942 ( .A(n8460), .B(n8459), .S(n8547), .Z(n8461) );
  MUX2_X1 U9943 ( .A(n8464), .B(n8463), .S(n8547), .Z(n8465) );
  NAND2_X1 U9944 ( .A1(n8466), .A2(n8465), .ZN(n8467) );
  INV_X1 U9945 ( .A(n8930), .ZN(n8937) );
  NAND2_X1 U9946 ( .A1(n8467), .A2(n8937), .ZN(n8470) );
  NAND3_X1 U9947 ( .A1(n8468), .A2(n8866), .A3(n8540), .ZN(n8469) );
  NAND2_X1 U9948 ( .A1(n8470), .A2(n8469), .ZN(n8477) );
  NAND2_X1 U9949 ( .A1(n8477), .A2(n8863), .ZN(n8472) );
  NAND3_X1 U9950 ( .A1(n8472), .A2(n8480), .A3(n8471), .ZN(n8474) );
  INV_X1 U9951 ( .A(n8475), .ZN(n8476) );
  OAI21_X1 U9952 ( .B1(n8477), .B2(n8476), .A(n8863), .ZN(n8479) );
  NAND2_X1 U9953 ( .A1(n8479), .A2(n8478), .ZN(n8481) );
  AND2_X1 U9954 ( .A1(n8492), .A2(n8484), .ZN(n8486) );
  INV_X1 U9955 ( .A(n8488), .ZN(n8485) );
  AOI21_X1 U9956 ( .B1(n8491), .B2(n8486), .A(n8485), .ZN(n8499) );
  NAND2_X1 U9957 ( .A1(n8488), .A2(n8487), .ZN(n8489) );
  NAND2_X1 U9958 ( .A1(n8489), .A2(n8540), .ZN(n8490) );
  INV_X1 U9959 ( .A(n8490), .ZN(n8498) );
  NAND2_X1 U9960 ( .A1(n8491), .A2(n8490), .ZN(n8494) );
  NAND3_X1 U9961 ( .A1(n8494), .A2(n8493), .A3(n8492), .ZN(n8495) );
  NAND2_X1 U9962 ( .A1(n8495), .A2(n8540), .ZN(n8497) );
  OAI211_X1 U9963 ( .C1(n8499), .C2(n8498), .A(n8497), .B(n8496), .ZN(n8500)
         );
  INV_X1 U9964 ( .A(n8500), .ZN(n8504) );
  MUX2_X1 U9965 ( .A(n8502), .B(n8501), .S(n8547), .Z(n8503) );
  OAI211_X1 U9966 ( .C1(n8505), .C2(n8504), .A(n4290), .B(n8503), .ZN(n8510)
         );
  NAND2_X1 U9967 ( .A1(n8513), .A2(n8506), .ZN(n8508) );
  MUX2_X1 U9968 ( .A(n8508), .B(n8507), .S(n8547), .Z(n8509) );
  MUX2_X1 U9969 ( .A(n8513), .B(n8512), .S(n8540), .Z(n8514) );
  NAND2_X1 U9970 ( .A1(n8732), .A2(n8514), .ZN(n8518) );
  MUX2_X1 U9971 ( .A(n8516), .B(n8515), .S(n8547), .Z(n8517) );
  MUX2_X1 U9972 ( .A(n8520), .B(n8519), .S(n8540), .Z(n8521) );
  MUX2_X1 U9973 ( .A(n8524), .B(n8523), .S(n8547), .Z(n8525) );
  INV_X1 U9974 ( .A(n8531), .ZN(n8532) );
  INV_X1 U9975 ( .A(n8533), .ZN(n8536) );
  INV_X1 U9976 ( .A(n8534), .ZN(n8535) );
  NAND2_X1 U9977 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  NAND2_X1 U9978 ( .A1(n8538), .A2(n8537), .ZN(n8546) );
  INV_X1 U9979 ( .A(n8539), .ZN(n8541) );
  INV_X1 U9980 ( .A(n8549), .ZN(n8550) );
  OAI21_X1 U9981 ( .B1(n8552), .B2(n5819), .A(n8551), .ZN(n8553) );
  NAND3_X1 U9982 ( .A1(n8557), .A2(n8556), .A3(n8072), .ZN(n8558) );
  OAI211_X1 U9983 ( .C1(n8559), .C2(n8561), .A(n8558), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8560) );
  OAI21_X1 U9984 ( .B1(n8562), .B2(n8561), .A(n8560), .ZN(P2_U3296) );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8563), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9986 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8564), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9987 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8565), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8566), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9989 ( .A(n8567), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8687), .Z(
        P2_U3517) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8766), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9991 ( .A(n8780), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8687), .Z(
        P2_U3514) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8792), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8779), .S(P2_U3893), .Z(
        P2_U3512) );
  INV_X1 U9994 ( .A(n8568), .ZN(n8810) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8810), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8569), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8838), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8570), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8837), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n5118), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10001 ( .A(n8933), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8687), .Z(
        P2_U3504) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8571), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10003 ( .A(n8572), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8687), .Z(
        P2_U3502) );
  MUX2_X1 U10004 ( .A(n8573), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8687), .Z(
        P2_U3501) );
  MUX2_X1 U10005 ( .A(n8574), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8687), .Z(
        P2_U3500) );
  MUX2_X1 U10006 ( .A(n8575), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8687), .Z(
        P2_U3499) );
  MUX2_X1 U10007 ( .A(n8576), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8687), .Z(
        P2_U3498) );
  MUX2_X1 U10008 ( .A(n8577), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8687), .Z(
        P2_U3497) );
  MUX2_X1 U10009 ( .A(n8578), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8687), .Z(
        P2_U3496) );
  MUX2_X1 U10010 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8579), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10011 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8580), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10012 ( .A(n8581), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8687), .Z(
        P2_U3493) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8582), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10014 ( .A(n7113), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8687), .Z(
        P2_U3491) );
  OAI21_X1 U10015 ( .B1(n8585), .B2(n8584), .A(n8583), .ZN(n8586) );
  NAND2_X1 U10016 ( .A1(n8586), .A2(n8665), .ZN(n8607) );
  INV_X1 U10017 ( .A(n8587), .ZN(n8591) );
  INV_X1 U10018 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n8589) );
  OAI21_X1 U10019 ( .B1(n8695), .B2(n8589), .A(n8588), .ZN(n8590) );
  AOI21_X1 U10020 ( .B1(n8674), .B2(n8591), .A(n8590), .ZN(n8606) );
  AND3_X1 U10021 ( .A1(n8594), .A2(n8593), .A3(n8592), .ZN(n8595) );
  OAI21_X1 U10022 ( .B1(n8596), .B2(n8595), .A(n8697), .ZN(n8605) );
  INV_X1 U10023 ( .A(n8597), .ZN(n8598) );
  NOR3_X1 U10024 ( .A1(n8600), .A2(n8599), .A3(n8598), .ZN(n8603) );
  OAI21_X1 U10025 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(n8604) );
  NAND4_X1 U10026 ( .A1(n8607), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(
        P2_U3190) );
  AOI21_X1 U10027 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8624) );
  INV_X1 U10028 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9714) );
  OAI21_X1 U10029 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8614) );
  NAND2_X1 U10030 ( .A1(n8665), .A2(n8614), .ZN(n8615) );
  OAI211_X1 U10031 ( .C1(n8695), .C2(n9714), .A(n8616), .B(n8615), .ZN(n8621)
         );
  AOI21_X1 U10032 ( .B1(n4342), .B2(n8618), .A(n8617), .ZN(n8619) );
  NOR2_X1 U10033 ( .A1(n8619), .A2(n8675), .ZN(n8620) );
  AOI211_X1 U10034 ( .C1(n8674), .C2(n8622), .A(n8621), .B(n8620), .ZN(n8623)
         );
  OAI21_X1 U10035 ( .B1(n8624), .B2(n8698), .A(n8623), .ZN(P2_U3196) );
  AOI21_X1 U10036 ( .B1(n8872), .B2(n8626), .A(n8625), .ZN(n8639) );
  OAI21_X1 U10037 ( .B1(n8629), .B2(n8628), .A(n8627), .ZN(n8637) );
  INV_X1 U10038 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9718) );
  INV_X1 U10039 ( .A(n8630), .ZN(n8631) );
  OAI21_X1 U10040 ( .B1(n8695), .B2(n9718), .A(n8631), .ZN(n8636) );
  AOI21_X1 U10041 ( .B1(n8633), .B2(n8923), .A(n8632), .ZN(n8634) );
  OAI22_X1 U10042 ( .A1(n8634), .A2(n8675), .B1(n8686), .B2(n5505), .ZN(n8635)
         );
  AOI211_X1 U10043 ( .C1(n8665), .C2(n8637), .A(n8636), .B(n8635), .ZN(n8638)
         );
  OAI21_X1 U10044 ( .B1(n8639), .B2(n8698), .A(n8638), .ZN(P2_U3197) );
  INV_X1 U10045 ( .A(n8640), .ZN(n8641) );
  AOI21_X1 U10046 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n8659) );
  INV_X1 U10047 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9722) );
  INV_X1 U10048 ( .A(n8644), .ZN(n8650) );
  OAI21_X1 U10049 ( .B1(n8647), .B2(n8646), .A(n8645), .ZN(n8648) );
  NAND2_X1 U10050 ( .A1(n8665), .A2(n8648), .ZN(n8649) );
  OAI211_X1 U10051 ( .C1(n8695), .C2(n9722), .A(n8650), .B(n8649), .ZN(n8656)
         );
  NAND2_X1 U10052 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  AOI21_X1 U10053 ( .B1(n8654), .B2(n8653), .A(n8675), .ZN(n8655) );
  AOI211_X1 U10054 ( .C1(n8674), .C2(n8657), .A(n8656), .B(n8655), .ZN(n8658)
         );
  OAI21_X1 U10055 ( .B1(n8659), .B2(n8698), .A(n8658), .ZN(P2_U3198) );
  AOI21_X1 U10056 ( .B1(n8661), .B2(n8917), .A(n8660), .ZN(n8676) );
  INV_X1 U10057 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9726) );
  OAI21_X1 U10058 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8666) );
  NAND2_X1 U10059 ( .A1(n8666), .A2(n8665), .ZN(n8668) );
  OAI211_X1 U10060 ( .C1(n9726), .C2(n8695), .A(n8668), .B(n8667), .ZN(n8672)
         );
  AOI21_X1 U10061 ( .B1(n8679), .B2(n8678), .A(n8677), .ZN(n8699) );
  NOR2_X1 U10062 ( .A1(n8685), .A2(n8684), .ZN(n8690) );
  INV_X1 U10063 ( .A(n8690), .ZN(n8688) );
  OAI21_X1 U10064 ( .B1(n8688), .B2(n8687), .A(n8686), .ZN(n8693) );
  NOR2_X1 U10065 ( .A1(n8690), .A2(n8689), .ZN(n8692) );
  INV_X1 U10066 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10069) );
  OAI21_X1 U10067 ( .B1(n8695), .B2(n10069), .A(n8694), .ZN(n8696) );
  OR2_X1 U10068 ( .A1(n8701), .A2(n8700), .ZN(n8946) );
  OAI21_X1 U10069 ( .B1(n10034), .B2(n8946), .A(n8702), .ZN(n8704) );
  AOI21_X1 U10070 ( .B1(n10034), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8704), .ZN(
        n8703) );
  OAI21_X1 U10071 ( .B1(n8884), .B2(n10020), .A(n8703), .ZN(P2_U3202) );
  AOI21_X1 U10072 ( .B1(n10034), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8704), .ZN(
        n8705) );
  OAI21_X1 U10073 ( .B1(n8367), .B2(n10020), .A(n8705), .ZN(P2_U3203) );
  NAND2_X1 U10074 ( .A1(n8706), .A2(n4275), .ZN(n8713) );
  INV_X1 U10075 ( .A(n8707), .ZN(n8709) );
  OAI22_X1 U10076 ( .A1(n8709), .A2(n10017), .B1(n4275), .B2(n8708), .ZN(n8710) );
  AOI21_X1 U10077 ( .B1(n8711), .B2(n10026), .A(n8710), .ZN(n8712) );
  OAI211_X1 U10078 ( .C1(n8714), .C2(n10025), .A(n8713), .B(n8712), .ZN(
        P2_U3206) );
  XOR2_X1 U10079 ( .A(n8719), .B(n8715), .Z(n8957) );
  INV_X1 U10080 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U10081 ( .A1(n8731), .A2(n8716), .ZN(n8718) );
  INV_X1 U10082 ( .A(n8887), .ZN(n8952) );
  MUX2_X1 U10083 ( .A(n8725), .B(n8952), .S(n4275), .Z(n8728) );
  AOI22_X1 U10084 ( .A1(n8954), .A2(n10026), .B1(n10028), .B2(n8726), .ZN(
        n8727) );
  OAI211_X1 U10085 ( .C1(n8957), .C2(n10025), .A(n8728), .B(n8727), .ZN(
        P2_U3207) );
  XNOR2_X1 U10086 ( .A(n8729), .B(n8732), .ZN(n8960) );
  NAND2_X1 U10087 ( .A1(n8731), .A2(n8730), .ZN(n8733) );
  XNOR2_X1 U10088 ( .A(n8733), .B(n8732), .ZN(n8734) );
  OAI222_X1 U10089 ( .A1(n8867), .A2(n8736), .B1(n8865), .B2(n8735), .C1(n8862), .C2(n8734), .ZN(n8958) );
  NOR2_X1 U10090 ( .A1(n8959), .A2(n9738), .ZN(n8737) );
  OAI21_X1 U10091 ( .B1(n8958), .B2(n8737), .A(n4275), .ZN(n8740) );
  AOI22_X1 U10092 ( .A1(n8738), .A2(n10028), .B1(n10034), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8739) );
  OAI211_X1 U10093 ( .C1(n8960), .C2(n10025), .A(n8740), .B(n8739), .ZN(
        P2_U3208) );
  XOR2_X1 U10094 ( .A(n8751), .B(n8741), .Z(n8742) );
  OAI222_X1 U10095 ( .A1(n8867), .A2(n8744), .B1(n8865), .B2(n8743), .C1(n8862), .C2(n8742), .ZN(n8963) );
  INV_X1 U10096 ( .A(n8745), .ZN(n8746) );
  OAI22_X1 U10097 ( .A1(n8964), .A2(n9738), .B1(n8746), .B2(n10017), .ZN(n8747) );
  OAI21_X1 U10098 ( .B1(n8963), .B2(n8747), .A(n4275), .ZN(n8754) );
  INV_X1 U10099 ( .A(n8748), .ZN(n8749) );
  OR2_X1 U10100 ( .A1(n8965), .A2(n10025), .ZN(n8753) );
  OAI211_X1 U10101 ( .C1(n4275), .C2(n8755), .A(n8754), .B(n8753), .ZN(
        P2_U3209) );
  XNOR2_X1 U10102 ( .A(n8757), .B(n8756), .ZN(n8973) );
  OR2_X1 U10103 ( .A1(n8758), .A2(n8759), .ZN(n8761) );
  NAND3_X1 U10104 ( .A1(n8778), .A2(n8763), .A3(n8762), .ZN(n8764) );
  NAND2_X1 U10105 ( .A1(n8765), .A2(n8764), .ZN(n8767) );
  AOI222_X1 U10106 ( .A1(n8928), .A2(n8767), .B1(n8766), .B2(n8932), .C1(n8792), .C2(n8934), .ZN(n8968) );
  MUX2_X1 U10107 ( .A(n8768), .B(n8968), .S(n4275), .Z(n8771) );
  AOI22_X1 U10108 ( .A1(n8970), .A2(n10026), .B1(n10028), .B2(n8769), .ZN(
        n8770) );
  OAI211_X1 U10109 ( .C1(n8973), .C2(n10025), .A(n8771), .B(n8770), .ZN(
        P2_U3210) );
  XNOR2_X1 U10110 ( .A(n8772), .B(n4290), .ZN(n8979) );
  INV_X1 U10111 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8782) );
  OR2_X1 U10112 ( .A1(n8758), .A2(n8773), .ZN(n8775) );
  NAND3_X1 U10113 ( .A1(n8791), .A2(n4290), .A3(n8776), .ZN(n8777) );
  NAND2_X1 U10114 ( .A1(n8778), .A2(n8777), .ZN(n8781) );
  AOI222_X1 U10115 ( .A1(n8928), .A2(n8781), .B1(n8780), .B2(n8932), .C1(n8779), .C2(n8934), .ZN(n8974) );
  MUX2_X1 U10116 ( .A(n8782), .B(n8974), .S(n4275), .Z(n8785) );
  AOI22_X1 U10117 ( .A1(n8976), .A2(n10026), .B1(n10028), .B2(n8783), .ZN(
        n8784) );
  OAI211_X1 U10118 ( .C1(n8979), .C2(n10025), .A(n8785), .B(n8784), .ZN(
        P2_U3211) );
  XNOR2_X1 U10119 ( .A(n8787), .B(n8786), .ZN(n8985) );
  OR2_X1 U10120 ( .A1(n8758), .A2(n8803), .ZN(n8798) );
  NAND3_X1 U10121 ( .A1(n8798), .A2(n8789), .A3(n8788), .ZN(n8790) );
  NAND2_X1 U10122 ( .A1(n8791), .A2(n8790), .ZN(n8793) );
  AOI222_X1 U10123 ( .A1(n8928), .A2(n8793), .B1(n8792), .B2(n8932), .C1(n8810), .C2(n8934), .ZN(n8980) );
  MUX2_X1 U10124 ( .A(n8794), .B(n8980), .S(n4275), .Z(n8797) );
  AOI22_X1 U10125 ( .A1(n8982), .A2(n10026), .B1(n10028), .B2(n8795), .ZN(
        n8796) );
  OAI211_X1 U10126 ( .C1(n8985), .C2(n10025), .A(n8797), .B(n8796), .ZN(
        P2_U3212) );
  INV_X1 U10127 ( .A(n8798), .ZN(n8799) );
  AOI21_X1 U10128 ( .B1(n8803), .B2(n8758), .A(n8799), .ZN(n8800) );
  OAI222_X1 U10129 ( .A1(n8867), .A2(n8801), .B1(n8865), .B2(n8826), .C1(n8862), .C2(n8800), .ZN(n8903) );
  AOI21_X1 U10130 ( .B1(n10028), .B2(n8802), .A(n8903), .ZN(n8808) );
  XOR2_X1 U10131 ( .A(n8804), .B(n8803), .Z(n8904) );
  OAI22_X1 U10132 ( .A1(n8990), .A2(n10020), .B1(n4275), .B2(n8805), .ZN(n8806) );
  AOI21_X1 U10133 ( .B1(n8904), .B2(n10030), .A(n8806), .ZN(n8807) );
  OAI21_X1 U10134 ( .B1(n8808), .B2(n10034), .A(n8807), .ZN(P2_U3213) );
  XNOR2_X1 U10135 ( .A(n8809), .B(n8816), .ZN(n8811) );
  AOI222_X1 U10136 ( .A1(n8928), .A2(n8811), .B1(n8810), .B2(n8932), .C1(n8838), .C2(n8934), .ZN(n8911) );
  INV_X1 U10137 ( .A(n8812), .ZN(n8813) );
  OAI22_X1 U10138 ( .A1(n4275), .A2(n8814), .B1(n8813), .B2(n10017), .ZN(n8819) );
  OAI21_X1 U10139 ( .B1(n8817), .B2(n8816), .A(n8815), .ZN(n8912) );
  NOR2_X1 U10140 ( .A1(n8912), .A2(n10025), .ZN(n8818) );
  AOI211_X1 U10141 ( .C1(n10026), .C2(n8909), .A(n8819), .B(n8818), .ZN(n8820)
         );
  OAI21_X1 U10142 ( .B1(n8911), .B2(n10034), .A(n8820), .ZN(P2_U3214) );
  OAI21_X1 U10143 ( .B1(n8822), .B2(n5428), .A(n8821), .ZN(n8995) );
  XNOR2_X1 U10144 ( .A(n8823), .B(n8824), .ZN(n8825) );
  OAI222_X1 U10145 ( .A1(n8867), .A2(n8826), .B1(n8865), .B2(n8851), .C1(n8825), .C2(n8862), .ZN(n8913) );
  NAND2_X1 U10146 ( .A1(n8913), .A2(n4275), .ZN(n8832) );
  INV_X1 U10147 ( .A(n8827), .ZN(n8828) );
  OAI22_X1 U10148 ( .A1(n4275), .A2(n8829), .B1(n8828), .B2(n10017), .ZN(n8830) );
  AOI21_X1 U10149 ( .B1(n8914), .B2(n10026), .A(n8830), .ZN(n8831) );
  OAI211_X1 U10150 ( .C1(n8995), .C2(n10025), .A(n8832), .B(n8831), .ZN(
        P2_U3215) );
  XNOR2_X1 U10151 ( .A(n8833), .B(n8835), .ZN(n9001) );
  OAI211_X1 U10152 ( .C1(n8836), .C2(n8835), .A(n8834), .B(n8928), .ZN(n8840)
         );
  AOI22_X1 U10153 ( .A1(n8838), .A2(n8932), .B1(n8837), .B2(n8934), .ZN(n8839)
         );
  MUX2_X1 U10154 ( .A(n8671), .B(n8996), .S(n4275), .Z(n8843) );
  AOI22_X1 U10155 ( .A1(n8998), .A2(n10026), .B1(n10028), .B2(n8841), .ZN(
        n8842) );
  OAI211_X1 U10156 ( .C1(n9001), .C2(n10025), .A(n8843), .B(n8842), .ZN(
        P2_U3216) );
  NAND2_X1 U10157 ( .A1(n8844), .A2(n8845), .ZN(n8846) );
  XNOR2_X1 U10158 ( .A(n8846), .B(n8848), .ZN(n9007) );
  INV_X1 U10159 ( .A(n8847), .ZN(n8849) );
  AOI21_X1 U10160 ( .B1(n8849), .B2(n8848), .A(n8862), .ZN(n8854) );
  OAI22_X1 U10161 ( .A1(n8851), .A2(n8867), .B1(n8850), .B2(n8865), .ZN(n8852)
         );
  AOI21_X1 U10162 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n9002) );
  MUX2_X1 U10163 ( .A(n8855), .B(n9002), .S(n4275), .Z(n8858) );
  AOI22_X1 U10164 ( .A1(n9004), .A2(n10026), .B1(n10028), .B2(n8856), .ZN(
        n8857) );
  OAI211_X1 U10165 ( .C1(n9007), .C2(n10025), .A(n8858), .B(n8857), .ZN(
        P2_U3217) );
  XNOR2_X1 U10166 ( .A(n8860), .B(n8859), .ZN(n9015) );
  INV_X1 U10167 ( .A(n8861), .ZN(n8864) );
  AOI21_X1 U10168 ( .B1(n8864), .B2(n8863), .A(n8862), .ZN(n8871) );
  OAI22_X1 U10169 ( .A1(n8868), .A2(n8867), .B1(n8866), .B2(n8865), .ZN(n8869)
         );
  AOI21_X1 U10170 ( .B1(n8871), .B2(n8870), .A(n8869), .ZN(n9008) );
  MUX2_X1 U10171 ( .A(n8872), .B(n9008), .S(n4275), .Z(n8875) );
  AOI22_X1 U10172 ( .A1(n9011), .A2(n10026), .B1(n10028), .B2(n8873), .ZN(
        n8874) );
  OAI211_X1 U10173 ( .C1(n9015), .C2(n10025), .A(n8875), .B(n8874), .ZN(
        P2_U3218) );
  OAI22_X1 U10174 ( .A1(n8877), .A2(n9738), .B1(n8876), .B2(n10017), .ZN(n8878) );
  OAI21_X1 U10175 ( .B1(n8879), .B2(n8878), .A(n4275), .ZN(n8881) );
  NAND2_X1 U10176 ( .A1(n10034), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8880) );
  OAI211_X1 U10177 ( .C1(n8882), .C2(n10025), .A(n8881), .B(n8880), .ZN(
        P2_U3220) );
  NOR2_X1 U10178 ( .A1(n8946), .A2(n8944), .ZN(n8885) );
  AOI21_X1 U10179 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n8944), .A(n8885), .ZN(
        n8883) );
  OAI21_X1 U10180 ( .B1(n8884), .B2(n8908), .A(n8883), .ZN(P2_U3490) );
  AOI21_X1 U10181 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n8944), .A(n8885), .ZN(
        n8886) );
  OAI21_X1 U10182 ( .B1(n8367), .B2(n8908), .A(n8886), .ZN(P2_U3489) );
  MUX2_X1 U10183 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8887), .S(n8942), .Z(n8890) );
  INV_X1 U10184 ( .A(n8954), .ZN(n8888) );
  OAI22_X1 U10185 ( .A1(n8957), .A2(n8927), .B1(n8888), .B2(n8908), .ZN(n8889)
         );
  OR2_X1 U10186 ( .A1(n8890), .A2(n8889), .ZN(P2_U3485) );
  MUX2_X1 U10187 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8958), .S(n8942), .Z(n8892) );
  OAI22_X1 U10188 ( .A1(n8960), .A2(n8927), .B1(n8959), .B2(n8908), .ZN(n8891)
         );
  OR2_X1 U10189 ( .A1(n8892), .A2(n8891), .ZN(P2_U3484) );
  MUX2_X1 U10190 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8963), .S(n8942), .Z(n8894) );
  OAI22_X1 U10191 ( .A1(n8965), .A2(n8927), .B1(n8964), .B2(n8908), .ZN(n8893)
         );
  OR2_X1 U10192 ( .A1(n8894), .A2(n8893), .ZN(P2_U3483) );
  INV_X1 U10193 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U10194 ( .A(n8895), .B(n8968), .S(n8942), .Z(n8897) );
  INV_X1 U10195 ( .A(n8908), .ZN(n8924) );
  NAND2_X1 U10196 ( .A1(n8970), .A2(n8924), .ZN(n8896) );
  OAI211_X1 U10197 ( .C1(n8973), .C2(n8927), .A(n8897), .B(n8896), .ZN(
        P2_U3482) );
  MUX2_X1 U10198 ( .A(n9534), .B(n8974), .S(n8942), .Z(n8899) );
  NAND2_X1 U10199 ( .A1(n8976), .A2(n8924), .ZN(n8898) );
  OAI211_X1 U10200 ( .C1(n8979), .C2(n8927), .A(n8899), .B(n8898), .ZN(
        P2_U3481) );
  INV_X1 U10201 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U10202 ( .A(n8900), .B(n8980), .S(n8942), .Z(n8902) );
  NAND2_X1 U10203 ( .A1(n8982), .A2(n8924), .ZN(n8901) );
  OAI211_X1 U10204 ( .C1(n8927), .C2(n8985), .A(n8902), .B(n8901), .ZN(
        P2_U3480) );
  INV_X1 U10205 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8906) );
  AOI21_X1 U10206 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8986) );
  MUX2_X1 U10207 ( .A(n8906), .B(n8986), .S(n8942), .Z(n8907) );
  OAI21_X1 U10208 ( .B1(n8990), .B2(n8908), .A(n8907), .ZN(P2_U3479) );
  NAND2_X1 U10209 ( .A1(n8909), .A2(n8915), .ZN(n8910) );
  OAI211_X1 U10210 ( .C1(n8940), .C2(n8912), .A(n8911), .B(n8910), .ZN(n8991)
         );
  MUX2_X1 U10211 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8991), .S(n8942), .Z(
        P2_U3478) );
  INV_X1 U10212 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9602) );
  AOI21_X1 U10213 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n8992) );
  MUX2_X1 U10214 ( .A(n9602), .B(n8992), .S(n8942), .Z(n8916) );
  OAI21_X1 U10215 ( .B1(n8927), .B2(n8995), .A(n8916), .ZN(P2_U3477) );
  MUX2_X1 U10216 ( .A(n8917), .B(n8996), .S(n8942), .Z(n8919) );
  NAND2_X1 U10217 ( .A1(n8998), .A2(n8924), .ZN(n8918) );
  OAI211_X1 U10218 ( .C1(n8927), .C2(n9001), .A(n8919), .B(n8918), .ZN(
        P2_U3476) );
  MUX2_X1 U10219 ( .A(n8920), .B(n9002), .S(n8942), .Z(n8922) );
  NAND2_X1 U10220 ( .A1(n9004), .A2(n8924), .ZN(n8921) );
  OAI211_X1 U10221 ( .C1(n9007), .C2(n8927), .A(n8922), .B(n8921), .ZN(
        P2_U3475) );
  MUX2_X1 U10222 ( .A(n8923), .B(n9008), .S(n8942), .Z(n8926) );
  NAND2_X1 U10223 ( .A1(n9011), .A2(n8924), .ZN(n8925) );
  OAI211_X1 U10224 ( .C1(n8927), .C2(n9015), .A(n8926), .B(n8925), .ZN(
        P2_U3474) );
  OAI211_X1 U10225 ( .C1(n8931), .C2(n8930), .A(n8929), .B(n8928), .ZN(n8936)
         );
  AOI22_X1 U10226 ( .A1(n8934), .A2(n8933), .B1(n5118), .B2(n8932), .ZN(n8935)
         );
  NAND2_X1 U10227 ( .A1(n8936), .A2(n8935), .ZN(n9741) );
  XNOR2_X1 U10228 ( .A(n8938), .B(n8937), .ZN(n9734) );
  OAI22_X1 U10229 ( .A1(n9734), .A2(n8940), .B1(n9739), .B2(n8939), .ZN(n8941)
         );
  NOR2_X1 U10230 ( .A1(n9741), .A2(n8941), .ZN(n9744) );
  OR2_X1 U10231 ( .A1(n8942), .A2(n5095), .ZN(n8943) );
  OAI21_X1 U10232 ( .B1(n9744), .B2(n8944), .A(n8943), .ZN(P2_U3473) );
  INV_X1 U10233 ( .A(n8989), .ZN(n9010) );
  NAND2_X1 U10234 ( .A1(n8945), .A2(n9010), .ZN(n8948) );
  INV_X1 U10235 ( .A(n8946), .ZN(n8947) );
  NAND2_X1 U10236 ( .A1(n8947), .A2(n10057), .ZN(n8949) );
  OAI211_X1 U10237 ( .C1(n8317), .C2(n10057), .A(n8948), .B(n8949), .ZN(
        P2_U3458) );
  INV_X1 U10238 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U10239 ( .A1(n8366), .A2(n9010), .ZN(n8950) );
  OAI211_X1 U10240 ( .C1(n8951), .C2(n10057), .A(n8950), .B(n8949), .ZN(
        P2_U3457) );
  MUX2_X1 U10241 ( .A(n8953), .B(n8952), .S(n10057), .Z(n8956) );
  NAND2_X1 U10242 ( .A1(n8954), .A2(n9010), .ZN(n8955) );
  OAI211_X1 U10243 ( .C1(n8957), .C2(n9014), .A(n8956), .B(n8955), .ZN(
        P2_U3453) );
  MUX2_X1 U10244 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8958), .S(n10057), .Z(
        n8962) );
  OAI22_X1 U10245 ( .A1(n8960), .A2(n9014), .B1(n8959), .B2(n8989), .ZN(n8961)
         );
  OR2_X1 U10246 ( .A1(n8962), .A2(n8961), .ZN(P2_U3452) );
  MUX2_X1 U10247 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8963), .S(n10057), .Z(
        n8967) );
  OAI22_X1 U10248 ( .A1(n8965), .A2(n9014), .B1(n8964), .B2(n8989), .ZN(n8966)
         );
  OR2_X1 U10249 ( .A1(n8967), .A2(n8966), .ZN(P2_U3451) );
  INV_X1 U10250 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8969) );
  MUX2_X1 U10251 ( .A(n8969), .B(n8968), .S(n10057), .Z(n8972) );
  NAND2_X1 U10252 ( .A1(n8970), .A2(n9010), .ZN(n8971) );
  OAI211_X1 U10253 ( .C1(n8973), .C2(n9014), .A(n8972), .B(n8971), .ZN(
        P2_U3450) );
  INV_X1 U10254 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8975) );
  MUX2_X1 U10255 ( .A(n8975), .B(n8974), .S(n10057), .Z(n8978) );
  NAND2_X1 U10256 ( .A1(n8976), .A2(n9010), .ZN(n8977) );
  OAI211_X1 U10257 ( .C1(n8979), .C2(n9014), .A(n8978), .B(n8977), .ZN(
        P2_U3449) );
  INV_X1 U10258 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U10259 ( .A(n8981), .B(n8980), .S(n10057), .Z(n8984) );
  NAND2_X1 U10260 ( .A1(n8982), .A2(n9010), .ZN(n8983) );
  OAI211_X1 U10261 ( .C1(n8985), .C2(n9014), .A(n8984), .B(n8983), .ZN(
        P2_U3448) );
  INV_X1 U10262 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8987) );
  MUX2_X1 U10263 ( .A(n8987), .B(n8986), .S(n10057), .Z(n8988) );
  OAI21_X1 U10264 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(P2_U3447) );
  MUX2_X1 U10265 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8991), .S(n10057), .Z(
        P2_U3446) );
  INV_X1 U10266 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8993) );
  MUX2_X1 U10267 ( .A(n8993), .B(n8992), .S(n10057), .Z(n8994) );
  OAI21_X1 U10268 ( .B1(n8995), .B2(n9014), .A(n8994), .ZN(P2_U3444) );
  INV_X1 U10269 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8997) );
  MUX2_X1 U10270 ( .A(n8997), .B(n8996), .S(n10057), .Z(n9000) );
  NAND2_X1 U10271 ( .A1(n8998), .A2(n9010), .ZN(n8999) );
  OAI211_X1 U10272 ( .C1(n9001), .C2(n9014), .A(n9000), .B(n8999), .ZN(
        P2_U3441) );
  INV_X1 U10273 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U10274 ( .A(n9003), .B(n9002), .S(n10057), .Z(n9006) );
  NAND2_X1 U10275 ( .A1(n9004), .A2(n9010), .ZN(n9005) );
  OAI211_X1 U10276 ( .C1(n9007), .C2(n9014), .A(n9006), .B(n9005), .ZN(
        P2_U3438) );
  MUX2_X1 U10277 ( .A(n9009), .B(n9008), .S(n10057), .Z(n9013) );
  NAND2_X1 U10278 ( .A1(n9011), .A2(n9010), .ZN(n9012) );
  OAI211_X1 U10279 ( .C1(n9015), .C2(n9014), .A(n9013), .B(n9012), .ZN(
        P2_U3435) );
  INV_X1 U10280 ( .A(n9016), .ZN(n9676) );
  NAND3_X1 U10281 ( .A1(n9017), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9018) );
  OAI22_X1 U10282 ( .A1(n4806), .A2(n9018), .B1(n6509), .B2(n9021), .ZN(n9019)
         );
  INV_X1 U10283 ( .A(n9019), .ZN(n9020) );
  OAI21_X1 U10284 ( .B1(n9676), .B2(n9024), .A(n9020), .ZN(P2_U3264) );
  OAI222_X1 U10285 ( .A1(n4809), .A2(P2_U3151), .B1(n9024), .B2(n9023), .C1(
        n9022), .C2(n9021), .ZN(P2_U3265) );
  NAND2_X1 U10286 ( .A1(n4743), .A2(n9026), .ZN(n9028) );
  XNOR2_X1 U10287 ( .A(n9028), .B(n9027), .ZN(n9035) );
  AOI22_X1 U10288 ( .A1(n9029), .A2(n9753), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n9030) );
  OAI21_X1 U10289 ( .B1(n9760), .B2(n9031), .A(n9030), .ZN(n9032) );
  AOI21_X1 U10290 ( .B1(n9033), .B2(n9141), .A(n9032), .ZN(n9034) );
  OAI21_X1 U10291 ( .B1(n9035), .B2(n9755), .A(n9034), .ZN(P1_U3215) );
  AOI21_X1 U10292 ( .B1(n9041), .B2(n9040), .A(n9039), .ZN(n9042) );
  NAND2_X1 U10293 ( .A1(n9156), .A2(n9086), .ZN(n9045) );
  OR2_X1 U10294 ( .A1(n9053), .A2(n9117), .ZN(n9044) );
  NAND2_X1 U10295 ( .A1(n9045), .A2(n9044), .ZN(n9340) );
  AOI22_X1 U10296 ( .A1(n9340), .A2(n9753), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9046) );
  OAI21_X1 U10297 ( .B1(n9760), .B2(n9047), .A(n9046), .ZN(n9048) );
  AOI21_X1 U10298 ( .B1(n9463), .B2(n9141), .A(n9048), .ZN(n9049) );
  OAI21_X1 U10299 ( .B1(n9050), .B2(n9755), .A(n9049), .ZN(P1_U3216) );
  XOR2_X1 U10300 ( .A(n9052), .B(n9051), .Z(n9059) );
  OR2_X1 U10301 ( .A1(n9053), .A2(n9129), .ZN(n9055) );
  NAND2_X1 U10302 ( .A1(n9160), .A2(n9131), .ZN(n9054) );
  NAND2_X1 U10303 ( .A1(n9055), .A2(n9054), .ZN(n9369) );
  AOI22_X1 U10304 ( .A1(n9369), .A2(n9753), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9056) );
  OAI21_X1 U10305 ( .B1(n9760), .B2(n9376), .A(n9056), .ZN(n9057) );
  AOI21_X1 U10306 ( .B1(n9375), .B2(n9141), .A(n9057), .ZN(n9058) );
  OAI21_X1 U10307 ( .B1(n9059), .B2(n9755), .A(n9058), .ZN(P1_U3223) );
  NAND2_X1 U10308 ( .A1(n9060), .A2(n9061), .ZN(n9062) );
  NAND2_X1 U10309 ( .A1(n9062), .A2(n9063), .ZN(n9072) );
  OAI21_X1 U10310 ( .B1(n9063), .B2(n9062), .A(n9072), .ZN(n9064) );
  NAND2_X1 U10311 ( .A1(n9064), .A2(n9148), .ZN(n9070) );
  NOR2_X1 U10312 ( .A1(n9065), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9195) );
  NOR2_X1 U10313 ( .A1(n9760), .A2(n9066), .ZN(n9067) );
  AOI211_X1 U10314 ( .C1(n9753), .C2(n9068), .A(n9195), .B(n9067), .ZN(n9069)
         );
  OAI211_X1 U10315 ( .C1(n9668), .C2(n9749), .A(n9070), .B(n9069), .ZN(
        P1_U3226) );
  NAND2_X1 U10316 ( .A1(n9072), .A2(n9071), .ZN(n9074) );
  OAI21_X1 U10317 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9076) );
  NAND2_X1 U10318 ( .A1(n9076), .A2(n9148), .ZN(n9081) );
  AND2_X1 U10319 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9209) );
  NOR2_X1 U10320 ( .A1(n9760), .A2(n9077), .ZN(n9078) );
  AOI211_X1 U10321 ( .C1(n9753), .C2(n9079), .A(n9209), .B(n9078), .ZN(n9080)
         );
  OAI211_X1 U10322 ( .C1(n9082), .C2(n9749), .A(n9081), .B(n9080), .ZN(
        P1_U3228) );
  OAI21_X1 U10323 ( .B1(n9084), .B2(n6460), .A(n9083), .ZN(n9085) );
  NAND2_X1 U10324 ( .A1(n9085), .A2(n9148), .ZN(n9093) );
  NAND2_X1 U10325 ( .A1(n9155), .A2(n9086), .ZN(n9088) );
  NAND2_X1 U10326 ( .A1(n9157), .A2(n9131), .ZN(n9087) );
  AND2_X1 U10327 ( .A1(n9088), .A2(n9087), .ZN(n9323) );
  OAI22_X1 U10328 ( .A1(n9323), .A2(n9090), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9089), .ZN(n9091) );
  AOI21_X1 U10329 ( .B1(n9327), .B2(n9097), .A(n9091), .ZN(n9092) );
  OAI211_X1 U10330 ( .C1(n9644), .C2(n9749), .A(n9093), .B(n9092), .ZN(
        P1_U3229) );
  OAI21_X1 U10331 ( .B1(n9096), .B2(n9094), .A(n9095), .ZN(n9101) );
  OAI22_X1 U10332 ( .A1(n9106), .A2(n9129), .B1(n9119), .B2(n9117), .ZN(n9386)
         );
  AOI22_X1 U10333 ( .A1(n9386), .A2(n9753), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9099) );
  NAND2_X1 U10334 ( .A1(n9097), .A2(n9392), .ZN(n9098) );
  OAI211_X1 U10335 ( .C1(n9657), .C2(n9749), .A(n9099), .B(n9098), .ZN(n9100)
         );
  AOI21_X1 U10336 ( .B1(n9101), .B2(n9148), .A(n9100), .ZN(n9102) );
  INV_X1 U10337 ( .A(n9102), .ZN(P1_U3233) );
  AOI21_X1 U10338 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9112) );
  INV_X1 U10339 ( .A(n9357), .ZN(n9109) );
  OAI22_X1 U10340 ( .A1(n9107), .A2(n9129), .B1(n9106), .B2(n9117), .ZN(n9351)
         );
  AOI22_X1 U10341 ( .A1(n9351), .A2(n9753), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9108) );
  OAI21_X1 U10342 ( .B1(n9135), .B2(n9109), .A(n9108), .ZN(n9110) );
  AOI21_X1 U10343 ( .B1(n9356), .B2(n9141), .A(n9110), .ZN(n9111) );
  OAI21_X1 U10344 ( .B1(n9112), .B2(n9755), .A(n9111), .ZN(P1_U3235) );
  NAND2_X1 U10345 ( .A1(n9113), .A2(n9114), .ZN(n9116) );
  XNOR2_X1 U10346 ( .A(n9116), .B(n9115), .ZN(n9123) );
  OAI22_X1 U10347 ( .A1(n9119), .A2(n9129), .B1(n9118), .B2(n9117), .ZN(n9417)
         );
  AOI22_X1 U10348 ( .A1(n9417), .A2(n9753), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9120) );
  OAI21_X1 U10349 ( .B1(n9135), .B2(n9428), .A(n9120), .ZN(n9121) );
  AOI21_X1 U10350 ( .B1(n9426), .B2(n9141), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10351 ( .B1(n9123), .B2(n9755), .A(n9122), .ZN(P1_U3238) );
  AND2_X1 U10352 ( .A1(n9125), .A2(n9124), .ZN(n9128) );
  OAI211_X1 U10353 ( .C1(n9128), .C2(n9127), .A(n9126), .B(n9148), .ZN(n9138)
         );
  OR2_X1 U10354 ( .A1(n9130), .A2(n9129), .ZN(n9133) );
  NAND2_X1 U10355 ( .A1(n9155), .A2(n9131), .ZN(n9132) );
  NAND2_X1 U10356 ( .A1(n9133), .A2(n9132), .ZN(n9289) );
  OAI22_X1 U10357 ( .A1(n9135), .A2(n9294), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9134), .ZN(n9136) );
  AOI21_X1 U10358 ( .B1(n9289), .B2(n9753), .A(n9136), .ZN(n9137) );
  OAI211_X1 U10359 ( .C1(n9639), .C2(n9749), .A(n9138), .B(n9137), .ZN(
        P1_U3240) );
  OAI21_X1 U10360 ( .B1(n9139), .B2(n9140), .A(n9060), .ZN(n9149) );
  NAND2_X1 U10361 ( .A1(n9142), .A2(n9141), .ZN(n9145) );
  AOI22_X1 U10362 ( .A1(n9143), .A2(n9753), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9144) );
  OAI211_X1 U10363 ( .C1(n9760), .C2(n9146), .A(n9145), .B(n9144), .ZN(n9147)
         );
  AOI21_X1 U10364 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(n9150) );
  INV_X1 U10365 ( .A(n9150), .ZN(P1_U3241) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9151), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9152), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9153), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10369 ( .A(n9154), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9177), .Z(
        P1_U3580) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9155), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10371 ( .A(n9156), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9177), .Z(
        P1_U3578) );
  MUX2_X1 U10372 ( .A(n9157), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9177), .Z(
        P1_U3577) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9158), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10374 ( .A(n9159), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9177), .Z(
        P1_U3575) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9160), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9161), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9162), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9163), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n6096), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9164), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10381 ( .A(n9165), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9177), .Z(
        P1_U3567) );
  MUX2_X1 U10382 ( .A(n9166), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9177), .Z(
        P1_U3566) );
  MUX2_X1 U10383 ( .A(n9167), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9177), .Z(
        P1_U3565) );
  MUX2_X1 U10384 ( .A(n9168), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9177), .Z(
        P1_U3564) );
  MUX2_X1 U10385 ( .A(n9169), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9177), .Z(
        P1_U3563) );
  MUX2_X1 U10386 ( .A(n9170), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9177), .Z(
        P1_U3562) );
  MUX2_X1 U10387 ( .A(n9171), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9177), .Z(
        P1_U3561) );
  MUX2_X1 U10388 ( .A(n9172), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9177), .Z(
        P1_U3560) );
  MUX2_X1 U10389 ( .A(n9173), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9177), .Z(
        P1_U3559) );
  MUX2_X1 U10390 ( .A(n9174), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9177), .Z(
        P1_U3558) );
  MUX2_X1 U10391 ( .A(n9175), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9177), .Z(
        P1_U3557) );
  MUX2_X1 U10392 ( .A(n9176), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9177), .Z(
        P1_U3556) );
  MUX2_X1 U10393 ( .A(n6268), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9177), .Z(
        P1_U3555) );
  MUX2_X1 U10394 ( .A(n6275), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9177), .Z(
        P1_U3554) );
  NAND2_X1 U10395 ( .A1(n9196), .A2(n9179), .ZN(n9178) );
  OAI21_X1 U10396 ( .B1(n9196), .B2(n9179), .A(n9178), .ZN(n9180) );
  INV_X1 U10397 ( .A(n9180), .ZN(n9186) );
  NAND2_X1 U10398 ( .A1(n9182), .A2(n9181), .ZN(n9184) );
  NAND2_X1 U10399 ( .A1(n9184), .A2(n9183), .ZN(n9185) );
  NOR2_X1 U10400 ( .A1(n9185), .A2(n9186), .ZN(n9203) );
  AOI21_X1 U10401 ( .B1(n9186), .B2(n9185), .A(n9203), .ZN(n9199) );
  NOR2_X1 U10402 ( .A1(n9188), .A2(n9187), .ZN(n9190) );
  NAND2_X1 U10403 ( .A1(n9196), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9200) );
  OAI21_X1 U10404 ( .B1(n9196), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9200), .ZN(
        n9192) );
  INV_X1 U10405 ( .A(n9201), .ZN(n9191) );
  AOI211_X1 U10406 ( .C1(n9193), .C2(n9192), .A(n9191), .B(n9784), .ZN(n9194)
         );
  AOI211_X1 U10407 ( .C1(n9794), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9195), .B(
        n9194), .ZN(n9198) );
  NAND2_X1 U10408 ( .A1(n9776), .A2(n9196), .ZN(n9197) );
  OAI211_X1 U10409 ( .C1(n9199), .C2(n9242), .A(n9198), .B(n9197), .ZN(
        P1_U3259) );
  INV_X1 U10410 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9570) );
  AOI22_X1 U10411 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9222), .B1(n9211), .B2(
        n9570), .ZN(n9202) );
  OAI21_X1 U10412 ( .B1(n4341), .B2(n9202), .A(n9223), .ZN(n9215) );
  AOI21_X1 U10413 ( .B1(n9179), .B2(n9204), .A(n9203), .ZN(n9207) );
  AOI22_X1 U10414 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(n9211), .B1(n9222), .B2(
        n9205), .ZN(n9206) );
  NOR2_X1 U10415 ( .A1(n9207), .A2(n9206), .ZN(n9217) );
  AOI21_X1 U10416 ( .B1(n9207), .B2(n9206), .A(n9217), .ZN(n9208) );
  NOR2_X1 U10417 ( .A1(n9208), .A2(n9242), .ZN(n9213) );
  AOI21_X1 U10418 ( .B1(n9794), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9209), .ZN(
        n9210) );
  OAI21_X1 U10419 ( .B1(n9798), .B2(n9211), .A(n9210), .ZN(n9212) );
  AOI211_X1 U10420 ( .C1(n9215), .C2(n9214), .A(n9213), .B(n9212), .ZN(n9216)
         );
  INV_X1 U10421 ( .A(n9216), .ZN(P1_U3260) );
  INV_X1 U10422 ( .A(n9235), .ZN(n9230) );
  INV_X1 U10423 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9621) );
  XNOR2_X1 U10424 ( .A(n9235), .B(n9621), .ZN(n9221) );
  OR2_X1 U10425 ( .A1(n9222), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9219) );
  INV_X1 U10426 ( .A(n9217), .ZN(n9218) );
  AND2_X1 U10427 ( .A1(n9219), .A2(n9218), .ZN(n9220) );
  NAND2_X1 U10428 ( .A1(n9221), .A2(n9220), .ZN(n9237) );
  OAI211_X1 U10429 ( .C1(n9221), .C2(n9220), .A(n9789), .B(n9237), .ZN(n9229)
         );
  AND2_X1 U10430 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9227) );
  INV_X1 U10431 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9429) );
  MUX2_X1 U10432 ( .A(n9429), .B(P1_REG2_REG_18__SCAN_IN), .S(n9235), .Z(n9224) );
  NOR2_X1 U10433 ( .A1(n9224), .A2(n9225), .ZN(n9232) );
  AOI211_X1 U10434 ( .C1(n9225), .C2(n9224), .A(n9232), .B(n9784), .ZN(n9226)
         );
  AOI211_X1 U10435 ( .C1(n9794), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9227), .B(
        n9226), .ZN(n9228) );
  OAI211_X1 U10436 ( .C1(n9798), .C2(n9230), .A(n9229), .B(n9228), .ZN(
        P1_U3261) );
  AND2_X1 U10437 ( .A1(n9235), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9231) );
  XNOR2_X1 U10438 ( .A(n9234), .B(n9233), .ZN(n9240) );
  NAND2_X1 U10439 ( .A1(n9235), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U10440 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  XNOR2_X1 U10441 ( .A(n9238), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U10442 ( .A1(n9789), .A2(n9241), .ZN(n9239) );
  INV_X1 U10443 ( .A(n9240), .ZN(n9243) );
  NAND2_X1 U10444 ( .A1(n9794), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9245) );
  NAND2_X1 U10445 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9244) );
  NAND2_X1 U10446 ( .A1(n9245), .A2(n9244), .ZN(n9246) );
  NOR2_X1 U10447 ( .A1(n5759), .A2(n9427), .ZN(n9247) );
  AOI211_X1 U10448 ( .C1(n9898), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9248), .B(
        n9247), .ZN(n9249) );
  OAI21_X1 U10449 ( .B1(n9831), .B2(n9250), .A(n9249), .ZN(P1_U3264) );
  OAI21_X1 U10450 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9256) );
  INV_X1 U10451 ( .A(n9254), .ZN(n9255) );
  AOI21_X1 U10452 ( .B1(n9256), .B2(n9868), .A(n9255), .ZN(n9441) );
  OR2_X1 U10453 ( .A1(n9258), .A2(n9257), .ZN(n9438) );
  NAND3_X1 U10454 ( .A1(n9438), .A2(n9259), .A3(n9874), .ZN(n9266) );
  AOI211_X1 U10455 ( .C1(n9261), .C2(n9268), .A(n9425), .B(n9260), .ZN(n9439)
         );
  AOI22_X1 U10456 ( .A1(n9262), .A2(n9899), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9898), .ZN(n9263) );
  OAI21_X1 U10457 ( .B1(n4614), .B2(n9427), .A(n9263), .ZN(n9264) );
  AOI21_X1 U10458 ( .B1(n9439), .B2(n9905), .A(n9264), .ZN(n9265) );
  OAI211_X1 U10459 ( .C1(n9898), .C2(n9441), .A(n9266), .B(n9265), .ZN(
        P1_U3265) );
  XNOR2_X1 U10460 ( .A(n9267), .B(n9275), .ZN(n9446) );
  INV_X1 U10461 ( .A(n9268), .ZN(n9269) );
  AOI211_X1 U10462 ( .C1(n6199), .C2(n4618), .A(n9425), .B(n9269), .ZN(n9443)
         );
  AOI22_X1 U10463 ( .A1(n9270), .A2(n9899), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9898), .ZN(n9271) );
  OAI21_X1 U10464 ( .B1(n9272), .B2(n9427), .A(n9271), .ZN(n9280) );
  OAI21_X1 U10465 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9278) );
  INV_X1 U10466 ( .A(n9276), .ZN(n9277) );
  AOI21_X1 U10467 ( .B1(n9278), .B2(n9868), .A(n9277), .ZN(n9445) );
  NOR2_X1 U10468 ( .A1(n9445), .A2(n9898), .ZN(n9279) );
  AOI211_X1 U10469 ( .C1(n9443), .C2(n9905), .A(n9280), .B(n9279), .ZN(n9281)
         );
  OAI21_X1 U10470 ( .B1(n9446), .B2(n9412), .A(n9281), .ZN(P1_U3266) );
  XNOR2_X1 U10471 ( .A(n9282), .B(n9284), .ZN(n9449) );
  INV_X1 U10472 ( .A(n9449), .ZN(n9300) );
  NAND2_X1 U10473 ( .A1(n9303), .A2(n9283), .ZN(n9285) );
  NAND2_X1 U10474 ( .A1(n9285), .A2(n9284), .ZN(n9287) );
  NAND2_X1 U10475 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  NAND2_X1 U10476 ( .A1(n9288), .A2(n9868), .ZN(n9291) );
  INV_X1 U10477 ( .A(n9289), .ZN(n9290) );
  NAND2_X1 U10478 ( .A1(n9291), .A2(n9290), .ZN(n9447) );
  AOI211_X1 U10479 ( .C1(n9293), .C2(n9309), .A(n9425), .B(n9292), .ZN(n9448)
         );
  NAND2_X1 U10480 ( .A1(n9448), .A2(n9905), .ZN(n9297) );
  INV_X1 U10481 ( .A(n9294), .ZN(n9295) );
  AOI22_X1 U10482 ( .A1(n9295), .A2(n9899), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9898), .ZN(n9296) );
  OAI211_X1 U10483 ( .C1(n9639), .C2(n9427), .A(n9297), .B(n9296), .ZN(n9298)
         );
  AOI21_X1 U10484 ( .B1(n9836), .B2(n9447), .A(n9298), .ZN(n9299) );
  OAI21_X1 U10485 ( .B1(n9300), .B2(n9412), .A(n9299), .ZN(P1_U3267) );
  XNOR2_X1 U10486 ( .A(n9301), .B(n9302), .ZN(n9456) );
  OAI211_X1 U10487 ( .C1(n9305), .C2(n9304), .A(n9303), .B(n9868), .ZN(n9308)
         );
  INV_X1 U10488 ( .A(n9306), .ZN(n9307) );
  NAND2_X1 U10489 ( .A1(n9308), .A2(n9307), .ZN(n9452) );
  INV_X1 U10490 ( .A(n9325), .ZN(n9311) );
  INV_X1 U10491 ( .A(n9309), .ZN(n9310) );
  AOI211_X1 U10492 ( .C1(n9454), .C2(n9311), .A(n9425), .B(n9310), .ZN(n9453)
         );
  NAND2_X1 U10493 ( .A1(n9453), .A2(n9905), .ZN(n9314) );
  AOI22_X1 U10494 ( .A1(n9312), .A2(n9899), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9898), .ZN(n9313) );
  OAI211_X1 U10495 ( .C1(n9315), .C2(n9427), .A(n9314), .B(n9313), .ZN(n9316)
         );
  AOI21_X1 U10496 ( .B1(n9836), .B2(n9452), .A(n9316), .ZN(n9317) );
  OAI21_X1 U10497 ( .B1(n9456), .B2(n9412), .A(n9317), .ZN(P1_U3268) );
  XNOR2_X1 U10498 ( .A(n9318), .B(n9319), .ZN(n9459) );
  INV_X1 U10499 ( .A(n9459), .ZN(n9332) );
  OAI211_X1 U10500 ( .C1(n9322), .C2(n9321), .A(n9320), .B(n9868), .ZN(n9324)
         );
  NAND2_X1 U10501 ( .A1(n9324), .A2(n9323), .ZN(n9457) );
  AOI211_X1 U10502 ( .C1(n9326), .C2(n9336), .A(n9425), .B(n9325), .ZN(n9458)
         );
  NAND2_X1 U10503 ( .A1(n9458), .A2(n9905), .ZN(n9329) );
  AOI22_X1 U10504 ( .A1(n9327), .A2(n9899), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9898), .ZN(n9328) );
  OAI211_X1 U10505 ( .C1(n9644), .C2(n9427), .A(n9329), .B(n9328), .ZN(n9330)
         );
  AOI21_X1 U10506 ( .B1(n9836), .B2(n9457), .A(n9330), .ZN(n9331) );
  OAI21_X1 U10507 ( .B1(n9332), .B2(n9412), .A(n9331), .ZN(P1_U3269) );
  XNOR2_X1 U10508 ( .A(n9333), .B(n9334), .ZN(n9466) );
  AOI21_X1 U10509 ( .B1(n9463), .B2(n9354), .A(n9425), .ZN(n9335) );
  AND2_X1 U10510 ( .A1(n9336), .A2(n9335), .ZN(n9462) );
  INV_X1 U10511 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9337) );
  OAI22_X1 U10512 ( .A1(n4619), .A2(n9427), .B1(n9337), .B2(n9836), .ZN(n9345)
         );
  OAI21_X1 U10513 ( .B1(n4788), .B2(n9339), .A(n9338), .ZN(n9341) );
  AOI21_X1 U10514 ( .B1(n9341), .B2(n9868), .A(n9340), .ZN(n9465) );
  NAND2_X1 U10515 ( .A1(n9342), .A2(n9899), .ZN(n9343) );
  AOI21_X1 U10516 ( .B1(n9465), .B2(n9343), .A(n9898), .ZN(n9344) );
  AOI211_X1 U10517 ( .C1(n9462), .C2(n9905), .A(n9345), .B(n9344), .ZN(n9346)
         );
  OAI21_X1 U10518 ( .B1(n9466), .B2(n9412), .A(n9346), .ZN(P1_U3270) );
  XOR2_X1 U10519 ( .A(n9347), .B(n9349), .Z(n9469) );
  INV_X1 U10520 ( .A(n9469), .ZN(n9362) );
  OAI211_X1 U10521 ( .C1(n9350), .C2(n9349), .A(n9348), .B(n9868), .ZN(n9353)
         );
  INV_X1 U10522 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U10523 ( .A1(n9353), .A2(n9352), .ZN(n9467) );
  INV_X1 U10524 ( .A(n9354), .ZN(n9355) );
  AOI211_X1 U10525 ( .C1(n9356), .C2(n9372), .A(n9425), .B(n9355), .ZN(n9468)
         );
  NAND2_X1 U10526 ( .A1(n9468), .A2(n9905), .ZN(n9359) );
  AOI22_X1 U10527 ( .A1(n9898), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9357), .B2(
        n9899), .ZN(n9358) );
  OAI211_X1 U10528 ( .C1(n9649), .C2(n9427), .A(n9359), .B(n9358), .ZN(n9360)
         );
  AOI21_X1 U10529 ( .B1(n9836), .B2(n9467), .A(n9360), .ZN(n9361) );
  OAI21_X1 U10530 ( .B1(n9362), .B2(n9412), .A(n9361), .ZN(P1_U3271) );
  XNOR2_X1 U10531 ( .A(n9363), .B(n9367), .ZN(n9474) );
  INV_X1 U10532 ( .A(n9474), .ZN(n9382) );
  INV_X1 U10533 ( .A(n9365), .ZN(n9385) );
  NAND2_X1 U10534 ( .A1(n9364), .A2(n9385), .ZN(n9384) );
  NAND2_X1 U10535 ( .A1(n9384), .A2(n9366), .ZN(n9368) );
  XNOR2_X1 U10536 ( .A(n9368), .B(n9367), .ZN(n9371) );
  INV_X1 U10537 ( .A(n9369), .ZN(n9370) );
  OAI21_X1 U10538 ( .B1(n9371), .B2(n9895), .A(n9370), .ZN(n9472) );
  INV_X1 U10539 ( .A(n9389), .ZN(n9374) );
  INV_X1 U10540 ( .A(n9372), .ZN(n9373) );
  AOI211_X1 U10541 ( .C1(n9375), .C2(n9374), .A(n9425), .B(n9373), .ZN(n9473)
         );
  NAND2_X1 U10542 ( .A1(n9473), .A2(n9905), .ZN(n9379) );
  INV_X1 U10543 ( .A(n9376), .ZN(n9377) );
  AOI22_X1 U10544 ( .A1(n9898), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9377), .B2(
        n9899), .ZN(n9378) );
  OAI211_X1 U10545 ( .C1(n9653), .C2(n9427), .A(n9379), .B(n9378), .ZN(n9380)
         );
  AOI21_X1 U10546 ( .B1(n9836), .B2(n9472), .A(n9380), .ZN(n9381) );
  OAI21_X1 U10547 ( .B1(n9382), .B2(n9412), .A(n9381), .ZN(P1_U3272) );
  XNOR2_X1 U10548 ( .A(n9383), .B(n9385), .ZN(n9479) );
  INV_X1 U10549 ( .A(n9479), .ZN(n9397) );
  OAI211_X1 U10550 ( .C1(n9364), .C2(n9385), .A(n9384), .B(n9868), .ZN(n9388)
         );
  INV_X1 U10551 ( .A(n9386), .ZN(n9387) );
  NAND2_X1 U10552 ( .A1(n9388), .A2(n9387), .ZN(n9477) );
  INV_X1 U10553 ( .A(n9399), .ZN(n9390) );
  AOI211_X1 U10554 ( .C1(n9391), .C2(n9390), .A(n9425), .B(n9389), .ZN(n9478)
         );
  NAND2_X1 U10555 ( .A1(n9478), .A2(n9905), .ZN(n9394) );
  AOI22_X1 U10556 ( .A1(n9898), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9392), .B2(
        n9899), .ZN(n9393) );
  OAI211_X1 U10557 ( .C1(n9657), .C2(n9427), .A(n9394), .B(n9393), .ZN(n9395)
         );
  AOI21_X1 U10558 ( .B1(n9836), .B2(n9477), .A(n9395), .ZN(n9396) );
  OAI21_X1 U10559 ( .B1(n9397), .B2(n9412), .A(n9396), .ZN(P1_U3273) );
  XOR2_X1 U10560 ( .A(n9398), .B(n9405), .Z(n9486) );
  AOI211_X1 U10561 ( .C1(n9483), .C2(n9423), .A(n9425), .B(n9399), .ZN(n9482)
         );
  INV_X1 U10562 ( .A(n9400), .ZN(n9401) );
  AOI22_X1 U10563 ( .A1(n9898), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9401), .B2(
        n9899), .ZN(n9402) );
  OAI21_X1 U10564 ( .B1(n9403), .B2(n9427), .A(n9402), .ZN(n9410) );
  NAND2_X1 U10565 ( .A1(n9415), .A2(n9404), .ZN(n9406) );
  XOR2_X1 U10566 ( .A(n9406), .B(n9405), .Z(n9408) );
  AOI21_X1 U10567 ( .B1(n9408), .B2(n9868), .A(n9407), .ZN(n9485) );
  NOR2_X1 U10568 ( .A1(n9485), .A2(n9898), .ZN(n9409) );
  AOI211_X1 U10569 ( .C1(n9482), .C2(n9905), .A(n9410), .B(n9409), .ZN(n9411)
         );
  OAI21_X1 U10570 ( .B1(n9486), .B2(n9412), .A(n9411), .ZN(P1_U3274) );
  NAND2_X1 U10571 ( .A1(n9413), .A2(n9421), .ZN(n9414) );
  NAND2_X1 U10572 ( .A1(n9415), .A2(n9414), .ZN(n9416) );
  NAND2_X1 U10573 ( .A1(n9416), .A2(n9868), .ZN(n9419) );
  INV_X1 U10574 ( .A(n9417), .ZN(n9418) );
  NAND2_X1 U10575 ( .A1(n9419), .A2(n9418), .ZN(n9618) );
  INV_X1 U10576 ( .A(n9618), .ZN(n9434) );
  OAI21_X1 U10577 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9620) );
  NAND2_X1 U10578 ( .A1(n9620), .A2(n9874), .ZN(n9433) );
  INV_X1 U10579 ( .A(n9423), .ZN(n9424) );
  AOI211_X1 U10580 ( .C1(n9426), .C2(n8139), .A(n9425), .B(n9424), .ZN(n9619)
         );
  NOR2_X1 U10581 ( .A1(n9662), .A2(n9427), .ZN(n9431) );
  OAI22_X1 U10582 ( .A1(n9836), .A2(n9429), .B1(n9428), .B2(n9878), .ZN(n9430)
         );
  AOI211_X1 U10583 ( .C1(n9619), .C2(n9905), .A(n9431), .B(n9430), .ZN(n9432)
         );
  OAI211_X1 U10584 ( .C1(n9898), .C2(n9434), .A(n9433), .B(n9432), .ZN(
        P1_U3275) );
  NAND2_X1 U10585 ( .A1(n9436), .A2(n4781), .ZN(n9437) );
  OAI21_X1 U10586 ( .B1(n5759), .B2(n9633), .A(n9437), .ZN(P1_U3552) );
  NAND3_X1 U10587 ( .A1(n9438), .A2(n9259), .A3(n9987), .ZN(n9442) );
  AOI21_X1 U10588 ( .B1(n9977), .B2(n9261), .A(n9439), .ZN(n9440) );
  NAND3_X1 U10589 ( .A1(n9442), .A2(n9441), .A3(n9440), .ZN(n9634) );
  MUX2_X1 U10590 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9634), .S(n10015), .Z(
        P1_U3550) );
  AOI21_X1 U10591 ( .B1(n9977), .B2(n6199), .A(n9443), .ZN(n9444) );
  OAI211_X1 U10592 ( .C1(n9446), .C2(n9941), .A(n9445), .B(n9444), .ZN(n9635)
         );
  MUX2_X1 U10593 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9635), .S(n10015), .Z(
        P1_U3549) );
  AOI211_X1 U10594 ( .C1(n9449), .C2(n9987), .A(n9448), .B(n9447), .ZN(n9636)
         );
  MUX2_X1 U10595 ( .A(n9450), .B(n9636), .S(n10015), .Z(n9451) );
  OAI21_X1 U10596 ( .B1(n9639), .B2(n9633), .A(n9451), .ZN(P1_U3548) );
  AOI211_X1 U10597 ( .C1(n9977), .C2(n9454), .A(n9453), .B(n9452), .ZN(n9455)
         );
  OAI21_X1 U10598 ( .B1(n9456), .B2(n9941), .A(n9455), .ZN(n9640) );
  MUX2_X1 U10599 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9640), .S(n10015), .Z(
        P1_U3547) );
  INV_X1 U10600 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9460) );
  AOI211_X1 U10601 ( .C1(n9459), .C2(n9987), .A(n9458), .B(n9457), .ZN(n9641)
         );
  MUX2_X1 U10602 ( .A(n9460), .B(n9641), .S(n10015), .Z(n9461) );
  OAI21_X1 U10603 ( .B1(n9644), .B2(n9633), .A(n9461), .ZN(P1_U3546) );
  AOI21_X1 U10604 ( .B1(n9977), .B2(n9463), .A(n9462), .ZN(n9464) );
  OAI211_X1 U10605 ( .C1(n9466), .C2(n9941), .A(n9465), .B(n9464), .ZN(n9645)
         );
  MUX2_X1 U10606 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9645), .S(n10015), .Z(
        P1_U3545) );
  INV_X1 U10607 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9470) );
  AOI211_X1 U10608 ( .C1(n9469), .C2(n9987), .A(n9468), .B(n9467), .ZN(n9646)
         );
  MUX2_X1 U10609 ( .A(n9470), .B(n9646), .S(n10015), .Z(n9471) );
  OAI21_X1 U10610 ( .B1(n9649), .B2(n9633), .A(n9471), .ZN(P1_U3544) );
  INV_X1 U10611 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9475) );
  AOI211_X1 U10612 ( .C1(n9474), .C2(n9987), .A(n9473), .B(n9472), .ZN(n9650)
         );
  MUX2_X1 U10613 ( .A(n9475), .B(n9650), .S(n10015), .Z(n9476) );
  OAI21_X1 U10614 ( .B1(n9653), .B2(n9633), .A(n9476), .ZN(P1_U3543) );
  INV_X1 U10615 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9480) );
  AOI211_X1 U10616 ( .C1(n9479), .C2(n9987), .A(n9478), .B(n9477), .ZN(n9654)
         );
  MUX2_X1 U10617 ( .A(n9480), .B(n9654), .S(n10015), .Z(n9481) );
  OAI21_X1 U10618 ( .B1(n9657), .B2(n9633), .A(n9481), .ZN(P1_U3542) );
  AOI21_X1 U10619 ( .B1(n9977), .B2(n9483), .A(n9482), .ZN(n9484) );
  OAI211_X1 U10620 ( .C1(n9486), .C2(n9941), .A(n9485), .B(n9484), .ZN(n9658)
         );
  MUX2_X1 U10621 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9658), .S(n10015), .Z(
        n9617) );
  NAND3_X1 U10622 ( .A1(keyinput0), .A2(keyinput16), .A3(keyinput54), .ZN(
        n9488) );
  NAND3_X1 U10623 ( .A1(keyinput44), .A2(keyinput5), .A3(keyinput32), .ZN(
        n9487) );
  OR4_X1 U10624 ( .A1(n9488), .A2(n9487), .A3(keyinput30), .A4(keyinput12), 
        .ZN(n9499) );
  NAND2_X1 U10625 ( .A1(keyinput48), .A2(keyinput22), .ZN(n9489) );
  NOR3_X1 U10626 ( .A1(keyinput23), .A2(keyinput37), .A3(n9489), .ZN(n9492) );
  NOR3_X1 U10627 ( .A1(keyinput24), .A2(keyinput29), .A3(keyinput27), .ZN(
        n9491) );
  NOR4_X1 U10628 ( .A1(keyinput36), .A2(keyinput8), .A3(keyinput46), .A4(
        keyinput25), .ZN(n9490) );
  NAND4_X1 U10629 ( .A1(n9492), .A2(keyinput13), .A3(n9491), .A4(n9490), .ZN(
        n9498) );
  NOR3_X1 U10630 ( .A1(keyinput26), .A2(keyinput60), .A3(keyinput38), .ZN(
        n9494) );
  NOR3_X1 U10631 ( .A1(keyinput33), .A2(keyinput17), .A3(keyinput20), .ZN(
        n9493) );
  NAND4_X1 U10632 ( .A1(keyinput41), .A2(n9494), .A3(keyinput55), .A4(n9493), 
        .ZN(n9497) );
  NOR2_X1 U10633 ( .A1(keyinput31), .A2(keyinput11), .ZN(n9495) );
  NAND3_X1 U10634 ( .A1(keyinput53), .A2(keyinput52), .A3(n9495), .ZN(n9496)
         );
  OR4_X1 U10635 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n9588)
         );
  NOR4_X1 U10636 ( .A1(keyinput9), .A2(keyinput1), .A3(keyinput21), .A4(
        keyinput4), .ZN(n9509) );
  NOR4_X1 U10637 ( .A1(keyinput28), .A2(keyinput42), .A3(keyinput39), .A4(
        keyinput58), .ZN(n9508) );
  OR4_X1 U10638 ( .A1(keyinput59), .A2(keyinput63), .A3(keyinput51), .A4(
        keyinput15), .ZN(n9501) );
  NAND2_X1 U10639 ( .A1(keyinput45), .A2(keyinput49), .ZN(n9500) );
  NOR4_X1 U10640 ( .A1(keyinput19), .A2(keyinput18), .A3(n9501), .A4(n9500), 
        .ZN(n9507) );
  NAND4_X1 U10641 ( .A1(keyinput57), .A2(keyinput61), .A3(keyinput40), .A4(
        keyinput56), .ZN(n9505) );
  NAND4_X1 U10642 ( .A1(keyinput47), .A2(keyinput43), .A3(keyinput34), .A4(
        keyinput35), .ZN(n9504) );
  NAND4_X1 U10643 ( .A1(keyinput50), .A2(keyinput62), .A3(keyinput14), .A4(
        keyinput10), .ZN(n9503) );
  NAND4_X1 U10644 ( .A1(keyinput3), .A2(keyinput2), .A3(keyinput6), .A4(
        keyinput7), .ZN(n9502) );
  NOR4_X1 U10645 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n9506)
         );
  NAND4_X1 U10646 ( .A1(n9509), .A2(n9508), .A3(n9507), .A4(n9506), .ZN(n9587)
         );
  AOI22_X1 U10647 ( .A1(n9511), .A2(keyinput30), .B1(keyinput32), .B2(n8794), 
        .ZN(n9510) );
  OAI221_X1 U10648 ( .B1(n9511), .B2(keyinput30), .C1(n8794), .C2(keyinput32), 
        .A(n9510), .ZN(n9521) );
  INV_X1 U10649 ( .A(keyinput44), .ZN(n9513) );
  AOI22_X1 U10650 ( .A1(n9514), .A2(keyinput5), .B1(P2_ADDR_REG_0__SCAN_IN), 
        .B2(n9513), .ZN(n9512) );
  OAI221_X1 U10651 ( .B1(n9514), .B2(keyinput5), .C1(n9513), .C2(
        P2_ADDR_REG_0__SCAN_IN), .A(n9512), .ZN(n9520) );
  INV_X1 U10652 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9913) );
  AOI22_X1 U10653 ( .A1(n7363), .A2(keyinput28), .B1(n9913), .B2(keyinput51), 
        .ZN(n9515) );
  OAI221_X1 U10654 ( .B1(n7363), .B2(keyinput28), .C1(n9913), .C2(keyinput51), 
        .A(n9515), .ZN(n9519) );
  AOI22_X1 U10655 ( .A1(n9914), .A2(keyinput43), .B1(keyinput35), .B2(n9517), 
        .ZN(n9516) );
  OAI221_X1 U10656 ( .B1(n9914), .B2(keyinput43), .C1(n9517), .C2(keyinput35), 
        .A(n9516), .ZN(n9518) );
  OR4_X1 U10657 ( .A1(n9521), .A2(n9520), .A3(n9519), .A4(n9518), .ZN(n9532)
         );
  AOI22_X1 U10658 ( .A1(n9911), .A2(keyinput20), .B1(keyinput55), .B2(n9523), 
        .ZN(n9522) );
  OAI221_X1 U10659 ( .B1(n9911), .B2(keyinput20), .C1(n9523), .C2(keyinput55), 
        .A(n9522), .ZN(n9531) );
  XNOR2_X1 U10660 ( .A(n9912), .B(keyinput38), .ZN(n9530) );
  XOR2_X1 U10661 ( .A(n6924), .B(keyinput9), .Z(n9528) );
  XOR2_X1 U10662 ( .A(n9524), .B(keyinput29), .Z(n9527) );
  XOR2_X1 U10663 ( .A(n6072), .B(keyinput31), .Z(n9526) );
  XNOR2_X1 U10664 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput4), .ZN(n9525) );
  NAND4_X1 U10665 ( .A1(n9528), .A2(n9527), .A3(n9526), .A4(n9525), .ZN(n9529)
         );
  NOR4_X1 U10666 ( .A1(n9532), .A2(n9531), .A3(n9530), .A4(n9529), .ZN(n9586)
         );
  AOI22_X1 U10667 ( .A1(n8768), .A2(keyinput10), .B1(keyinput6), .B2(n9534), 
        .ZN(n9533) );
  OAI221_X1 U10668 ( .B1(n8768), .B2(keyinput10), .C1(n9534), .C2(keyinput6), 
        .A(n9533), .ZN(n9538) );
  AOI22_X1 U10669 ( .A1(n8782), .A2(keyinput48), .B1(n9536), .B2(keyinput37), 
        .ZN(n9535) );
  OAI221_X1 U10670 ( .B1(n8782), .B2(keyinput48), .C1(n9536), .C2(keyinput37), 
        .A(n9535), .ZN(n9537) );
  NOR2_X1 U10671 ( .A1(n9538), .A2(n9537), .ZN(n9567) );
  AOI22_X1 U10672 ( .A1(n5070), .A2(keyinput0), .B1(n9540), .B2(keyinput12), 
        .ZN(n9539) );
  OAI221_X1 U10673 ( .B1(n5070), .B2(keyinput0), .C1(n9540), .C2(keyinput12), 
        .A(n9539), .ZN(n9543) );
  INV_X1 U10674 ( .A(keyinput17), .ZN(n9541) );
  XNOR2_X1 U10675 ( .A(n9541), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(n9542) );
  NOR2_X1 U10676 ( .A1(n9543), .A2(n9542), .ZN(n9566) );
  XNOR2_X1 U10677 ( .A(SI_0_), .B(keyinput41), .ZN(n9547) );
  XNOR2_X1 U10678 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput22), .ZN(n9546) );
  XNOR2_X1 U10679 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput33), .ZN(n9545) );
  XNOR2_X1 U10680 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput23), .ZN(n9544)
         );
  NAND4_X1 U10681 ( .A1(n9547), .A2(n9546), .A3(n9545), .A4(n9544), .ZN(n9553)
         );
  XNOR2_X1 U10682 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput13), .ZN(n9551) );
  XNOR2_X1 U10683 ( .A(P1_REG3_REG_17__SCAN_IN), .B(keyinput11), .ZN(n9550) );
  XNOR2_X1 U10684 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput36), .ZN(n9549) );
  XNOR2_X1 U10685 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput52), .ZN(n9548) );
  NAND4_X1 U10686 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(n9552)
         );
  NOR2_X1 U10687 ( .A1(n9553), .A2(n9552), .ZN(n9565) );
  XNOR2_X1 U10688 ( .A(P2_REG0_REG_17__SCAN_IN), .B(keyinput8), .ZN(n9557) );
  XNOR2_X1 U10689 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput53), .ZN(n9556) );
  XNOR2_X1 U10690 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput27), .ZN(n9555) );
  XNOR2_X1 U10691 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput24), .ZN(n9554) );
  NAND4_X1 U10692 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n9563)
         );
  XNOR2_X1 U10693 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput50), .ZN(n9561) );
  XNOR2_X1 U10694 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput18), .ZN(n9560) );
  XNOR2_X1 U10695 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput14), .ZN(n9559) );
  XNOR2_X1 U10696 ( .A(P2_REG0_REG_26__SCAN_IN), .B(keyinput61), .ZN(n9558) );
  NAND4_X1 U10697 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(n9562)
         );
  NOR2_X1 U10698 ( .A1(n9563), .A2(n9562), .ZN(n9564) );
  NAND4_X1 U10699 ( .A1(n9567), .A2(n9566), .A3(n9565), .A4(n9564), .ZN(n9584)
         );
  INV_X1 U10700 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9569) );
  AOI22_X1 U10701 ( .A1(n9570), .A2(keyinput59), .B1(keyinput49), .B2(n9569), 
        .ZN(n9568) );
  OAI221_X1 U10702 ( .B1(n9570), .B2(keyinput59), .C1(n9569), .C2(keyinput49), 
        .A(n9568), .ZN(n9583) );
  AOI22_X1 U10703 ( .A1(n5529), .A2(keyinput19), .B1(n9910), .B2(keyinput45), 
        .ZN(n9571) );
  OAI221_X1 U10704 ( .B1(n5529), .B2(keyinput19), .C1(n9910), .C2(keyinput45), 
        .A(n9571), .ZN(n9582) );
  AOI22_X1 U10705 ( .A1(n9573), .A2(keyinput16), .B1(keyinput54), .B2(n5020), 
        .ZN(n9572) );
  OAI221_X1 U10706 ( .B1(n9573), .B2(keyinput16), .C1(n5020), .C2(keyinput54), 
        .A(n9572), .ZN(n9580) );
  AOI22_X1 U10707 ( .A1(n9576), .A2(keyinput46), .B1(keyinput25), .B2(n9575), 
        .ZN(n9574) );
  OAI221_X1 U10708 ( .B1(n9576), .B2(keyinput46), .C1(n9575), .C2(keyinput25), 
        .A(n9574), .ZN(n9579) );
  AOI22_X1 U10709 ( .A1(n9777), .A2(keyinput26), .B1(n4843), .B2(keyinput60), 
        .ZN(n9577) );
  OAI221_X1 U10710 ( .B1(n9777), .B2(keyinput26), .C1(n4843), .C2(keyinput60), 
        .A(n9577), .ZN(n9578) );
  OR3_X1 U10711 ( .A1(n9580), .A2(n9579), .A3(n9578), .ZN(n9581) );
  NOR4_X1 U10712 ( .A1(n9584), .A2(n9583), .A3(n9582), .A4(n9581), .ZN(n9585)
         );
  OAI211_X1 U10713 ( .C1(n9588), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9589)
         );
  INV_X1 U10714 ( .A(n9589), .ZN(n9615) );
  AOI22_X1 U10715 ( .A1(n6047), .A2(keyinput39), .B1(n9591), .B2(keyinput3), 
        .ZN(n9590) );
  OAI221_X1 U10716 ( .B1(n6047), .B2(keyinput39), .C1(n9591), .C2(keyinput3), 
        .A(n9590), .ZN(n9600) );
  AOI22_X1 U10717 ( .A1(n6042), .A2(keyinput1), .B1(keyinput63), .B2(n5127), 
        .ZN(n9592) );
  OAI221_X1 U10718 ( .B1(n6042), .B2(keyinput1), .C1(n5127), .C2(keyinput63), 
        .A(n9592), .ZN(n9599) );
  INV_X1 U10719 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U10720 ( .A1(n9594), .A2(keyinput57), .B1(n9983), .B2(keyinput7), 
        .ZN(n9593) );
  OAI221_X1 U10721 ( .B1(n9594), .B2(keyinput57), .C1(n9983), .C2(keyinput7), 
        .A(n9593), .ZN(n9598) );
  AOI22_X1 U10722 ( .A1(n4933), .A2(keyinput56), .B1(P2_U3151), .B2(keyinput62), .ZN(n9595) );
  OAI221_X1 U10723 ( .B1(n4933), .B2(keyinput56), .C1(P2_U3151), .C2(
        keyinput62), .A(n9595), .ZN(n9597) );
  NOR4_X1 U10724 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9614)
         );
  AOI22_X1 U10725 ( .A1(n5305), .A2(keyinput15), .B1(keyinput2), .B2(n9602), 
        .ZN(n9601) );
  OAI221_X1 U10726 ( .B1(n5305), .B2(keyinput15), .C1(n9602), .C2(keyinput2), 
        .A(n9601), .ZN(n9612) );
  AOI22_X1 U10727 ( .A1(n9604), .A2(keyinput21), .B1(keyinput40), .B2(n9642), 
        .ZN(n9603) );
  OAI221_X1 U10728 ( .B1(n9604), .B2(keyinput21), .C1(n9642), .C2(keyinput40), 
        .A(n9603), .ZN(n9611) );
  INV_X1 U10729 ( .A(keyinput47), .ZN(n9606) );
  AOI22_X1 U10730 ( .A1(n9607), .A2(keyinput42), .B1(P2_ADDR_REG_14__SCAN_IN), 
        .B2(n9606), .ZN(n9605) );
  OAI221_X1 U10731 ( .B1(n9607), .B2(keyinput42), .C1(n9606), .C2(
        P2_ADDR_REG_14__SCAN_IN), .A(n9605), .ZN(n9610) );
  INV_X1 U10732 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10052) );
  INV_X1 U10733 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U10734 ( .A1(n10052), .A2(keyinput58), .B1(n9909), .B2(keyinput34), 
        .ZN(n9608) );
  OAI221_X1 U10735 ( .B1(n10052), .B2(keyinput58), .C1(n9909), .C2(keyinput34), 
        .A(n9608), .ZN(n9609) );
  NOR4_X1 U10736 ( .A1(n9612), .A2(n9611), .A3(n9610), .A4(n9609), .ZN(n9613)
         );
  NAND3_X1 U10737 ( .A1(n9615), .A2(n9614), .A3(n9613), .ZN(n9616) );
  XNOR2_X1 U10738 ( .A(n9617), .B(n9616), .ZN(P1_U3541) );
  AOI211_X1 U10739 ( .C1(n9620), .C2(n9987), .A(n9619), .B(n9618), .ZN(n9659)
         );
  MUX2_X1 U10740 ( .A(n9621), .B(n9659), .S(n10015), .Z(n9622) );
  OAI21_X1 U10741 ( .B1(n9662), .B2(n9633), .A(n9622), .ZN(P1_U3540) );
  AOI21_X1 U10742 ( .B1(n9977), .B2(n9624), .A(n9623), .ZN(n9625) );
  OAI211_X1 U10743 ( .C1(n9627), .C2(n9941), .A(n9626), .B(n9625), .ZN(n9663)
         );
  MUX2_X1 U10744 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9663), .S(n10015), .Z(
        P1_U3539) );
  OAI211_X1 U10745 ( .C1(n9630), .C2(n9941), .A(n9629), .B(n9628), .ZN(n9631)
         );
  INV_X1 U10746 ( .A(n9631), .ZN(n9664) );
  MUX2_X1 U10747 ( .A(n9179), .B(n9664), .S(n10015), .Z(n9632) );
  OAI21_X1 U10748 ( .B1(n9668), .B2(n9633), .A(n9632), .ZN(P1_U3538) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9634), .S(n10000), .Z(
        P1_U3518) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9635), .S(n10000), .Z(
        P1_U3517) );
  INV_X1 U10751 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9637) );
  MUX2_X1 U10752 ( .A(n9637), .B(n9636), .S(n10000), .Z(n9638) );
  OAI21_X1 U10753 ( .B1(n9639), .B2(n9667), .A(n9638), .ZN(P1_U3516) );
  MUX2_X1 U10754 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9640), .S(n10000), .Z(
        P1_U3515) );
  MUX2_X1 U10755 ( .A(n9642), .B(n9641), .S(n10000), .Z(n9643) );
  OAI21_X1 U10756 ( .B1(n9644), .B2(n9667), .A(n9643), .ZN(P1_U3514) );
  MUX2_X1 U10757 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9645), .S(n10000), .Z(
        P1_U3513) );
  INV_X1 U10758 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9647) );
  MUX2_X1 U10759 ( .A(n9647), .B(n9646), .S(n10000), .Z(n9648) );
  OAI21_X1 U10760 ( .B1(n9649), .B2(n9667), .A(n9648), .ZN(P1_U3512) );
  INV_X1 U10761 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9651) );
  MUX2_X1 U10762 ( .A(n9651), .B(n9650), .S(n10000), .Z(n9652) );
  OAI21_X1 U10763 ( .B1(n9653), .B2(n9667), .A(n9652), .ZN(P1_U3511) );
  INV_X1 U10764 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9655) );
  MUX2_X1 U10765 ( .A(n9655), .B(n9654), .S(n10000), .Z(n9656) );
  OAI21_X1 U10766 ( .B1(n9657), .B2(n9667), .A(n9656), .ZN(P1_U3510) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9658), .S(n10000), .Z(
        P1_U3509) );
  INV_X1 U10768 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9660) );
  MUX2_X1 U10769 ( .A(n9660), .B(n9659), .S(n10000), .Z(n9661) );
  OAI21_X1 U10770 ( .B1(n9662), .B2(n9667), .A(n9661), .ZN(P1_U3507) );
  MUX2_X1 U10771 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9663), .S(n10000), .Z(
        P1_U3504) );
  INV_X1 U10772 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9665) );
  MUX2_X1 U10773 ( .A(n9665), .B(n9664), .S(n10000), .Z(n9666) );
  OAI21_X1 U10774 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(P1_U3501) );
  MUX2_X1 U10775 ( .A(P1_D_REG_1__SCAN_IN), .B(n9669), .S(n9915), .Z(P1_U3440)
         );
  NOR4_X1 U10776 ( .A1(n4736), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9670), .ZN(n9672) );
  AOI21_X1 U10777 ( .B1(n9673), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9672), .ZN(
        n9674) );
  OAI21_X1 U10778 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(P1_U3324) );
  NOR2_X1 U10779 ( .A1(n9677), .A2(n9678), .ZN(n9733) );
  NOR2_X1 U10780 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9729) );
  NOR2_X1 U10781 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9725) );
  NOR2_X1 U10782 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9721) );
  NOR2_X1 U10783 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9717) );
  NOR2_X1 U10784 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9713) );
  NOR2_X1 U10785 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9709) );
  NOR2_X1 U10786 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9705) );
  NOR2_X1 U10787 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9701) );
  NOR2_X1 U10788 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9697) );
  NOR2_X1 U10789 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9693) );
  NOR2_X1 U10790 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9691) );
  NOR2_X1 U10791 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9689) );
  NOR2_X1 U10792 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9687) );
  NOR2_X1 U10793 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9685) );
  NAND2_X1 U10794 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9683) );
  XOR2_X1 U10795 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10100) );
  NAND2_X1 U10796 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9681) );
  AOI21_X1 U10797 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10062) );
  INV_X1 U10798 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10066) );
  INV_X1 U10799 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10065) );
  NOR2_X1 U10800 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  AND2_X1 U10801 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10064), .ZN(n10061) );
  NOR2_X1 U10802 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10061), .ZN(n9679) );
  NOR2_X1 U10803 ( .A1(n10062), .A2(n9679), .ZN(n10098) );
  XOR2_X1 U10804 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10097) );
  NAND2_X1 U10805 ( .A1(n10098), .A2(n10097), .ZN(n9680) );
  NAND2_X1 U10806 ( .A1(n9681), .A2(n9680), .ZN(n10099) );
  NAND2_X1 U10807 ( .A1(n10100), .A2(n10099), .ZN(n9682) );
  NAND2_X1 U10808 ( .A1(n9683), .A2(n9682), .ZN(n10102) );
  XNOR2_X1 U10809 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10101) );
  NOR2_X1 U10810 ( .A1(n10102), .A2(n10101), .ZN(n9684) );
  NOR2_X1 U10811 ( .A1(n9685), .A2(n9684), .ZN(n10090) );
  XNOR2_X1 U10812 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10089) );
  NOR2_X1 U10813 ( .A1(n10090), .A2(n10089), .ZN(n9686) );
  NOR2_X1 U10814 ( .A1(n9687), .A2(n9686), .ZN(n10088) );
  XNOR2_X1 U10815 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10087) );
  NOR2_X1 U10816 ( .A1(n10088), .A2(n10087), .ZN(n9688) );
  NOR2_X1 U10817 ( .A1(n9689), .A2(n9688), .ZN(n10094) );
  XNOR2_X1 U10818 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10093) );
  NOR2_X1 U10819 ( .A1(n10094), .A2(n10093), .ZN(n9690) );
  NOR2_X1 U10820 ( .A1(n9691), .A2(n9690), .ZN(n10096) );
  XNOR2_X1 U10821 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10095) );
  NOR2_X1 U10822 ( .A1(n10096), .A2(n10095), .ZN(n9692) );
  NOR2_X1 U10823 ( .A1(n9693), .A2(n9692), .ZN(n10092) );
  INV_X1 U10824 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U10825 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9695), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n9694), .ZN(n10091) );
  NOR2_X1 U10826 ( .A1(n10092), .A2(n10091), .ZN(n9696) );
  NOR2_X1 U10827 ( .A1(n9697), .A2(n9696), .ZN(n10086) );
  INV_X1 U10828 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U10829 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9699), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n9698), .ZN(n10085) );
  NOR2_X1 U10830 ( .A1(n10086), .A2(n10085), .ZN(n9700) );
  NOR2_X1 U10831 ( .A1(n9701), .A2(n9700), .ZN(n10084) );
  INV_X1 U10832 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9703) );
  AOI22_X1 U10833 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9703), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n9702), .ZN(n10083) );
  NOR2_X1 U10834 ( .A1(n10084), .A2(n10083), .ZN(n9704) );
  NOR2_X1 U10835 ( .A1(n9705), .A2(n9704), .ZN(n10082) );
  INV_X1 U10836 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U10837 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n9707), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n9706), .ZN(n10081) );
  NOR2_X1 U10838 ( .A1(n10082), .A2(n10081), .ZN(n9708) );
  NOR2_X1 U10839 ( .A1(n9709), .A2(n9708), .ZN(n10080) );
  INV_X1 U10840 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9711) );
  AOI22_X1 U10841 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9711), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n9710), .ZN(n10079) );
  NOR2_X1 U10842 ( .A1(n10080), .A2(n10079), .ZN(n9712) );
  NOR2_X1 U10843 ( .A1(n9713), .A2(n9712), .ZN(n10078) );
  INV_X1 U10844 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9715) );
  AOI22_X1 U10845 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9715), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n9714), .ZN(n10077) );
  NOR2_X1 U10846 ( .A1(n10078), .A2(n10077), .ZN(n9716) );
  NOR2_X1 U10847 ( .A1(n9717), .A2(n9716), .ZN(n10076) );
  INV_X1 U10848 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9719) );
  AOI22_X1 U10849 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9719), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n9718), .ZN(n10075) );
  NOR2_X1 U10850 ( .A1(n10076), .A2(n10075), .ZN(n9720) );
  NOR2_X1 U10851 ( .A1(n9721), .A2(n9720), .ZN(n10074) );
  INV_X1 U10852 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9723) );
  AOI22_X1 U10853 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9723), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n9722), .ZN(n10073) );
  NOR2_X1 U10854 ( .A1(n10074), .A2(n10073), .ZN(n9724) );
  NOR2_X1 U10855 ( .A1(n9725), .A2(n9724), .ZN(n10072) );
  INV_X1 U10856 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9727) );
  AOI22_X1 U10857 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9727), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n9726), .ZN(n10071) );
  NOR2_X1 U10858 ( .A1(n10072), .A2(n10071), .ZN(n9728) );
  NOR2_X1 U10859 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  NOR2_X1 U10860 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9730), .ZN(n10067) );
  AND2_X1 U10861 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9730), .ZN(n10068) );
  NOR2_X1 U10862 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10068), .ZN(n9731) );
  NOR2_X1 U10863 ( .A1(n10067), .A2(n9731), .ZN(n9732) );
  XOR2_X1 U10864 ( .A(n9733), .B(n9732), .Z(ADD_1068_U4) );
  INV_X1 U10865 ( .A(n9734), .ZN(n9736) );
  NAND2_X1 U10866 ( .A1(n9736), .A2(n9735), .ZN(n9737) );
  OAI211_X1 U10867 ( .C1(n9739), .C2(n9738), .A(n9737), .B(n4275), .ZN(n9740)
         );
  OAI22_X1 U10868 ( .A1(n9741), .A2(n9740), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n4275), .ZN(n9742) );
  OAI21_X1 U10869 ( .B1(n9743), .B2(n10017), .A(n9742), .ZN(P2_U3219) );
  AOI22_X1 U10870 ( .A1(n10060), .A2(n5098), .B1(n9744), .B2(n10057), .ZN(
        P2_U3432) );
  INV_X1 U10871 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U10872 ( .A1(n10060), .A2(n9746), .B1(n9745), .B2(n10057), .ZN(
        P2_U3429) );
  AOI21_X1 U10873 ( .B1(n9748), .B2(n9747), .A(n4331), .ZN(n9756) );
  NOR2_X1 U10874 ( .A1(n5674), .A2(n9749), .ZN(n9750) );
  AOI211_X1 U10875 ( .C1(n9753), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9754)
         );
  OAI21_X1 U10876 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  INV_X1 U10877 ( .A(n9757), .ZN(n9758) );
  OAI21_X1 U10878 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(P1_U3217) );
  XNOR2_X1 U10879 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NOR2_X1 U10880 ( .A1(n9761), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9763) );
  OR2_X1 U10881 ( .A1(n9762), .A2(n9763), .ZN(n9765) );
  INV_X1 U10882 ( .A(n9763), .ZN(n9764) );
  MUX2_X1 U10883 ( .A(n9765), .B(n9764), .S(n5599), .Z(n9767) );
  NAND2_X1 U10884 ( .A1(n9767), .A2(n9766), .ZN(n9769) );
  AOI22_X1 U10885 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9794), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9768) );
  OAI21_X1 U10886 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(P1_U3243) );
  AOI22_X1 U10887 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9794), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9783) );
  AOI211_X1 U10888 ( .C1(n9773), .C2(n9772), .A(n9771), .B(n9784), .ZN(n9774)
         );
  AOI21_X1 U10889 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9782) );
  NOR2_X1 U10890 ( .A1(n5599), .A2(n9777), .ZN(n9780) );
  OAI211_X1 U10891 ( .C1(n9780), .C2(n9779), .A(n9789), .B(n9778), .ZN(n9781)
         );
  NAND3_X1 U10892 ( .A1(n9783), .A2(n9782), .A3(n9781), .ZN(P1_U3244) );
  AOI211_X1 U10893 ( .C1(n9787), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9800)
         );
  OAI211_X1 U10894 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9796)
         );
  INV_X1 U10895 ( .A(n9792), .ZN(n9793) );
  AOI21_X1 U10896 ( .B1(n9794), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9793), .ZN(
        n9795) );
  OAI211_X1 U10897 ( .C1(n9798), .C2(n9797), .A(n9796), .B(n9795), .ZN(n9799)
         );
  OR3_X1 U10898 ( .A1(n9801), .A2(n9800), .A3(n9799), .ZN(P1_U3247) );
  XNOR2_X1 U10899 ( .A(n9802), .B(n9804), .ZN(n9996) );
  NAND2_X1 U10900 ( .A1(n7678), .A2(n9803), .ZN(n9805) );
  XNOR2_X1 U10901 ( .A(n9805), .B(n9804), .ZN(n9806) );
  NOR2_X1 U10902 ( .A1(n9806), .A2(n9895), .ZN(n9808) );
  AOI211_X1 U10903 ( .C1(n9996), .C2(n9973), .A(n9808), .B(n9807), .ZN(n9993)
         );
  INV_X1 U10904 ( .A(n9809), .ZN(n9810) );
  AOI222_X1 U10905 ( .A1(n9811), .A2(n9906), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9898), .C1(n9899), .C2(n9810), .ZN(n9816) );
  AND2_X1 U10906 ( .A1(n9836), .A2(n9812), .ZN(n9903) );
  OAI211_X1 U10907 ( .C1(n9992), .C2(n4611), .A(n4343), .B(n9901), .ZN(n9990)
         );
  INV_X1 U10908 ( .A(n9990), .ZN(n9814) );
  AOI22_X1 U10909 ( .A1(n9996), .A2(n9903), .B1(n9905), .B2(n9814), .ZN(n9815)
         );
  OAI211_X1 U10910 ( .C1(n9898), .C2(n9993), .A(n9816), .B(n9815), .ZN(
        P1_U3282) );
  XNOR2_X1 U10911 ( .A(n9817), .B(n9820), .ZN(n9982) );
  NAND2_X1 U10912 ( .A1(n9819), .A2(n9818), .ZN(n9821) );
  XNOR2_X1 U10913 ( .A(n9821), .B(n9820), .ZN(n9822) );
  NAND2_X1 U10914 ( .A1(n9822), .A2(n9868), .ZN(n9980) );
  INV_X1 U10915 ( .A(n9823), .ZN(n9826) );
  INV_X1 U10916 ( .A(n9824), .ZN(n9825) );
  AOI21_X1 U10917 ( .B1(n9899), .B2(n9826), .A(n9825), .ZN(n9827) );
  OAI211_X1 U10918 ( .C1(n9830), .C2(n9880), .A(n9980), .B(n9827), .ZN(n9828)
         );
  AOI22_X1 U10919 ( .A1(n9982), .A2(n9874), .B1(n9828), .B2(n9836), .ZN(n9835)
         );
  OAI211_X1 U10920 ( .C1(n7563), .C2(n9830), .A(n9901), .B(n9829), .ZN(n9978)
         );
  AOI21_X1 U10921 ( .B1(n9978), .B2(n9832), .A(n9831), .ZN(n9833) );
  INV_X1 U10922 ( .A(n9833), .ZN(n9834) );
  OAI211_X1 U10923 ( .C1(n9836), .C2(n6042), .A(n9835), .B(n9834), .ZN(
        P1_U3284) );
  XNOR2_X1 U10924 ( .A(n9837), .B(n9838), .ZN(n9963) );
  XNOR2_X1 U10925 ( .A(n9839), .B(n9838), .ZN(n9840) );
  NOR2_X1 U10926 ( .A1(n9840), .A2(n9895), .ZN(n9841) );
  AOI211_X1 U10927 ( .C1(n9973), .C2(n9963), .A(n9842), .B(n9841), .ZN(n9960)
         );
  INV_X1 U10928 ( .A(n9843), .ZN(n9844) );
  AOI222_X1 U10929 ( .A1(n9845), .A2(n9906), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9898), .C1(n9844), .C2(n9899), .ZN(n9850) );
  INV_X1 U10930 ( .A(n9846), .ZN(n9847) );
  OAI211_X1 U10931 ( .C1(n9959), .C2(n4604), .A(n9847), .B(n9901), .ZN(n9958)
         );
  INV_X1 U10932 ( .A(n9958), .ZN(n9848) );
  AOI22_X1 U10933 ( .A1(n9963), .A2(n9903), .B1(n9905), .B2(n9848), .ZN(n9849)
         );
  OAI211_X1 U10934 ( .C1(n9898), .C2(n9960), .A(n9850), .B(n9849), .ZN(
        P1_U3286) );
  NAND2_X1 U10935 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  XOR2_X1 U10936 ( .A(n9861), .B(n9853), .Z(n9856) );
  INV_X1 U10937 ( .A(n9854), .ZN(n9855) );
  AOI21_X1 U10938 ( .B1(n9856), .B2(n9868), .A(n9855), .ZN(n9946) );
  INV_X1 U10939 ( .A(n9857), .ZN(n9858) );
  AOI222_X1 U10940 ( .A1(n9859), .A2(n9906), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n9898), .C1(n9858), .C2(n9899), .ZN(n9866) );
  XNOR2_X1 U10941 ( .A(n9860), .B(n9861), .ZN(n9949) );
  OAI211_X1 U10942 ( .C1(n9863), .C2(n9945), .A(n9862), .B(n9901), .ZN(n9944)
         );
  INV_X1 U10943 ( .A(n9944), .ZN(n9864) );
  AOI22_X1 U10944 ( .A1(n9949), .A2(n9874), .B1(n9905), .B2(n9864), .ZN(n9865)
         );
  OAI211_X1 U10945 ( .C1(n9898), .C2(n9946), .A(n9866), .B(n9865), .ZN(
        P1_U3288) );
  XNOR2_X1 U10946 ( .A(n6538), .B(n6007), .ZN(n9869) );
  AOI21_X1 U10947 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9931) );
  INV_X1 U10948 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9871) );
  AOI222_X1 U10949 ( .A1(n9871), .A2(n9899), .B1(n9898), .B2(
        P1_REG2_REG_3__SCAN_IN), .C1(n9870), .C2(n9906), .ZN(n9876) );
  XNOR2_X1 U10950 ( .A(n7347), .B(n6007), .ZN(n9934) );
  OAI211_X1 U10951 ( .C1(n4602), .C2(n9930), .A(n9901), .B(n9872), .ZN(n9929)
         );
  INV_X1 U10952 ( .A(n9929), .ZN(n9873) );
  AOI22_X1 U10953 ( .A1(n9934), .A2(n9874), .B1(n9905), .B2(n9873), .ZN(n9875)
         );
  OAI211_X1 U10954 ( .C1(n9898), .C2(n9931), .A(n9876), .B(n9875), .ZN(
        P1_U3290) );
  XNOR2_X1 U10955 ( .A(n9877), .B(n9881), .ZN(n9927) );
  INV_X1 U10956 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9879) );
  OAI22_X1 U10957 ( .A1(n9924), .A2(n9880), .B1(n9879), .B2(n9878), .ZN(n9885)
         );
  XNOR2_X1 U10958 ( .A(n9882), .B(n9881), .ZN(n9884) );
  OAI21_X1 U10959 ( .B1(n9884), .B2(n9895), .A(n9883), .ZN(n9925) );
  AOI211_X1 U10960 ( .C1(n9973), .C2(n9927), .A(n9885), .B(n9925), .ZN(n9890)
         );
  OAI211_X1 U10961 ( .C1(n5630), .C2(n9924), .A(n9901), .B(n9886), .ZN(n9923)
         );
  INV_X1 U10962 ( .A(n9923), .ZN(n9887) );
  AOI22_X1 U10963 ( .A1(n9927), .A2(n9903), .B1(n9905), .B2(n9887), .ZN(n9888)
         );
  OAI221_X1 U10964 ( .B1(n9898), .B2(n9890), .C1(n9836), .C2(n9889), .A(n9888), 
        .ZN(P1_U3291) );
  XNOR2_X1 U10965 ( .A(n9892), .B(n9891), .ZN(n9921) );
  XOR2_X1 U10966 ( .A(n9893), .B(n9892), .Z(n9896) );
  OAI21_X1 U10967 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9897) );
  AOI21_X1 U10968 ( .B1(n9973), .B2(n9921), .A(n9897), .ZN(n9918) );
  AOI22_X1 U10969 ( .A1(n9899), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n9898), .ZN(n9908) );
  OAI211_X1 U10970 ( .C1(n6701), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9917)
         );
  INV_X1 U10971 ( .A(n9917), .ZN(n9904) );
  AOI222_X1 U10972 ( .A1(n4278), .A2(n9906), .B1(n9905), .B2(n9904), .C1(n9921), .C2(n9903), .ZN(n9907) );
  OAI211_X1 U10973 ( .C1(n9898), .C2(n9918), .A(n9908), .B(n9907), .ZN(
        P1_U3292) );
  NOR2_X1 U10974 ( .A1(n9915), .A2(n9909), .ZN(P1_U3294) );
  AND2_X1 U10975 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9916), .ZN(P1_U3295) );
  AND2_X1 U10976 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9916), .ZN(P1_U3296) );
  AND2_X1 U10977 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9916), .ZN(P1_U3297) );
  AND2_X1 U10978 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9916), .ZN(P1_U3298) );
  AND2_X1 U10979 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9916), .ZN(P1_U3299) );
  AND2_X1 U10980 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9916), .ZN(P1_U3300) );
  NOR2_X1 U10981 ( .A1(n9915), .A2(n9910), .ZN(P1_U3301) );
  AND2_X1 U10982 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9916), .ZN(P1_U3302) );
  AND2_X1 U10983 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9916), .ZN(P1_U3303) );
  AND2_X1 U10984 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9916), .ZN(P1_U3304) );
  AND2_X1 U10985 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9916), .ZN(P1_U3305) );
  NOR2_X1 U10986 ( .A1(n9915), .A2(n9911), .ZN(P1_U3306) );
  AND2_X1 U10987 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9916), .ZN(P1_U3307) );
  NOR2_X1 U10988 ( .A1(n9915), .A2(n9912), .ZN(P1_U3308) );
  AND2_X1 U10989 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9916), .ZN(P1_U3309) );
  AND2_X1 U10990 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9916), .ZN(P1_U3310) );
  AND2_X1 U10991 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9916), .ZN(P1_U3311) );
  NOR2_X1 U10992 ( .A1(n9915), .A2(n9913), .ZN(P1_U3312) );
  NOR2_X1 U10993 ( .A1(n9915), .A2(n9914), .ZN(P1_U3313) );
  AND2_X1 U10994 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9916), .ZN(P1_U3314) );
  AND2_X1 U10995 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9916), .ZN(P1_U3315) );
  AND2_X1 U10996 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9916), .ZN(P1_U3316) );
  AND2_X1 U10997 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9916), .ZN(P1_U3317) );
  AND2_X1 U10998 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9916), .ZN(P1_U3318) );
  AND2_X1 U10999 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9916), .ZN(P1_U3319) );
  AND2_X1 U11000 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9916), .ZN(P1_U3320) );
  AND2_X1 U11001 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9916), .ZN(P1_U3321) );
  AND2_X1 U11002 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9916), .ZN(P1_U3322) );
  AND2_X1 U11003 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9916), .ZN(P1_U3323) );
  INV_X1 U11004 ( .A(n9969), .ZN(n9997) );
  OAI21_X1 U11005 ( .B1(n6701), .B2(n9991), .A(n9917), .ZN(n9920) );
  INV_X1 U11006 ( .A(n9918), .ZN(n9919) );
  AOI211_X1 U11007 ( .C1(n9997), .C2(n9921), .A(n9920), .B(n9919), .ZN(n10001)
         );
  INV_X1 U11008 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U11009 ( .A1(n10000), .A2(n10001), .B1(n9922), .B2(n9998), .ZN(
        P1_U3456) );
  OAI21_X1 U11010 ( .B1(n9924), .B2(n9991), .A(n9923), .ZN(n9926) );
  AOI211_X1 U11011 ( .C1(n9987), .C2(n9927), .A(n9926), .B(n9925), .ZN(n10003)
         );
  INV_X1 U11012 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9928) );
  AOI22_X1 U11013 ( .A1(n10000), .A2(n10003), .B1(n9928), .B2(n9998), .ZN(
        P1_U3459) );
  OAI21_X1 U11014 ( .B1(n9930), .B2(n9991), .A(n9929), .ZN(n9933) );
  INV_X1 U11015 ( .A(n9931), .ZN(n9932) );
  AOI211_X1 U11016 ( .C1(n9987), .C2(n9934), .A(n9933), .B(n9932), .ZN(n10004)
         );
  INV_X1 U11017 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U11018 ( .A1(n10000), .A2(n10004), .B1(n9935), .B2(n9998), .ZN(
        P1_U3462) );
  AOI21_X1 U11019 ( .B1(n9977), .B2(n9937), .A(n9936), .ZN(n9939) );
  OAI211_X1 U11020 ( .C1(n9941), .C2(n9940), .A(n9939), .B(n9938), .ZN(n9942)
         );
  INV_X1 U11021 ( .A(n9942), .ZN(n10006) );
  INV_X1 U11022 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U11023 ( .A1(n10000), .A2(n10006), .B1(n9943), .B2(n9998), .ZN(
        P1_U3465) );
  OAI21_X1 U11024 ( .B1(n9945), .B2(n9991), .A(n9944), .ZN(n9948) );
  INV_X1 U11025 ( .A(n9946), .ZN(n9947) );
  AOI211_X1 U11026 ( .C1(n9987), .C2(n9949), .A(n9948), .B(n9947), .ZN(n10007)
         );
  INV_X1 U11027 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U11028 ( .A1(n10000), .A2(n10007), .B1(n9950), .B2(n9998), .ZN(
        P1_U3468) );
  AND2_X1 U11029 ( .A1(n9951), .A2(n9987), .ZN(n9955) );
  OAI21_X1 U11030 ( .B1(n9953), .B2(n9991), .A(n9952), .ZN(n9954) );
  NOR3_X1 U11031 ( .A1(n9956), .A2(n9955), .A3(n9954), .ZN(n10008) );
  INV_X1 U11032 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11033 ( .A1(n10000), .A2(n10008), .B1(n9957), .B2(n9998), .ZN(
        P1_U3471) );
  OAI21_X1 U11034 ( .B1(n9959), .B2(n9991), .A(n9958), .ZN(n9962) );
  INV_X1 U11035 ( .A(n9960), .ZN(n9961) );
  AOI211_X1 U11036 ( .C1(n9997), .C2(n9963), .A(n9962), .B(n9961), .ZN(n10009)
         );
  INV_X1 U11037 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11038 ( .A1(n10000), .A2(n10009), .B1(n9964), .B2(n9998), .ZN(
        P1_U3474) );
  INV_X1 U11039 ( .A(n9970), .ZN(n9972) );
  AOI211_X1 U11040 ( .C1(n9977), .C2(n9967), .A(n9966), .B(n9965), .ZN(n9968)
         );
  OAI21_X1 U11041 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9971) );
  AOI21_X1 U11042 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(n10010) );
  INV_X1 U11043 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11044 ( .A1(n10000), .A2(n10010), .B1(n9974), .B2(n9998), .ZN(
        P1_U3477) );
  AOI21_X1 U11045 ( .B1(n9977), .B2(n9976), .A(n9975), .ZN(n9979) );
  NAND3_X1 U11046 ( .A1(n9980), .A2(n9979), .A3(n9978), .ZN(n9981) );
  AOI21_X1 U11047 ( .B1(n9982), .B2(n9987), .A(n9981), .ZN(n10011) );
  AOI22_X1 U11048 ( .A1(n10000), .A2(n10011), .B1(n9983), .B2(n9998), .ZN(
        P1_U3480) );
  OAI211_X1 U11049 ( .C1(n5674), .C2(n9991), .A(n9985), .B(n9984), .ZN(n9986)
         );
  AOI21_X1 U11050 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n10012) );
  INV_X1 U11051 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9989) );
  AOI22_X1 U11052 ( .A1(n10000), .A2(n10012), .B1(n9989), .B2(n9998), .ZN(
        P1_U3483) );
  OAI21_X1 U11053 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(n9995) );
  INV_X1 U11054 ( .A(n9993), .ZN(n9994) );
  AOI211_X1 U11055 ( .C1(n9997), .C2(n9996), .A(n9995), .B(n9994), .ZN(n10014)
         );
  INV_X1 U11056 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9999) );
  AOI22_X1 U11057 ( .A1(n10000), .A2(n10014), .B1(n9999), .B2(n9998), .ZN(
        P1_U3486) );
  AOI22_X1 U11058 ( .A1(n10015), .A2(n10001), .B1(n6925), .B2(n10013), .ZN(
        P1_U3523) );
  AOI22_X1 U11059 ( .A1(n10015), .A2(n10003), .B1(n10002), .B2(n10013), .ZN(
        P1_U3524) );
  AOI22_X1 U11060 ( .A1(n10015), .A2(n10004), .B1(n6924), .B2(n10013), .ZN(
        P1_U3525) );
  AOI22_X1 U11061 ( .A1(n10015), .A2(n10006), .B1(n10005), .B2(n10013), .ZN(
        P1_U3526) );
  AOI22_X1 U11062 ( .A1(n10015), .A2(n10007), .B1(n6013), .B2(n10013), .ZN(
        P1_U3527) );
  AOI22_X1 U11063 ( .A1(n10015), .A2(n10008), .B1(n6992), .B2(n10013), .ZN(
        P1_U3528) );
  AOI22_X1 U11064 ( .A1(n10015), .A2(n10009), .B1(n7006), .B2(n10013), .ZN(
        P1_U3529) );
  AOI22_X1 U11065 ( .A1(n10015), .A2(n10010), .B1(n7102), .B2(n10013), .ZN(
        P1_U3530) );
  AOI22_X1 U11066 ( .A1(n10015), .A2(n10011), .B1(n6041), .B2(n10013), .ZN(
        P1_U3531) );
  AOI22_X1 U11067 ( .A1(n10015), .A2(n10012), .B1(n7294), .B2(n10013), .ZN(
        P1_U3532) );
  AOI22_X1 U11068 ( .A1(n10015), .A2(n10014), .B1(n7435), .B2(n10013), .ZN(
        P1_U3533) );
  MUX2_X1 U11069 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10016), .S(n4275), .Z(
        n10022) );
  OAI22_X1 U11070 ( .A1(n10020), .A2(n10019), .B1(n10018), .B2(n10017), .ZN(
        n10021) );
  NOR2_X1 U11071 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  OAI21_X1 U11072 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(P2_U3227) );
  AOI222_X1 U11073 ( .A1(n10031), .A2(n10030), .B1(n10029), .B2(n10028), .C1(
        n10027), .C2(n10026), .ZN(n10032) );
  OAI221_X1 U11074 ( .B1(n10034), .B2(n10033), .C1(n4275), .C2(n5446), .A(
        n10032), .ZN(P2_U3229) );
  INV_X1 U11075 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U11076 ( .A1(n10060), .A2(n10036), .B1(n10035), .B2(n10057), .ZN(
        P2_U3390) );
  AOI22_X1 U11077 ( .A1(n10060), .A2(n4921), .B1(n10037), .B2(n10057), .ZN(
        P2_U3393) );
  AOI22_X1 U11078 ( .A1(n10060), .A2(n4953), .B1(n10038), .B2(n10057), .ZN(
        P2_U3396) );
  INV_X1 U11079 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11080 ( .A1(n10060), .A2(n10040), .B1(n10039), .B2(n10057), .ZN(
        P2_U3399) );
  INV_X1 U11081 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U11082 ( .A1(n10060), .A2(n10042), .B1(n10041), .B2(n10057), .ZN(
        P2_U3402) );
  INV_X1 U11083 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U11084 ( .A1(n10060), .A2(n10044), .B1(n10043), .B2(n10057), .ZN(
        P2_U3405) );
  INV_X1 U11085 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U11086 ( .A1(n10060), .A2(n10046), .B1(n10045), .B2(n10057), .ZN(
        P2_U3408) );
  INV_X1 U11087 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10048) );
  AOI22_X1 U11088 ( .A1(n10060), .A2(n10048), .B1(n10047), .B2(n10057), .ZN(
        P2_U3411) );
  INV_X1 U11089 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U11090 ( .A1(n10060), .A2(n10050), .B1(n10049), .B2(n10057), .ZN(
        P2_U3414) );
  AOI22_X1 U11091 ( .A1(n10060), .A2(n10052), .B1(n10051), .B2(n10057), .ZN(
        P2_U3417) );
  INV_X1 U11092 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10054) );
  AOI22_X1 U11093 ( .A1(n10060), .A2(n10054), .B1(n10053), .B2(n10057), .ZN(
        P2_U3420) );
  INV_X1 U11094 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11095 ( .A1(n10060), .A2(n10056), .B1(n10055), .B2(n10057), .ZN(
        P2_U3423) );
  INV_X1 U11096 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U11097 ( .A1(n10060), .A2(n10059), .B1(n10058), .B2(n10057), .ZN(
        P2_U3426) );
  NOR2_X1 U11098 ( .A1(n10062), .A2(n10061), .ZN(n10063) );
  XOR2_X1 U11099 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10063), .Z(ADD_1068_U5) );
  AOI21_X1 U11100 ( .B1(n10066), .B2(n10065), .A(n10064), .ZN(ADD_1068_U46) );
  NOR2_X1 U11101 ( .A1(n10068), .A2(n10067), .ZN(n10070) );
  XNOR2_X1 U11102 ( .A(n10070), .B(n10069), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11103 ( .A(n10072), .B(n10071), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11104 ( .A(n10074), .B(n10073), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11105 ( .A(n10076), .B(n10075), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11106 ( .A(n10078), .B(n10077), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11107 ( .A(n10080), .B(n10079), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11108 ( .A(n10082), .B(n10081), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11109 ( .A(n10084), .B(n10083), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11110 ( .A(n10086), .B(n10085), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11111 ( .A(n10088), .B(n10087), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11112 ( .A(n10090), .B(n10089), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11113 ( .A(n10092), .B(n10091), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11114 ( .A(n10094), .B(n10093), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11115 ( .A(n10096), .B(n10095), .ZN(ADD_1068_U48) );
  XOR2_X1 U11116 ( .A(n10098), .B(n10097), .Z(ADD_1068_U54) );
  XOR2_X1 U11117 ( .A(n10100), .B(n10099), .Z(ADD_1068_U53) );
  XNOR2_X1 U11118 ( .A(n10102), .B(n10101), .ZN(ADD_1068_U52) );
  INV_X2 U4786 ( .A(n8318), .ZN(n4959) );
  CLKBUF_X1 U4784 ( .A(n5994), .Z(n6249) );
endmodule

