

module b22_C_SARLock_k_128_1 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6559, n6560, n6561, n6562, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473;

  AND3_X1 U7308 ( .A1(n12297), .A2(n12339), .A3(n12296), .ZN(n12344) );
  INV_X1 U7309 ( .A(n6627), .ZN(n7025) );
  INV_X4 U7310 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  OR2_X1 U7311 ( .A1(n12953), .A2(n12958), .ZN(n12955) );
  NAND2_X1 U7312 ( .A1(n9008), .A2(n9007), .ZN(n13586) );
  CLKBUF_X2 U7313 ( .A(n12877), .Z(n6973) );
  AND2_X1 U7314 ( .A1(n9652), .A2(n9653), .ZN(n11716) );
  INV_X1 U7315 ( .A(n7887), .ZN(n8247) );
  CLKBUF_X2 U7316 ( .A(n9433), .Z(n12259) );
  INV_X1 U7317 ( .A(n12264), .ZN(n9631) );
  AND3_X1 U7318 ( .A1(n8979), .A2(n8343), .A3(n8342), .ZN(n9993) );
  NOR2_X1 U7319 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9265) );
  AOI21_X1 U7320 ( .B1(n7293), .B2(n7298), .A(n12012), .ZN(n7291) );
  INV_X1 U7321 ( .A(n12256), .ZN(n12293) );
  AND2_X1 U7322 ( .A1(n7295), .A2(n6704), .ZN(n7293) );
  NAND2_X1 U7323 ( .A1(n9732), .A2(n11185), .ZN(n6567) );
  INV_X1 U7324 ( .A(n12396), .ZN(n12464) );
  INV_X1 U7325 ( .A(n7841), .ZN(n8222) );
  AND2_X1 U7326 ( .A1(n12761), .A2(n12630), .ZN(n12746) );
  INV_X1 U7327 ( .A(n8214), .ZN(n8191) );
  INV_X1 U7328 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8285) );
  AOI22_X1 U7329 ( .A1(n13826), .A2(n13827), .B1(n12384), .B2(n12383), .ZN(
        n13755) );
  NAND2_X1 U7330 ( .A1(n14364), .A2(n9284), .ZN(n12266) );
  INV_X1 U7331 ( .A(n12266), .ZN(n9718) );
  INV_X1 U7332 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9411) );
  AND2_X1 U7333 ( .A1(n6756), .A2(n9134), .ZN(n10335) );
  XNOR2_X1 U7334 ( .A(n7315), .B(n14986), .ZN(n14977) );
  AND2_X1 U7335 ( .A1(n11896), .A2(n11716), .ZN(n9655) );
  NAND2_X1 U7336 ( .A1(n7167), .A2(n9611), .ZN(n14265) );
  NAND2_X1 U7337 ( .A1(n12440), .A2(n12439), .ZN(n13746) );
  AND2_X1 U7338 ( .A1(n9432), .A2(n9431), .ZN(n14530) );
  OR2_X1 U7339 ( .A1(n6785), .A2(n6783), .ZN(n13860) );
  INV_X1 U7340 ( .A(n9926), .ZN(n6559) );
  OR2_X4 U7341 ( .A1(n8194), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n6599) );
  AND2_X2 U7342 ( .A1(n12900), .A2(n13138), .ZN(n8280) );
  OR2_X2 U7343 ( .A1(n14922), .A2(n7305), .ZN(n7304) );
  OAI21_X2 U7344 ( .B1(n8613), .B2(n7095), .A(n7092), .ZN(n8731) );
  NAND2_X2 U7345 ( .A1(n7516), .A2(n7518), .ZN(n8613) );
  OAI211_X2 U7346 ( .C1(n12039), .C2(n12038), .A(n6908), .B(n6907), .ZN(n13585) );
  OAI22_X2 U7347 ( .A1(n10974), .A2(n10973), .B1(n10972), .B2(n14796), .ZN(
        n11139) );
  NOR2_X2 U7348 ( .A1(n11255), .A2(n13667), .ZN(n11431) );
  XNOR2_X1 U7349 ( .A(n11007), .B(n11039), .ZN(n14906) );
  NAND2_X1 U7350 ( .A1(n11006), .A2(n11005), .ZN(n11007) );
  XNOR2_X2 U7351 ( .A(n6802), .B(n9279), .ZN(n9282) );
  AND2_X4 U7352 ( .A1(n8373), .A2(n12067), .ZN(n9931) );
  INV_X1 U7353 ( .A(n14831), .ZN(n10776) );
  NAND2_X2 U7354 ( .A1(n9132), .A2(n9131), .ZN(n9139) );
  AND2_X2 U7355 ( .A1(n9251), .A2(n9130), .ZN(n9131) );
  XNOR2_X2 U7356 ( .A(n8372), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8383) );
  NOR2_X4 U7357 ( .A1(n7591), .A2(n7592), .ZN(n9506) );
  NAND2_X1 U7358 ( .A1(n10350), .A2(n6987), .ZN(n10439) );
  XNOR2_X2 U7359 ( .A(n7436), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8377) );
  NAND2_X2 U7360 ( .A1(n14955), .A2(n11012), .ZN(n7315) );
  CLKBUF_X2 U7362 ( .A(n9740), .Z(n6560) );
  OAI211_X1 U7363 ( .C1(n8821), .C2(n10051), .A(n8369), .B(n8368), .ZN(n9740)
         );
  NAND2_X1 U7364 ( .A1(n7730), .A2(n13207), .ZN(n6561) );
  NOR2_X2 U7365 ( .A1(n11640), .A2(n11641), .ZN(n11643) );
  NOR2_X2 U7366 ( .A1(n11457), .A2(n7982), .ZN(n11640) );
  AOI21_X2 U7367 ( .B1(n14106), .B2(n14105), .A(n9706), .ZN(n14083) );
  NAND2_X2 U7368 ( .A1(n14124), .A2(n9705), .ZN(n14106) );
  INV_X1 U7369 ( .A(n11022), .ZN(n6562) );
  INV_X1 U7371 ( .A(n6562), .ZN(n6564) );
  AOI21_X2 U7372 ( .B1(n14544), .B2(n9082), .A(n14541), .ZN(n14547) );
  XNOR2_X2 U7373 ( .A(n9067), .B(n9068), .ZN(n14393) );
  NAND2_X2 U7374 ( .A1(n7080), .A2(n9066), .ZN(n9067) );
  AOI21_X1 U7375 ( .B1(n7023), .B2(n7025), .A(n7022), .ZN(n7021) );
  AND2_X1 U7376 ( .A1(n7024), .A2(n15130), .ZN(n7023) );
  OR2_X1 U7377 ( .A1(n7025), .A2(n13138), .ZN(n7024) );
  NAND2_X1 U7378 ( .A1(n7090), .A2(n7089), .ZN(n12014) );
  CLKBUF_X1 U7379 ( .A(n13289), .Z(n6977) );
  OAI21_X1 U7380 ( .B1(n8871), .B2(n7420), .A(n8893), .ZN(n7419) );
  OR2_X1 U7381 ( .A1(n13496), .A2(n13495), .ZN(n13620) );
  XNOR2_X1 U7382 ( .A(n9628), .B(n9627), .ZN(n12048) );
  AND2_X1 U7383 ( .A1(n7317), .A2(n6752), .ZN(n14460) );
  NAND2_X1 U7384 ( .A1(n8898), .A2(n8897), .ZN(n13603) );
  NAND2_X1 U7385 ( .A1(n10895), .A2(n7917), .ZN(n11114) );
  NAND2_X1 U7386 ( .A1(n6803), .A2(n10439), .ZN(n6804) );
  NAND2_X1 U7387 ( .A1(n9437), .A2(n9436), .ZN(n14401) );
  INV_X1 U7388 ( .A(n12394), .ZN(n12462) );
  NAND2_X1 U7389 ( .A1(n13859), .A2(n10441), .ZN(n12106) );
  INV_X1 U7390 ( .A(n13856), .ZN(n11204) );
  INV_X1 U7391 ( .A(n13860), .ZN(n7583) );
  INV_X1 U7392 ( .A(n14837), .ZN(n10795) );
  INV_X1 U7393 ( .A(n13321), .ZN(n10659) );
  INV_X1 U7394 ( .A(n13323), .ZN(n10801) );
  INV_X4 U7395 ( .A(n9749), .ZN(n9880) );
  INV_X4 U7396 ( .A(n9749), .ZN(n9937) );
  AND4_X1 U7397 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(n10596)
         );
  INV_X4 U7398 ( .A(n9743), .ZN(n9906) );
  CLKBUF_X1 U7399 ( .A(n7836), .Z(n7489) );
  NOR2_X2 U7400 ( .A1(n10644), .A2(n9993), .ZN(n9743) );
  INV_X4 U7401 ( .A(n12746), .ZN(n12750) );
  INV_X4 U7402 ( .A(n8463), .ZN(n6565) );
  AND2_X1 U7403 ( .A1(n12273), .A2(n12275), .ZN(n12288) );
  XNOR2_X1 U7404 ( .A(n9291), .B(n9290), .ZN(n14370) );
  INV_X2 U7405 ( .A(n8417), .ZN(n6566) );
  OAI21_X1 U7406 ( .B1(n12753), .B2(n12752), .A(n12751), .ZN(n7158) );
  AND2_X1 U7407 ( .A1(n13588), .A2(n13587), .ZN(n6990) );
  OAI21_X1 U7408 ( .B1(n7066), .B2(n13063), .A(n8255), .ZN(n12901) );
  AOI21_X1 U7409 ( .B1(n9856), .B2(n6636), .A(n7676), .ZN(n9866) );
  OR2_X1 U7410 ( .A1(n9951), .A2(n6663), .ZN(n6579) );
  NAND2_X1 U7411 ( .A1(n7035), .A2(n7375), .ZN(n12909) );
  NAND2_X1 U7412 ( .A1(n7378), .A2(n7377), .ZN(n12926) );
  AND2_X1 U7413 ( .A1(n7294), .A2(n7293), .ZN(n13427) );
  NOR2_X1 U7414 ( .A1(n7150), .A2(n7380), .ZN(n7374) );
  NAND2_X1 U7415 ( .A1(n13458), .A2(n12033), .ZN(n13440) );
  NAND2_X1 U7416 ( .A1(n13796), .A2(n13797), .ZN(n13795) );
  INV_X1 U7417 ( .A(n6993), .ZN(n6761) );
  AND2_X1 U7418 ( .A1(n12843), .A2(n12857), .ZN(n6993) );
  XNOR2_X1 U7419 ( .A(n12842), .B(n14466), .ZN(n14475) );
  OR2_X1 U7420 ( .A1(n13084), .A2(n8228), .ZN(n12747) );
  NOR2_X1 U7421 ( .A1(n6608), .A2(n7389), .ZN(n7388) );
  NAND2_X1 U7422 ( .A1(n8193), .A2(n8192), .ZN(n12960) );
  OR2_X1 U7423 ( .A1(n12994), .A2(n7012), .ZN(n7006) );
  NAND2_X1 U7424 ( .A1(n8178), .A2(n8177), .ZN(n12531) );
  NAND2_X1 U7425 ( .A1(n7303), .A2(n12000), .ZN(n13566) );
  NAND2_X1 U7426 ( .A1(n7318), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U7427 ( .A1(n7628), .A2(n7627), .ZN(n12076) );
  AOI21_X1 U7428 ( .B1(n6603), .B2(n12321), .A(n7350), .ZN(n7349) );
  AND2_X1 U7429 ( .A1(n6899), .A2(n12026), .ZN(n6898) );
  NAND2_X1 U7430 ( .A1(n8696), .A2(n8695), .ZN(n11937) );
  NAND2_X1 U7431 ( .A1(n11630), .A2(n12773), .ZN(n6772) );
  NAND2_X1 U7432 ( .A1(n11780), .A2(n12700), .ZN(n11930) );
  AOI21_X1 U7433 ( .B1(n11429), .B2(n11428), .A(n11427), .ZN(n11686) );
  OAI21_X1 U7434 ( .B1(n6835), .B2(n6834), .A(n6833), .ZN(n9796) );
  OAI21_X1 U7435 ( .B1(n11248), .B2(n11247), .A(n11249), .ZN(n11429) );
  OAI21_X1 U7436 ( .B1(n11346), .B2(n7508), .A(n7505), .ZN(n11588) );
  OR2_X1 U7437 ( .A1(n11859), .A2(n11884), .ZN(n11889) );
  NAND2_X1 U7438 ( .A1(n11281), .A2(n7961), .ZN(n11282) );
  NAND2_X1 U7439 ( .A1(n11114), .A2(n12596), .ZN(n11113) );
  NAND2_X1 U7440 ( .A1(n7550), .A2(n6628), .ZN(n10932) );
  NAND2_X1 U7441 ( .A1(n6804), .A2(n7547), .ZN(n7550) );
  AND2_X1 U7442 ( .A1(n11560), .A2(n11561), .ZN(n7560) );
  AND2_X1 U7443 ( .A1(n10690), .A2(n7903), .ZN(n10897) );
  NAND4_X1 U7444 ( .A1(n8227), .A2(n8226), .A3(n8225), .A4(n8224), .ZN(n12913)
         );
  NOR2_X1 U7445 ( .A1(n11550), .A2(n7557), .ZN(n7556) );
  NAND2_X1 U7446 ( .A1(n7004), .A2(n12654), .ZN(n10894) );
  NAND2_X1 U7447 ( .A1(n10860), .A2(n10859), .ZN(n10858) );
  NOR2_X1 U7448 ( .A1(n6615), .A2(n6992), .ZN(n11016) );
  NAND2_X1 U7449 ( .A1(n10871), .A2(n7868), .ZN(n10860) );
  OAI21_X2 U7450 ( .B1(n9011), .B2(n10712), .A(n13571), .ZN(n13302) );
  NAND2_X1 U7451 ( .A1(n7440), .A2(n7439), .ZN(n14620) );
  AND2_X1 U7452 ( .A1(n12654), .A2(n12649), .ZN(n12652) );
  OR2_X1 U7453 ( .A1(n14958), .A2(n14957), .ZN(n14955) );
  INV_X1 U7454 ( .A(n10771), .ZN(n10768) );
  INV_X1 U7455 ( .A(n14684), .ZN(n12115) );
  AND2_X1 U7456 ( .A1(n6989), .A2(n10492), .ZN(n15060) );
  INV_X1 U7457 ( .A(n10708), .ZN(n10441) );
  NOR2_X1 U7458 ( .A1(n9058), .A2(n9059), .ZN(n9060) );
  INV_X2 U7459 ( .A(n8410), .ZN(n8964) );
  NAND2_X1 U7460 ( .A1(n6666), .A2(n7845), .ZN(n15063) );
  INV_X1 U7461 ( .A(n14672), .ZN(n12100) );
  AND4_X1 U7462 ( .A1(n7306), .A2(n8426), .A3(n8424), .A4(n8425), .ZN(n10610)
         );
  NAND2_X1 U7463 ( .A1(n8421), .A2(n8420), .ZN(n14837) );
  AOI21_X1 U7464 ( .B1(n6949), .B2(n6948), .A(n9032), .ZN(n9061) );
  NAND2_X1 U7465 ( .A1(n10344), .A2(n14014), .ZN(n14631) );
  INV_X2 U7466 ( .A(n7489), .ZN(n8113) );
  AND4_X1 U7467 ( .A1(n9301), .A2(n9300), .A3(n9299), .A4(n9298), .ZN(n10741)
         );
  NAND2_X1 U7468 ( .A1(n12883), .A2(n10577), .ZN(n9251) );
  NAND2_X1 U7469 ( .A1(n10647), .A2(n11176), .ZN(n8811) );
  XNOR2_X1 U7470 ( .A(n9732), .B(n9993), .ZN(n13402) );
  OR2_X2 U7471 ( .A1(n12286), .A2(n12273), .ZN(n14242) );
  NAND2_X1 U7472 ( .A1(n9653), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U7473 ( .A1(n6825), .A2(n6824), .ZN(n10723) );
  NAND2_X1 U7474 ( .A1(n12759), .A2(n12877), .ZN(n7836) );
  NAND2_X1 U7475 ( .A1(n8112), .A2(n8242), .ZN(n12883) );
  NAND2_X2 U7476 ( .A1(n9284), .A2(n9283), .ZN(n9598) );
  OAI21_X1 U7477 ( .B1(n7747), .B2(n6609), .A(n7224), .ZN(n7942) );
  NAND2_X1 U7478 ( .A1(n9282), .A2(n9283), .ZN(n12264) );
  NAND2_X1 U7479 ( .A1(n8394), .A2(n10006), .ZN(n8821) );
  AND2_X1 U7480 ( .A1(n12067), .A2(n13696), .ZN(n8576) );
  INV_X1 U7481 ( .A(n9283), .ZN(n14364) );
  INV_X2 U7482 ( .A(n8394), .ZN(n10141) );
  XNOR2_X1 U7483 ( .A(n6881), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U7484 ( .A1(n7807), .A2(n7806), .ZN(n12759) );
  XNOR2_X1 U7485 ( .A(n8288), .B(n8287), .ZN(n11422) );
  NAND2_X1 U7486 ( .A1(n9012), .A2(n12050), .ZN(n8394) );
  AND2_X1 U7487 ( .A1(n7723), .A2(n7395), .ZN(n7729) );
  NAND2_X1 U7488 ( .A1(n9529), .A2(n9641), .ZN(n14014) );
  NOR2_X1 U7489 ( .A1(n9049), .A2(n14378), .ZN(n15469) );
  OAI21_X1 U7490 ( .B1(n8290), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8291) );
  XNOR2_X1 U7491 ( .A(n8244), .B(n8243), .ZN(n10577) );
  OR2_X1 U7492 ( .A1(n9012), .A2(n10006), .ZN(n6889) );
  XNOR2_X1 U7493 ( .A(n9639), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14371) );
  XNOR2_X1 U7494 ( .A(n9640), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12273) );
  XNOR2_X1 U7495 ( .A(n7280), .B(n8371), .ZN(n13696) );
  NOR2_X1 U7496 ( .A1(n8337), .A2(n8345), .ZN(n8967) );
  OR2_X1 U7497 ( .A1(n8009), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U7498 ( .A1(n8337), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7436) );
  XNOR2_X1 U7499 ( .A(n7721), .B(n7720), .ZN(n12365) );
  NAND2_X1 U7500 ( .A1(n14358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6802) );
  OR2_X1 U7501 ( .A1(n8286), .A2(n8285), .ZN(n8288) );
  NAND2_X1 U7502 ( .A1(n8370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6965) );
  OR2_X1 U7503 ( .A1(n8240), .A2(n7645), .ZN(n8317) );
  NAND2_X2 U7504 ( .A1(n10025), .A2(P1_U3086), .ZN(n14366) );
  AOI21_X1 U7505 ( .B1(n8971), .B2(n8359), .A(n8358), .ZN(n8363) );
  OAI21_X1 U7506 ( .B1(n9050), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6673), .ZN(
        n7072) );
  NOR2_X1 U7507 ( .A1(n8240), .A2(n7642), .ZN(n8286) );
  XNOR2_X1 U7508 ( .A(n8341), .B(n8334), .ZN(n11176) );
  NAND2_X1 U7509 ( .A1(n13691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8372) );
  OAI21_X1 U7510 ( .B1(n9643), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U7511 ( .A1(n7281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7280) );
  INV_X4 U7512 ( .A(n6566), .ZN(n10006) );
  NAND2_X1 U7513 ( .A1(n8971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U7514 ( .A1(n8352), .A2(n8348), .ZN(n8971) );
  NOR2_X1 U7515 ( .A1(n8970), .A2(n8350), .ZN(n8351) );
  AND2_X1 U7516 ( .A1(n7713), .A2(n8110), .ZN(n7716) );
  NAND2_X1 U7517 ( .A1(n7169), .A2(n7168), .ZN(n8417) );
  AOI21_X1 U7518 ( .B1(n9043), .B2(n7257), .A(n7254), .ZN(n9040) );
  NAND2_X1 U7519 ( .A1(n7834), .A2(n7835), .ZN(n6940) );
  AND2_X1 U7520 ( .A1(n9274), .A2(n9504), .ZN(n9505) );
  AND2_X1 U7521 ( .A1(n7711), .A2(n7972), .ZN(n7976) );
  INV_X1 U7522 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7972) );
  INV_X1 U7523 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7812) );
  INV_X1 U7524 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n15400) );
  INV_X1 U7525 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n15399) );
  INV_X1 U7526 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9406) );
  NOR2_X1 U7527 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6807) );
  INV_X1 U7528 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8592) );
  NOR2_X1 U7529 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8329) );
  INV_X1 U7530 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7878) );
  INV_X1 U7531 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6809) );
  INV_X1 U7532 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9263) );
  INV_X1 U7533 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8340) );
  INV_X1 U7534 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7814) );
  INV_X4 U7535 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7536 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7649) );
  INV_X1 U7537 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7815) );
  NOR2_X1 U7538 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8331) );
  INV_X1 U7539 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9267) );
  XNOR2_X1 U7540 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7875) );
  INV_X4 U7541 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7542 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8287) );
  INV_X1 U7543 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7995) );
  INV_X1 U7544 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n15406) );
  NOR2_X1 U7545 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7707) );
  NOR2_X4 U7546 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7833) );
  NAND2_X4 U7547 ( .A1(n12464), .A2(n14631), .ZN(n12394) );
  OAI21_X2 U7548 ( .B1(n10563), .B2(n7622), .A(n7618), .ZN(n10888) );
  NAND2_X1 U7549 ( .A1(n10474), .A2(n9146), .ZN(n10563) );
  AOI21_X2 U7550 ( .B1(n14048), .B2(n14047), .A(n9708), .ZN(n14032) );
  AOI22_X2 U7551 ( .A1(n13470), .A2(n13478), .B1(n13475), .B2(n13484), .ZN(
        n13455) );
  OAI22_X2 U7552 ( .A1(n12031), .A2(n13482), .B1(n13237), .B2(n13621), .ZN(
        n13470) );
  XNOR2_X2 U7553 ( .A(n12382), .B(n12383), .ZN(n13826) );
  NOR2_X2 U7554 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7885) );
  INV_X1 U7555 ( .A(n12352), .ZN(n6568) );
  NAND2_X1 U7556 ( .A1(n10647), .A2(n11176), .ZN(n6569) );
  INV_X2 U7557 ( .A(n10442), .ZN(n12455) );
  NOR2_X2 U7558 ( .A1(n7918), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7934) );
  OR2_X2 U7559 ( .A1(n7904), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7918) );
  NOR2_X2 U7560 ( .A1(n8066), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8081) );
  OR2_X2 U7561 ( .A1(n8045), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8066) );
  OR2_X2 U7562 ( .A1(n7841), .A2(n12946), .ZN(n8209) );
  NOR2_X4 U7563 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n6599), .ZN(n8218) );
  NAND2_X1 U7564 ( .A1(n7151), .A2(n12968), .ZN(n7149) );
  INV_X1 U7565 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9269) );
  AOI21_X1 U7566 ( .B1(n7050), .B2(n7048), .A(n7047), .ZN(n7046) );
  INV_X1 U7567 ( .A(n7052), .ZN(n7048) );
  NAND2_X1 U7568 ( .A1(n13242), .A2(n6646), .ZN(n13289) );
  INV_X1 U7569 ( .A(n13292), .ZN(n6872) );
  INV_X1 U7570 ( .A(n8821), .ZN(n8434) );
  OAI21_X1 U7571 ( .B1(n8815), .B2(n8817), .A(n6854), .ZN(n7531) );
  INV_X1 U7572 ( .A(n6855), .ZN(n6854) );
  OAI21_X1 U7573 ( .B1(n8814), .B2(n8817), .A(n7532), .ZN(n6855) );
  AND2_X1 U7574 ( .A1(n7542), .A2(n6853), .ZN(n6852) );
  NAND2_X1 U7575 ( .A1(n8752), .A2(n10407), .ZN(n8753) );
  AOI21_X1 U7576 ( .B1(n6859), .B2(n6857), .A(n6856), .ZN(n8752) );
  NOR2_X1 U7577 ( .A1(n8750), .A2(n10382), .ZN(n6856) );
  AND2_X1 U7578 ( .A1(n8710), .A2(n6858), .ZN(n6857) );
  NAND2_X1 U7579 ( .A1(n8750), .A2(n10382), .ZN(n6858) );
  AOI21_X1 U7580 ( .B1(n7177), .B2(n7094), .A(n7093), .ZN(n7092) );
  INV_X1 U7581 ( .A(n7525), .ZN(n7093) );
  AND2_X1 U7582 ( .A1(n8710), .A2(n8709), .ZN(n8732) );
  NAND2_X1 U7583 ( .A1(n6782), .A2(n7268), .ZN(n7271) );
  AND2_X1 U7584 ( .A1(n7267), .A2(n6597), .ZN(n6782) );
  AND2_X1 U7585 ( .A1(n6618), .A2(n7488), .ZN(n7396) );
  INV_X1 U7586 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7488) );
  INV_X1 U7587 ( .A(n9545), .ZN(n9433) );
  NAND2_X1 U7588 ( .A1(n9305), .A2(n6566), .ZN(n9545) );
  OR2_X1 U7589 ( .A1(n9771), .A2(n9772), .ZN(n7669) );
  NAND2_X1 U7590 ( .A1(n6831), .A2(n9831), .ZN(n9834) );
  NAND2_X1 U7591 ( .A1(n6828), .A2(n6826), .ZN(n6831) );
  AOI21_X1 U7592 ( .B1(n9850), .B2(n9849), .A(n9847), .ZN(n9848) );
  INV_X1 U7593 ( .A(n7681), .ZN(n7680) );
  OAI21_X1 U7594 ( .B1(n7682), .B2(n7684), .A(n9861), .ZN(n7681) );
  NAND2_X1 U7595 ( .A1(n12258), .A2(n7115), .ZN(n7114) );
  INV_X1 U7596 ( .A(n7145), .ZN(n7142) );
  AND2_X1 U7597 ( .A1(n11046), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7305) );
  AOI21_X1 U7598 ( .B1(n7376), .B2(n12934), .A(n6656), .ZN(n7375) );
  NAND2_X1 U7599 ( .A1(n12955), .A2(n7374), .ZN(n7035) );
  OR2_X1 U7600 ( .A1(n12986), .A2(n8173), .ZN(n12736) );
  NOR2_X1 U7601 ( .A1(n12592), .A2(n7514), .ZN(n7513) );
  INV_X1 U7602 ( .A(n12691), .ZN(n7514) );
  AOI21_X1 U7603 ( .B1(n7371), .B2(n7373), .A(n7369), .ZN(n7368) );
  OAI21_X1 U7604 ( .B1(n8261), .B2(n7947), .A(n6741), .ZN(n11279) );
  AOI21_X1 U7605 ( .B1(n12665), .B2(n6743), .A(n6742), .ZN(n6741) );
  INV_X1 U7606 ( .A(n12662), .ZN(n6743) );
  INV_X1 U7607 ( .A(n12666), .ZN(n6742) );
  OR2_X1 U7608 ( .A1(n12905), .A2(n12765), .ZN(n12612) );
  INV_X1 U7609 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7709) );
  AND2_X1 U7610 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  INV_X1 U7611 ( .A(n7993), .ZN(n7239) );
  INV_X1 U7612 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U7613 ( .A1(n7742), .A2(n7743), .ZN(n7223) );
  NAND2_X1 U7614 ( .A1(n6821), .A2(n6818), .ZN(n9883) );
  INV_X1 U7615 ( .A(n7293), .ZN(n7292) );
  NOR2_X1 U7616 ( .A1(n13488), .A2(n13621), .ZN(n6891) );
  NOR2_X1 U7617 ( .A1(n13635), .A2(n7133), .ZN(n7131) );
  INV_X1 U7618 ( .A(n13565), .ZN(n7353) );
  NAND2_X1 U7619 ( .A1(n14837), .A2(n10610), .ZN(n10622) );
  INV_X1 U7620 ( .A(n11812), .ZN(n6798) );
  NAND2_X1 U7621 ( .A1(n7325), .A2(n6614), .ZN(n7189) );
  AOI21_X1 U7622 ( .B1(n7602), .B2(n14174), .A(n6581), .ZN(n7600) );
  OR2_X1 U7623 ( .A1(n14165), .A2(n7601), .ZN(n6887) );
  INV_X1 U7624 ( .A(n7602), .ZN(n7601) );
  NAND2_X1 U7625 ( .A1(n6873), .A2(n7605), .ZN(n14229) );
  AOI21_X1 U7626 ( .B1(n7606), .B2(n14517), .A(n6660), .ZN(n7605) );
  NAND2_X1 U7627 ( .A1(n14516), .A2(n7606), .ZN(n6873) );
  AOI21_X1 U7628 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(n10354) );
  NAND2_X1 U7629 ( .A1(n6880), .A2(n6648), .ZN(n9280) );
  INV_X1 U7630 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9270) );
  AND4_X1 U7631 ( .A1(n9313), .A2(n9268), .A3(n9504), .A4(n9267), .ZN(n7437)
         );
  NAND2_X1 U7632 ( .A1(n8545), .A2(n8544), .ZN(n8565) );
  NAND2_X1 U7633 ( .A1(n7165), .A2(n8478), .ZN(n8499) );
  NAND2_X1 U7634 ( .A1(n8476), .A2(n8475), .ZN(n7165) );
  AND2_X1 U7635 ( .A1(n9218), .A2(n7617), .ZN(n7616) );
  OR2_X1 U7636 ( .A1(n12568), .A2(n9217), .ZN(n7617) );
  NAND2_X1 U7637 ( .A1(n6758), .A2(n6757), .ZN(n6756) );
  INV_X1 U7638 ( .A(n12351), .ZN(n6758) );
  NAND2_X1 U7639 ( .A1(n9137), .A2(n9136), .ZN(n6757) );
  XNOR2_X1 U7640 ( .A(n7304), .B(n11053), .ZN(n14943) );
  NOR2_X1 U7641 ( .A1(n14943), .A2(n11051), .ZN(n14942) );
  INV_X1 U7642 ( .A(n14997), .ZN(n6773) );
  XNOR2_X1 U7643 ( .A(n11016), .B(n15022), .ZN(n15018) );
  NOR2_X1 U7644 ( .A1(n15018), .A2(n11077), .ZN(n15017) );
  NAND2_X1 U7645 ( .A1(n7302), .A2(n7301), .ZN(n7300) );
  NAND2_X1 U7646 ( .A1(n11462), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7301) );
  NAND2_X1 U7647 ( .A1(n6964), .A2(n6737), .ZN(n7268) );
  INV_X1 U7648 ( .A(n11905), .ZN(n6964) );
  NAND2_X1 U7649 ( .A1(n12793), .A2(n12804), .ZN(n12827) );
  NAND2_X1 U7650 ( .A1(n13018), .A2(n13017), .ZN(n7387) );
  AND2_X1 U7651 ( .A1(n7043), .A2(n6690), .ZN(n7042) );
  NAND2_X1 U7652 ( .A1(n13067), .A2(n7051), .ZN(n8268) );
  NAND2_X1 U7653 ( .A1(n8052), .A2(n6711), .ZN(n7391) );
  NAND2_X1 U7654 ( .A1(n7038), .A2(n7382), .ZN(n7037) );
  NOR2_X1 U7655 ( .A1(n12685), .A2(n7383), .ZN(n7382) );
  NAND2_X1 U7656 ( .A1(n6602), .A2(n7040), .ZN(n7038) );
  NAND2_X1 U7657 ( .A1(n11113), .A2(n7393), .ZN(n11281) );
  AND2_X1 U7658 ( .A1(n7947), .A2(n7933), .ZN(n7393) );
  NOR2_X1 U7659 ( .A1(n10532), .A2(n15124), .ZN(n10489) );
  NAND2_X1 U7660 ( .A1(n10492), .A2(n15062), .ZN(n15065) );
  INV_X1 U7661 ( .A(n15050), .ZN(n15064) );
  AND3_X1 U7662 ( .A1(n10554), .A2(n7489), .A3(n12746), .ZN(n15061) );
  NAND2_X1 U7663 ( .A1(n7806), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U7664 ( .A1(n8150), .A2(n7786), .ZN(n8163) );
  AOI21_X1 U7665 ( .B1(n8135), .B2(n7206), .A(n7205), .ZN(n7204) );
  INV_X1 U7666 ( .A(n7783), .ZN(n7205) );
  INV_X1 U7667 ( .A(n7781), .ZN(n7206) );
  INV_X1 U7668 ( .A(n8135), .ZN(n7207) );
  NAND2_X1 U7669 ( .A1(n8055), .A2(n8054), .ZN(n8057) );
  OAI21_X1 U7670 ( .B1(n7956), .B2(n6669), .A(n7753), .ZN(n7971) );
  AND2_X1 U7671 ( .A1(n7957), .A2(n7976), .ZN(n8111) );
  XNOR2_X1 U7672 ( .A(n10049), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U7673 ( .A1(n13289), .A2(n7428), .ZN(n13212) );
  AND2_X1 U7674 ( .A1(n8952), .A2(n8926), .ZN(n7428) );
  XNOR2_X1 U7675 ( .A(n6567), .B(n10812), .ZN(n8378) );
  NAND2_X1 U7676 ( .A1(n9928), .A2(n9927), .ZN(n13382) );
  NAND2_X1 U7677 ( .A1(n13418), .A2(n6895), .ZN(n13383) );
  NOR2_X1 U7678 ( .A1(n13586), .A2(n13583), .ZN(n6895) );
  OR2_X1 U7679 ( .A1(n13430), .A2(n12037), .ZN(n7358) );
  NOR2_X1 U7680 ( .A1(n11854), .A2(n6919), .ZN(n6918) );
  INV_X1 U7681 ( .A(n11688), .ZN(n6919) );
  AOI21_X1 U7682 ( .B1(n7312), .B2(n7311), .A(n6658), .ZN(n7310) );
  AOI21_X1 U7683 ( .B1(n7554), .B2(n7560), .A(n6685), .ZN(n7553) );
  INV_X1 U7684 ( .A(n7556), .ZN(n7554) );
  INV_X1 U7685 ( .A(n11674), .ZN(n7559) );
  AND2_X1 U7686 ( .A1(n10377), .A2(n12450), .ZN(n7546) );
  NAND2_X1 U7687 ( .A1(n13785), .A2(n6649), .ZN(n13736) );
  NAND2_X1 U7688 ( .A1(n11574), .A2(n6796), .ZN(n6794) );
  NOR2_X1 U7689 ( .A1(n6799), .A2(n6798), .ZN(n6796) );
  INV_X1 U7690 ( .A(n7551), .ZN(n6799) );
  OR2_X1 U7691 ( .A1(n7553), .A2(n6798), .ZN(n6795) );
  OAI21_X1 U7692 ( .B1(n14100), .B2(n7599), .A(n7596), .ZN(n14057) );
  AOI21_X1 U7693 ( .B1(n7598), .B2(n7597), .A(n6633), .ZN(n7596) );
  INV_X1 U7694 ( .A(n9584), .ZN(n7597) );
  NAND2_X1 U7695 ( .A1(n14198), .A2(n7445), .ZN(n14133) );
  NOR2_X1 U7696 ( .A1(n14299), .A2(n7446), .ZN(n7445) );
  INV_X1 U7697 ( .A(n7447), .ZN(n7446) );
  NAND2_X1 U7698 ( .A1(n14165), .A2(n12321), .ZN(n7604) );
  INV_X1 U7699 ( .A(n7335), .ZN(n7334) );
  OAI21_X1 U7700 ( .B1(n6610), .B2(n7336), .A(n9701), .ZN(n7335) );
  NAND2_X1 U7701 ( .A1(n14238), .A2(n6610), .ZN(n7338) );
  OR2_X1 U7702 ( .A1(n14334), .A2(n14217), .ZN(n12181) );
  NAND2_X1 U7703 ( .A1(n11262), .A2(n7347), .ZN(n11399) );
  AND2_X1 U7704 ( .A1(n12312), .A2(n9690), .ZN(n7347) );
  OR2_X1 U7705 ( .A1(n10343), .A2(n10069), .ZN(n10363) );
  AOI21_X1 U7706 ( .B1(n9676), .B2(n9672), .A(n9671), .ZN(n10353) );
  NOR2_X1 U7707 ( .A1(n6574), .A2(n14032), .ZN(n7176) );
  INV_X1 U7708 ( .A(n9289), .ZN(n6880) );
  NOR2_X1 U7709 ( .A1(n9289), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n9288) );
  XNOR2_X1 U7710 ( .A(n8837), .B(SI_22_), .ZN(n9556) );
  NAND3_X1 U7711 ( .A1(n9506), .A2(n7483), .A3(n7481), .ZN(n9643) );
  INV_X1 U7712 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7483) );
  INV_X1 U7713 ( .A(n8799), .ZN(n8797) );
  NAND2_X1 U7714 ( .A1(n9506), .A2(n7481), .ZN(n9641) );
  NAND2_X1 U7715 ( .A1(n8773), .A2(n7542), .ZN(n8793) );
  NAND2_X1 U7716 ( .A1(n6859), .A2(n8710), .ZN(n8751) );
  NAND2_X1 U7717 ( .A1(n6947), .A2(n6946), .ZN(n7243) );
  NAND2_X1 U7718 ( .A1(n7249), .A2(n7244), .ZN(n6946) );
  INV_X1 U7719 ( .A(n14393), .ZN(n6947) );
  NAND2_X1 U7720 ( .A1(n7246), .A2(n7245), .ZN(n7244) );
  NAND2_X1 U7721 ( .A1(n6687), .A2(n7246), .ZN(n7078) );
  NAND2_X1 U7722 ( .A1(n7252), .A2(n15321), .ZN(n7074) );
  NAND2_X1 U7723 ( .A1(n12076), .A2(n9181), .ZN(n14436) );
  NAND2_X1 U7724 ( .A1(n12757), .A2(n12758), .ZN(n7486) );
  NAND2_X1 U7725 ( .A1(n6655), .A2(n7195), .ZN(n7194) );
  OR2_X1 U7726 ( .A1(n11020), .A2(n11019), .ZN(n7302) );
  NAND2_X1 U7727 ( .A1(n6748), .A2(n6930), .ZN(n6747) );
  INV_X1 U7728 ( .A(n12889), .ZN(n6930) );
  NAND2_X1 U7729 ( .A1(n12890), .A2(n15031), .ZN(n6748) );
  NAND2_X1 U7730 ( .A1(n6861), .A2(n13569), .ZN(n6860) );
  AOI21_X1 U7731 ( .B1(n6864), .B2(n7288), .A(n12018), .ZN(n6863) );
  NAND2_X1 U7732 ( .A1(n9605), .A2(n9604), .ZN(n14270) );
  NAND4_X1 U7733 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n13840)
         );
  XNOR2_X1 U7734 ( .A(n9638), .B(n9710), .ZN(n14263) );
  OR2_X1 U7735 ( .A1(n9067), .A2(n9068), .ZN(n7250) );
  NAND2_X1 U7736 ( .A1(n10807), .A2(n9743), .ZN(n6970) );
  NAND2_X1 U7737 ( .A1(n9906), .A2(n9734), .ZN(n6971) );
  NAND2_X1 U7738 ( .A1(n7470), .A2(n12121), .ZN(n7469) );
  OR2_X1 U7739 ( .A1(n7470), .A2(n12121), .ZN(n7468) );
  INV_X1 U7740 ( .A(n9778), .ZN(n6988) );
  NAND2_X1 U7741 ( .A1(n7668), .A2(n9778), .ZN(n7667) );
  NAND2_X1 U7742 ( .A1(n7670), .A2(n7669), .ZN(n7668) );
  INV_X1 U7743 ( .A(n9777), .ZN(n6983) );
  AND2_X1 U7744 ( .A1(n9771), .A2(n9772), .ZN(n7670) );
  NAND2_X1 U7745 ( .A1(n12181), .A2(n12171), .ZN(n12177) );
  INV_X1 U7746 ( .A(n9790), .ZN(n6834) );
  NAND2_X1 U7747 ( .A1(n7692), .A2(n7691), .ZN(n7690) );
  INV_X1 U7748 ( .A(n9795), .ZN(n7691) );
  OR2_X1 U7749 ( .A1(n9801), .A2(n6577), .ZN(n7689) );
  NAND2_X1 U7750 ( .A1(n9801), .A2(n6577), .ZN(n7692) );
  AOI21_X1 U7751 ( .B1(n7104), .B2(n7103), .A(n6683), .ZN(n7102) );
  NAND2_X1 U7752 ( .A1(n7451), .A2(n7100), .ZN(n7101) );
  INV_X1 U7753 ( .A(n9818), .ZN(n7675) );
  NAND2_X1 U7754 ( .A1(n9824), .A2(n9825), .ZN(n6830) );
  NAND2_X1 U7755 ( .A1(n7098), .A2(n7459), .ZN(n12223) );
  NAND2_X1 U7756 ( .A1(n7460), .A2(n7457), .ZN(n7098) );
  INV_X1 U7757 ( .A(n7461), .ZN(n7457) );
  NOR2_X1 U7758 ( .A1(n7461), .A2(n7459), .ZN(n7458) );
  NAND2_X1 U7759 ( .A1(n12226), .A2(n7474), .ZN(n7473) );
  INV_X1 U7760 ( .A(n12225), .ZN(n7474) );
  AND2_X1 U7761 ( .A1(n9854), .A2(n9855), .ZN(n7687) );
  NAND2_X1 U7762 ( .A1(n7683), .A2(n9860), .ZN(n7682) );
  NAND2_X1 U7763 ( .A1(n7687), .A2(n7684), .ZN(n7683) );
  AOI22_X1 U7764 ( .A1(n7680), .A2(n7682), .B1(n7678), .B2(n7687), .ZN(n7677)
         );
  NOR2_X1 U7765 ( .A1(n9860), .A2(n7679), .ZN(n7678) );
  INV_X1 U7766 ( .A(n7684), .ZN(n7679) );
  OAI22_X1 U7767 ( .A1(n12237), .A2(n7117), .B1(n7116), .B2(n12238), .ZN(
        n12242) );
  INV_X1 U7768 ( .A(n12236), .ZN(n7116) );
  NOR2_X1 U7769 ( .A1(n12239), .A2(n12236), .ZN(n7117) );
  NAND2_X1 U7770 ( .A1(n7464), .A2(n7465), .ZN(n12237) );
  INV_X1 U7771 ( .A(n12249), .ZN(n7480) );
  AOI21_X1 U7772 ( .B1(n7145), .B2(n7148), .A(n12934), .ZN(n7144) );
  OAI21_X1 U7773 ( .B1(n7700), .B2(n7529), .A(n8699), .ZN(n7528) );
  NOR2_X1 U7774 ( .A1(n7136), .A2(n7135), .ZN(n12729) );
  NOR2_X1 U7775 ( .A1(n7501), .A2(n12752), .ZN(n7499) );
  INV_X1 U7776 ( .A(n12687), .ZN(n7017) );
  INV_X1 U7777 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7398) );
  INV_X1 U7778 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8325) );
  AOI21_X1 U7779 ( .B1(n7178), .B2(n7181), .A(n7528), .ZN(n7177) );
  AND2_X1 U7780 ( .A1(n7184), .A2(n7699), .ZN(n7183) );
  NAND2_X1 U7781 ( .A1(n8612), .A2(n6866), .ZN(n7184) );
  OAI21_X1 U7782 ( .B1(n10006), .B2(P2_DATAO_REG_11__SCAN_IN), .A(n6968), .ZN(
        n8589) );
  NAND2_X1 U7783 ( .A1(n10006), .A2(n10138), .ZN(n6968) );
  NOR2_X1 U7784 ( .A1(n8585), .A2(n8563), .ZN(n7517) );
  INV_X1 U7785 ( .A(n8567), .ZN(n7519) );
  INV_X1 U7786 ( .A(n8501), .ZN(n7523) );
  INV_X1 U7787 ( .A(n8416), .ZN(n7084) );
  INV_X1 U7788 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9028) );
  AND2_X1 U7789 ( .A1(n7233), .A2(n7232), .ZN(n12615) );
  NAND2_X1 U7790 ( .A1(n13147), .A2(n12588), .ZN(n7232) );
  NAND2_X1 U7791 ( .A1(n12896), .A2(n12892), .ZN(n7233) );
  NAND2_X1 U7792 ( .A1(n14959), .A2(n11027), .ZN(n11028) );
  OAI21_X1 U7793 ( .B1(n11908), .B2(n14496), .A(n11907), .ZN(n12789) );
  NAND2_X1 U7794 ( .A1(n12823), .A2(n12822), .ZN(n6754) );
  NAND2_X1 U7795 ( .A1(n12624), .A2(n12623), .ZN(n7013) );
  OR2_X1 U7796 ( .A1(n13113), .A2(n13003), .ZN(n12722) );
  NAND2_X1 U7797 ( .A1(n8269), .A2(n7493), .ZN(n7490) );
  AND2_X1 U7798 ( .A1(n8264), .A2(n12674), .ZN(n7510) );
  INV_X1 U7799 ( .A(n12679), .ZN(n7506) );
  INV_X1 U7800 ( .A(n12674), .ZN(n7507) );
  NAND2_X1 U7801 ( .A1(n9137), .A2(n12634), .ZN(n15042) );
  INV_X1 U7802 ( .A(n10577), .ZN(n9250) );
  INV_X1 U7803 ( .A(n12913), .ZN(n8228) );
  INV_X1 U7804 ( .A(SI_12_), .ZN(n8614) );
  AND2_X1 U7805 ( .A1(n7716), .A2(n6618), .ZN(n6932) );
  INV_X1 U7806 ( .A(n8162), .ZN(n7199) );
  NAND2_X1 U7807 ( .A1(n7646), .A2(n8282), .ZN(n7645) );
  INV_X1 U7808 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8282) );
  INV_X1 U7809 ( .A(n7647), .ZN(n7646) );
  INV_X1 U7810 ( .A(n7212), .ZN(n7211) );
  OAI21_X1 U7811 ( .B1(n8054), .B2(n7213), .A(n7774), .ZN(n7212) );
  INV_X1 U7812 ( .A(n7772), .ZN(n7213) );
  INV_X1 U7813 ( .A(n7750), .ZN(n7226) );
  INV_X1 U7814 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7896) );
  INV_X1 U7815 ( .A(n8562), .ZN(n7427) );
  OR2_X1 U7816 ( .A1(n9944), .A2(n9910), .ZN(n9951) );
  INV_X1 U7817 ( .A(n13696), .ZN(n8373) );
  NAND2_X1 U7818 ( .A1(n9009), .A2(n13414), .ZN(n7287) );
  NOR2_X1 U7819 ( .A1(n7286), .A2(n7285), .ZN(n7284) );
  INV_X1 U7820 ( .A(n7287), .ZN(n7286) );
  AND2_X1 U7821 ( .A1(n8939), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8954) );
  XNOR2_X1 U7822 ( .A(n13603), .B(n13456), .ZN(n7299) );
  NAND2_X1 U7823 ( .A1(n13620), .A2(n7365), .ZN(n7364) );
  NOR2_X1 U7824 ( .A1(n13478), .A2(n7366), .ZN(n7365) );
  INV_X1 U7825 ( .A(n12032), .ZN(n7366) );
  INV_X1 U7826 ( .A(n12008), .ZN(n7262) );
  NAND2_X1 U7827 ( .A1(n13500), .A2(n7266), .ZN(n7265) );
  INV_X1 U7828 ( .A(n12005), .ZN(n7266) );
  INV_X1 U7829 ( .A(n13640), .ZN(n7134) );
  AND2_X1 U7830 ( .A1(n11144), .A2(n6917), .ZN(n6916) );
  INV_X1 U7831 ( .A(n11135), .ZN(n6917) );
  INV_X1 U7832 ( .A(n9733), .ZN(n9732) );
  NAND3_X1 U7833 ( .A1(n6943), .A2(n8347), .A3(n8346), .ZN(n8970) );
  INV_X1 U7834 ( .A(n8345), .ZN(n6943) );
  INV_X1 U7835 ( .A(n12447), .ZN(n7570) );
  OR2_X1 U7836 ( .A1(n11823), .A2(n7564), .ZN(n7563) );
  INV_X1 U7837 ( .A(n12450), .ZN(n6937) );
  NAND2_X1 U7838 ( .A1(n12257), .A2(n7113), .ZN(n7112) );
  NAND2_X1 U7839 ( .A1(n12255), .A2(n7110), .ZN(n7109) );
  AND2_X1 U7840 ( .A1(n9705), .A2(n9565), .ZN(n12324) );
  NAND2_X1 U7841 ( .A1(n14135), .A2(n9555), .ZN(n14115) );
  INV_X1 U7842 ( .A(n14228), .ZN(n7341) );
  AND2_X1 U7843 ( .A1(n7585), .A2(n11600), .ZN(n7584) );
  NOR2_X1 U7844 ( .A1(n7443), .A2(n14401), .ZN(n7442) );
  INV_X1 U7845 ( .A(n7444), .ZN(n7443) );
  NAND2_X1 U7846 ( .A1(n7594), .A2(n6637), .ZN(n11980) );
  OR2_X1 U7847 ( .A1(n14619), .A2(n6885), .ZN(n7594) );
  INV_X1 U7848 ( .A(n12300), .ZN(n6885) );
  NAND2_X1 U7849 ( .A1(n9306), .A2(n9307), .ZN(n10410) );
  NAND2_X1 U7850 ( .A1(n9318), .A2(n10708), .ZN(n12107) );
  INV_X1 U7851 ( .A(n6783), .ZN(n7581) );
  INV_X1 U7852 ( .A(n6785), .ZN(n7582) );
  NAND2_X1 U7853 ( .A1(n10741), .A2(n14632), .ZN(n12093) );
  NAND2_X1 U7854 ( .A1(n7188), .A2(n7189), .ZN(n7322) );
  AND2_X1 U7855 ( .A1(n7187), .A2(n7190), .ZN(n7186) );
  AOI21_X1 U7856 ( .B1(n7327), .B2(n6570), .A(n12328), .ZN(n7190) );
  NAND2_X1 U7857 ( .A1(n12062), .A2(n6570), .ZN(n7187) );
  NAND2_X1 U7858 ( .A1(n6887), .A2(n6886), .ZN(n14135) );
  AND2_X1 U7859 ( .A1(n7600), .A2(n9554), .ZN(n6886) );
  NAND2_X1 U7860 ( .A1(n7535), .A2(n7537), .ZN(n9885) );
  INV_X1 U7861 ( .A(n7538), .ZN(n7537) );
  OAI21_X1 U7862 ( .B1(n8934), .B2(n7539), .A(n9626), .ZN(n7538) );
  OAI21_X1 U7863 ( .B1(n7096), .B2(n6730), .A(n8913), .ZN(n8928) );
  NAND2_X1 U7864 ( .A1(n8894), .A2(n8895), .ZN(n7096) );
  AND2_X1 U7865 ( .A1(n6587), .A2(n7482), .ZN(n7481) );
  INV_X1 U7866 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7482) );
  OAI21_X1 U7867 ( .B1(n8613), .B2(n7119), .A(n7118), .ZN(n8700) );
  INV_X1 U7868 ( .A(n7120), .ZN(n7119) );
  AOI21_X1 U7869 ( .B1(n7120), .B2(n7094), .A(n7529), .ZN(n7118) );
  AOI21_X1 U7870 ( .B1(n7178), .B2(n7181), .A(n7121), .ZN(n7120) );
  OR2_X1 U7871 ( .A1(n9434), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9435) );
  NAND2_X1 U7872 ( .A1(n8589), .A2(n15455), .ZN(n6866) );
  NAND2_X1 U7873 ( .A1(n8454), .A2(n8453), .ZN(n8476) );
  XNOR2_X1 U7874 ( .A(n8432), .B(n6966), .ZN(n8430) );
  NAND2_X1 U7875 ( .A1(n6967), .A2(n6640), .ZN(n8413) );
  NAND2_X1 U7876 ( .A1(n7171), .A2(n7813), .ZN(n7169) );
  AND2_X1 U7877 ( .A1(n13863), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U7878 ( .A1(n15382), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n7257) );
  XNOR2_X1 U7879 ( .A(n7072), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n9038) );
  OAI22_X1 U7880 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n15353), .B1(n9088), .B2(
        n9087), .ZN(n9092) );
  NAND2_X1 U7881 ( .A1(n7621), .A2(n9150), .ZN(n7620) );
  INV_X1 U7882 ( .A(n10562), .ZN(n7621) );
  AOI21_X1 U7883 ( .B1(n7616), .B2(n9217), .A(n6672), .ZN(n7613) );
  OR2_X1 U7884 ( .A1(n12568), .A2(n9217), .ZN(n7614) );
  INV_X1 U7885 ( .A(n15063), .ZN(n12355) );
  NAND2_X1 U7886 ( .A1(n9182), .A2(n13066), .ZN(n9183) );
  NAND2_X1 U7887 ( .A1(n7948), .A2(n15369), .ZN(n7963) );
  AOI21_X1 U7888 ( .B1(n7633), .B2(n7631), .A(n7630), .ZN(n7629) );
  INV_X1 U7889 ( .A(n7633), .ZN(n7632) );
  INV_X1 U7890 ( .A(n9196), .ZN(n7630) );
  NOR2_X1 U7891 ( .A1(n12522), .A2(n7637), .ZN(n7636) );
  INV_X1 U7892 ( .A(n9183), .ZN(n7637) );
  NOR2_X1 U7893 ( .A1(n10993), .A2(n7624), .ZN(n7623) );
  NAND3_X1 U7894 ( .A1(n11629), .A2(n9168), .A3(n6772), .ZN(n7628) );
  NAND2_X1 U7895 ( .A1(n7155), .A2(n15071), .ZN(n7154) );
  AND4_X1 U7896 ( .A1(n12582), .A2(n8237), .A3(n8236), .A4(n8235), .ZN(n12765)
         );
  INV_X1 U7897 ( .A(n7856), .ZN(n7887) );
  OAI21_X1 U7898 ( .B1(n6940), .B2(n6751), .A(n10664), .ZN(n10553) );
  NOR2_X1 U7899 ( .A1(n6922), .A2(n10552), .ZN(n6751) );
  NOR2_X1 U7900 ( .A1(n14906), .A2(n11037), .ZN(n14905) );
  NAND2_X1 U7901 ( .A1(n14944), .A2(n11026), .ZN(n14961) );
  INV_X1 U7902 ( .A(n7304), .ZN(n11009) );
  NAND2_X1 U7903 ( .A1(n11056), .A2(n14937), .ZN(n14968) );
  XNOR2_X1 U7904 ( .A(n11028), .B(n11065), .ZN(n14992) );
  NAND2_X1 U7905 ( .A1(n14992), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n14991) );
  OR2_X1 U7906 ( .A1(n14976), .A2(n11014), .ZN(n6774) );
  INV_X1 U7907 ( .A(n7315), .ZN(n11013) );
  NAND2_X1 U7908 ( .A1(n15019), .A2(n11032), .ZN(n11033) );
  NAND2_X1 U7909 ( .A1(n11033), .A2(n11034), .ZN(n11463) );
  NAND2_X1 U7910 ( .A1(n6928), .A2(n11087), .ZN(n11459) );
  NAND2_X1 U7911 ( .A1(n12784), .A2(n7271), .ZN(n6939) );
  NAND2_X1 U7912 ( .A1(n12847), .A2(n12848), .ZN(n14450) );
  NAND2_X1 U7913 ( .A1(n14450), .A2(n14451), .ZN(n14449) );
  NOR2_X1 U7914 ( .A1(n12934), .A2(n7034), .ZN(n7033) );
  NAND2_X1 U7915 ( .A1(n12955), .A2(n7379), .ZN(n7378) );
  OR2_X1 U7916 ( .A1(n8211), .A2(n8210), .ZN(n7377) );
  NAND2_X1 U7917 ( .A1(n7060), .A2(n7058), .ZN(n7390) );
  AOI21_X1 U7918 ( .B1(n7061), .B2(n6572), .A(n7059), .ZN(n7058) );
  NOR2_X1 U7919 ( .A1(n12590), .A2(n7386), .ZN(n7385) );
  INV_X1 U7920 ( .A(n8134), .ZN(n7386) );
  AND2_X1 U7921 ( .A1(n12591), .A2(n12623), .ZN(n12993) );
  OR2_X1 U7922 ( .A1(n7063), .A2(n12590), .ZN(n13005) );
  OR2_X1 U7923 ( .A1(n13184), .A2(n13049), .ZN(n13013) );
  OR2_X1 U7924 ( .A1(n13056), .A2(n13065), .ZN(n13039) );
  NAND2_X1 U7925 ( .A1(n7051), .A2(n7054), .ZN(n7050) );
  NAND2_X1 U7926 ( .A1(n7041), .A2(n7046), .ZN(n13047) );
  OR2_X1 U7927 ( .A1(n8074), .A2(n7049), .ZN(n7041) );
  NOR2_X1 U7928 ( .A1(n8087), .A2(n7053), .ZN(n7052) );
  INV_X1 U7929 ( .A(n8073), .ZN(n7053) );
  NAND2_X1 U7930 ( .A1(n8268), .A2(n7492), .ZN(n13052) );
  INV_X1 U7931 ( .A(n13035), .ZN(n13065) );
  NAND2_X1 U7932 ( .A1(n6744), .A2(n12701), .ZN(n13067) );
  NAND2_X1 U7933 ( .A1(n11930), .A2(n12606), .ZN(n6744) );
  AND2_X1 U7934 ( .A1(n12702), .A2(n12701), .ZN(n12606) );
  AOI21_X1 U7935 ( .B1(n6580), .B2(n7018), .A(n11777), .ZN(n7015) );
  INV_X1 U7936 ( .A(n7513), .ZN(n7018) );
  OR2_X1 U7937 ( .A1(n11799), .A2(n8266), .ZN(n7515) );
  NAND2_X1 U7938 ( .A1(n7515), .A2(n7513), .ZN(n11778) );
  NAND2_X1 U7939 ( .A1(n8265), .A2(n12687), .ZN(n11799) );
  OR2_X1 U7940 ( .A1(n7368), .A2(n7040), .ZN(n7039) );
  INV_X1 U7941 ( .A(n7992), .ZN(n7040) );
  OAI21_X1 U7942 ( .B1(n11279), .B2(n8262), .A(n8263), .ZN(n11346) );
  AOI21_X1 U7943 ( .B1(n11348), .B2(n7372), .A(n6622), .ZN(n7371) );
  INV_X1 U7944 ( .A(n7962), .ZN(n7372) );
  NAND2_X1 U7945 ( .A1(n7370), .A2(n7368), .ZN(n11446) );
  NAND2_X1 U7946 ( .A1(n11282), .A2(n7962), .ZN(n11349) );
  INV_X1 U7947 ( .A(n12659), .ZN(n12596) );
  OAI211_X1 U7948 ( .C1(n12585), .C2(SI_2_), .A(n7852), .B(n7851), .ZN(n15043)
         );
  INV_X1 U7949 ( .A(n15062), .ZN(n6989) );
  INV_X1 U7950 ( .A(n9133), .ZN(n15059) );
  NAND2_X1 U7951 ( .A1(n12959), .A2(n12958), .ZN(n12957) );
  INV_X1 U7952 ( .A(n7033), .ZN(n7032) );
  OR2_X1 U7953 ( .A1(n10851), .A2(n8191), .ZN(n8152) );
  NAND2_X1 U7954 ( .A1(n8044), .A2(n8043), .ZN(n13137) );
  OR2_X1 U7955 ( .A1(n10251), .A2(n8191), .ZN(n8044) );
  NAND2_X1 U7956 ( .A1(n10554), .A2(n7489), .ZN(n8251) );
  OAI21_X1 U7957 ( .B1(n8176), .B2(n11740), .A(n7790), .ZN(n8188) );
  NAND2_X1 U7958 ( .A1(n7203), .A2(n7201), .ZN(n8150) );
  AOI21_X1 U7959 ( .B1(n7204), .B2(n7207), .A(n7202), .ZN(n7201) );
  INV_X1 U7960 ( .A(n8147), .ZN(n7202) );
  NAND2_X1 U7961 ( .A1(n8107), .A2(n7779), .ZN(n8125) );
  NAND2_X1 U7962 ( .A1(n8125), .A2(n8124), .ZN(n8127) );
  NAND2_X1 U7963 ( .A1(n8091), .A2(n7777), .ZN(n8105) );
  NAND2_X1 U7964 ( .A1(n8105), .A2(n8104), .ZN(n8107) );
  NAND2_X1 U7965 ( .A1(n8089), .A2(n8088), .ZN(n8091) );
  NAND2_X1 U7966 ( .A1(n8037), .A2(n7770), .ZN(n8055) );
  NAND2_X1 U7967 ( .A1(n7761), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7191) );
  INV_X1 U7968 ( .A(n7761), .ZN(n7762) );
  NOR2_X1 U7969 ( .A1(n7756), .A2(n7238), .ZN(n7237) );
  AND2_X1 U7970 ( .A1(n10136), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7756) );
  INV_X1 U7971 ( .A(n7754), .ZN(n7238) );
  OAI21_X1 U7972 ( .B1(n7942), .B2(n7751), .A(n7752), .ZN(n7956) );
  NOR2_X1 U7973 ( .A1(n7749), .A2(n7229), .ZN(n7228) );
  INV_X1 U7974 ( .A(n7746), .ZN(n7229) );
  NAND2_X1 U7975 ( .A1(n7223), .A2(n7875), .ZN(n7220) );
  XNOR2_X1 U7976 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7893) );
  NOR2_X1 U7977 ( .A1(n7877), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7897) );
  OR2_X1 U7978 ( .A1(n7850), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n7877) );
  OR3_X1 U7979 ( .A1(n11924), .A2(n11973), .A3(n11742), .ZN(n9997) );
  NAND2_X1 U7980 ( .A1(n6592), .A2(n8654), .ZN(n7430) );
  NAND2_X1 U7981 ( .A1(n7409), .A2(n7407), .ZN(n7406) );
  INV_X1 U7982 ( .A(n11965), .ZN(n7409) );
  NOR2_X1 U7983 ( .A1(n7411), .A2(n7408), .ZN(n7407) );
  NOR2_X1 U7984 ( .A1(n7405), .A2(n7414), .ZN(n7399) );
  OR2_X1 U7985 ( .A1(n11965), .A2(n7408), .ZN(n7405) );
  OR2_X1 U7986 ( .A1(n7406), .A2(n8744), .ZN(n7401) );
  AND2_X1 U7987 ( .A1(n13586), .A2(n11948), .ZN(n7397) );
  AOI21_X1 U7988 ( .B1(n10910), .B2(n10909), .A(n8517), .ZN(n10880) );
  NAND2_X1 U7989 ( .A1(n10880), .A2(n10879), .ZN(n10878) );
  NAND2_X1 U7990 ( .A1(n11362), .A2(n8611), .ZN(n11412) );
  NAND2_X1 U7991 ( .A1(n8870), .A2(n8869), .ZN(n8871) );
  NAND2_X1 U7992 ( .A1(n13219), .A2(n13218), .ZN(n13217) );
  OR2_X1 U7993 ( .A1(n10658), .A2(n10657), .ZN(n6890) );
  NAND3_X1 U7994 ( .A1(n6890), .A2(n6616), .A3(n10505), .ZN(n10504) );
  NAND2_X1 U7995 ( .A1(n13226), .A2(n13225), .ZN(n8792) );
  NAND2_X1 U7996 ( .A1(n7423), .A2(n7421), .ZN(n11362) );
  AND2_X1 U7997 ( .A1(n7424), .A2(n7422), .ZN(n7421) );
  INV_X1 U7998 ( .A(n11364), .ZN(n7422) );
  NAND2_X1 U7999 ( .A1(n9952), .A2(n6847), .ZN(n6846) );
  NAND2_X1 U8000 ( .A1(n8373), .A2(n8383), .ZN(n8422) );
  INV_X1 U8001 ( .A(n8422), .ZN(n8386) );
  NOR2_X1 U8002 ( .A1(n13382), .A2(n13583), .ZN(n7128) );
  NOR2_X1 U8003 ( .A1(n12014), .A2(n6865), .ZN(n6864) );
  NAND2_X1 U8004 ( .A1(n13418), .A2(n9009), .ZN(n13396) );
  OR2_X1 U8005 ( .A1(n13598), .A2(n13448), .ZN(n7359) );
  NAND2_X1 U8006 ( .A1(n7123), .A2(n7122), .ZN(n13432) );
  NAND2_X1 U8007 ( .A1(n7290), .A2(n7091), .ZN(n13413) );
  AOI21_X1 U8008 ( .B1(n7291), .B2(n7292), .A(n7289), .ZN(n7091) );
  INV_X1 U8009 ( .A(n12011), .ZN(n7289) );
  INV_X1 U8010 ( .A(n12013), .ZN(n13423) );
  NAND2_X1 U8011 ( .A1(n12036), .A2(n12035), .ZN(n13430) );
  NAND2_X1 U8012 ( .A1(n7364), .A2(n7363), .ZN(n13458) );
  AND2_X1 U8013 ( .A1(n13459), .A2(n6620), .ZN(n7363) );
  NAND2_X1 U8014 ( .A1(n12020), .A2(n6901), .ZN(n6900) );
  NOR2_X1 U8015 ( .A1(n7352), .A2(n6902), .ZN(n6901) );
  NAND2_X1 U8016 ( .A1(n12025), .A2(n12019), .ZN(n6902) );
  NAND2_X1 U8017 ( .A1(n7351), .A2(n12025), .ZN(n6899) );
  NAND2_X1 U8018 ( .A1(n12022), .A2(n6578), .ZN(n13554) );
  NAND2_X1 U8019 ( .A1(n7360), .A2(n6642), .ZN(n11882) );
  NAND2_X1 U8020 ( .A1(n6912), .A2(n11687), .ZN(n11726) );
  NAND2_X1 U8021 ( .A1(n11686), .A2(n11685), .ZN(n6912) );
  XNOR2_X1 U8022 ( .A(n13661), .B(n11758), .ZN(n11725) );
  NOR2_X1 U8023 ( .A1(n7308), .A2(n11689), .ZN(n7307) );
  AND2_X1 U8024 ( .A1(n11253), .A2(n11251), .ZN(n7312) );
  NAND2_X1 U8025 ( .A1(n6921), .A2(n11137), .ZN(n11248) );
  NAND2_X1 U8026 ( .A1(n10969), .A2(n10975), .ZN(n11136) );
  OAI21_X1 U8027 ( .B1(n10915), .B2(n10615), .A(n10616), .ZN(n10618) );
  NAND2_X1 U8028 ( .A1(n6914), .A2(n6913), .ZN(n10829) );
  INV_X1 U8029 ( .A(n10832), .ZN(n6913) );
  INV_X1 U8030 ( .A(n10618), .ZN(n6914) );
  NAND2_X1 U8031 ( .A1(n10812), .A2(n10723), .ZN(n10808) );
  NAND2_X1 U8032 ( .A1(n8620), .A2(n8619), .ZN(n13667) );
  AND2_X1 U8033 ( .A1(n8984), .A2(n8983), .ZN(n14810) );
  OR2_X1 U8034 ( .A1(n8971), .A2(n8970), .ZN(n8973) );
  AND2_X1 U8035 ( .A1(n13819), .A2(n7569), .ZN(n7568) );
  OR2_X1 U8036 ( .A1(n13747), .A2(n7570), .ZN(n7569) );
  INV_X1 U8037 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n15429) );
  NOR2_X1 U8038 ( .A1(n9416), .A2(n15303), .ZN(n9424) );
  AND2_X1 U8039 ( .A1(n11208), .A2(n11207), .ZN(n11209) );
  NAND2_X1 U8040 ( .A1(n13755), .A2(n13756), .ZN(n13754) );
  INV_X1 U8041 ( .A(n6801), .ZN(n6800) );
  OAI21_X1 U8042 ( .B1(n13756), .B2(n12388), .A(n13769), .ZN(n6801) );
  INV_X1 U8043 ( .A(n11580), .ZN(n7557) );
  AOI21_X1 U8044 ( .B1(n10342), .B2(n12463), .A(n7576), .ZN(n10377) );
  INV_X1 U8045 ( .A(n10346), .ZN(n10347) );
  INV_X1 U8046 ( .A(n13808), .ZN(n7572) );
  NOR2_X1 U8047 ( .A1(n13726), .A2(n7575), .ZN(n7574) );
  INV_X1 U8048 ( .A(n12400), .ZN(n7575) );
  NAND2_X1 U8049 ( .A1(n13736), .A2(n12417), .ZN(n13796) );
  INV_X1 U8050 ( .A(n7548), .ZN(n7547) );
  NAND2_X1 U8051 ( .A1(n13766), .A2(n13768), .ZN(n13807) );
  NAND2_X1 U8052 ( .A1(n13807), .A2(n13808), .ZN(n13806) );
  AND4_X1 U8053 ( .A1(n9459), .A2(n9458), .A3(n9457), .A4(n9456), .ZN(n12166)
         );
  INV_X1 U8054 ( .A(n13875), .ZN(n13878) );
  AND2_X1 U8055 ( .A1(n12062), .A2(n9610), .ZN(n7590) );
  AOI21_X1 U8056 ( .B1(n7346), .B2(n7344), .A(n6593), .ZN(n7343) );
  INV_X1 U8057 ( .A(n7346), .ZN(n7345) );
  AND2_X1 U8058 ( .A1(n14372), .A2(n9305), .ZN(n14128) );
  NOR2_X1 U8059 ( .A1(n14161), .A2(n7603), .ZN(n7602) );
  INV_X1 U8060 ( .A(n9538), .ZN(n7603) );
  OR2_X1 U8061 ( .A1(n14172), .A2(n12321), .ZN(n14173) );
  NAND2_X1 U8062 ( .A1(n9527), .A2(n12209), .ZN(n14165) );
  NOR2_X1 U8063 ( .A1(n14203), .A2(n7340), .ZN(n7337) );
  INV_X1 U8064 ( .A(n9477), .ZN(n7607) );
  INV_X1 U8065 ( .A(n14236), .ZN(n9700) );
  NAND2_X1 U8066 ( .A1(n9476), .A2(n9475), .ZN(n14514) );
  INV_X1 U8067 ( .A(n14516), .ZN(n9476) );
  AOI21_X1 U8068 ( .B1(n7589), .B2(n14530), .A(n7587), .ZN(n7586) );
  NOR2_X1 U8069 ( .A1(n9422), .A2(n13850), .ZN(n7587) );
  NOR2_X1 U8070 ( .A1(n14530), .A2(n12158), .ZN(n7588) );
  NAND2_X1 U8071 ( .A1(n11267), .A2(n9404), .ZN(n11398) );
  NAND2_X1 U8072 ( .A1(n11398), .A2(n11397), .ZN(n11396) );
  NAND2_X1 U8073 ( .A1(n7330), .A2(n7329), .ZN(n11264) );
  NAND2_X1 U8074 ( .A1(n7332), .A2(n9689), .ZN(n7329) );
  OR2_X1 U8075 ( .A1(n12287), .A2(n13878), .ZN(n14221) );
  NAND2_X1 U8076 ( .A1(n9679), .A2(n12093), .ZN(n12086) );
  NAND2_X1 U8077 ( .A1(n12106), .A2(n12107), .ZN(n10411) );
  NOR2_X1 U8078 ( .A1(n10054), .A2(n9545), .ZN(n6961) );
  INV_X1 U8079 ( .A(n14221), .ZN(n14207) );
  INV_X1 U8080 ( .A(n14029), .ZN(n14257) );
  NAND2_X1 U8081 ( .A1(n9493), .A2(n9492), .ZN(n14330) );
  XNOR2_X1 U8082 ( .A(n9925), .B(n9924), .ZN(n12260) );
  NAND2_X1 U8083 ( .A1(n9280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6881) );
  NOR2_X1 U8084 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6995) );
  NOR2_X1 U8085 ( .A1(n9645), .A2(n9276), .ZN(n9277) );
  XNOR2_X1 U8086 ( .A(n7096), .B(n6730), .ZN(n11895) );
  NAND2_X1 U8087 ( .A1(n9649), .A2(n9647), .ZN(n9653) );
  INV_X1 U8088 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U8089 ( .A1(n7531), .A2(n6718), .ZN(n8873) );
  INV_X1 U8090 ( .A(n8857), .ZN(n7530) );
  NAND2_X1 U8091 ( .A1(n7173), .A2(n7172), .ZN(n8814) );
  NOR2_X1 U8092 ( .A1(n6716), .A2(n10576), .ZN(n7172) );
  NAND2_X1 U8093 ( .A1(n6852), .A2(n8773), .ZN(n7173) );
  OAI21_X1 U8094 ( .B1(n6852), .B2(n6716), .A(n6850), .ZN(n7544) );
  NOR2_X1 U8095 ( .A1(n6851), .A2(SI_20_), .ZN(n6850) );
  NOR2_X1 U8096 ( .A1(n8773), .A2(n6716), .ZN(n6851) );
  NAND2_X1 U8097 ( .A1(n8753), .A2(n7543), .ZN(n7542) );
  NAND2_X1 U8098 ( .A1(n8753), .A2(n8773), .ZN(n8755) );
  OR2_X1 U8099 ( .A1(n8752), .A2(n10407), .ZN(n8773) );
  NAND2_X1 U8100 ( .A1(n7593), .A2(n9266), .ZN(n7592) );
  NAND2_X1 U8101 ( .A1(n6963), .A2(n9268), .ZN(n7591) );
  NAND2_X1 U8102 ( .A1(n7520), .A2(n8567), .ZN(n8587) );
  NAND2_X1 U8103 ( .A1(n8565), .A2(n8564), .ZN(n7520) );
  NAND2_X1 U8104 ( .A1(n9304), .A2(n8392), .ZN(n8397) );
  XNOR2_X1 U8105 ( .A(n8396), .B(SI_1_), .ZN(n8398) );
  INV_X2 U8106 ( .A(n6566), .ZN(n10025) );
  XNOR2_X1 U8107 ( .A(n9029), .B(n14916), .ZN(n9050) );
  NAND2_X1 U8108 ( .A1(n15466), .A2(n15467), .ZN(n7080) );
  AOI21_X1 U8109 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15016), .A(n9071), .ZN(
        n9072) );
  NAND2_X1 U8110 ( .A1(n9080), .A2(n9079), .ZN(n9084) );
  AND2_X1 U8111 ( .A1(n7076), .A2(n7075), .ZN(n9109) );
  OR2_X1 U8112 ( .A1(n12364), .A2(n8191), .ZN(n7817) );
  NAND2_X1 U8113 ( .A1(n6770), .A2(n7616), .ZN(n6769) );
  NOR2_X1 U8114 ( .A1(n9217), .A2(n6767), .ZN(n6766) );
  INV_X1 U8115 ( .A(n9215), .ZN(n6767) );
  NAND2_X1 U8116 ( .A1(n6759), .A2(n6756), .ZN(n6755) );
  NAND2_X1 U8117 ( .A1(n12351), .A2(n12354), .ZN(n6759) );
  NAND2_X1 U8118 ( .A1(n8140), .A2(n8139), .ZN(n13006) );
  OR2_X1 U8119 ( .A1(n10825), .A2(n8191), .ZN(n8140) );
  OR2_X1 U8120 ( .A1(n11423), .A2(n8191), .ZN(n8193) );
  INV_X1 U8121 ( .A(n12520), .ZN(n6976) );
  NAND2_X1 U8122 ( .A1(n8065), .A2(n8064), .ZN(n14442) );
  OR2_X1 U8123 ( .A1(n10295), .A2(n8191), .ZN(n8065) );
  OAI22_X1 U8124 ( .A1(n12845), .A2(n7489), .B1(n12585), .B2(n10294), .ZN(
        n8063) );
  NAND2_X1 U8125 ( .A1(n7003), .A2(n7002), .ZN(n14438) );
  INV_X1 U8126 ( .A(n12773), .ZN(n11631) );
  AND2_X1 U8127 ( .A1(n9221), .A2(n9242), .ZN(n14439) );
  NAND2_X1 U8128 ( .A1(n9222), .A2(n10489), .ZN(n12574) );
  CLKBUF_X1 U8129 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n6922) );
  XNOR2_X1 U8130 ( .A(n11022), .B(n10669), .ZN(n10667) );
  NAND2_X1 U8131 ( .A1(n10666), .A2(n10667), .ZN(n11006) );
  NOR2_X1 U8132 ( .A1(n14977), .A2(n11117), .ZN(n14976) );
  NOR2_X1 U8133 ( .A1(n15017), .A2(n11017), .ZN(n11020) );
  XNOR2_X1 U8134 ( .A(n7300), .B(n15454), .ZN(n11457) );
  OAI211_X1 U8135 ( .C1(n6993), .C2(P3_REG2_REG_17__SCAN_IN), .A(n6760), .B(
        n6763), .ZN(n6762) );
  INV_X1 U8136 ( .A(n12844), .ZN(n6763) );
  NAND2_X1 U8137 ( .A1(n6761), .A2(n14475), .ZN(n6760) );
  NAND2_X1 U8138 ( .A1(n7500), .A2(n7498), .ZN(n12613) );
  INV_X1 U8139 ( .A(n7501), .ZN(n7498) );
  NAND2_X1 U8140 ( .A1(n12933), .A2(n7504), .ZN(n7500) );
  NAND2_X1 U8141 ( .A1(n8234), .A2(n8233), .ZN(n12905) );
  NAND2_X1 U8142 ( .A1(n8217), .A2(n8216), .ZN(n13084) );
  NAND2_X1 U8143 ( .A1(n7057), .A2(n7061), .ZN(n12977) );
  AOI21_X1 U8144 ( .B1(n10140), .B2(n8214), .A(n8011), .ZN(n14490) );
  OAI22_X1 U8145 ( .A1(n12585), .A2(SI_13_), .B1(n7489), .B2(n12801), .ZN(
        n8011) );
  AND3_X1 U8146 ( .A1(n7932), .A2(n7931), .A3(n7930), .ZN(n12661) );
  NAND2_X1 U8147 ( .A1(n7067), .A2(n15144), .ZN(n7068) );
  INV_X1 U8148 ( .A(n8280), .ZN(n7067) );
  XNOR2_X1 U8149 ( .A(n8238), .B(n12611), .ZN(n7066) );
  INV_X1 U8150 ( .A(n12949), .ZN(n13157) );
  INV_X1 U8151 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7394) );
  MUX2_X1 U8152 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7805), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7807) );
  NAND2_X1 U8153 ( .A1(n7809), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7805) );
  XNOR2_X1 U8154 ( .A(n8239), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12761) );
  MUX2_X1 U8155 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8109), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8112) );
  NAND2_X1 U8156 ( .A1(n7978), .A2(n7977), .ZN(n11462) );
  NAND2_X1 U8157 ( .A1(n8938), .A2(n8937), .ZN(n13591) );
  INV_X1 U8158 ( .A(n7397), .ZN(n6879) );
  NAND2_X1 U8159 ( .A1(n13212), .A2(n8953), .ZN(n8966) );
  INV_X1 U8160 ( .A(n8379), .ZN(n6979) );
  NAND2_X1 U8161 ( .A1(n8716), .A2(n8715), .ZN(n13651) );
  NAND2_X1 U8162 ( .A1(n8881), .A2(n8880), .ZN(n13607) );
  INV_X1 U8163 ( .A(n10723), .ZN(n10807) );
  NAND2_X1 U8164 ( .A1(n8802), .A2(n8801), .ZN(n13635) );
  NAND2_X1 U8165 ( .A1(n8839), .A2(n8838), .ZN(n13621) );
  NAND2_X1 U8166 ( .A1(n8597), .A2(n8596), .ZN(n11389) );
  NAND2_X1 U8167 ( .A1(n8760), .A2(n8759), .ZN(n13645) );
  NAND2_X1 U8168 ( .A1(n8344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7650) );
  INV_X1 U8169 ( .A(n13382), .ZN(n13581) );
  AND2_X1 U8170 ( .A1(n6623), .A2(n13584), .ZN(n6924) );
  NOR2_X1 U8171 ( .A1(n7285), .A2(n6910), .ZN(n6909) );
  OR2_X1 U8172 ( .A1(n13589), .A2(n14840), .ZN(n6991) );
  INV_X1 U8173 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10573) );
  NAND2_X1 U8174 ( .A1(n6792), .A2(n6605), .ZN(n6791) );
  OAI21_X1 U8175 ( .B1(n13746), .B2(n6790), .A(n6787), .ZN(n6792) );
  AND2_X1 U8176 ( .A1(n11841), .A2(n6624), .ZN(n6793) );
  INV_X1 U8177 ( .A(n14206), .ZN(n13774) );
  NAND2_X1 U8178 ( .A1(n9540), .A2(n9539), .ZN(n14304) );
  AND2_X1 U8179 ( .A1(n9520), .A2(n9519), .ZN(n14318) );
  NAND2_X1 U8180 ( .A1(n7097), .A2(n9482), .ZN(n14334) );
  OR2_X1 U8181 ( .A1(n10361), .A2(n10358), .ZN(n13836) );
  AND2_X1 U8182 ( .A1(n9713), .A2(n13878), .ZN(n14209) );
  NOR2_X1 U8183 ( .A1(n7176), .A2(n6884), .ZN(n14262) );
  NAND2_X1 U8184 ( .A1(n14059), .A2(n9603), .ZN(n14044) );
  NAND2_X1 U8185 ( .A1(n9567), .A2(n9566), .ZN(n14291) );
  OAI211_X1 U8186 ( .C1(n14263), .C2(n14404), .A(n6883), .B(n6882), .ZN(n14340) );
  AND3_X1 U8187 ( .A1(n7319), .A2(n7320), .A3(n14261), .ZN(n6883) );
  AOI211_X1 U8188 ( .C1(n14697), .C2(n14260), .A(n14259), .B(n14258), .ZN(
        n14261) );
  OR2_X1 U8189 ( .A1(n14393), .A2(n7249), .ZN(n7242) );
  OR2_X1 U8190 ( .A1(n14393), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7247) );
  AND2_X1 U8191 ( .A1(n9076), .A2(n9077), .ZN(n14399) );
  NOR2_X1 U8192 ( .A1(n14554), .A2(n9099), .ZN(n14558) );
  OR2_X1 U8193 ( .A1(n14558), .A2(n14557), .ZN(n7251) );
  OAI21_X1 U8194 ( .B1(n12097), .B2(n12096), .A(n12095), .ZN(n12099) );
  OAI21_X1 U8195 ( .B1(n12118), .B2(n12117), .A(n12116), .ZN(n12120) );
  NAND2_X1 U8196 ( .A1(n12130), .A2(n7477), .ZN(n7476) );
  AND2_X1 U8197 ( .A1(n7655), .A2(n7656), .ZN(n7654) );
  INV_X1 U8198 ( .A(n6696), .ZN(n7655) );
  OAI21_X1 U8199 ( .B1(n9773), .B2(n7670), .A(n6674), .ZN(n9779) );
  NAND2_X1 U8200 ( .A1(n7652), .A2(n9788), .ZN(n7651) );
  NAND2_X1 U8201 ( .A1(n7654), .A2(n7653), .ZN(n7652) );
  NAND2_X1 U8202 ( .A1(n9783), .A2(n6696), .ZN(n7653) );
  NAND2_X1 U8203 ( .A1(n12147), .A2(n12146), .ZN(n12148) );
  AND2_X1 U8204 ( .A1(n12161), .A2(n7454), .ZN(n7453) );
  NAND2_X1 U8205 ( .A1(n12151), .A2(n7455), .ZN(n7454) );
  AND2_X1 U8206 ( .A1(n12162), .A2(n12160), .ZN(n12161) );
  INV_X1 U8207 ( .A(n12164), .ZN(n7107) );
  INV_X1 U8208 ( .A(n12163), .ZN(n7106) );
  NAND2_X1 U8209 ( .A1(n6841), .A2(n6840), .ZN(n6839) );
  INV_X1 U8210 ( .A(n7688), .ZN(n6841) );
  NAND2_X1 U8211 ( .A1(n9794), .A2(n7692), .ZN(n6840) );
  AOI21_X1 U8212 ( .B1(n7453), .B2(n7456), .A(n7452), .ZN(n7451) );
  NOR2_X1 U8213 ( .A1(n7455), .A2(n12151), .ZN(n7456) );
  NAND2_X1 U8214 ( .A1(n7108), .A2(n7105), .ZN(n7452) );
  INV_X1 U8215 ( .A(n12178), .ZN(n7108) );
  AOI21_X1 U8216 ( .B1(n7661), .B2(n7660), .A(n6722), .ZN(n7658) );
  NAND2_X1 U8217 ( .A1(n6836), .A2(n6837), .ZN(n9808) );
  OAI21_X1 U8218 ( .B1(n6839), .B2(n6712), .A(n6838), .ZN(n6836) );
  NAND2_X1 U8219 ( .A1(n6839), .A2(n6712), .ZN(n6837) );
  INV_X1 U8220 ( .A(n9804), .ZN(n6838) );
  NOR2_X1 U8221 ( .A1(n6611), .A2(n7662), .ZN(n7661) );
  NAND2_X1 U8222 ( .A1(n6611), .A2(n7662), .ZN(n7660) );
  AOI21_X1 U8223 ( .B1(n12657), .B2(n12656), .A(n12750), .ZN(n7159) );
  OAI21_X1 U8224 ( .B1(n12658), .B2(n12746), .A(n6582), .ZN(n7160) );
  NAND2_X1 U8225 ( .A1(n6832), .A2(n6829), .ZN(n6828) );
  AND2_X1 U8226 ( .A1(n7674), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U8227 ( .A1(n7675), .A2(n6632), .ZN(n7674) );
  INV_X1 U8228 ( .A(n6827), .ZN(n6826) );
  OAI22_X1 U8229 ( .A1(n9825), .A2(n9824), .B1(n9828), .B2(n9829), .ZN(n6827)
         );
  NOR2_X1 U8230 ( .A1(n12219), .A2(n12218), .ZN(n7461) );
  NAND2_X1 U8231 ( .A1(n7099), .A2(n7462), .ZN(n7460) );
  AOI21_X1 U8232 ( .B1(n12219), .B2(n12218), .A(n7463), .ZN(n7462) );
  INV_X1 U8233 ( .A(n12216), .ZN(n7463) );
  NOR2_X1 U8234 ( .A1(n7665), .A2(n6717), .ZN(n7663) );
  NOR2_X1 U8235 ( .A1(n9840), .A2(n9838), .ZN(n7665) );
  NAND2_X1 U8236 ( .A1(n12227), .A2(n12225), .ZN(n7472) );
  NAND2_X1 U8237 ( .A1(n7686), .A2(n7685), .ZN(n7684) );
  INV_X1 U8238 ( .A(n9855), .ZN(n7685) );
  INV_X1 U8239 ( .A(n9854), .ZN(n7686) );
  NAND2_X1 U8240 ( .A1(n7466), .A2(n12234), .ZN(n7465) );
  AOI21_X1 U8241 ( .B1(n7162), .B2(n7161), .A(n12699), .ZN(n12704) );
  INV_X1 U8242 ( .A(n12697), .ZN(n7161) );
  INV_X1 U8243 ( .A(n7677), .ZN(n7676) );
  NAND2_X1 U8244 ( .A1(n13005), .A2(n12724), .ZN(n7137) );
  OAI22_X1 U8245 ( .A1(n12718), .A2(n13055), .B1(n12717), .B2(n12716), .ZN(
        n7138) );
  NAND2_X1 U8246 ( .A1(n12728), .A2(n12993), .ZN(n7135) );
  INV_X1 U8247 ( .A(n15047), .ZN(n12600) );
  NAND2_X1 U8248 ( .A1(n7480), .A2(n12248), .ZN(n7479) );
  INV_X1 U8249 ( .A(n10411), .ZN(n12301) );
  INV_X1 U8250 ( .A(n7144), .ZN(n7143) );
  INV_X1 U8251 ( .A(n7377), .ZN(n7376) );
  NOR2_X1 U8252 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7715) );
  NOR2_X1 U8253 ( .A1(n8551), .A2(n8550), .ZN(n8572) );
  NAND2_X1 U8254 ( .A1(n8336), .A2(n8340), .ZN(n8345) );
  INV_X1 U8255 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8336) );
  AND2_X1 U8256 ( .A1(n7114), .A2(n12254), .ZN(n7110) );
  INV_X1 U8257 ( .A(n12258), .ZN(n7113) );
  OR2_X1 U8258 ( .A1(n14371), .A2(n14014), .ZN(n12087) );
  NAND2_X1 U8259 ( .A1(n7586), .A2(n7588), .ZN(n7585) );
  OAI21_X1 U8260 ( .B1(n11267), .B2(n12312), .A(n6868), .ZN(n6871) );
  AND2_X1 U8261 ( .A1(n7586), .A2(n6869), .ZN(n6868) );
  NAND2_X1 U8262 ( .A1(n11397), .A2(n6870), .ZN(n6869) );
  INV_X1 U8263 ( .A(n9404), .ZN(n6870) );
  INV_X1 U8264 ( .A(n14140), .ZN(n7350) );
  NAND2_X1 U8265 ( .A1(n9005), .A2(n7540), .ZN(n7539) );
  INV_X1 U8266 ( .A(n9627), .ZN(n7540) );
  INV_X1 U8267 ( .A(n7539), .ZN(n7536) );
  AOI21_X1 U8268 ( .B1(n7527), .B2(n7529), .A(n7526), .ZN(n7525) );
  INV_X1 U8269 ( .A(n8706), .ZN(n7526) );
  INV_X1 U8270 ( .A(n7528), .ZN(n7527) );
  INV_X1 U8271 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9504) );
  INV_X1 U8272 ( .A(n7700), .ZN(n7121) );
  OAI21_X1 U8273 ( .B1(n10025), .B2(n7744), .A(n6982), .ZN(n8452) );
  NAND2_X1 U8274 ( .A1(n10025), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6982) );
  INV_X1 U8275 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7811) );
  NAND2_X1 U8276 ( .A1(n6952), .A2(n6950), .ZN(n9074) );
  NAND2_X1 U8277 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n6951), .ZN(n6950) );
  NAND2_X1 U8278 ( .A1(n9072), .A2(n9073), .ZN(n6952) );
  NAND2_X1 U8279 ( .A1(n10317), .A2(n15062), .ZN(n12629) );
  INV_X1 U8280 ( .A(n12541), .ZN(n7631) );
  AOI21_X1 U8281 ( .B1(n7640), .B2(n11196), .A(n6650), .ZN(n7638) );
  NOR2_X1 U8282 ( .A1(n7497), .A2(n7034), .ZN(n7495) );
  INV_X1 U8283 ( .A(n7499), .ZN(n7497) );
  AOI21_X1 U8284 ( .B1(n7499), .B2(n12622), .A(n6594), .ZN(n7496) );
  NAND2_X1 U8285 ( .A1(n14925), .A2(n11024), .ZN(n11025) );
  OR2_X1 U8286 ( .A1(n14972), .A2(n11058), .ZN(n11012) );
  NAND2_X1 U8287 ( .A1(n14999), .A2(n11030), .ZN(n11031) );
  NAND2_X1 U8288 ( .A1(n11463), .A2(n11464), .ZN(n11644) );
  INV_X1 U8289 ( .A(n6731), .ZN(n7270) );
  NAND2_X1 U8290 ( .A1(n12827), .A2(n12828), .ZN(n12846) );
  OR2_X1 U8291 ( .A1(n14468), .A2(n6739), .ZN(n6927) );
  INV_X1 U8292 ( .A(n6927), .ZN(n12875) );
  OR2_X1 U8293 ( .A1(n12920), .A2(n8245), .ZN(n12621) );
  INV_X1 U8294 ( .A(n8201), .ZN(n7381) );
  INV_X1 U8295 ( .A(n8175), .ZN(n7389) );
  OR2_X1 U8296 ( .A1(n8116), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8130) );
  NOR2_X1 U8297 ( .A1(n8130), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U8298 ( .A1(n7046), .A2(n7049), .ZN(n7043) );
  INV_X1 U8299 ( .A(n7050), .ZN(n7049) );
  AOI21_X1 U8300 ( .B1(n7513), .B2(n8266), .A(n7512), .ZN(n7511) );
  NAND2_X1 U8301 ( .A1(n7513), .A2(n7017), .ZN(n7016) );
  INV_X1 U8302 ( .A(n12694), .ZN(n7512) );
  INV_X1 U8303 ( .A(n8007), .ZN(n7383) );
  INV_X1 U8304 ( .A(n12652), .ZN(n7902) );
  INV_X1 U8305 ( .A(n7218), .ZN(n7217) );
  OAI21_X1 U8306 ( .B1(n8187), .B2(n7219), .A(n7794), .ZN(n7218) );
  INV_X1 U8307 ( .A(n7792), .ZN(n7219) );
  NOR2_X1 U8308 ( .A1(n7197), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U8309 ( .A1(n8281), .A2(n7648), .ZN(n7647) );
  INV_X1 U8310 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15353) );
  INV_X1 U8311 ( .A(n7743), .ZN(n7222) );
  INV_X1 U8312 ( .A(n8633), .ZN(n7431) );
  INV_X1 U8313 ( .A(n13263), .ZN(n7420) );
  NOR2_X1 U8314 ( .A1(n7420), .A2(n7417), .ZN(n7416) );
  INV_X1 U8315 ( .A(n13218), .ZN(n7417) );
  AND2_X1 U8316 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8460) );
  NAND2_X1 U8317 ( .A1(n13232), .A2(n8836), .ZN(n8848) );
  NOR2_X1 U8318 ( .A1(n8761), .A2(n15363), .ZN(n8777) );
  INV_X1 U8319 ( .A(n12023), .ZN(n7352) );
  NAND2_X1 U8320 ( .A1(n11695), .A2(n11696), .ZN(n7277) );
  INV_X1 U8321 ( .A(n11696), .ZN(n7273) );
  NOR2_X1 U8322 ( .A1(n8665), .A2(n8664), .ZN(n8686) );
  NAND2_X1 U8323 ( .A1(n7126), .A2(n7125), .ZN(n11859) );
  OR2_X1 U8324 ( .A1(n8644), .A2(n8643), .ZN(n8665) );
  INV_X1 U8325 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8550) );
  AND2_X1 U8326 ( .A1(n10917), .A2(n14858), .ZN(n10632) );
  INV_X1 U8327 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8328) );
  INV_X1 U8328 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8354) );
  INV_X1 U8329 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8980) );
  OR2_X1 U8330 ( .A1(n8733), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8757) );
  INV_X1 U8331 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8326) );
  OR2_X1 U8332 ( .A1(n8502), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8522) );
  INV_X1 U8333 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U8334 ( .A1(n14371), .A2(n14014), .ZN(n12088) );
  INV_X1 U8335 ( .A(n12463), .ZN(n10442) );
  AND2_X1 U8336 ( .A1(n14072), .A2(n9707), .ZN(n7346) );
  OR2_X1 U8337 ( .A1(n14298), .A2(n13843), .ZN(n9705) );
  NOR2_X1 U8338 ( .A1(n14304), .A2(n7448), .ZN(n7447) );
  INV_X1 U8339 ( .A(n7449), .ZN(n7448) );
  AND2_X1 U8340 ( .A1(n7450), .A2(n14318), .ZN(n7449) );
  INV_X1 U8341 ( .A(n7337), .ZN(n7336) );
  AND2_X1 U8342 ( .A1(n9424), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9438) );
  NOR2_X1 U8343 ( .A1(n12159), .A2(n12150), .ZN(n7444) );
  NAND2_X1 U8344 ( .A1(n11980), .A2(n9355), .ZN(n11100) );
  NOR2_X2 U8345 ( .A1(n14620), .A2(n12115), .ZN(n14621) );
  INV_X1 U8346 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9273) );
  INV_X1 U8347 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9274) );
  INV_X1 U8348 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9657) );
  INV_X1 U8349 ( .A(n9645), .ZN(n7579) );
  NAND2_X1 U8350 ( .A1(n8873), .A2(n8872), .ZN(n7166) );
  NAND2_X1 U8351 ( .A1(n8707), .A2(n10294), .ZN(n8710) );
  INV_X1 U8352 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9262) );
  INV_X1 U8353 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9407) );
  INV_X1 U8354 ( .A(n6866), .ZN(n7180) );
  INV_X1 U8355 ( .A(n8635), .ZN(n7179) );
  INV_X1 U8356 ( .A(n7183), .ZN(n7181) );
  NAND2_X1 U8357 ( .A1(n8591), .A2(n6866), .ZN(n8612) );
  AOI21_X1 U8358 ( .B1(n8586), .B2(n7519), .A(n6677), .ZN(n7518) );
  OR2_X1 U8359 ( .A1(n9370), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9409) );
  AOI21_X1 U8360 ( .B1(n8519), .B2(n7523), .A(n6678), .ZN(n7521) );
  NAND3_X1 U8361 ( .A1(n7082), .A2(n8433), .A3(n7081), .ZN(n8451) );
  NAND2_X1 U8362 ( .A1(n8430), .A2(n7084), .ZN(n7081) );
  NAND2_X1 U8363 ( .A1(n8417), .A2(n10005), .ZN(n8360) );
  NAND2_X1 U8364 ( .A1(n9028), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7256) );
  INV_X1 U8365 ( .A(n6955), .ZN(n9031) );
  OAI21_X1 U8366 ( .B1(n9038), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6613), .ZN(
        n6955) );
  XNOR2_X1 U8367 ( .A(n9031), .B(n14954), .ZN(n9055) );
  NOR2_X1 U8368 ( .A1(n9037), .A2(n9036), .ZN(n9070) );
  INV_X1 U8369 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7245) );
  OR2_X1 U8370 ( .A1(n10215), .A2(n9074), .ZN(n9078) );
  NAND2_X1 U8371 ( .A1(n9205), .A2(n8173), .ZN(n6749) );
  NOR2_X1 U8372 ( .A1(n11530), .A2(n7641), .ZN(n7640) );
  INV_X1 U8373 ( .A(n9161), .ZN(n7641) );
  NOR2_X1 U8374 ( .A1(n12502), .A2(n7634), .ZN(n7633) );
  INV_X1 U8375 ( .A(n9194), .ZN(n7634) );
  NAND2_X1 U8376 ( .A1(n12542), .A2(n12541), .ZN(n7635) );
  INV_X1 U8377 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10564) );
  OR2_X1 U8378 ( .A1(n8166), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8179) );
  OR2_X1 U8379 ( .A1(n11195), .A2(n11196), .ZN(n11193) );
  AND2_X1 U8380 ( .A1(n7934), .A2(n10959), .ZN(n7948) );
  INV_X1 U8381 ( .A(n12629), .ZN(n12627) );
  INV_X1 U8382 ( .A(n12550), .ZN(n7000) );
  XNOR2_X1 U8383 ( .A(n9139), .B(n9133), .ZN(n9138) );
  NAND2_X1 U8384 ( .A1(n10563), .A2(n10562), .ZN(n7625) );
  INV_X1 U8385 ( .A(n7157), .ZN(n7156) );
  OAI21_X1 U8386 ( .B1(n12755), .B2(n12892), .A(n12754), .ZN(n7157) );
  INV_X1 U8387 ( .A(n12619), .ZN(n7195) );
  INV_X1 U8388 ( .A(n12611), .ZN(n7231) );
  OR2_X1 U8389 ( .A1(n8314), .A2(n11628), .ZN(n9998) );
  AND2_X1 U8390 ( .A1(n10681), .A2(n10680), .ZN(n10682) );
  NOR2_X1 U8391 ( .A1(n10682), .A2(n10683), .ZN(n11021) );
  NAND2_X1 U8392 ( .A1(n10549), .A2(n14895), .ZN(n10678) );
  NOR2_X1 U8393 ( .A1(n14905), .A2(n11008), .ZN(n14924) );
  NOR2_X1 U8394 ( .A1(n14924), .A2(n14923), .ZN(n14922) );
  NAND2_X1 U8395 ( .A1(n11042), .A2(n14900), .ZN(n14920) );
  XNOR2_X1 U8396 ( .A(n11025), .B(n14951), .ZN(n14945) );
  NAND2_X1 U8397 ( .A1(n14945), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n14944) );
  NAND2_X1 U8398 ( .A1(n11063), .A2(n14965), .ZN(n14983) );
  NAND2_X1 U8399 ( .A1(n14991), .A2(n11029), .ZN(n15000) );
  NAND2_X1 U8400 ( .A1(n11075), .A2(n15006), .ZN(n15025) );
  XNOR2_X1 U8401 ( .A(n11031), .B(n15022), .ZN(n15020) );
  NAND2_X1 U8402 ( .A1(n15020), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15019) );
  NOR2_X1 U8403 ( .A1(n15002), .A2(n11070), .ZN(n6992) );
  NAND2_X1 U8404 ( .A1(n7270), .A2(n12790), .ZN(n7269) );
  INV_X1 U8405 ( .A(n12806), .ZN(n6938) );
  NAND2_X1 U8406 ( .A1(n12791), .A2(n12792), .ZN(n12793) );
  NAND2_X1 U8407 ( .A1(n12824), .A2(n12853), .ZN(n7318) );
  INV_X1 U8408 ( .A(n6754), .ZN(n12824) );
  INV_X1 U8409 ( .A(n6752), .ZN(n12839) );
  XNOR2_X1 U8410 ( .A(n12846), .B(n12853), .ZN(n12829) );
  NAND2_X1 U8411 ( .A1(n6754), .A2(n6753), .ZN(n6752) );
  AOI21_X1 U8412 ( .B1(n12854), .B2(n12853), .A(n12852), .ZN(n14456) );
  NAND2_X1 U8413 ( .A1(n14449), .A2(n12849), .ZN(n12850) );
  XNOR2_X1 U8414 ( .A(n12850), .B(n14466), .ZN(n14467) );
  NOR2_X1 U8415 ( .A1(n14475), .A2(n14476), .ZN(n14473) );
  XNOR2_X1 U8416 ( .A(n6927), .B(n6926), .ZN(n12859) );
  NAND2_X1 U8417 ( .A1(n7502), .A2(n12621), .ZN(n7501) );
  NAND2_X1 U8418 ( .A1(n7504), .A2(n12934), .ZN(n7502) );
  NAND2_X1 U8419 ( .A1(n12941), .A2(n12743), .ZN(n12933) );
  OR2_X1 U8420 ( .A1(n8179), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8194) );
  AOI21_X1 U8421 ( .B1(n7011), .B2(n7009), .A(n7008), .ZN(n7007) );
  INV_X1 U8422 ( .A(n12736), .ZN(n7008) );
  OR2_X1 U8423 ( .A1(n7387), .A2(n6572), .ZN(n7057) );
  INV_X1 U8424 ( .A(n7062), .ZN(n7061) );
  OAI21_X1 U8425 ( .B1(n7385), .B2(n6572), .A(n7065), .ZN(n7062) );
  NAND2_X1 U8426 ( .A1(n9197), .A2(n12551), .ZN(n7065) );
  AND3_X1 U8427 ( .A1(n8146), .A2(n8145), .A3(n8144), .ZN(n13021) );
  INV_X1 U8428 ( .A(n8269), .ZN(n7491) );
  INV_X1 U8429 ( .A(n13032), .ZN(n8122) );
  NAND2_X1 U8430 ( .A1(n13052), .A2(n8269), .ZN(n13041) );
  AND2_X1 U8431 ( .A1(n13013), .A2(n12719), .ZN(n13032) );
  NAND2_X1 U8432 ( .A1(n13047), .A2(n8103), .ZN(n13033) );
  AND2_X1 U8433 ( .A1(n8081), .A2(n8080), .ZN(n8096) );
  INV_X1 U8434 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n12559) );
  NAND2_X1 U8435 ( .A1(n8096), .A2(n12559), .ZN(n8116) );
  OR2_X1 U8436 ( .A1(n7999), .A2(n7724), .ZN(n8012) );
  NOR2_X1 U8437 ( .A1(n8012), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8025) );
  INV_X1 U8438 ( .A(n7509), .ZN(n7508) );
  AOI21_X1 U8439 ( .B1(n7509), .B2(n7507), .A(n7506), .ZN(n7505) );
  NOR2_X1 U8440 ( .A1(n12676), .A2(n7510), .ZN(n7509) );
  AND2_X1 U8441 ( .A1(n7980), .A2(n7979), .ZN(n11353) );
  NAND2_X1 U8442 ( .A1(n10858), .A2(n7884), .ZN(n10692) );
  INV_X1 U8443 ( .A(n15042), .ZN(n6745) );
  NOR2_X1 U8444 ( .A1(n7503), .A2(n12893), .ZN(n13144) );
  INV_X1 U8445 ( .A(n13138), .ZN(n14498) );
  AND2_X1 U8446 ( .A1(n9998), .A2(n10066), .ZN(n9242) );
  AND2_X1 U8447 ( .A1(n12746), .A2(n12756), .ZN(n10286) );
  NAND2_X1 U8448 ( .A1(n8277), .A2(n10827), .ZN(n15124) );
  NAND2_X1 U8449 ( .A1(n8297), .A2(n8296), .ZN(n10485) );
  AOI22_X1 U8450 ( .A1(n12367), .A2(n12366), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(n14363), .ZN(n12575) );
  NAND2_X1 U8451 ( .A1(n7216), .A2(n7214), .ZN(n8213) );
  AOI21_X1 U8452 ( .B1(n7217), .B2(n7219), .A(n7215), .ZN(n7214) );
  NAND2_X1 U8453 ( .A1(n8188), .A2(n7217), .ZN(n7216) );
  INV_X1 U8454 ( .A(n7795), .ZN(n7215) );
  NAND2_X1 U8455 ( .A1(n7810), .A2(n7809), .ZN(n12877) );
  MUX2_X1 U8456 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7808), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n7810) );
  NAND2_X1 U8457 ( .A1(n7957), .A2(n6932), .ZN(n6931) );
  NAND2_X1 U8458 ( .A1(n7644), .A2(n7643), .ZN(n7642) );
  INV_X1 U8459 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7643) );
  INV_X1 U8460 ( .A(n7645), .ZN(n7644) );
  XNOR2_X1 U8461 ( .A(n8241), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12630) );
  AND2_X1 U8462 ( .A1(n7781), .A2(n7780), .ZN(n8124) );
  AND2_X1 U8463 ( .A1(n7779), .A2(n7778), .ZN(n8104) );
  INV_X1 U8464 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7706) );
  INV_X1 U8465 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7705) );
  AOI21_X1 U8466 ( .B1(n7211), .B2(n7213), .A(n7209), .ZN(n7208) );
  INV_X1 U8467 ( .A(n7775), .ZN(n7209) );
  AND2_X1 U8468 ( .A1(n7777), .A2(n7776), .ZN(n8088) );
  OR2_X1 U8469 ( .A1(n8041), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8059) );
  AND2_X1 U8470 ( .A1(n7770), .A2(n7769), .ZN(n8034) );
  NAND2_X1 U8471 ( .A1(n8035), .A2(n8034), .ZN(n8037) );
  INV_X1 U8472 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U8473 ( .A1(n7755), .A2(n7754), .ZN(n7988) );
  INV_X1 U8474 ( .A(n7225), .ZN(n7224) );
  OAI22_X1 U8475 ( .A1(n7228), .A2(n6609), .B1(n10045), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n7225) );
  AND2_X1 U8476 ( .A1(n7750), .A2(n7748), .ZN(n7911) );
  AND2_X1 U8477 ( .A1(n10033), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U8478 ( .A1(n6709), .A2(n11755), .ZN(n11938) );
  NAND2_X1 U8479 ( .A1(n10878), .A2(n8539), .ZN(n10944) );
  NAND2_X1 U8480 ( .A1(n10944), .A2(n10945), .ZN(n10943) );
  NAND2_X1 U8481 ( .A1(n11412), .A2(n11413), .ZN(n11411) );
  XNOR2_X1 U8482 ( .A(n8848), .B(n8846), .ZN(n13281) );
  NAND2_X1 U8483 ( .A1(n13281), .A2(n13280), .ZN(n13279) );
  AOI21_X1 U8484 ( .B1(n7425), .B2(n7426), .A(n6682), .ZN(n7424) );
  INV_X1 U8485 ( .A(n10945), .ZN(n7425) );
  NAND2_X1 U8486 ( .A1(n10878), .A2(n6645), .ZN(n7423) );
  INV_X1 U8487 ( .A(n8749), .ZN(n7408) );
  INV_X1 U8488 ( .A(n6612), .ZN(n7411) );
  AND2_X1 U8489 ( .A1(n11937), .A2(n8744), .ZN(n7412) );
  NOR2_X1 U8490 ( .A1(n9916), .A2(n6579), .ZN(n6849) );
  INV_X1 U8491 ( .A(n7534), .ZN(n7533) );
  OAI211_X1 U8492 ( .C1(n9951), .C2(n9950), .A(n9949), .B(n9948), .ZN(n7534)
         );
  AND2_X1 U8493 ( .A1(n8380), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8385) );
  AOI21_X1 U8494 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n10174), .A(n10252), .ZN(
        n10194) );
  AOI21_X1 U8495 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n10176), .A(n14725), .ZN(
        n10180) );
  AOI21_X1 U8496 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n10276), .A(n14743), .ZN(
        n10279) );
  NAND2_X1 U8497 ( .A1(n10423), .A2(n10422), .ZN(n11476) );
  NAND2_X1 U8498 ( .A1(n14789), .A2(n11484), .ZN(n11608) );
  NAND2_X1 U8499 ( .A1(n12017), .A2(n12016), .ZN(n12018) );
  NAND2_X1 U8500 ( .A1(n13591), .A2(n13298), .ZN(n7089) );
  NAND2_X1 U8501 ( .A1(n6862), .A2(n6621), .ZN(n6861) );
  NAND2_X1 U8502 ( .A1(n7284), .A2(n13398), .ZN(n6862) );
  AND2_X1 U8503 ( .A1(n8954), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12041) );
  NAND2_X1 U8504 ( .A1(n7355), .A2(n7354), .ZN(n13399) );
  AOI21_X1 U8505 ( .B1(n7356), .B2(n12037), .A(n6630), .ZN(n7354) );
  NOR2_X1 U8506 ( .A1(n13423), .A2(n7357), .ZN(n7356) );
  INV_X1 U8507 ( .A(n7359), .ZN(n7357) );
  AND2_X1 U8508 ( .A1(n12010), .A2(n12011), .ZN(n13431) );
  NAND2_X1 U8509 ( .A1(n7299), .A2(n7296), .ZN(n7295) );
  INV_X1 U8510 ( .A(n13445), .ZN(n7296) );
  INV_X1 U8511 ( .A(n7299), .ZN(n13446) );
  NAND2_X1 U8512 ( .A1(n6573), .A2(n13462), .ZN(n13461) );
  NAND2_X1 U8513 ( .A1(n13455), .A2(n13454), .ZN(n13453) );
  NOR2_X1 U8514 ( .A1(n13629), .A2(n7130), .ZN(n7129) );
  INV_X1 U8515 ( .A(n7131), .ZN(n7130) );
  INV_X1 U8516 ( .A(n6891), .ZN(n13489) );
  AND2_X1 U8517 ( .A1(n13500), .A2(n12008), .ZN(n7263) );
  OAI21_X1 U8518 ( .B1(n6680), .B2(n7262), .A(n6584), .ZN(n7261) );
  AND2_X1 U8519 ( .A1(n8777), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U8520 ( .A1(n12006), .A2(n12005), .ZN(n13517) );
  NAND2_X1 U8521 ( .A1(n13557), .A2(n7132), .ZN(n13545) );
  NAND2_X1 U8522 ( .A1(n13557), .A2(n13563), .ZN(n13558) );
  NOR2_X2 U8523 ( .A1(n11889), .A2(n13651), .ZN(n13557) );
  NAND2_X1 U8524 ( .A1(n8736), .A2(n8735), .ZN(n11884) );
  OAI21_X1 U8525 ( .B1(n11718), .B2(n7274), .A(n7272), .ZN(n11887) );
  INV_X1 U8526 ( .A(n7276), .ZN(n7274) );
  AOI21_X1 U8527 ( .B1(n7276), .B2(n7273), .A(n6657), .ZN(n7272) );
  AND2_X1 U8528 ( .A1(n11854), .A2(n7277), .ZN(n7276) );
  NAND2_X1 U8529 ( .A1(n8686), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8737) );
  NOR2_X1 U8530 ( .A1(n13661), .A2(n11692), .ZN(n6894) );
  NAND2_X1 U8531 ( .A1(n11431), .A2(n11506), .ZN(n11721) );
  NOR2_X1 U8532 ( .A1(n6916), .A2(n6607), .ZN(n6915) );
  AND3_X1 U8533 ( .A1(n10632), .A2(n7124), .A3(n6892), .ZN(n11238) );
  NOR2_X1 U8534 ( .A1(n10835), .A2(n11141), .ZN(n6892) );
  AND2_X1 U8535 ( .A1(n11238), .A2(n11239), .ZN(n11236) );
  NAND2_X1 U8536 ( .A1(n10829), .A2(n10828), .ZN(n10831) );
  NAND2_X1 U8537 ( .A1(n10632), .A2(n10715), .ZN(n10843) );
  AND2_X1 U8538 ( .A1(n10762), .A2(n10794), .ZN(n10917) );
  NAND2_X1 U8539 ( .A1(n10614), .A2(n10613), .ZN(n10915) );
  NAND2_X1 U8540 ( .A1(n6893), .A2(n10776), .ZN(n10791) );
  INV_X1 U8541 ( .A(n10808), .ZN(n6893) );
  NOR2_X1 U8542 ( .A1(n10791), .A2(n14837), .ZN(n10794) );
  AND2_X1 U8543 ( .A1(n14877), .A2(n11360), .ZN(n10603) );
  NOR2_X1 U8544 ( .A1(n9993), .A2(n8377), .ZN(n10647) );
  AND2_X1 U8545 ( .A1(n12040), .A2(n13383), .ZN(n13582) );
  INV_X1 U8546 ( .A(n12038), .ZN(n6910) );
  NAND2_X1 U8547 ( .A1(n7275), .A2(n11696), .ZN(n11849) );
  OR2_X1 U8548 ( .A1(n11718), .A2(n11695), .ZN(n7275) );
  INV_X1 U8549 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8371) );
  AOI21_X1 U8550 ( .B1(n7568), .B2(n7570), .A(n6651), .ZN(n7566) );
  NAND2_X1 U8551 ( .A1(n7565), .A2(n11953), .ZN(n7562) );
  INV_X1 U8552 ( .A(n9568), .ZN(n9569) );
  NOR2_X1 U8553 ( .A1(n7555), .A2(n7552), .ZN(n7551) );
  INV_X1 U8554 ( .A(n11573), .ZN(n7552) );
  INV_X1 U8555 ( .A(n7560), .ZN(n7555) );
  INV_X1 U8556 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n15303) );
  NOR2_X1 U8557 ( .A1(n9533), .A2(n13732), .ZN(n9541) );
  INV_X1 U8558 ( .A(n7566), .ZN(n6790) );
  AOI21_X1 U8559 ( .B1(n7566), .B2(n6789), .A(n6788), .ZN(n6787) );
  INV_X1 U8560 ( .A(n7568), .ZN(n6789) );
  INV_X1 U8561 ( .A(n13704), .ZN(n6788) );
  INV_X1 U8562 ( .A(n10440), .ZN(n6803) );
  AND3_X1 U8563 ( .A1(n12270), .A2(n12269), .A3(n12268), .ZN(n12291) );
  INV_X1 U8564 ( .A(n9598), .ZN(n9633) );
  NAND2_X1 U8565 ( .A1(n6784), .A2(n6606), .ZN(n6783) );
  NAND2_X1 U8566 ( .A1(n9719), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U8567 ( .A1(n12285), .A2(n12284), .ZN(n12292) );
  NAND2_X1 U8568 ( .A1(n14059), .A2(n6647), .ZN(n14042) );
  NAND2_X1 U8569 ( .A1(n14057), .A2(n14056), .ZN(n14059) );
  NAND2_X1 U8570 ( .A1(n14092), .A2(n9707), .ZN(n14064) );
  NAND2_X1 U8571 ( .A1(n14092), .A2(n7346), .ZN(n14066) );
  INV_X1 U8572 ( .A(n9577), .ZN(n9578) );
  NAND2_X1 U8573 ( .A1(n14083), .A2(n14085), .ZN(n14092) );
  NAND2_X1 U8574 ( .A1(n14100), .A2(n9584), .ZN(n14088) );
  AOI21_X1 U8575 ( .B1(n14115), .B2(n14118), .A(n6659), .ZN(n7701) );
  NAND2_X1 U8576 ( .A1(n7701), .A2(n14101), .ZN(n14100) );
  NAND2_X1 U8577 ( .A1(n14198), .A2(n7449), .ZN(n14166) );
  NAND2_X1 U8578 ( .A1(n14198), .A2(n14318), .ZN(n14181) );
  NAND2_X1 U8579 ( .A1(n7595), .A2(n9516), .ZN(n14182) );
  NOR2_X1 U8580 ( .A1(n9496), .A2(n9495), .ZN(n9510) );
  OR2_X1 U8581 ( .A1(n9468), .A2(n15429), .ZN(n9496) );
  NAND2_X1 U8582 ( .A1(n9698), .A2(n9697), .ZN(n14507) );
  NAND2_X1 U8583 ( .A1(n6874), .A2(n9460), .ZN(n14516) );
  NAND2_X1 U8584 ( .A1(n11785), .A2(n12317), .ZN(n6874) );
  NAND2_X1 U8585 ( .A1(n9438), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9454) );
  OR2_X1 U8586 ( .A1(n9454), .A2(n9453), .ZN(n9468) );
  AND2_X1 U8587 ( .A1(n12170), .A2(n7442), .ZN(n7441) );
  AND4_X1 U8588 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), .ZN(n13829)
         );
  NAND2_X1 U8589 ( .A1(n11403), .A2(n7444), .ZN(n11597) );
  NAND2_X1 U8590 ( .A1(n11399), .A2(n9691), .ZN(n11373) );
  NAND2_X1 U8591 ( .A1(n11403), .A2(n14603), .ZN(n11402) );
  OR2_X1 U8592 ( .A1(n9398), .A2(n9397), .ZN(n9416) );
  NAND2_X1 U8593 ( .A1(n7594), .A2(n12299), .ZN(n11978) );
  INV_X1 U8594 ( .A(n14242), .ZN(n14622) );
  OR2_X1 U8595 ( .A1(n12264), .A2(n9296), .ZN(n9299) );
  NAND2_X1 U8596 ( .A1(n14032), .A2(n6585), .ZN(n7319) );
  AOI21_X1 U8597 ( .B1(n7321), .B2(n14611), .A(n7326), .ZN(n7320) );
  AND2_X1 U8598 ( .A1(n14034), .A2(n14209), .ZN(n7326) );
  NAND2_X1 U8599 ( .A1(n9630), .A2(n9629), .ZN(n14260) );
  AND2_X1 U8600 ( .A1(n6887), .A2(n7600), .ZN(n14136) );
  INV_X1 U8601 ( .A(n10822), .ZN(n7439) );
  OR2_X1 U8602 ( .A1(n10356), .A2(n14371), .ZN(n14702) );
  AND2_X1 U8603 ( .A1(n10246), .A2(n9673), .ZN(n10235) );
  XNOR2_X1 U8604 ( .A(n9885), .B(n9884), .ZN(n13694) );
  AND2_X1 U8605 ( .A1(n9006), .A2(n8936), .ZN(n12049) );
  OR2_X1 U8606 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NOR2_X2 U8607 ( .A1(n9656), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U8608 ( .A1(n8815), .A2(n8814), .ZN(n8819) );
  NAND2_X1 U8609 ( .A1(n8819), .A2(n8818), .ZN(n8852) );
  CLKBUF_X1 U8610 ( .A(n9479), .Z(n9490) );
  INV_X1 U8611 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9446) );
  XNOR2_X1 U8612 ( .A(n8634), .B(n7699), .ZN(n10201) );
  NAND2_X1 U8613 ( .A1(n7182), .A2(n6866), .ZN(n8634) );
  OR2_X1 U8614 ( .A1(n8613), .A2(n8612), .ZN(n7182) );
  NAND2_X1 U8615 ( .A1(n7524), .A2(n8501), .ZN(n8520) );
  NAND2_X1 U8616 ( .A1(n8499), .A2(n8498), .ZN(n7524) );
  NAND2_X1 U8617 ( .A1(n6963), .A2(n9268), .ZN(n9340) );
  INV_X1 U8618 ( .A(n8430), .ZN(n8429) );
  INV_X1 U8619 ( .A(n8413), .ZN(n8411) );
  AND2_X1 U8620 ( .A1(n6942), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9043) );
  INV_X1 U8621 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6942) );
  XNOR2_X1 U8622 ( .A(n9038), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U8623 ( .A1(n7259), .A2(n9063), .ZN(n9065) );
  NAND2_X1 U8624 ( .A1(n14392), .A2(n14391), .ZN(n7259) );
  AOI22_X1 U8625 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n15351), .B1(n9084), .B2(
        n9083), .ZN(n9088) );
  INV_X1 U8626 ( .A(n14551), .ZN(n7240) );
  INV_X1 U8627 ( .A(n7623), .ZN(n7622) );
  INV_X1 U8628 ( .A(n7619), .ZN(n7618) );
  OAI21_X1 U8629 ( .B1(n10993), .B2(n7620), .A(n6676), .ZN(n7619) );
  AND2_X1 U8630 ( .A1(n7613), .A2(n7611), .ZN(n7610) );
  INV_X1 U8631 ( .A(n7616), .ZN(n7611) );
  NAND2_X1 U8632 ( .A1(n7613), .A2(n7615), .ZN(n7612) );
  OR2_X1 U8633 ( .A1(n9218), .A2(n9217), .ZN(n7615) );
  NAND2_X1 U8634 ( .A1(n9205), .A2(n12532), .ZN(n12488) );
  NAND2_X1 U8635 ( .A1(n11193), .A2(n9161), .ZN(n11529) );
  NAND2_X1 U8636 ( .A1(n7866), .A2(n6601), .ZN(n15089) );
  NAND2_X1 U8637 ( .A1(n8215), .A2(n6966), .ZN(n7029) );
  NAND2_X1 U8638 ( .A1(n7635), .A2(n9194), .ZN(n12501) );
  INV_X1 U8639 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U8640 ( .A1(n14438), .A2(n9183), .ZN(n12523) );
  NAND2_X1 U8641 ( .A1(n14438), .A2(n7636), .ZN(n12524) );
  INV_X1 U8642 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15369) );
  NAND2_X1 U8643 ( .A1(n6775), .A2(n9200), .ZN(n12550) );
  NAND2_X1 U8644 ( .A1(n6777), .A2(n6776), .ZN(n6775) );
  INV_X1 U8645 ( .A(n9198), .ZN(n6776) );
  INV_X1 U8646 ( .A(n9199), .ZN(n6777) );
  OAI21_X1 U8647 ( .B1(n7003), .B2(n6765), .A(n6764), .ZN(n12558) );
  INV_X1 U8648 ( .A(n7636), .ZN(n6765) );
  AOI21_X1 U8649 ( .B1(n7636), .B2(n14435), .A(n6671), .ZN(n6764) );
  NAND2_X1 U8650 ( .A1(n8095), .A2(n8094), .ZN(n13056) );
  OR2_X1 U8651 ( .A1(n10408), .A2(n8191), .ZN(n8095) );
  NAND2_X1 U8652 ( .A1(n7625), .A2(n9150), .ZN(n10992) );
  AND2_X1 U8653 ( .A1(n9177), .A2(n9178), .ZN(n7627) );
  INV_X1 U8654 ( .A(n14433), .ZN(n14444) );
  INV_X1 U8655 ( .A(n12764), .ZN(n7485) );
  INV_X1 U8656 ( .A(n12783), .ZN(n10942) );
  NAND2_X1 U8657 ( .A1(n7887), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n6746) );
  INV_X1 U8658 ( .A(n7838), .ZN(n12782) );
  NOR2_X2 U8659 ( .A1(n9998), .A2(n13200), .ZN(n12783) );
  INV_X1 U8660 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14899) );
  NAND2_X1 U8661 ( .A1(n6750), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10665) );
  AOI21_X1 U8662 ( .B1(n10545), .B2(n10538), .A(n10537), .ZN(n10539) );
  NAND2_X1 U8663 ( .A1(n10539), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10681) );
  INV_X1 U8664 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14916) );
  INV_X1 U8665 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14954) );
  INV_X1 U8666 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14975) );
  INV_X1 U8667 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15016) );
  INV_X1 U8668 ( .A(n6774), .ZN(n14998) );
  NAND2_X1 U8669 ( .A1(n11461), .A2(n11460), .ZN(n11657) );
  INV_X1 U8670 ( .A(n7300), .ZN(n11639) );
  INV_X1 U8671 ( .A(n12823), .ZN(n12821) );
  INV_X1 U8672 ( .A(n6939), .ZN(n12786) );
  NOR2_X1 U8673 ( .A1(n12839), .A2(n7317), .ZN(n12838) );
  AND2_X1 U8674 ( .A1(n10556), .A2(n10555), .ZN(n14474) );
  AND2_X1 U8675 ( .A1(n7235), .A2(n7234), .ZN(n12896) );
  NAND2_X1 U8676 ( .A1(n8215), .A2(SI_31_), .ZN(n7234) );
  NAND2_X1 U8677 ( .A1(n12926), .A2(n12934), .ZN(n12925) );
  NAND2_X1 U8678 ( .A1(n7390), .A2(n8175), .ZN(n12965) );
  NAND2_X1 U8679 ( .A1(n7010), .A2(n12623), .ZN(n12975) );
  OR2_X1 U8680 ( .A1(n12994), .A2(n12624), .ZN(n7010) );
  NAND2_X1 U8681 ( .A1(n8165), .A2(n8164), .ZN(n12986) );
  NAND2_X1 U8682 ( .A1(n7064), .A2(n12589), .ZN(n12990) );
  NAND2_X1 U8683 ( .A1(n7387), .A2(n7385), .ZN(n7064) );
  NAND2_X1 U8684 ( .A1(n7387), .A2(n8134), .ZN(n13000) );
  NAND2_X1 U8685 ( .A1(n8129), .A2(n8128), .ZN(n13113) );
  OR2_X1 U8686 ( .A1(n10575), .A2(n8191), .ZN(n8129) );
  NAND2_X1 U8687 ( .A1(n7045), .A2(n7050), .ZN(n13048) );
  NAND2_X1 U8688 ( .A1(n8074), .A2(n7052), .ZN(n7045) );
  NAND2_X1 U8689 ( .A1(n8268), .A2(n12705), .ZN(n13054) );
  NAND2_X1 U8690 ( .A1(n8074), .A2(n8073), .ZN(n13062) );
  NAND2_X1 U8691 ( .A1(n7391), .A2(n8053), .ZN(n11926) );
  INV_X1 U8692 ( .A(n13029), .ZN(n13073) );
  NAND2_X1 U8693 ( .A1(n7515), .A2(n12691), .ZN(n11744) );
  NAND2_X1 U8694 ( .A1(n8024), .A2(n8023), .ZN(n14481) );
  NAND2_X1 U8695 ( .A1(n7384), .A2(n8007), .ZN(n11801) );
  OAI21_X1 U8696 ( .B1(n7370), .B2(n7040), .A(n6602), .ZN(n7384) );
  NAND2_X1 U8697 ( .A1(n11446), .A2(n7992), .ZN(n11589) );
  OAI21_X1 U8698 ( .B1(n11282), .B2(n7373), .A(n7371), .ZN(n11447) );
  NAND2_X1 U8699 ( .A1(n11349), .A2(n11348), .ZN(n11347) );
  INV_X1 U8700 ( .A(n13026), .ZN(n13071) );
  NAND2_X1 U8701 ( .A1(n8261), .A2(n12662), .ZN(n11226) );
  NAND2_X1 U8702 ( .A1(n11113), .A2(n7933), .ZN(n11228) );
  NOR2_X1 U8703 ( .A1(n7056), .A2(n6589), .ZN(n7055) );
  NOR2_X1 U8704 ( .A1(n7489), .A2(n10536), .ZN(n7056) );
  INV_X1 U8705 ( .A(n15072), .ZN(n13069) );
  OR2_X1 U8706 ( .A1(n15118), .A2(n15129), .ZN(n13138) );
  OAI21_X1 U8707 ( .B1(n12957), .B2(n7032), .A(n7030), .ZN(n12919) );
  INV_X1 U8708 ( .A(n7031), .ZN(n7030) );
  OAI21_X1 U8709 ( .B1(n8272), .B2(n7032), .A(n12917), .ZN(n7031) );
  INV_X1 U8710 ( .A(n7026), .ZN(n7022) );
  AOI21_X1 U8711 ( .B1(n12920), .B2(n7028), .A(n7027), .ZN(n7026) );
  NOR2_X1 U8712 ( .A1(n15130), .A2(n13152), .ZN(n7027) );
  INV_X1 U8713 ( .A(n12531), .ZN(n13165) );
  NAND2_X1 U8714 ( .A1(n8115), .A2(n8114), .ZN(n13184) );
  INV_X1 U8715 ( .A(n10492), .ZN(n10317) );
  OR2_X1 U8716 ( .A1(n8293), .A2(n6781), .ZN(n6780) );
  INV_X1 U8717 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8718 ( .A1(n10533), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13200) );
  NAND2_X1 U8719 ( .A1(n7395), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7721) );
  INV_X1 U8720 ( .A(n7729), .ZN(n13207) );
  NAND2_X1 U8721 ( .A1(n8190), .A2(n7792), .ZN(n8203) );
  OAI21_X1 U8722 ( .B1(n8127), .B2(n7207), .A(n7204), .ZN(n8148) );
  INV_X1 U8723 ( .A(n12630), .ZN(n10827) );
  NAND2_X1 U8724 ( .A1(n8136), .A2(n8135), .ZN(n8138) );
  NAND2_X1 U8725 ( .A1(n8127), .A2(n7781), .ZN(n8136) );
  INV_X1 U8726 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8243) );
  INV_X1 U8727 ( .A(SI_19_), .ZN(n10530) );
  INV_X1 U8728 ( .A(SI_18_), .ZN(n10407) );
  NAND2_X1 U8729 ( .A1(n8057), .A2(n7772), .ZN(n8076) );
  INV_X1 U8730 ( .A(SI_17_), .ZN(n10382) );
  INV_X1 U8731 ( .A(SI_16_), .ZN(n10294) );
  INV_X1 U8732 ( .A(SI_15_), .ZN(n10250) );
  INV_X1 U8733 ( .A(SI_14_), .ZN(n10232) );
  NAND2_X1 U8734 ( .A1(n7763), .A2(n7191), .ZN(n8008) );
  NAND2_X1 U8735 ( .A1(n7236), .A2(n7757), .ZN(n7994) );
  NAND2_X1 U8736 ( .A1(n7227), .A2(n7750), .ZN(n7926) );
  NAND2_X1 U8737 ( .A1(n7747), .A2(n7228), .ZN(n7227) );
  OR2_X1 U8738 ( .A1(n7899), .A2(n7898), .ZN(n11053) );
  OR2_X1 U8739 ( .A1(n7833), .A2(n6936), .ZN(n6935) );
  NAND2_X1 U8740 ( .A1(n8285), .A2(n7279), .ZN(n7278) );
  NAND2_X1 U8741 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6936) );
  NOR2_X1 U8742 ( .A1(n9997), .A2(n9996), .ZN(n10145) );
  AND2_X1 U8743 ( .A1(n8956), .A2(n8942), .ZN(n13419) );
  NAND2_X1 U8744 ( .A1(n6977), .A2(n8926), .ZN(n13210) );
  NAND2_X1 U8745 ( .A1(n10943), .A2(n8562), .ZN(n10999) );
  AND2_X1 U8746 ( .A1(n7401), .A2(n8772), .ZN(n7400) );
  NAND2_X1 U8747 ( .A1(n11705), .A2(n6643), .ZN(n6875) );
  NAND2_X1 U8748 ( .A1(n8776), .A2(n8775), .ZN(n13640) );
  INV_X1 U8749 ( .A(n13316), .ZN(n11181) );
  OR2_X1 U8750 ( .A1(n8394), .A2(n10331), .ZN(n8368) );
  NAND2_X1 U8751 ( .A1(n9926), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U8752 ( .A1(n7433), .A2(n7432), .ZN(n13232) );
  AND2_X1 U8753 ( .A1(n13233), .A2(n6586), .ZN(n7432) );
  AND2_X1 U8754 ( .A1(n7433), .A2(n6586), .ZN(n13234) );
  NAND2_X1 U8755 ( .A1(n7402), .A2(n7410), .ZN(n13257) );
  OR2_X1 U8756 ( .A1(n7412), .A2(n7411), .ZN(n7402) );
  NAND2_X1 U8757 ( .A1(n13264), .A2(n13263), .ZN(n13262) );
  NAND2_X1 U8758 ( .A1(n13217), .A2(n8871), .ZN(n13264) );
  AND2_X1 U8759 ( .A1(n6890), .A2(n6616), .ZN(n10506) );
  NAND2_X1 U8760 ( .A1(n13701), .A2(n8394), .ZN(n6825) );
  OR2_X1 U8761 ( .A1(n8394), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6824) );
  INV_X1 U8762 ( .A(n7433), .ZN(n13269) );
  NAND2_X1 U8763 ( .A1(n11411), .A2(n8633), .ZN(n11438) );
  NOR2_X1 U8764 ( .A1(n13252), .A2(n13524), .ZN(n13284) );
  AND2_X1 U8765 ( .A1(n9019), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13283) );
  NAND2_X1 U8766 ( .A1(n7423), .A2(n7424), .ZN(n11365) );
  NAND2_X1 U8767 ( .A1(n9020), .A2(n8423), .ZN(n7306) );
  OR2_X1 U8768 ( .A1(n9011), .A2(n9990), .ZN(n13252) );
  NAND2_X1 U8769 ( .A1(n7404), .A2(n7403), .ZN(n11966) );
  NAND2_X1 U8770 ( .A1(n7412), .A2(n7410), .ZN(n7403) );
  AOI21_X1 U8771 ( .B1(n7410), .B2(n7411), .A(n7408), .ZN(n7404) );
  NAND2_X1 U8772 ( .A1(n13242), .A2(n8911), .ZN(n13291) );
  AND2_X1 U8773 ( .A1(n8402), .A2(n8404), .ZN(n6923) );
  NAND2_X1 U8774 ( .A1(n9931), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6925) );
  OAI21_X1 U8775 ( .B1(n13334), .B2(n13329), .A(n10172), .ZN(n13332) );
  INV_X1 U8776 ( .A(n11476), .ZN(n14753) );
  XNOR2_X1 U8777 ( .A(n11608), .B(n11497), .ZN(n11485) );
  AND2_X1 U8778 ( .A1(n10178), .A2(n12050), .ZN(n14782) );
  INV_X1 U8779 ( .A(n13384), .ZN(n13385) );
  AND2_X1 U8780 ( .A1(n13397), .A2(n13396), .ZN(n7087) );
  NAND2_X1 U8781 ( .A1(n13401), .A2(n13400), .ZN(n13589) );
  OR2_X1 U8782 ( .A1(n13399), .A2(n13398), .ZN(n13400) );
  NAND2_X1 U8783 ( .A1(n7358), .A2(n7356), .ZN(n13593) );
  NAND2_X1 U8784 ( .A1(n7358), .A2(n7359), .ZN(n13424) );
  AND2_X1 U8785 ( .A1(n7362), .A2(n6620), .ZN(n13460) );
  NAND2_X1 U8786 ( .A1(n13620), .A2(n12032), .ZN(n13477) );
  INV_X1 U8787 ( .A(n7362), .ZN(n13476) );
  NOR2_X1 U8788 ( .A1(n6897), .A2(n6896), .ZN(n13514) );
  INV_X1 U8789 ( .A(n6899), .ZN(n6896) );
  INV_X1 U8790 ( .A(n6900), .ZN(n6897) );
  NAND2_X1 U8791 ( .A1(n13554), .A2(n12023), .ZN(n13534) );
  NAND2_X1 U8792 ( .A1(n12022), .A2(n12021), .ZN(n13556) );
  NAND2_X1 U8793 ( .A1(n7360), .A2(n11856), .ZN(n11858) );
  NAND2_X1 U8794 ( .A1(n6920), .A2(n11688), .ZN(n11855) );
  NAND2_X1 U8795 ( .A1(n7309), .A2(n7310), .ZN(n11690) );
  NAND2_X1 U8796 ( .A1(n7313), .A2(n7312), .ZN(n11425) );
  NAND2_X1 U8797 ( .A1(n8571), .A2(n8570), .ZN(n11190) );
  INV_X1 U8798 ( .A(n14803), .ZN(n13547) );
  NAND2_X1 U8799 ( .A1(n11136), .A2(n11135), .ZN(n11235) );
  NOR2_X1 U8800 ( .A1(n13469), .A2(n10711), .ZN(n14806) );
  INV_X1 U8801 ( .A(n6560), .ZN(n10812) );
  NAND2_X1 U8802 ( .A1(n14818), .A2(n10603), .ZN(n13571) );
  INV_X2 U8803 ( .A(n14888), .ZN(n14891) );
  INV_X1 U8804 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6911) );
  AND2_X1 U8805 ( .A1(n9017), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14818) );
  INV_X1 U8806 ( .A(n14814), .ZN(n14811) );
  NAND3_X1 U8807 ( .A1(n8352), .A2(n7367), .A3(n8351), .ZN(n13691) );
  AND2_X1 U8808 ( .A1(n8353), .A2(n8371), .ZN(n7367) );
  NAND2_X1 U8809 ( .A1(n8363), .A2(n8370), .ZN(n12050) );
  NAND2_X1 U8810 ( .A1(n8975), .A2(n8974), .ZN(n11973) );
  XNOR2_X1 U8811 ( .A(n8969), .B(n8968), .ZN(n11924) );
  INV_X1 U8812 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8968) );
  XNOR2_X1 U8813 ( .A(n8978), .B(n8977), .ZN(n11742) );
  INV_X1 U8814 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8977) );
  INV_X1 U8815 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10333) );
  INV_X1 U8816 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n15428) );
  INV_X1 U8817 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10245) );
  INV_X1 U8818 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10204) );
  INV_X1 U8819 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10138) );
  INV_X1 U8820 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10065) );
  INV_X1 U8821 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10058) );
  INV_X1 U8822 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10045) );
  INV_X1 U8823 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10039) );
  INV_X1 U8824 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10033) );
  INV_X1 U8825 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10034) );
  AND2_X2 U8826 ( .A1(n10075), .A2(n9655), .ZN(n10343) );
  NAND2_X1 U8827 ( .A1(n6786), .A2(n7566), .ZN(n13703) );
  NAND2_X1 U8828 ( .A1(n13746), .A2(n7568), .ZN(n6786) );
  NAND2_X1 U8829 ( .A1(n13795), .A2(n12424), .ZN(n13719) );
  NAND2_X1 U8830 ( .A1(n6797), .A2(n7553), .ZN(n11813) );
  NAND2_X1 U8831 ( .A1(n11574), .A2(n7551), .ZN(n6797) );
  AND4_X1 U8832 ( .A1(n9338), .A2(n9337), .A3(n9336), .A4(n9335), .ZN(n12114)
         );
  NAND2_X1 U8833 ( .A1(n13806), .A2(n12400), .ZN(n13727) );
  NAND2_X1 U8834 ( .A1(n13806), .A2(n7574), .ZN(n13728) );
  AND2_X1 U8835 ( .A1(n7558), .A2(n7561), .ZN(n11579) );
  NAND2_X1 U8836 ( .A1(n13785), .A2(n12412), .ZN(n13738) );
  NAND2_X1 U8837 ( .A1(n11824), .A2(n11823), .ZN(n11954) );
  NAND2_X1 U8838 ( .A1(n13754), .A2(n12389), .ZN(n13767) );
  NAND2_X1 U8839 ( .A1(n11559), .A2(n7560), .ZN(n11673) );
  OR2_X1 U8840 ( .A1(n10361), .A2(n10359), .ZN(n13811) );
  OAI21_X1 U8841 ( .B1(n13807), .B2(n7573), .A(n7571), .ZN(n13787) );
  AOI21_X1 U8842 ( .B1(n7572), .B2(n7574), .A(n6724), .ZN(n7571) );
  INV_X1 U8843 ( .A(n7574), .ZN(n7573) );
  NAND2_X1 U8844 ( .A1(n13787), .A2(n13786), .ZN(n13785) );
  NAND2_X1 U8845 ( .A1(n11954), .A2(n11953), .ZN(n12373) );
  AND3_X1 U8846 ( .A1(n6794), .A2(n6795), .A3(n6624), .ZN(n11840) );
  XNOR2_X1 U8847 ( .A(n10591), .B(n10590), .ZN(n7548) );
  INV_X1 U8848 ( .A(n7550), .ZN(n10594) );
  AND2_X1 U8849 ( .A1(n11302), .A2(n11300), .ZN(n7001) );
  INV_X1 U8850 ( .A(n13836), .ZN(n13809) );
  NAND2_X1 U8851 ( .A1(n7567), .A2(n12447), .ZN(n13818) );
  NAND2_X1 U8852 ( .A1(n13746), .A2(n13747), .ZN(n7567) );
  NAND2_X1 U8853 ( .A1(n9595), .A2(n9594), .ZN(n14275) );
  AND2_X1 U8854 ( .A1(n10586), .A2(n10072), .ZN(n12346) );
  OR2_X1 U8855 ( .A1(n9525), .A2(n9524), .ZN(n14206) );
  NAND4_X1 U8856 ( .A1(n9350), .A2(n9349), .A3(n9348), .A4(n9347), .ZN(n13856)
         );
  INV_X1 U8857 ( .A(n9318), .ZN(n13859) );
  INV_X1 U8858 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7813) );
  INV_X1 U8859 ( .A(n12292), .ZN(n14254) );
  NAND2_X1 U8860 ( .A1(n12262), .A2(n12261), .ZN(n14029) );
  NAND2_X1 U8861 ( .A1(n9587), .A2(n9586), .ZN(n14077) );
  NAND2_X1 U8862 ( .A1(n9576), .A2(n9575), .ZN(n14097) );
  NAND2_X1 U8863 ( .A1(n7604), .A2(n9538), .ZN(n14162) );
  NAND2_X1 U8864 ( .A1(n7604), .A2(n7602), .ZN(n14306) );
  AND2_X1 U8865 ( .A1(n14173), .A2(n12215), .ZN(n14150) );
  INV_X1 U8866 ( .A(n14318), .ZN(n14193) );
  NAND2_X1 U8867 ( .A1(n7338), .A2(n7337), .ZN(n14204) );
  AND2_X1 U8868 ( .A1(n9509), .A2(n9508), .ZN(n14202) );
  NAND2_X1 U8869 ( .A1(n14238), .A2(n12181), .ZN(n14216) );
  NAND2_X1 U8870 ( .A1(n14514), .A2(n9477), .ZN(n14247) );
  NAND2_X1 U8871 ( .A1(n9466), .A2(n9465), .ZN(n14513) );
  OAI21_X1 U8872 ( .B1(n11396), .B2(n7588), .A(n7586), .ZN(n11596) );
  INV_X1 U8873 ( .A(n14530), .ZN(n12159) );
  NAND2_X1 U8874 ( .A1(n11396), .A2(n9422), .ZN(n11377) );
  AND2_X1 U8875 ( .A1(n11262), .A2(n9690), .ZN(n11400) );
  NAND2_X1 U8876 ( .A1(n7333), .A2(n9688), .ZN(n11124) );
  NAND2_X1 U8877 ( .A1(n11162), .A2(n9686), .ZN(n7333) );
  AND2_X1 U8878 ( .A1(n12086), .A2(n12098), .ZN(n10409) );
  OR2_X1 U8879 ( .A1(n9715), .A2(n14143), .ZN(n14196) );
  NAND2_X1 U8880 ( .A1(n9317), .A2(n6960), .ZN(n10708) );
  NOR2_X1 U8881 ( .A1(n6617), .A2(n6961), .ZN(n6960) );
  INV_X1 U8882 ( .A(n14616), .ZN(n14512) );
  AND3_X2 U8883 ( .A1(n9294), .A2(n9295), .A3(n9293), .ZN(n14672) );
  INV_X1 U8884 ( .A(n14249), .ZN(n14627) );
  AND2_X1 U8885 ( .A1(n10081), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10072) );
  NAND2_X1 U8886 ( .A1(n6880), .A2(n6653), .ZN(n14358) );
  AND2_X1 U8887 ( .A1(n6998), .A2(n9281), .ZN(n7608) );
  OR2_X1 U8888 ( .A1(n9288), .A2(n6959), .ZN(n6997) );
  NAND2_X1 U8889 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n6959) );
  XNOR2_X1 U8890 ( .A(n8859), .B(SI_23_), .ZN(n11669) );
  OR2_X1 U8891 ( .A1(n9556), .A2(n10025), .ZN(n9557) );
  NAND2_X1 U8892 ( .A1(n9644), .A2(n9643), .ZN(n12275) );
  NAND2_X1 U8893 ( .A1(n7544), .A2(n8814), .ZN(n8798) );
  NAND2_X1 U8894 ( .A1(n8773), .A2(n7541), .ZN(n8774) );
  INV_X1 U8895 ( .A(n7542), .ZN(n7541) );
  INV_X1 U8896 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10390) );
  INV_X1 U8897 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n15293) );
  INV_X1 U8898 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10385) );
  INV_X1 U8899 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n15357) );
  INV_X1 U8900 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10243) );
  INV_X1 U8901 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10078) );
  INV_X1 U8902 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10063) );
  INV_X1 U8903 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10060) );
  INV_X1 U8904 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10049) );
  INV_X1 U8905 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10047) );
  INV_X1 U8906 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10028) );
  INV_X1 U8907 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10053) );
  CLKBUF_X1 U8908 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14566) );
  AND2_X1 U8909 ( .A1(n9048), .A2(n9047), .ZN(n14377) );
  XNOR2_X1 U8910 ( .A(n9039), .B(n7253), .ZN(n15462) );
  INV_X1 U8911 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7253) );
  OAI21_X1 U8912 ( .B1(n9052), .B2(n9051), .A(n15468), .ZN(n15461) );
  XNOR2_X1 U8913 ( .A(n9060), .B(n7260), .ZN(n14392) );
  INV_X1 U8914 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7260) );
  XNOR2_X1 U8915 ( .A(n9065), .B(n7258), .ZN(n15466) );
  INV_X1 U8916 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7258) );
  AND4_X1 U8917 ( .A1(n7243), .A2(n7078), .A3(n7248), .A4(n7077), .ZN(n14398)
         );
  NOR2_X1 U8918 ( .A1(n14547), .A2(n14548), .ZN(n14546) );
  NOR2_X1 U8919 ( .A1(n9091), .A2(n9090), .ZN(n14550) );
  AND2_X1 U8920 ( .A1(n9091), .A2(n9090), .ZN(n14551) );
  NOR2_X1 U8921 ( .A1(n6954), .A2(n6953), .ZN(n14553) );
  INV_X1 U8922 ( .A(n9097), .ZN(n6953) );
  INV_X1 U8923 ( .A(n9107), .ZN(n7073) );
  AND2_X1 U8924 ( .A1(n9108), .A2(n9107), .ZN(n14561) );
  AND2_X1 U8925 ( .A1(n9114), .A2(n9113), .ZN(n14411) );
  NAND2_X1 U8926 ( .A1(n6769), .A2(n6715), .ZN(n6768) );
  NOR2_X1 U8927 ( .A1(n6755), .A2(n12353), .ZN(n12360) );
  NAND2_X1 U8928 ( .A1(n6976), .A2(n6975), .ZN(n6974) );
  NAND2_X1 U8929 ( .A1(n12960), .A2(n14441), .ZN(n6975) );
  AND2_X1 U8930 ( .A1(n12573), .A2(n6725), .ZN(n6944) );
  OR2_X1 U8931 ( .A1(n12763), .A2(n12762), .ZN(n7484) );
  INV_X1 U8932 ( .A(n7302), .ZN(n11456) );
  AOI21_X1 U8933 ( .B1(n6588), .B2(n15023), .A(n6747), .ZN(n6929) );
  NAND2_X1 U8934 ( .A1(n15141), .A2(n9259), .ZN(n7069) );
  OAI21_X1 U8935 ( .B1(n12901), .B2(n8280), .A(n15130), .ZN(n8324) );
  NAND2_X1 U8936 ( .A1(n6878), .A2(n6879), .ZN(n6877) );
  NAND2_X1 U8937 ( .A1(n6986), .A2(n6984), .ZN(P2_U3233) );
  AOI21_X1 U8938 ( .B1(n13374), .B2(n13373), .A(n6985), .ZN(n6984) );
  NAND2_X1 U8939 ( .A1(n13375), .A2(n10646), .ZN(n6986) );
  OAI21_X1 U8940 ( .B1(n14767), .B2(n7812), .A(n13376), .ZN(n6985) );
  OAI21_X1 U8941 ( .B1(n13585), .B2(n14840), .A(n6924), .ZN(n13672) );
  OAI21_X1 U8942 ( .B1(n13585), .B2(n6906), .A(n6904), .ZN(P2_U3496) );
  NAND2_X1 U8943 ( .A1(n14880), .A2(n13618), .ZN(n6906) );
  INV_X1 U8944 ( .A(n6905), .ZN(n6904) );
  OAI21_X1 U8945 ( .B1(n6924), .B2(n14878), .A(n6732), .ZN(n6905) );
  NAND2_X1 U8946 ( .A1(n7086), .A2(n6733), .ZN(P2_U3495) );
  NAND2_X1 U8947 ( .A1(n13673), .A2(n14880), .ZN(n7086) );
  INV_X1 U8948 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7085) );
  XNOR2_X1 U8949 ( .A(n6791), .B(n6619), .ZN(n12473) );
  OAI21_X1 U8950 ( .B1(n14262), .B2(n14642), .A(n9729), .ZN(n9730) );
  AOI211_X1 U8951 ( .C1(n14626), .C2(n14264), .A(n12065), .B(n12064), .ZN(
        n12066) );
  AND2_X1 U8952 ( .A1(n6934), .A2(n6933), .ZN(n14046) );
  AOI21_X1 U8953 ( .B1(n14269), .B2(n14626), .A(n14045), .ZN(n6934) );
  OR2_X1 U8954 ( .A1(n14273), .A2(n14249), .ZN(n6933) );
  OR2_X1 U8955 ( .A1(n14720), .A2(n6957), .ZN(n6956) );
  INV_X1 U8956 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8957 ( .A1(n14708), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U8958 ( .A1(n14340), .A2(n14710), .ZN(n7175) );
  AND2_X1 U8959 ( .A1(n7247), .A2(n7250), .ZN(n14396) );
  NAND2_X1 U8960 ( .A1(n7248), .A2(n7242), .ZN(n14394) );
  INV_X1 U8961 ( .A(n7251), .ZN(n14556) );
  INV_X1 U8962 ( .A(n14517), .ZN(n9475) );
  AND2_X1 U8963 ( .A1(n12179), .A2(n12180), .ZN(n14517) );
  NAND2_X1 U8964 ( .A1(n14265), .A2(n9709), .ZN(n6570) );
  INV_X2 U8965 ( .A(n9743), .ZN(n9749) );
  MUX2_X2 U8966 ( .A(n12090), .B(n12089), .S(n12271), .Z(n12165) );
  NAND2_X1 U8967 ( .A1(n6709), .A2(n7413), .ZN(n7410) );
  NAND3_X1 U8968 ( .A1(n6935), .A2(n7278), .A3(n7850), .ZN(n11022) );
  OR2_X1 U8969 ( .A1(n7063), .A2(n8161), .ZN(n6572) );
  INV_X1 U8970 ( .A(n11348), .ZN(n7373) );
  AOI21_X1 U8971 ( .B1(n7183), .B2(n7180), .A(n7179), .ZN(n7178) );
  INV_X1 U8972 ( .A(n7178), .ZN(n7094) );
  AND2_X1 U8973 ( .A1(n6891), .A2(n13475), .ZN(n6573) );
  OR2_X1 U8974 ( .A1(n6634), .A2(n14234), .ZN(n6574) );
  NAND2_X1 U8975 ( .A1(n9623), .A2(n9622), .ZN(n12326) );
  OAI22_X1 U8976 ( .A1(n12587), .A2(n8191), .B1(n12586), .B2(n12585), .ZN(
        n13147) );
  NOR3_X1 U8977 ( .A1(n12193), .A2(n12192), .A3(n12198), .ZN(n6575) );
  INV_X1 U8978 ( .A(n9197), .ZN(n13172) );
  NAND2_X1 U8979 ( .A1(n8152), .A2(n8151), .ZN(n9197) );
  OAI22_X1 U8980 ( .A1(n12896), .A2(n12892), .B1(n13147), .B2(n12588), .ZN(
        n12620) );
  AND2_X1 U8981 ( .A1(n7821), .A2(n7820), .ZN(n6576) );
  INV_X1 U8982 ( .A(n12328), .ZN(n9710) );
  XNOR2_X1 U8983 ( .A(n14270), .B(n13840), .ZN(n7328) );
  INV_X1 U8984 ( .A(n7328), .ZN(n7325) );
  AND2_X1 U8985 ( .A1(n9798), .A2(n9797), .ZN(n6577) );
  AND2_X1 U8986 ( .A1(n7353), .A2(n12021), .ZN(n6578) );
  AND2_X1 U8987 ( .A1(n7511), .A2(n7016), .ZN(n6580) );
  AND2_X1 U8988 ( .A1(n14304), .A2(n13844), .ZN(n6581) );
  AND2_X1 U8989 ( .A1(n12659), .A2(n6631), .ZN(n6582) );
  OR2_X1 U8990 ( .A1(n12186), .A2(n12165), .ZN(n6583) );
  OR2_X1 U8991 ( .A1(n13629), .A2(n13523), .ZN(n6584) );
  AND2_X1 U8992 ( .A1(n6686), .A2(n14611), .ZN(n6585) );
  INV_X1 U8993 ( .A(n14796), .ZN(n7124) );
  NAND2_X1 U8994 ( .A1(n8813), .A2(n8812), .ZN(n6586) );
  OAI211_X1 U8995 ( .C1(n9449), .C2(n10028), .A(n9326), .B(n9325), .ZN(n10822)
         );
  AND2_X1 U8996 ( .A1(n6681), .A2(n9505), .ZN(n6587) );
  INV_X1 U8997 ( .A(n14435), .ZN(n7002) );
  XOR2_X1 U8998 ( .A(n12888), .B(n12887), .Z(n6588) );
  AND2_X1 U8999 ( .A1(n8215), .A2(SI_0_), .ZN(n6589) );
  AND2_X1 U9000 ( .A1(n7563), .A2(n12372), .ZN(n6590) );
  AND2_X1 U9001 ( .A1(n12152), .A2(n7453), .ZN(n6591) );
  OR2_X1 U9002 ( .A1(n11437), .A2(n7431), .ZN(n6592) );
  NAND2_X1 U9003 ( .A1(n12747), .A2(n12917), .ZN(n12934) );
  INV_X1 U9004 ( .A(n12934), .ZN(n7150) );
  NOR2_X1 U9005 ( .A1(n14282), .A2(n13841), .ZN(n6593) );
  INV_X1 U9006 ( .A(n9783), .ZN(n7656) );
  AND2_X1 U9007 ( .A1(n13147), .A2(n7503), .ZN(n6594) );
  AND2_X1 U9008 ( .A1(n7007), .A2(n7005), .ZN(n6595) );
  NAND2_X1 U9009 ( .A1(n11574), .A2(n11573), .ZN(n7558) );
  NAND2_X1 U9010 ( .A1(n7817), .A2(n7816), .ZN(n12920) );
  INV_X1 U9011 ( .A(n11150), .ZN(n7311) );
  INV_X2 U9012 ( .A(n14878), .ZN(n14880) );
  NAND2_X1 U9013 ( .A1(n8683), .A2(n8682), .ZN(n13656) );
  INV_X1 U9014 ( .A(n13656), .ZN(n7125) );
  AND2_X1 U9015 ( .A1(n10533), .A2(n12746), .ZN(n6596) );
  AND2_X1 U9016 ( .A1(n7269), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6597) );
  INV_X1 U9017 ( .A(n12463), .ZN(n12395) );
  INV_X1 U9018 ( .A(n8215), .ZN(n12585) );
  NAND2_X1 U9019 ( .A1(n9905), .A2(n9904), .ZN(n13583) );
  OR2_X1 U9020 ( .A1(n14082), .A2(n14077), .ZN(n6598) );
  NAND2_X1 U9021 ( .A1(n9918), .A2(n9917), .ZN(n6600) );
  AND2_X1 U9022 ( .A1(n7865), .A2(n7029), .ZN(n6601) );
  NAND2_X1 U9023 ( .A1(n6566), .A2(n7836), .ZN(n7847) );
  INV_X1 U9024 ( .A(n12039), .ZN(n7285) );
  NAND2_X1 U9025 ( .A1(n8205), .A2(n8204), .ZN(n12949) );
  AND2_X1 U9026 ( .A1(n7039), .A2(n8006), .ZN(n6602) );
  INV_X1 U9027 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6998) );
  AND2_X1 U9028 ( .A1(n14161), .A2(n12215), .ZN(n6603) );
  INV_X1 U9029 ( .A(n7842), .ZN(n12584) );
  AND2_X1 U9030 ( .A1(n12365), .A2(n7729), .ZN(n7842) );
  NAND2_X1 U9031 ( .A1(n7730), .A2(n7729), .ZN(n7841) );
  AND4_X1 U9032 ( .A1(n7829), .A2(n7828), .A3(n7827), .A4(n7826), .ZN(n7838)
         );
  NAND2_X1 U9033 ( .A1(n14088), .A2(n7598), .ZN(n14073) );
  AND2_X1 U9034 ( .A1(n7626), .A2(n12532), .ZN(n6604) );
  NAND2_X1 U9035 ( .A1(n12461), .A2(n12460), .ZN(n6605) );
  OR2_X1 U9036 ( .A1(n12264), .A2(n10084), .ZN(n6606) );
  AND2_X1 U9037 ( .A1(n11334), .A2(n13316), .ZN(n6607) );
  AND2_X1 U9038 ( .A1(n12531), .A2(n12767), .ZN(n6608) );
  OR2_X1 U9039 ( .A1(n7925), .A2(n7226), .ZN(n6609) );
  AND2_X1 U9040 ( .A1(n12181), .A2(n7341), .ZN(n6610) );
  AND2_X1 U9041 ( .A1(n9806), .A2(n9805), .ZN(n6611) );
  NOR2_X1 U9042 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8365) );
  NAND2_X1 U9043 ( .A1(n7762), .A2(n10243), .ZN(n7763) );
  OR2_X1 U9044 ( .A1(n13255), .A2(n13254), .ZN(n6612) );
  OR2_X1 U9045 ( .A1(n9030), .A2(n14936), .ZN(n6613) );
  INV_X1 U9046 ( .A(n14632), .ZN(n7578) );
  INV_X1 U9047 ( .A(n10741), .ZN(n10342) );
  AND2_X1 U9048 ( .A1(n6570), .A2(n7327), .ZN(n6614) );
  NOR2_X1 U9049 ( .A1(n10998), .A2(n7427), .ZN(n7426) );
  INV_X1 U9050 ( .A(n13055), .ZN(n7047) );
  AND2_X1 U9051 ( .A1(n6774), .A2(n6773), .ZN(n6615) );
  NAND2_X1 U9052 ( .A1(n8428), .A2(n8427), .ZN(n6616) );
  AND2_X1 U9053 ( .A1(n9530), .A2(n13890), .ZN(n6617) );
  INV_X1 U9054 ( .A(n12676), .ZN(n7369) );
  INV_X1 U9055 ( .A(n12019), .ZN(n6903) );
  NAND2_X1 U9056 ( .A1(n9313), .A2(n9267), .ZN(n9315) );
  OR2_X1 U9057 ( .A1(n14041), .A2(n13840), .ZN(n7327) );
  AND2_X1 U9058 ( .A1(n12214), .A2(n12215), .ZN(n14174) );
  AND4_X1 U9059 ( .A1(n7718), .A2(n7717), .A3(n7648), .A4(n8287), .ZN(n6618)
         );
  OAI211_X2 U9060 ( .C1(n6559), .C2(n10034), .A(n8400), .B(n8401), .ZN(n14831)
         );
  XNOR2_X1 U9061 ( .A(n12467), .B(n12466), .ZN(n6619) );
  OR2_X1 U9062 ( .A1(n13614), .A2(n13484), .ZN(n6620) );
  OR2_X1 U9063 ( .A1(n7287), .A2(n12039), .ZN(n6621) );
  NAND2_X1 U9064 ( .A1(n8861), .A2(n8860), .ZN(n13614) );
  INV_X1 U9065 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14936) );
  INV_X1 U9066 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8348) );
  INV_X1 U9067 ( .A(n12589), .ZN(n7063) );
  AND2_X1 U9068 ( .A1(n12774), .A2(n11353), .ZN(n6622) );
  AND3_X1 U9069 ( .A1(n7282), .A2(n6863), .A3(n6860), .ZN(n6623) );
  NOR2_X1 U9070 ( .A1(n8108), .A2(n7710), .ZN(n8110) );
  INV_X1 U9071 ( .A(n12222), .ZN(n7459) );
  NAND2_X1 U9072 ( .A1(n11811), .A2(n11810), .ZN(n6624) );
  NAND2_X1 U9073 ( .A1(n14173), .A2(n6603), .ZN(n14139) );
  NOR2_X1 U9074 ( .A1(n12839), .A2(n7316), .ZN(n6625) );
  AND4_X1 U9075 ( .A1(n7715), .A2(n7896), .A3(n7878), .A4(n7714), .ZN(n6626)
         );
  OAI22_X1 U9076 ( .A1(n12394), .A2(n7583), .B1(n14672), .B2(n12391), .ZN(
        n10349) );
  NAND2_X1 U9077 ( .A1(n8642), .A2(n8641), .ZN(n11692) );
  AND2_X1 U9078 ( .A1(n12916), .A2(n12915), .ZN(n6627) );
  AND2_X1 U9079 ( .A1(n10597), .A2(n7549), .ZN(n6628) );
  AND2_X1 U9080 ( .A1(n9141), .A2(n12781), .ZN(n6629) );
  NAND2_X1 U9081 ( .A1(n8823), .A2(n8822), .ZN(n13629) );
  AND2_X1 U9082 ( .A1(n13591), .A2(n13428), .ZN(n6630) );
  OR2_X1 U9083 ( .A1(n12660), .A2(n12746), .ZN(n6631) );
  AND2_X1 U9084 ( .A1(n9817), .A2(n9816), .ZN(n6632) );
  AND2_X1 U9085 ( .A1(n14077), .A2(n13841), .ZN(n6633) );
  OR2_X1 U9086 ( .A1(n7323), .A2(n9710), .ZN(n6634) );
  NAND2_X1 U9087 ( .A1(n7649), .A2(n8365), .ZN(n8418) );
  AND4_X1 U9088 ( .A1(n12741), .A2(n7150), .A3(n12918), .A4(n12610), .ZN(n6635) );
  OR2_X1 U9089 ( .A1(n7680), .A2(n7678), .ZN(n6636) );
  INV_X1 U9090 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8353) );
  INV_X1 U9091 ( .A(n12622), .ZN(n7504) );
  AND2_X1 U9092 ( .A1(n12304), .A2(n12299), .ZN(n6637) );
  NOR2_X1 U9093 ( .A1(n14473), .A2(n6993), .ZN(n6638) );
  NOR2_X1 U9094 ( .A1(n14248), .A2(n7607), .ZN(n7606) );
  AND2_X1 U9095 ( .A1(n7006), .A2(n7007), .ZN(n6639) );
  OR2_X1 U9096 ( .A1(n8396), .A2(n10008), .ZN(n6640) );
  INV_X1 U9097 ( .A(n14299), .ZN(n14149) );
  NAND2_X1 U9098 ( .A1(n9547), .A2(n9546), .ZN(n14299) );
  AND2_X1 U9099 ( .A1(n12721), .A2(n12720), .ZN(n6641) );
  INV_X1 U9100 ( .A(n7123), .ZN(n13441) );
  NOR2_X1 U9101 ( .A1(n13461), .A2(n13603), .ZN(n7123) );
  AND2_X1 U9102 ( .A1(n11856), .A2(n11851), .ZN(n6642) );
  AND2_X1 U9103 ( .A1(n7399), .A2(n8685), .ZN(n6643) );
  INV_X1 U9104 ( .A(n9150), .ZN(n7624) );
  OR2_X1 U9105 ( .A1(n9850), .A2(n9849), .ZN(n6644) );
  AND2_X1 U9106 ( .A1(n7426), .A2(n8539), .ZN(n6645) );
  INV_X1 U9107 ( .A(n12235), .ZN(n7466) );
  AND2_X1 U9108 ( .A1(n6872), .A2(n8911), .ZN(n6646) );
  AND2_X1 U9109 ( .A1(n7325), .A2(n9603), .ZN(n6647) );
  INV_X1 U9110 ( .A(n11953), .ZN(n7564) );
  AND2_X1 U9111 ( .A1(n6998), .A2(n9290), .ZN(n6648) );
  NAND2_X1 U9112 ( .A1(n12736), .A2(n8174), .ZN(n12976) );
  INV_X1 U9113 ( .A(n12976), .ZN(n7059) );
  AND2_X1 U9114 ( .A1(n12414), .A2(n12412), .ZN(n6649) );
  INV_X1 U9115 ( .A(n7152), .ZN(n7151) );
  NAND2_X1 U9116 ( .A1(n12958), .A2(n7153), .ZN(n7152) );
  INV_X1 U9117 ( .A(n7298), .ZN(n7297) );
  NAND2_X1 U9118 ( .A1(n7299), .A2(n13454), .ZN(n7298) );
  AND2_X1 U9119 ( .A1(n12666), .A2(n12667), .ZN(n12665) );
  AND2_X1 U9120 ( .A1(n9163), .A2(n12774), .ZN(n6650) );
  AND2_X1 U9121 ( .A1(n12454), .A2(n12453), .ZN(n6651) );
  INV_X2 U9122 ( .A(n8598), .ZN(n8526) );
  AND2_X2 U9123 ( .A1(n8383), .A2(n13696), .ZN(n8380) );
  OR2_X1 U9124 ( .A1(n9747), .A2(n9746), .ZN(n6652) );
  INV_X1 U9125 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9290) );
  AND2_X1 U9126 ( .A1(n7608), .A2(n9290), .ZN(n6653) );
  AND2_X1 U9127 ( .A1(n8270), .A2(n7490), .ZN(n6654) );
  INV_X1 U9128 ( .A(n12685), .ZN(n8019) );
  AND2_X1 U9129 ( .A1(n12691), .A2(n12688), .ZN(n12685) );
  XOR2_X1 U9130 ( .A(n12618), .B(n12883), .Z(n6655) );
  INV_X1 U9131 ( .A(n7493), .ZN(n7492) );
  NAND2_X1 U9132 ( .A1(n7047), .A2(n12705), .ZN(n7493) );
  NOR2_X1 U9133 ( .A1(n13084), .A2(n12913), .ZN(n6656) );
  NOR2_X1 U9134 ( .A1(n13656), .A2(n11850), .ZN(n6657) );
  NOR2_X1 U9135 ( .A1(n13667), .A2(n11424), .ZN(n6658) );
  NOR2_X1 U9136 ( .A1(n14128), .A2(n13843), .ZN(n6659) );
  NOR2_X1 U9137 ( .A1(n14334), .A2(n13846), .ZN(n6660) );
  OR2_X1 U9138 ( .A1(n6972), .A2(n6983), .ZN(n6661) );
  NAND2_X1 U9139 ( .A1(n7744), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6662) );
  INV_X1 U9140 ( .A(n8087), .ZN(n7054) );
  INV_X1 U9141 ( .A(n7340), .ZN(n7339) );
  NOR2_X1 U9142 ( .A1(n14227), .A2(n14208), .ZN(n7340) );
  AND2_X1 U9143 ( .A1(n9915), .A2(n9914), .ZN(n6663) );
  XOR2_X1 U9144 ( .A(n9127), .B(n7815), .Z(n6664) );
  AND2_X1 U9145 ( .A1(n7294), .A2(n7295), .ZN(n6665) );
  AND2_X1 U9146 ( .A1(n12038), .A2(n9968), .ZN(n13398) );
  INV_X1 U9147 ( .A(n13398), .ZN(n7288) );
  AND3_X1 U9148 ( .A1(n7844), .A2(n7846), .A3(n6746), .ZN(n6666) );
  AND2_X1 U9149 ( .A1(n7653), .A2(n9787), .ZN(n6667) );
  INV_X1 U9150 ( .A(n12153), .ZN(n7455) );
  NAND2_X1 U9151 ( .A1(n8636), .A2(n10139), .ZN(n8656) );
  INV_X1 U9152 ( .A(n8656), .ZN(n7529) );
  AND2_X1 U9153 ( .A1(n12741), .A2(n12740), .ZN(n6668) );
  AND2_X1 U9154 ( .A1(n10065), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U9155 ( .A1(n9506), .A2(n6587), .ZN(n6670) );
  NOR2_X1 U9156 ( .A1(n9184), .A2(n12562), .ZN(n6671) );
  NOR2_X1 U9157 ( .A1(n7614), .A2(n9218), .ZN(n6672) );
  AND2_X1 U9158 ( .A1(n12370), .A2(n12369), .ZN(n12371) );
  OR2_X1 U9159 ( .A1(n9029), .A2(n14916), .ZN(n6673) );
  INV_X1 U9160 ( .A(n7414), .ZN(n7413) );
  NAND2_X1 U9161 ( .A1(n6612), .A2(n11755), .ZN(n7414) );
  INV_X1 U9162 ( .A(n6575), .ZN(n7103) );
  AND2_X1 U9163 ( .A1(n7669), .A2(n6988), .ZN(n6674) );
  NAND2_X1 U9164 ( .A1(n14088), .A2(n9585), .ZN(n6675) );
  INV_X1 U9165 ( .A(n7133), .ZN(n7132) );
  NAND2_X1 U9166 ( .A1(n13563), .A2(n7134), .ZN(n7133) );
  NAND2_X1 U9167 ( .A1(n9152), .A2(n12778), .ZN(n6676) );
  AND2_X1 U9168 ( .A1(n8588), .A2(SI_10_), .ZN(n6677) );
  AND2_X1 U9169 ( .A1(n8521), .A2(SI_7_), .ZN(n6678) );
  OR2_X1 U9170 ( .A1(n8240), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6679) );
  INV_X1 U9171 ( .A(n12131), .ZN(n7477) );
  INV_X1 U9172 ( .A(n7380), .ZN(n7379) );
  OR2_X1 U9173 ( .A1(n8210), .A2(n7381), .ZN(n7380) );
  AND2_X1 U9174 ( .A1(n12007), .A2(n7265), .ZN(n6680) );
  NOR2_X1 U9175 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6681) );
  INV_X1 U9176 ( .A(n7599), .ZN(n7598) );
  NAND2_X1 U9177 ( .A1(n14063), .A2(n9585), .ZN(n7599) );
  AND2_X1 U9178 ( .A1(n8584), .A2(n8583), .ZN(n6682) );
  NAND2_X1 U9179 ( .A1(n12207), .A2(n12206), .ZN(n6683) );
  NAND2_X1 U9180 ( .A1(n7842), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n6684) );
  INV_X1 U9181 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10136) );
  INV_X1 U9182 ( .A(n12309), .ZN(n11130) );
  INV_X1 U9183 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9287) );
  AND2_X1 U9184 ( .A1(n11672), .A2(n7559), .ZN(n6685) );
  NAND2_X1 U9185 ( .A1(n9422), .A2(n13850), .ZN(n7589) );
  INV_X1 U9186 ( .A(n12257), .ZN(n7115) );
  OAI21_X1 U9187 ( .B1(n6578), .B2(n7352), .A(n12024), .ZN(n7351) );
  OAI21_X1 U9188 ( .B1(n11905), .B2(n7270), .A(n12790), .ZN(n12784) );
  AND2_X1 U9189 ( .A1(n7322), .A2(n9710), .ZN(n6686) );
  NAND2_X1 U9190 ( .A1(n7250), .A2(n14395), .ZN(n6687) );
  INV_X1 U9191 ( .A(n7332), .ZN(n7331) );
  NAND2_X1 U9192 ( .A1(n12309), .A2(n9688), .ZN(n7332) );
  INV_X1 U9193 ( .A(n14072), .ZN(n14063) );
  INV_X1 U9194 ( .A(n9734), .ZN(n10619) );
  OR2_X1 U9195 ( .A1(n9121), .A2(n9120), .ZN(n6688) );
  OR2_X2 U9196 ( .A1(n10343), .A2(n12288), .ZN(n12396) );
  NAND2_X1 U9197 ( .A1(n9452), .A2(n9451), .ZN(n12171) );
  AND2_X1 U9198 ( .A1(n9686), .A2(n9689), .ZN(n6689) );
  INV_X1 U9199 ( .A(n12475), .ZN(n12918) );
  AND2_X1 U9200 ( .A1(n12739), .A2(n12938), .ZN(n12958) );
  AND2_X1 U9201 ( .A1(n8122), .A2(n8103), .ZN(n6690) );
  AND2_X1 U9202 ( .A1(n8654), .A2(n11413), .ZN(n6691) );
  AND2_X1 U9203 ( .A1(n7660), .A2(n6722), .ZN(n6692) );
  AND2_X1 U9204 ( .A1(n7221), .A2(n6662), .ZN(n6693) );
  NOR2_X1 U9205 ( .A1(n12747), .A2(n12746), .ZN(n6694) );
  AND2_X1 U9206 ( .A1(n12941), .A2(n7033), .ZN(n6695) );
  AND2_X1 U9207 ( .A1(n9781), .A2(n9780), .ZN(n6696) );
  OR2_X1 U9208 ( .A1(n7466), .A2(n12234), .ZN(n6697) );
  AND2_X1 U9209 ( .A1(n9526), .A2(n9516), .ZN(n6698) );
  OR2_X1 U9210 ( .A1(n12185), .A2(n6575), .ZN(n6699) );
  OR2_X1 U9211 ( .A1(n12248), .A2(n7480), .ZN(n6700) );
  OR2_X1 U9212 ( .A1(n7666), .A2(n9839), .ZN(n6701) );
  AND2_X1 U9213 ( .A1(n7114), .A2(n12250), .ZN(n6702) );
  OR2_X1 U9214 ( .A1(n12130), .A2(n7477), .ZN(n6703) );
  NAND2_X1 U9215 ( .A1(n13603), .A2(n13294), .ZN(n6704) );
  INV_X1 U9216 ( .A(n12122), .ZN(n7470) );
  AND2_X1 U9217 ( .A1(n7719), .A2(n7394), .ZN(n6705) );
  AND2_X1 U9218 ( .A1(n9009), .A2(n7128), .ZN(n6706) );
  INV_X1 U9219 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9281) );
  INV_X1 U9220 ( .A(n7012), .ZN(n7011) );
  NAND2_X1 U9221 ( .A1(n7059), .A2(n7013), .ZN(n7012) );
  OR2_X1 U9222 ( .A1(n6632), .A2(n7675), .ZN(n6707) );
  INV_X1 U9223 ( .A(n6848), .ZN(n6847) );
  OAI21_X1 U9224 ( .B1(n6579), .B2(n6600), .A(n7533), .ZN(n6848) );
  INV_X1 U9225 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7279) );
  INV_X1 U9226 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7719) );
  INV_X1 U9227 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U9228 ( .A1(n11144), .A2(n10975), .ZN(n6708) );
  INV_X1 U9229 ( .A(n13061), .ZN(n7051) );
  INV_X1 U9230 ( .A(n12892), .ZN(n7503) );
  INV_X1 U9231 ( .A(n14085), .ZN(n7344) );
  INV_X1 U9232 ( .A(n8576), .ZN(n8463) );
  AND2_X1 U9233 ( .A1(n11705), .A2(n8685), .ZN(n6709) );
  AND2_X1 U9234 ( .A1(n13557), .A2(n7131), .ZN(n6710) );
  NAND2_X1 U9235 ( .A1(n7558), .A2(n7556), .ZN(n11559) );
  INV_X1 U9236 ( .A(n8380), .ZN(n8598) );
  NAND2_X1 U9237 ( .A1(n13137), .A2(n14415), .ZN(n6711) );
  AND2_X1 U9238 ( .A1(n9803), .A2(n9802), .ZN(n6712) );
  AND2_X1 U9239 ( .A1(n9842), .A2(n9841), .ZN(n6713) );
  NAND4_X1 U9240 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(n14034)
         );
  AND2_X1 U9241 ( .A1(n14198), .A2(n7447), .ZN(n6714) );
  INV_X1 U9242 ( .A(n15002), .ZN(n11072) );
  INV_X1 U9243 ( .A(n12968), .ZN(n7005) );
  NOR2_X1 U9244 ( .A1(n6806), .A2(n6805), .ZN(n8546) );
  AND3_X1 U9245 ( .A1(n12483), .A2(n12478), .A3(n14439), .ZN(n6715) );
  NAND2_X1 U9246 ( .A1(n8916), .A2(n8915), .ZN(n13598) );
  INV_X1 U9247 ( .A(n13598), .ZN(n7122) );
  INV_X1 U9248 ( .A(n12551), .ZN(n13002) );
  NAND2_X1 U9249 ( .A1(n7628), .A2(n9177), .ZN(n12074) );
  AND2_X1 U9250 ( .A1(n8796), .A2(n10530), .ZN(n6716) );
  OR2_X1 U9251 ( .A1(n12949), .A2(n9234), .ZN(n12743) );
  INV_X1 U9252 ( .A(n12743), .ZN(n7034) );
  AND4_X1 U9253 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n12158)
         );
  INV_X1 U9254 ( .A(n12158), .ZN(n13850) );
  NAND2_X1 U9255 ( .A1(n7044), .A2(n7042), .ZN(n13031) );
  NOR2_X1 U9256 ( .A1(n9833), .A2(n9832), .ZN(n6717) );
  AND2_X1 U9257 ( .A1(n8856), .A2(n7530), .ZN(n6718) );
  AND2_X1 U9258 ( .A1(n7635), .A2(n7633), .ZN(n6719) );
  AND2_X1 U9259 ( .A1(n14514), .A2(n7606), .ZN(n6720) );
  AOI21_X1 U9260 ( .B1(n7370), .B2(n6602), .A(n7037), .ZN(n7036) );
  AND2_X1 U9261 ( .A1(n7313), .A2(n11251), .ZN(n6721) );
  INV_X1 U9262 ( .A(SI_3_), .ZN(n6966) );
  AND2_X1 U9263 ( .A1(n9810), .A2(n9809), .ZN(n6722) );
  AND2_X1 U9264 ( .A1(n7338), .A2(n7339), .ZN(n6723) );
  AND2_X1 U9265 ( .A1(n12405), .A2(n12404), .ZN(n6724) );
  OR2_X1 U9266 ( .A1(n9197), .A2(n13002), .ZN(n12623) );
  INV_X1 U9267 ( .A(n12623), .ZN(n7009) );
  INV_X1 U9268 ( .A(n13586), .ZN(n9009) );
  OR2_X1 U9269 ( .A1(n13157), .A2(n12574), .ZN(n6725) );
  NAND2_X1 U9270 ( .A1(n14202), .A2(n14220), .ZN(n6726) );
  AND2_X1 U9271 ( .A1(n7239), .A2(n7757), .ZN(n6727) );
  AND2_X1 U9272 ( .A1(n7703), .A2(n8053), .ZN(n6728) );
  INV_X1 U9273 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U9274 ( .A1(n15130), .A2(n15105), .ZN(n13196) );
  INV_X1 U9275 ( .A(n13196), .ZN(n7028) );
  INV_X1 U9276 ( .A(n11851), .ZN(n7361) );
  AND2_X1 U9277 ( .A1(n6780), .A2(n6778), .ZN(n9129) );
  NAND2_X1 U9278 ( .A1(n8661), .A2(n8660), .ZN(n13661) );
  INV_X1 U9279 ( .A(n13661), .ZN(n7127) );
  NOR2_X2 U9280 ( .A1(n9011), .A2(n9002), .ZN(n13278) );
  NAND2_X1 U9281 ( .A1(n8172), .A2(n8171), .ZN(n12731) );
  AND2_X1 U9282 ( .A1(n11403), .A2(n7442), .ZN(n6729) );
  XOR2_X1 U9283 ( .A(n8912), .B(SI_25_), .Z(n6730) );
  NAND2_X1 U9284 ( .A1(n9532), .A2(n9531), .ZN(n14313) );
  INV_X1 U9285 ( .A(n14313), .ZN(n7450) );
  NAND2_X1 U9286 ( .A1(n14390), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6731) );
  OR2_X1 U9287 ( .A1(n14880), .A2(n6911), .ZN(n6732) );
  OR2_X1 U9288 ( .A1(n14880), .A2(n7085), .ZN(n6733) );
  NAND2_X1 U9289 ( .A1(n11431), .A2(n6894), .ZN(n11720) );
  INV_X1 U9290 ( .A(n11720), .ZN(n7126) );
  NAND2_X1 U9291 ( .A1(n10858), .A2(n7392), .ZN(n10690) );
  AND2_X1 U9292 ( .A1(n11193), .A2(n7640), .ZN(n6734) );
  AND2_X1 U9293 ( .A1(n7625), .A2(n7623), .ZN(n6735) );
  AND2_X1 U9294 ( .A1(n7333), .A2(n7331), .ZN(n6736) );
  INV_X1 U9295 ( .A(n8877), .ZN(n8876) );
  AND2_X1 U9296 ( .A1(n12801), .A2(n6731), .ZN(n6737) );
  OR2_X1 U9297 ( .A1(n8240), .A2(n7647), .ZN(n6738) );
  INV_X1 U9298 ( .A(SI_20_), .ZN(n10576) );
  INV_X1 U9299 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15234) );
  AND2_X1 U9300 ( .A1(n12858), .A2(n12857), .ZN(n6739) );
  INV_X1 U9301 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7246) );
  INV_X1 U9302 ( .A(n12884), .ZN(n6926) );
  NAND2_X1 U9303 ( .A1(n13402), .A2(n13373), .ZN(n11185) );
  NAND2_X1 U9304 ( .A1(n6994), .A2(n6997), .ZN(n13875) );
  AND2_X2 U9305 ( .A1(n10235), .A2(n10247), .ZN(n14710) );
  NAND2_X1 U9306 ( .A1(n6867), .A2(n9319), .ZN(n10816) );
  AND2_X1 U9307 ( .A1(n8042), .A2(n8059), .ZN(n12853) );
  INV_X1 U9308 ( .A(n12853), .ZN(n6753) );
  AND2_X2 U9309 ( .A1(n10488), .A2(n9258), .ZN(n15144) );
  AND2_X1 U9310 ( .A1(n10351), .A2(n7545), .ZN(n6740) );
  INV_X1 U9311 ( .A(n6804), .ZN(n10444) );
  INV_X1 U9312 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6810) );
  INV_X1 U9313 ( .A(n10646), .ZN(n13373) );
  INV_X1 U9314 ( .A(n8383), .ZN(n12067) );
  INV_X1 U9315 ( .A(n12883), .ZN(n12872) );
  INV_X1 U9316 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15382) );
  INV_X1 U9317 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6948) );
  INV_X1 U9318 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U9319 ( .A1(n7285), .A2(n13569), .ZN(n6865) );
  AND2_X1 U9320 ( .A1(n7284), .A2(n13569), .ZN(n7283) );
  INV_X2 U9321 ( .A(n13520), .ZN(n13569) );
  OAI21_X1 U9322 ( .B1(n15047), .B2(n6745), .A(n12626), .ZN(n10867) );
  NAND2_X1 U9323 ( .A1(n12626), .A2(n12635), .ZN(n15047) );
  NAND2_X2 U9324 ( .A1(n12957), .A2(n8272), .ZN(n12941) );
  NAND3_X1 U9325 ( .A1(n7716), .A2(n7957), .A3(n7396), .ZN(n7809) );
  NAND4_X1 U9326 ( .A1(n7716), .A2(n7957), .A3(n7396), .A4(n7719), .ZN(n7806)
         );
  NOR2_X4 U9327 ( .A1(n7943), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U9328 ( .A1(n7019), .A2(n6626), .ZN(n7943) );
  INV_X1 U9329 ( .A(n6749), .ZN(n7626) );
  NAND2_X1 U9330 ( .A1(n6749), .A2(n12532), .ZN(n9209) );
  INV_X1 U9331 ( .A(n10553), .ZN(n6750) );
  NAND2_X1 U9332 ( .A1(n7833), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10664) );
  NOR2_X2 U9333 ( .A1(n14460), .A2(n14459), .ZN(n14461) );
  INV_X1 U9334 ( .A(n6762), .ZN(n12871) );
  NAND2_X1 U9335 ( .A1(n12558), .A2(n12557), .ZN(n9188) );
  NAND2_X2 U9336 ( .A1(n12518), .A2(n9215), .ZN(n12567) );
  NAND2_X1 U9337 ( .A1(n12518), .A2(n6766), .ZN(n6770) );
  OAI211_X1 U9338 ( .C1(n6769), .C2(n12487), .A(n6768), .B(n12486), .ZN(
        P3_U3160) );
  NOR2_X1 U9339 ( .A1(n6771), .A2(n9166), .ZN(n11730) );
  INV_X1 U9340 ( .A(n6772), .ZN(n6771) );
  OAI21_X2 U9341 ( .B1(n12542), .B2(n7632), .A(n7629), .ZN(n9199) );
  NAND2_X1 U9342 ( .A1(n8292), .A2(n8293), .ZN(n8295) );
  NAND3_X1 U9343 ( .A1(n8292), .A2(n8293), .A3(n6779), .ZN(n6778) );
  INV_X1 U9344 ( .A(n8293), .ZN(n11628) );
  INV_X1 U9345 ( .A(n8294), .ZN(n6781) );
  NOR2_X2 U9346 ( .A1(n9999), .A2(n6629), .ZN(n10475) );
  NOR2_X2 U9347 ( .A1(n10000), .A2(n10001), .ZN(n9999) );
  NAND2_X1 U9348 ( .A1(n13719), .A2(n13720), .ZN(n12432) );
  NAND2_X1 U9349 ( .A1(n9286), .A2(n9285), .ZN(n6785) );
  NAND3_X1 U9350 ( .A1(n6794), .A2(n6795), .A3(n6793), .ZN(n11824) );
  OAI21_X1 U9351 ( .B1(n13755), .B2(n12388), .A(n6800), .ZN(n13766) );
  NAND4_X1 U9352 ( .A1(n6810), .A2(n6808), .A3(n6809), .A4(n7649), .ZN(n8435)
         );
  NAND4_X1 U9353 ( .A1(n6809), .A2(n6808), .A3(n8326), .A4(n8325), .ZN(n6805)
         );
  NAND4_X1 U9354 ( .A1(n6807), .A2(n7398), .A3(n6810), .A4(n7649), .ZN(n6806)
         );
  NAND2_X1 U9355 ( .A1(n6812), .A2(n6811), .ZN(n9763) );
  OR2_X1 U9356 ( .A1(n6815), .A2(n9757), .ZN(n6811) );
  NAND2_X1 U9357 ( .A1(n6814), .A2(n6813), .ZN(n6812) );
  INV_X1 U9358 ( .A(n9756), .ZN(n6813) );
  NAND2_X1 U9359 ( .A1(n6815), .A2(n9757), .ZN(n6814) );
  NAND2_X1 U9360 ( .A1(n7672), .A2(n7671), .ZN(n6815) );
  NAND3_X1 U9361 ( .A1(n9995), .A2(n6816), .A3(n9994), .ZN(P2_U3328) );
  OAI211_X1 U9362 ( .C1(n9989), .C2(n9963), .A(n6817), .B(n9967), .ZN(n6816)
         );
  NAND2_X1 U9363 ( .A1(n9989), .A2(n9966), .ZN(n6817) );
  NAND2_X1 U9364 ( .A1(n6820), .A2(n6819), .ZN(n6818) );
  INV_X1 U9365 ( .A(n9874), .ZN(n6819) );
  INV_X1 U9366 ( .A(n6823), .ZN(n6820) );
  NAND2_X1 U9367 ( .A1(n6822), .A2(n9873), .ZN(n6821) );
  NAND2_X1 U9368 ( .A1(n6823), .A2(n9874), .ZN(n6822) );
  NAND2_X1 U9369 ( .A1(n9868), .A2(n9867), .ZN(n6823) );
  NAND3_X1 U9370 ( .A1(n9814), .A2(n6707), .A3(n9815), .ZN(n6832) );
  OAI21_X1 U9371 ( .B1(n9784), .B2(n7654), .A(n6667), .ZN(n6833) );
  AOI21_X1 U9372 ( .B1(n9784), .B2(n7653), .A(n7651), .ZN(n6835) );
  OR2_X1 U9373 ( .A1(n9808), .A2(n7661), .ZN(n7657) );
  NAND2_X1 U9374 ( .A1(n6843), .A2(n6842), .ZN(n9850) );
  NAND2_X1 U9375 ( .A1(n6713), .A2(n6845), .ZN(n6842) );
  OR2_X1 U9376 ( .A1(n9844), .A2(n6844), .ZN(n6843) );
  NOR2_X1 U9377 ( .A1(n6713), .A2(n6845), .ZN(n6844) );
  INV_X1 U9378 ( .A(n9843), .ZN(n6845) );
  OAI211_X1 U9379 ( .C1(n6849), .C2(n6848), .A(n6846), .B(n9955), .ZN(n9960)
         );
  INV_X1 U9380 ( .A(n8794), .ZN(n6853) );
  NAND2_X1 U9381 ( .A1(n8731), .A2(n8732), .ZN(n6859) );
  NAND2_X1 U9382 ( .A1(n10816), .A2(n9327), .ZN(n9329) );
  NAND2_X1 U9383 ( .A1(n10410), .A2(n10411), .ZN(n6867) );
  NAND2_X1 U9384 ( .A1(n6871), .A2(n7584), .ZN(n9445) );
  OAI211_X2 U9385 ( .C1(n7406), .C2(n11937), .A(n6875), .B(n7400), .ZN(n13226)
         );
  OAI211_X1 U9386 ( .C1(n9010), .C2(n6877), .A(n6876), .B(n9027), .ZN(P2_U3192) );
  NAND3_X1 U9387 ( .A1(n9010), .A2(n6878), .A3(n13586), .ZN(n6876) );
  AOI22_X1 U9388 ( .A1(n7397), .A2(n13304), .B1(n9009), .B2(n13304), .ZN(n6878) );
  NAND2_X1 U9389 ( .A1(n7319), .A2(n7320), .ZN(n6884) );
  INV_X1 U9390 ( .A(n7176), .ZN(n6882) );
  NAND2_X1 U9391 ( .A1(n14340), .A2(n14720), .ZN(n6958) );
  NAND2_X4 U9392 ( .A1(n6889), .A2(n6888), .ZN(n9926) );
  NAND3_X1 U9393 ( .A1(n8363), .A2(n6566), .A3(n8370), .ZN(n6888) );
  XNOR2_X2 U9394 ( .A(n6965), .B(n8353), .ZN(n9012) );
  NAND2_X1 U9395 ( .A1(n10504), .A2(n8448), .ZN(n10497) );
  NOR2_X1 U9396 ( .A1(n13860), .A2(n12100), .ZN(n12101) );
  NAND3_X1 U9397 ( .A1(n7124), .A2(n10632), .A3(n10715), .ZN(n10982) );
  NAND2_X1 U9398 ( .A1(n6900), .A2(n6898), .ZN(n12028) );
  NAND2_X1 U9399 ( .A1(n12020), .A2(n12019), .ZN(n12022) );
  NAND2_X1 U9400 ( .A1(n13401), .A2(n6909), .ZN(n6907) );
  OR2_X1 U9401 ( .A1(n13401), .A2(n12039), .ZN(n6908) );
  OAI21_X1 U9402 ( .B1(n10970), .B2(n6708), .A(n6915), .ZN(n11178) );
  NAND2_X1 U9403 ( .A1(n6920), .A2(n6918), .ZN(n7360) );
  NAND2_X1 U9404 ( .A1(n11726), .A2(n11725), .ZN(n6920) );
  NAND2_X1 U9405 ( .A1(n10831), .A2(n10830), .ZN(n10968) );
  NAND2_X1 U9406 ( .A1(n11178), .A2(n11179), .ZN(n6921) );
  OAI22_X1 U9407 ( .A1(n10803), .A2(n10802), .B1(n6560), .B2(n13325), .ZN(
        n10769) );
  NAND2_X1 U9408 ( .A1(n13399), .A2(n13398), .ZN(n13401) );
  NAND2_X1 U9409 ( .A1(n9734), .A2(n10807), .ZN(n10607) );
  NAND2_X1 U9410 ( .A1(n11882), .A2(n11881), .ZN(n12020) );
  NAND2_X1 U9411 ( .A1(n12030), .A2(n12029), .ZN(n13496) );
  NOR2_X2 U9412 ( .A1(n14461), .A2(n12841), .ZN(n12842) );
  NOR2_X1 U9413 ( .A1(n14942), .A2(n11010), .ZN(n14958) );
  OAI22_X2 U9414 ( .A1(n11824), .A2(n7562), .B1(n6590), .B2(n12371), .ZN(
        n13711) );
  AOI21_X2 U9415 ( .B1(n11211), .B2(n11210), .A(n11209), .ZN(n11212) );
  NOR2_X2 U9416 ( .A1(n7545), .A2(n10351), .ZN(n10440) );
  NOR2_X1 U9417 ( .A1(n7546), .A2(n10375), .ZN(n7545) );
  NAND2_X1 U9418 ( .A1(n12432), .A2(n12431), .ZN(n13778) );
  NAND2_X1 U9419 ( .A1(n10932), .A2(n10931), .ZN(n11208) );
  NAND2_X1 U9420 ( .A1(n11543), .A2(n11542), .ZN(n11574) );
  OAI22_X1 U9421 ( .A1(n12391), .A2(n7578), .B1(n10345), .B2(n13867), .ZN(
        n10346) );
  NAND2_X1 U9422 ( .A1(n11301), .A2(n7001), .ZN(n11543) );
  XNOR2_X1 U9423 ( .A(n10348), .B(n6937), .ZN(n10350) );
  NAND2_X1 U9424 ( .A1(n9970), .A2(n10782), .ZN(n10771) );
  NAND2_X1 U9425 ( .A1(n8434), .A2(n9312), .ZN(n8401) );
  NAND3_X2 U9426 ( .A1(n8405), .A2(n8403), .A3(n6923), .ZN(n13323) );
  NAND3_X1 U9427 ( .A1(n8413), .A2(n8430), .A3(n8412), .ZN(n7082) );
  NAND2_X1 U9428 ( .A1(n7531), .A2(n8856), .ZN(n8858) );
  NAND2_X1 U9429 ( .A1(n10622), .A2(n9972), .ZN(n10783) );
  NAND2_X2 U9430 ( .A1(n6941), .A2(n6925), .ZN(n13325) );
  NAND2_X1 U9431 ( .A1(n10612), .A2(n10611), .ZN(n10753) );
  XNOR2_X2 U9432 ( .A(n13325), .B(n9740), .ZN(n10803) );
  NAND2_X1 U9433 ( .A1(n9209), .A2(n12533), .ZN(n12513) );
  NAND2_X1 U9434 ( .A1(n10954), .A2(n9157), .ZN(n11195) );
  NAND2_X1 U9435 ( .A1(n9188), .A2(n9187), .ZN(n12495) );
  OAI22_X1 U9436 ( .A1(n10335), .A2(n10336), .B1(n9140), .B2(n15063), .ZN(
        n10000) );
  NAND2_X1 U9437 ( .A1(n7000), .A2(n13002), .ZN(n12548) );
  NAND2_X1 U9438 ( .A1(n15030), .A2(n11089), .ZN(n6928) );
  OAI21_X1 U9439 ( .B1(n12891), .B2(n15036), .A(n6929), .ZN(P3_U3201) );
  NAND2_X1 U9440 ( .A1(n6931), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U9441 ( .A1(n14104), .A2(n14288), .ZN(n14082) );
  NAND2_X1 U9442 ( .A1(n10738), .A2(n10441), .ZN(n10820) );
  INV_X1 U9443 ( .A(n10820), .ZN(n7440) );
  OR2_X1 U9444 ( .A1(n11161), .A2(n12129), .ZN(n11159) );
  OR2_X2 U9445 ( .A1(n14133), .A2(n14128), .ZN(n14125) );
  AND2_X2 U9446 ( .A1(n11274), .A2(n11500), .ZN(n11403) );
  NAND2_X1 U9447 ( .A1(n11164), .A2(n11165), .ZN(n11163) );
  NOR2_X1 U9448 ( .A1(n6996), .A2(n6995), .ZN(n6994) );
  NAND2_X2 U9449 ( .A1(n13875), .A2(n14370), .ZN(n9305) );
  NAND2_X1 U9450 ( .A1(n13860), .A2(n14672), .ZN(n12098) );
  NAND2_X1 U9451 ( .A1(n6999), .A2(n6726), .ZN(n7595) );
  NAND2_X1 U9452 ( .A1(n9503), .A2(n9502), .ZN(n14197) );
  INV_X1 U9453 ( .A(n9280), .ZN(n6996) );
  NAND2_X1 U9454 ( .A1(n13711), .A2(n13712), .ZN(n13710) );
  NAND2_X1 U9455 ( .A1(n9191), .A2(n9190), .ZN(n12542) );
  AND3_X1 U9456 ( .A1(n8374), .A2(n8376), .A3(n8375), .ZN(n6941) );
  NAND2_X1 U9457 ( .A1(n6939), .A2(n6938), .ZN(n12823) );
  NOR2_X2 U9458 ( .A1(n11643), .A2(n11642), .ZN(n11905) );
  NAND2_X1 U9459 ( .A1(n11905), .A2(n12790), .ZN(n7267) );
  NAND2_X1 U9460 ( .A1(n10665), .A2(n10664), .ZN(n10666) );
  NAND2_X1 U9461 ( .A1(n15472), .A2(n15473), .ZN(n9045) );
  XNOR2_X1 U9462 ( .A(n9044), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15472) );
  NOR2_X2 U9463 ( .A1(n14561), .A2(n9109), .ZN(n9113) );
  NOR2_X1 U9464 ( .A1(n15469), .A2(n15470), .ZN(n9052) );
  NOR2_X2 U9465 ( .A1(n7079), .A2(n14399), .ZN(n14542) );
  OAI21_X1 U9466 ( .B1(n6571), .B2(n8108), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8109) );
  XNOR2_X1 U9467 ( .A(n9121), .B(n9120), .ZN(n14374) );
  OAI21_X1 U9468 ( .B1(n10350), .B2(n6987), .A(n10439), .ZN(n10351) );
  NAND2_X1 U9469 ( .A1(n6945), .A2(n6944), .ZN(P3_U3180) );
  NAND2_X1 U9470 ( .A1(n12569), .A2(n14439), .ZN(n6945) );
  NAND2_X1 U9471 ( .A1(n7210), .A2(n7208), .ZN(n8089) );
  NAND2_X1 U9472 ( .A1(n7158), .A2(n7156), .ZN(n7155) );
  AOI21_X1 U9473 ( .B1(n7144), .B2(n7142), .A(n6694), .ZN(n7141) );
  NAND2_X1 U9474 ( .A1(n7200), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U9475 ( .A1(n7236), .A2(n6727), .ZN(n7760) );
  NAND2_X1 U9476 ( .A1(n7764), .A2(n7763), .ZN(n8021) );
  NAND2_X1 U9477 ( .A1(n6668), .A2(n7149), .ZN(n7148) );
  NAND2_X1 U9478 ( .A1(n7192), .A2(n7484), .ZN(P3_U3296) );
  NOR2_X1 U9479 ( .A1(n9115), .A2(n14412), .ZN(n9121) );
  INV_X1 U9480 ( .A(n7072), .ZN(n9030) );
  OAI22_X1 U9481 ( .A1(n9061), .A2(n9034), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14975), .ZN(n9035) );
  INV_X1 U9482 ( .A(n6954), .ZN(n9098) );
  INV_X1 U9483 ( .A(n14546), .ZN(n7071) );
  NOR2_X1 U9484 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  OAI21_X1 U9485 ( .B1(n9040), .B2(n9041), .A(n7256), .ZN(n7255) );
  NAND2_X1 U9486 ( .A1(n7241), .A2(n7240), .ZN(n6954) );
  OAI21_X1 U9487 ( .B1(n14374), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6688), .ZN(
        n6969) );
  NAND2_X1 U9488 ( .A1(n9086), .A2(n14768), .ZN(n7070) );
  NAND2_X1 U9489 ( .A1(n7070), .A2(n7071), .ZN(n9091) );
  INV_X1 U9490 ( .A(n9055), .ZN(n6949) );
  INV_X1 U9491 ( .A(n9077), .ZN(n7077) );
  XNOR2_X1 U9492 ( .A(n6969), .B(n6664), .ZN(SUB_1596_U4) );
  NOR2_X1 U9493 ( .A1(n9064), .A2(n13940), .ZN(n9036) );
  INV_X1 U9494 ( .A(n7419), .ZN(n7418) );
  NAND2_X1 U9495 ( .A1(n10578), .A2(n8409), .ZN(n10658) );
  OAI21_X2 U9496 ( .B1(n10465), .B2(n10464), .A(n8496), .ZN(n10910) );
  NAND2_X1 U9497 ( .A1(n6958), .A2(n6956), .ZN(P1_U3557) );
  AND2_X4 U9498 ( .A1(n9305), .A2(n10006), .ZN(n12283) );
  NAND2_X1 U9499 ( .A1(n9329), .A2(n9328), .ZN(n14619) );
  INV_X1 U9501 ( .A(n7696), .ZN(n7549) );
  INV_X1 U9502 ( .A(n9315), .ZN(n6963) );
  NAND2_X1 U9503 ( .A1(n13778), .A2(n13779), .ZN(n12440) );
  MUX2_X1 U9504 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7832), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n7835) );
  INV_X1 U9505 ( .A(n9129), .ZN(n8310) );
  NAND2_X1 U9506 ( .A1(n9129), .A2(n12758), .ZN(n9132) );
  NAND2_X1 U9507 ( .A1(n12028), .A2(n12027), .ZN(n13510) );
  NAND2_X1 U9508 ( .A1(n10968), .A2(n10967), .ZN(n10970) );
  NAND2_X1 U9509 ( .A1(n7716), .A2(n7957), .ZN(n8240) );
  NAND2_X1 U9510 ( .A1(n15060), .A2(n12638), .ZN(n9137) );
  NAND3_X1 U9511 ( .A1(n6576), .A2(n6684), .A3(n7822), .ZN(n15062) );
  NAND2_X1 U9512 ( .A1(n13413), .A2(n13423), .ZN(n7090) );
  NAND2_X1 U9513 ( .A1(n6991), .A2(n6990), .ZN(n13673) );
  INV_X1 U9514 ( .A(n12014), .ZN(n13391) );
  NAND2_X1 U9515 ( .A1(n8398), .A2(n8397), .ZN(n6967) );
  INV_X1 U9516 ( .A(n7310), .ZN(n7308) );
  NAND2_X1 U9517 ( .A1(n11998), .A2(n6903), .ZN(n7303) );
  INV_X1 U9518 ( .A(n12006), .ZN(n7264) );
  OR2_X1 U9519 ( .A1(n13395), .A2(n13394), .ZN(n7088) );
  NAND2_X1 U9520 ( .A1(n7088), .A2(n13393), .ZN(n13404) );
  NAND2_X1 U9521 ( .A1(n7309), .A2(n7307), .ZN(n11694) );
  NAND2_X1 U9522 ( .A1(n8858), .A2(n8857), .ZN(n8874) );
  NAND2_X1 U9523 ( .A1(n9006), .A2(n9005), .ZN(n9628) );
  NAND2_X1 U9524 ( .A1(n7175), .A2(n7174), .ZN(P1_U3525) );
  NAND2_X1 U9525 ( .A1(n8935), .A2(n8934), .ZN(n9006) );
  NAND2_X1 U9526 ( .A1(n7166), .A2(n8874), .ZN(n8878) );
  NAND2_X1 U9527 ( .A1(n8927), .A2(SI_26_), .ZN(n8933) );
  NAND2_X1 U9528 ( .A1(n6981), .A2(n8876), .ZN(n8894) );
  INV_X1 U9529 ( .A(n12463), .ZN(n12391) );
  AOI21_X1 U9530 ( .B1(n7325), .B2(n7327), .A(n12062), .ZN(n7324) );
  OR2_X1 U9531 ( .A1(n14550), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7241) );
  NAND3_X1 U9532 ( .A1(n7074), .A2(n7251), .A3(n7073), .ZN(n7076) );
  NAND2_X1 U9533 ( .A1(n14558), .A2(n14557), .ZN(n7252) );
  NOR2_X1 U9534 ( .A1(n14553), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n9099) );
  NOR2_X1 U9535 ( .A1(n14398), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7079) );
  NAND2_X1 U9536 ( .A1(n14927), .A2(n14926), .ZN(n14925) );
  NAND3_X1 U9537 ( .A1(n6971), .A2(n9971), .A3(n6970), .ZN(n9737) );
  NAND2_X1 U9538 ( .A1(n9739), .A2(n9738), .ZN(n9747) );
  NAND3_X1 U9539 ( .A1(n9748), .A2(n7673), .A3(n6652), .ZN(n7672) );
  AOI21_X1 U9540 ( .B1(n9773), .B2(n7669), .A(n7667), .ZN(n6972) );
  OR2_X1 U9541 ( .A1(n12519), .A2(n6974), .ZN(P3_U3165) );
  OR2_X1 U9542 ( .A1(n10730), .A2(n10731), .ZN(n10728) );
  NAND2_X1 U9543 ( .A1(n6978), .A2(n8395), .ZN(n10730) );
  NAND2_X1 U9544 ( .A1(n11707), .A2(n11706), .ZN(n11705) );
  NAND2_X1 U9545 ( .A1(n13244), .A2(n13243), .ZN(n13242) );
  NAND2_X1 U9546 ( .A1(n7415), .A2(n7418), .ZN(n13244) );
  NAND2_X2 U9547 ( .A1(n13279), .A2(n8849), .ZN(n8870) );
  XNOR2_X2 U9548 ( .A(n8870), .B(n8868), .ZN(n13219) );
  NAND2_X1 U9549 ( .A1(n10496), .A2(n8473), .ZN(n10465) );
  NAND2_X1 U9550 ( .A1(n6980), .A2(n6979), .ZN(n6978) );
  INV_X1 U9551 ( .A(n8378), .ZN(n6980) );
  INV_X1 U9552 ( .A(n8878), .ZN(n6981) );
  NAND2_X1 U9553 ( .A1(n7170), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7168) );
  INV_X1 U9554 ( .A(n7148), .ZN(n7147) );
  NAND2_X1 U9555 ( .A1(n8153), .A2(n12552), .ZN(n8166) );
  NAND2_X1 U9556 ( .A1(n7193), .A2(n7485), .ZN(n7192) );
  OAI21_X1 U9557 ( .B1(n7155), .B2(n12756), .A(n7154), .ZN(n7487) );
  NAND4_X2 U9558 ( .A1(n8209), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n12928)
         );
  AOI21_X1 U9559 ( .B1(n7141), .B2(n7143), .A(n12475), .ZN(n7139) );
  NAND2_X1 U9560 ( .A1(n7140), .A2(n7139), .ZN(n12748) );
  XNOR2_X1 U9561 ( .A(n14848), .B(n10659), .ZN(n10752) );
  XNOR2_X2 U9562 ( .A(n9654), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10075) );
  AND2_X4 U9563 ( .A1(n10345), .A2(n12288), .ZN(n12463) );
  NAND2_X1 U9564 ( .A1(n7659), .A2(n7658), .ZN(n9813) );
  NAND2_X1 U9565 ( .A1(n9960), .A2(n9959), .ZN(n9989) );
  INV_X1 U9566 ( .A(n13372), .ZN(n13369) );
  XNOR2_X1 U9567 ( .A(n13362), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13372) );
  NOR2_X1 U9568 ( .A1(n13347), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13360) );
  XNOR2_X1 U9569 ( .A(n13359), .B(n13364), .ZN(n13347) );
  INV_X1 U9570 ( .A(n10349), .ZN(n6987) );
  NAND2_X1 U9571 ( .A1(n7580), .A2(n7579), .ZN(n9656) );
  NOR2_X1 U9572 ( .A1(n10376), .A2(n10377), .ZN(n10375) );
  NAND2_X1 U9573 ( .A1(n13710), .A2(n12378), .ZN(n12382) );
  NAND2_X1 U9574 ( .A1(n9506), .A2(n9505), .ZN(n9646) );
  INV_X1 U9575 ( .A(n9646), .ZN(n7580) );
  NAND2_X1 U9576 ( .A1(n7657), .A2(n6692), .ZN(n9814) );
  NAND2_X1 U9577 ( .A1(n7055), .A2(n7824), .ZN(n10492) );
  NAND2_X2 U9578 ( .A1(n9214), .A2(n12514), .ZN(n12518) );
  INV_X1 U9579 ( .A(n14436), .ZN(n7003) );
  NAND2_X1 U9580 ( .A1(n9204), .A2(n9203), .ZN(n9205) );
  NAND2_X1 U9581 ( .A1(n10888), .A2(n10887), .ZN(n10886) );
  INV_X1 U9582 ( .A(n7850), .ZN(n7019) );
  INV_X1 U9583 ( .A(n7324), .ZN(n7323) );
  INV_X1 U9584 ( .A(n7177), .ZN(n7095) );
  INV_X1 U9585 ( .A(n9730), .ZN(n9731) );
  NAND3_X1 U9586 ( .A1(n7437), .A2(n7593), .A3(n9266), .ZN(n9479) );
  INV_X1 U9587 ( .A(n14197), .ZN(n6999) );
  NAND2_X1 U9588 ( .A1(n12061), .A2(n9623), .ZN(n9638) );
  NAND2_X1 U9589 ( .A1(n14042), .A2(n7590), .ZN(n12061) );
  NAND3_X1 U9590 ( .A1(n8352), .A2(n8353), .A3(n8351), .ZN(n7281) );
  NAND2_X1 U9591 ( .A1(n7664), .A2(n6701), .ZN(n9844) );
  OAI21_X1 U9592 ( .B1(n9866), .B2(n7693), .A(n9865), .ZN(n9868) );
  NAND2_X1 U9593 ( .A1(n9733), .A2(n10646), .ZN(n10644) );
  AND2_X2 U9594 ( .A1(n8377), .A2(n11176), .ZN(n9733) );
  NAND2_X1 U9595 ( .A1(n7639), .A2(n7638), .ZN(n9165) );
  NAND2_X1 U9596 ( .A1(n10894), .A2(n12594), .ZN(n8259) );
  NAND2_X1 U9597 ( .A1(n10693), .A2(n12652), .ZN(n7004) );
  NAND2_X1 U9598 ( .A1(n8258), .A2(n12648), .ZN(n10693) );
  NAND2_X1 U9599 ( .A1(n7006), .A2(n6595), .ZN(n12969) );
  NAND2_X1 U9600 ( .A1(n8265), .A2(n6580), .ZN(n7014) );
  NAND2_X1 U9601 ( .A1(n7014), .A2(n7015), .ZN(n11780) );
  NAND2_X1 U9602 ( .A1(n13081), .A2(n7023), .ZN(n7020) );
  NAND2_X1 U9603 ( .A1(n7020), .A2(n7021), .ZN(P3_U3455) );
  AOI21_X1 U9604 ( .B1(n13081), .B2(n13138), .A(n7025), .ZN(n13151) );
  AND2_X4 U9605 ( .A1(n7836), .A2(n10006), .ZN(n8215) );
  NAND2_X1 U9606 ( .A1(n7867), .A2(n8256), .ZN(n10871) );
  INV_X1 U9607 ( .A(n7036), .ZN(n11800) );
  NAND2_X1 U9608 ( .A1(n8074), .A2(n7046), .ZN(n7044) );
  NAND2_X1 U9609 ( .A1(n7387), .A2(n7061), .ZN(n7060) );
  OAI21_X1 U9610 ( .B1(n12901), .B2(n7068), .A(n7069), .ZN(n9261) );
  NAND2_X1 U9611 ( .A1(n7074), .A2(n7251), .ZN(n9108) );
  INV_X1 U9612 ( .A(n7076), .ZN(n14560) );
  INV_X1 U9613 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7075) );
  NAND3_X1 U9614 ( .A1(n7078), .A2(n7248), .A3(n7243), .ZN(n9076) );
  NAND3_X1 U9615 ( .A1(n7544), .A2(n8814), .A3(n8797), .ZN(n8815) );
  NAND2_X1 U9616 ( .A1(n7083), .A2(n8416), .ZN(n8431) );
  NAND2_X1 U9617 ( .A1(n8413), .A2(n8412), .ZN(n7083) );
  NOR2_X2 U9618 ( .A1(n13404), .A2(n7087), .ZN(n13588) );
  NAND2_X1 U9619 ( .A1(n10384), .A2(n12259), .ZN(n7097) );
  NAND3_X1 U9620 ( .A1(n12213), .A2(n12212), .A3(n14174), .ZN(n7099) );
  NOR2_X1 U9621 ( .A1(n6699), .A2(n6591), .ZN(n7100) );
  NAND2_X1 U9622 ( .A1(n7101), .A2(n7102), .ZN(n12211) );
  OAI21_X1 U9623 ( .B1(n12185), .B2(n14517), .A(n6583), .ZN(n7104) );
  NAND3_X1 U9624 ( .A1(n12162), .A2(n7107), .A3(n7106), .ZN(n7105) );
  NAND2_X1 U9625 ( .A1(n12251), .A2(n6702), .ZN(n7111) );
  NAND3_X1 U9626 ( .A1(n7111), .A2(n7109), .A3(n7112), .ZN(n12277) );
  NAND2_X1 U9627 ( .A1(n12242), .A2(n12243), .ZN(n12241) );
  OAI21_X1 U9628 ( .B1(n8613), .B2(n7181), .A(n7178), .ZN(n8655) );
  AND2_X1 U9629 ( .A1(n13418), .A2(n6706), .ZN(n13384) );
  NAND2_X1 U9630 ( .A1(n13557), .A2(n7129), .ZN(n13488) );
  AOI21_X1 U9631 ( .B1(n7138), .B2(n6641), .A(n7137), .ZN(n7136) );
  NAND2_X1 U9632 ( .A1(n12733), .A2(n7141), .ZN(n7140) );
  AOI21_X2 U9633 ( .B1(n7147), .B2(n7152), .A(n7146), .ZN(n7145) );
  INV_X1 U9634 ( .A(n12745), .ZN(n7146) );
  INV_X1 U9635 ( .A(n12742), .ZN(n7153) );
  OAI211_X1 U9636 ( .C1(n7160), .C2(n7159), .A(n12664), .B(n12665), .ZN(n12670) );
  NAND3_X1 U9637 ( .A1(n7164), .A2(n7163), .A3(n12698), .ZN(n7162) );
  NAND3_X1 U9638 ( .A1(n12690), .A2(n12689), .A3(n12750), .ZN(n7163) );
  NAND3_X1 U9639 ( .A1(n12695), .A2(n12746), .A3(n12694), .ZN(n7164) );
  NAND3_X1 U9640 ( .A1(n8499), .A2(n8519), .A3(n8498), .ZN(n7522) );
  NAND2_X1 U9641 ( .A1(n12060), .A2(n9709), .ZN(n9622) );
  NAND2_X1 U9642 ( .A1(n12048), .A2(n9433), .ZN(n7167) );
  NAND3_X1 U9643 ( .A1(n7815), .A2(n7814), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7170) );
  NAND3_X1 U9644 ( .A1(n7812), .A2(n7811), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7171) );
  NAND2_X1 U9645 ( .A1(n7323), .A2(n9710), .ZN(n7185) );
  AOI22_X1 U9646 ( .A1(n7185), .A2(n7322), .B1(n7186), .B2(n7189), .ZN(n7321)
         );
  OAI21_X1 U9647 ( .B1(n12062), .B2(n7327), .A(n6570), .ZN(n7188) );
  NAND3_X1 U9648 ( .A1(n7763), .A2(P1_DATAO_REG_13__SCAN_IN), .A3(n7191), .ZN(
        n7764) );
  NAND3_X1 U9649 ( .A1(n7487), .A2(n7486), .A3(n7194), .ZN(n7193) );
  NAND2_X1 U9650 ( .A1(n7789), .A2(n7790), .ZN(n8176) );
  NAND2_X1 U9651 ( .A1(n7198), .A2(n7196), .ZN(n7790) );
  NAND2_X1 U9652 ( .A1(n7198), .A2(n7787), .ZN(n7788) );
  INV_X1 U9653 ( .A(n7787), .ZN(n7197) );
  INV_X1 U9654 ( .A(n8163), .ZN(n7200) );
  NAND2_X1 U9655 ( .A1(n8127), .A2(n7204), .ZN(n7203) );
  NAND2_X1 U9656 ( .A1(n8055), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U9657 ( .A1(n8188), .A2(n8187), .ZN(n8190) );
  OAI21_X1 U9658 ( .B1(n7862), .B2(n7220), .A(n6693), .ZN(n7894) );
  NAND3_X1 U9659 ( .A1(n7223), .A2(n7875), .A3(n7222), .ZN(n7221) );
  OAI21_X1 U9660 ( .B1(n7862), .B2(n7742), .A(n7743), .ZN(n7876) );
  NAND2_X1 U9661 ( .A1(n7747), .A2(n7746), .ZN(n7912) );
  XNOR2_X1 U9662 ( .A(n7230), .B(n12872), .ZN(n12757) );
  NAND4_X1 U9663 ( .A1(n12755), .A2(n12615), .A3(n7231), .A4(n6635), .ZN(n7230) );
  NAND2_X1 U9664 ( .A1(n13201), .A2(n8214), .ZN(n7235) );
  NAND2_X1 U9665 ( .A1(n7755), .A2(n7237), .ZN(n7236) );
  OR2_X1 U9666 ( .A1(n7250), .A2(n14395), .ZN(n7248) );
  OR2_X1 U9667 ( .A1(n14395), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7249) );
  INV_X1 U9668 ( .A(n7255), .ZN(n9029) );
  AOI21_X2 U9669 ( .B1(n7264), .B2(n7263), .A(n7261), .ZN(n13482) );
  NAND3_X1 U9670 ( .A1(n7268), .A2(n7269), .A3(n7267), .ZN(n11906) );
  INV_X1 U9671 ( .A(n7271), .ZN(n12785) );
  AND2_X2 U9672 ( .A1(n8333), .A2(n8546), .ZN(n8352) );
  NAND2_X1 U9673 ( .A1(n12014), .A2(n7283), .ZN(n7282) );
  NOR2_X1 U9674 ( .A1(n12014), .A2(n13398), .ZN(n13394) );
  NAND2_X1 U9675 ( .A1(n13455), .A2(n7291), .ZN(n7290) );
  NAND2_X1 U9676 ( .A1(n13455), .A2(n7297), .ZN(n7294) );
  OAI21_X2 U9677 ( .B1(n13566), .B2(n12001), .A(n12003), .ZN(n13536) );
  INV_X2 U9678 ( .A(n10610), .ZN(n13322) );
  NAND2_X1 U9679 ( .A1(n11252), .A2(n7312), .ZN(n7309) );
  INV_X1 U9680 ( .A(n11252), .ZN(n7314) );
  NAND2_X1 U9681 ( .A1(n7314), .A2(n11150), .ZN(n7313) );
  INV_X1 U9682 ( .A(n7318), .ZN(n7316) );
  OAI21_X1 U9683 ( .B1(n14032), .B2(n7325), .A(n7327), .ZN(n12052) );
  NAND2_X1 U9684 ( .A1(n11162), .A2(n6689), .ZN(n7330) );
  OAI21_X1 U9685 ( .B1(n14238), .B2(n7336), .A(n7334), .ZN(n14186) );
  NAND2_X1 U9686 ( .A1(n7342), .A2(n12107), .ZN(n10817) );
  NAND4_X1 U9687 ( .A1(n12086), .A2(n12107), .A3(n12106), .A4(n12098), .ZN(
        n7342) );
  OAI21_X2 U9688 ( .B1(n14083), .B2(n7345), .A(n7343), .ZN(n14048) );
  NAND2_X1 U9689 ( .A1(n11373), .A2(n9692), .ZN(n9694) );
  NAND2_X1 U9690 ( .A1(n7348), .A2(n7349), .ZN(n9703) );
  NAND2_X1 U9691 ( .A1(n14172), .A2(n6603), .ZN(n7348) );
  OAI21_X2 U9692 ( .B1(n14507), .B2(n9699), .A(n12180), .ZN(n14236) );
  NAND2_X1 U9693 ( .A1(n11103), .A2(n9685), .ZN(n11162) );
  NAND2_X1 U9694 ( .A1(n11264), .A2(n11263), .ZN(n11262) );
  NAND2_X1 U9695 ( .A1(n14186), .A2(n14185), .ZN(n14184) );
  NAND2_X1 U9696 ( .A1(n11984), .A2(n9683), .ZN(n11104) );
  OAI21_X1 U9697 ( .B1(n14608), .B2(n9682), .A(n9681), .ZN(n11982) );
  NAND2_X1 U9698 ( .A1(n9700), .A2(n14248), .ZN(n14238) );
  NOR2_X2 U9699 ( .A1(n13591), .A2(n13432), .ZN(n13418) );
  NAND2_X1 U9700 ( .A1(n13430), .A2(n7356), .ZN(n7355) );
  CLKBUF_X1 U9701 ( .A(n7364), .Z(n7362) );
  NAND2_X1 U9702 ( .A1(n8352), .A2(n8351), .ZN(n8370) );
  NAND2_X1 U9703 ( .A1(n11282), .A2(n7371), .ZN(n7370) );
  NAND2_X1 U9704 ( .A1(n12955), .A2(n8201), .ZN(n12943) );
  NAND2_X1 U9705 ( .A1(n7390), .A2(n7388), .ZN(n8186) );
  NAND2_X1 U9706 ( .A1(n7391), .A2(n6728), .ZN(n8074) );
  AND2_X1 U9707 ( .A1(n7902), .A2(n7884), .ZN(n7392) );
  NAND4_X1 U9708 ( .A1(n7396), .A2(n7716), .A3(n6705), .A4(n7957), .ZN(n7395)
         );
  NAND2_X1 U9709 ( .A1(n13219), .A2(n7416), .ZN(n7415) );
  NAND2_X1 U9710 ( .A1(n11412), .A2(n6691), .ZN(n7429) );
  NAND2_X1 U9711 ( .A1(n7429), .A2(n7430), .ZN(n11707) );
  NAND2_X1 U9712 ( .A1(n8792), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U9713 ( .A1(n8792), .A2(n13224), .ZN(n13270) );
  NOR2_X1 U9714 ( .A1(n13271), .A2(n7435), .ZN(n7434) );
  INV_X1 U9715 ( .A(n13224), .ZN(n7435) );
  NOR2_X4 U9716 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9313) );
  AND4_X2 U9717 ( .A1(n7438), .A2(n9406), .A3(n9262), .A4(n9407), .ZN(n9266)
         );
  NOR2_X2 U9718 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7438) );
  NOR2_X2 U9719 ( .A1(n6598), .A2(n14275), .ZN(n14051) );
  NOR2_X2 U9720 ( .A1(n14125), .A2(n14291), .ZN(n14104) );
  NOR2_X2 U9721 ( .A1(n12100), .A2(n14632), .ZN(n10738) );
  NAND2_X1 U9722 ( .A1(n11403), .A2(n7441), .ZN(n14518) );
  NAND2_X1 U9723 ( .A1(n7460), .A2(n7458), .ZN(n12221) );
  NAND3_X1 U9724 ( .A1(n12232), .A2(n12233), .A3(n6697), .ZN(n7464) );
  NAND2_X1 U9725 ( .A1(n7467), .A2(n7469), .ZN(n12126) );
  NAND3_X1 U9726 ( .A1(n12120), .A2(n7468), .A3(n12119), .ZN(n7467) );
  NAND2_X1 U9727 ( .A1(n7471), .A2(n7472), .ZN(n12231) );
  NAND3_X1 U9728 ( .A1(n12224), .A2(n7473), .A3(n12223), .ZN(n7471) );
  NAND2_X1 U9729 ( .A1(n7475), .A2(n7476), .ZN(n12135) );
  NAND3_X1 U9730 ( .A1(n12128), .A2(n6703), .A3(n12127), .ZN(n7475) );
  NAND2_X1 U9731 ( .A1(n7478), .A2(n7479), .ZN(n12252) );
  NAND3_X1 U9732 ( .A1(n12247), .A2(n12246), .A3(n6700), .ZN(n7478) );
  NOR2_X1 U9733 ( .A1(n6596), .A2(n8113), .ZN(n10540) );
  OAI21_X2 U9734 ( .B1(n8268), .B2(n7491), .A(n6654), .ZN(n13015) );
  NAND2_X1 U9735 ( .A1(n7494), .A2(n7496), .ZN(n12617) );
  NAND2_X1 U9736 ( .A1(n12941), .A2(n7495), .ZN(n7494) );
  OAI21_X1 U9737 ( .B1(n11346), .B2(n8264), .A(n12674), .ZN(n11445) );
  OAI21_X2 U9738 ( .B1(n13004), .B2(n12725), .A(n12727), .ZN(n12994) );
  NAND2_X1 U9739 ( .A1(n8565), .A2(n7517), .ZN(n7516) );
  NAND2_X1 U9740 ( .A1(n7522), .A2(n7521), .ZN(n8542) );
  AND2_X1 U9741 ( .A1(n8850), .A2(n8851), .ZN(n7532) );
  NAND2_X1 U9742 ( .A1(n8932), .A2(n8933), .ZN(n8935) );
  NAND3_X1 U9743 ( .A1(n8932), .A2(n8933), .A3(n7536), .ZN(n7535) );
  INV_X1 U9744 ( .A(n8754), .ZN(n7543) );
  NOR2_X1 U9745 ( .A1(n10440), .A2(n6740), .ZN(n10367) );
  NOR2_X1 U9746 ( .A1(n10594), .A2(n7696), .ZN(n10598) );
  INV_X1 U9747 ( .A(n11550), .ZN(n7561) );
  INV_X1 U9748 ( .A(n12371), .ZN(n7565) );
  OAI21_X1 U9749 ( .B1(n12396), .B2(n7578), .A(n7577), .ZN(n7576) );
  NAND2_X1 U9750 ( .A1(n10343), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7577) );
  NAND3_X1 U9751 ( .A1(n7582), .A2(n7581), .A3(n12100), .ZN(n9679) );
  OAI22_X1 U9752 ( .A1(n10442), .A2(n7583), .B1(n14672), .B2(n12396), .ZN(
        n10348) );
  XNOR2_X1 U9753 ( .A(n10747), .B(n7583), .ZN(n10742) );
  OAI22_X1 U9754 ( .A1(n14218), .A2(n7583), .B1(n10596), .B2(n14221), .ZN(
        n10412) );
  AND2_X1 U9755 ( .A1(n14042), .A2(n9610), .ZN(n12063) );
  AND4_X2 U9756 ( .A1(n9265), .A2(n9264), .A3(n9411), .A4(n9263), .ZN(n7593)
         );
  NAND2_X1 U9757 ( .A1(n7595), .A2(n6698), .ZN(n9527) );
  NAND2_X1 U9758 ( .A1(n12567), .A2(n7610), .ZN(n7609) );
  OAI211_X1 U9759 ( .C1(n12567), .C2(n7612), .A(n7609), .B(n14439), .ZN(n9240)
         );
  NAND2_X1 U9760 ( .A1(n12567), .A2(n12568), .ZN(n12566) );
  NAND2_X1 U9761 ( .A1(n11195), .A2(n7640), .ZN(n7639) );
  XNOR2_X2 U9762 ( .A(n7650), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U9763 ( .A1(n9808), .A2(n7660), .ZN(n7659) );
  INV_X1 U9764 ( .A(n9807), .ZN(n7662) );
  NAND2_X1 U9765 ( .A1(n9834), .A2(n7663), .ZN(n7664) );
  INV_X1 U9766 ( .A(n9838), .ZN(n7666) );
  OR2_X1 U9767 ( .A1(n9752), .A2(n9753), .ZN(n7671) );
  NAND2_X1 U9768 ( .A1(n9753), .A2(n9752), .ZN(n7673) );
  OAI21_X1 U9769 ( .B1(n9796), .B2(n7690), .A(n7689), .ZN(n7688) );
  OR2_X1 U9770 ( .A1(n13696), .A2(n8381), .ZN(n8382) );
  CLKBUF_X1 U9771 ( .A(n11786), .Z(n11789) );
  OR2_X1 U9772 ( .A1(n8117), .A2(n10669), .ZN(n7844) );
  NOR2_X2 U9773 ( .A1(n14240), .A2(n14330), .ZN(n14225) );
  NAND2_X1 U9774 ( .A1(n12091), .A2(n12189), .ZN(n12097) );
  INV_X1 U9775 ( .A(n12365), .ZN(n7730) );
  OAI21_X1 U9776 ( .B1(n12394), .B2(n10741), .A(n10347), .ZN(n10376) );
  INV_X1 U9777 ( .A(n10075), .ZN(n11976) );
  AOI21_X1 U9778 ( .B1(n14258), .B2(n14626), .A(n9728), .ZN(n9729) );
  INV_X1 U9779 ( .A(n9282), .ZN(n9284) );
  AND2_X1 U9780 ( .A1(n8310), .A2(n10485), .ZN(n9245) );
  NAND2_X1 U9781 ( .A1(n9278), .A2(n9277), .ZN(n9289) );
  INV_X1 U9782 ( .A(n9479), .ZN(n9278) );
  AND2_X1 U9783 ( .A1(P3_U3897), .A2(n12759), .ZN(n15031) );
  NAND2_X1 U9784 ( .A1(n8317), .A2(n8316), .ZN(n10533) );
  XNOR2_X1 U9785 ( .A(n12052), .B(n12326), .ZN(n12055) );
  NAND2_X1 U9786 ( .A1(n9201), .A2(n9202), .ZN(n12532) );
  NAND2_X1 U9787 ( .A1(n9851), .A2(n6644), .ZN(n9856) );
  NAND2_X1 U9788 ( .A1(n8290), .A2(n8284), .ZN(n8294) );
  XNOR2_X1 U9789 ( .A(n8291), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8293) );
  AND2_X1 U9790 ( .A1(n9863), .A2(n9862), .ZN(n7693) );
  NAND2_X2 U9791 ( .A1(n10491), .A2(n15072), .ZN(n15077) );
  INV_X1 U9792 ( .A(n15077), .ZN(n15079) );
  NOR2_X1 U9793 ( .A1(n9173), .A2(n9172), .ZN(n7694) );
  OR2_X1 U9794 ( .A1(n12264), .A2(n9308), .ZN(n7695) );
  AND2_X1 U9795 ( .A1(n10593), .A2(n10592), .ZN(n7696) );
  OR2_X1 U9796 ( .A1(n9260), .A2(n13136), .ZN(n7697) );
  OR2_X1 U9797 ( .A1(n14263), .A2(n14249), .ZN(n7698) );
  NOR2_X1 U9798 ( .A1(n9260), .A2(n13196), .ZN(n8320) );
  INV_X1 U9799 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8080) );
  INV_X1 U9800 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8485) );
  AND2_X1 U9801 ( .A1(n8635), .A2(n8617), .ZN(n7699) );
  INV_X1 U9802 ( .A(n14134), .ZN(n9554) );
  AND2_X2 U9803 ( .A1(n8318), .A2(n9242), .ZN(n15130) );
  INV_X1 U9804 ( .A(n15130), .ZN(n8319) );
  AND2_X1 U9805 ( .A1(n8656), .A2(n8638), .ZN(n7700) );
  INV_X1 U9806 ( .A(n15061), .ZN(n15049) );
  INV_X1 U9807 ( .A(n12958), .ZN(n8200) );
  OR2_X1 U9808 ( .A1(n7836), .A2(n6940), .ZN(n7702) );
  INV_X2 U9809 ( .A(n14226), .ZN(n14642) );
  OR2_X1 U9810 ( .A1(n14442), .A2(n12769), .ZN(n7703) );
  OR2_X1 U9811 ( .A1(n12102), .A2(n12101), .ZN(n7704) );
  INV_X1 U9812 ( .A(n13540), .ZN(n13522) );
  AND2_X1 U9813 ( .A1(n13571), .A2(n10643), .ZN(n13469) );
  INV_X1 U9814 ( .A(n13469), .ZN(n13562) );
  AOI21_X1 U9815 ( .B1(n9747), .B2(n9746), .A(n9744), .ZN(n9745) );
  INV_X1 U9816 ( .A(n12086), .ZN(n12091) );
  NAND2_X1 U9817 ( .A1(n12094), .A2(n12256), .ZN(n12095) );
  OR2_X1 U9818 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  AOI21_X1 U9819 ( .B1(n9796), .B2(n9795), .A(n9793), .ZN(n9794) );
  INV_X1 U9820 ( .A(n14202), .ZN(n12204) );
  OR2_X1 U9821 ( .A1(n12231), .A2(n12230), .ZN(n12232) );
  NAND2_X1 U9822 ( .A1(n9921), .A2(n9749), .ZN(n9922) );
  INV_X1 U9823 ( .A(n7976), .ZN(n7712) );
  INV_X1 U9824 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8330) );
  NOR2_X1 U9825 ( .A1(n9175), .A2(n12770), .ZN(n9176) );
  INV_X1 U9826 ( .A(n12665), .ZN(n7947) );
  AND2_X1 U9827 ( .A1(n10060), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7751) );
  INV_X1 U9828 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8349) );
  INV_X1 U9829 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8327) );
  INV_X1 U9830 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9268) );
  INV_X1 U9831 ( .A(n12780), .ZN(n9144) );
  NOR2_X1 U9832 ( .A1(n7694), .A2(n9176), .ZN(n9177) );
  AND2_X1 U9833 ( .A1(n11007), .A2(n11039), .ZN(n11008) );
  INV_X1 U9834 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15291) );
  INV_X1 U9835 ( .A(n12927), .ZN(n8245) );
  INV_X1 U9836 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8281) );
  INV_X1 U9837 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7711) );
  AND2_X1 U9838 ( .A1(n8572), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8599) );
  INV_X1 U9839 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n15363) );
  INV_X1 U9840 ( .A(n11547), .ZN(n11549) );
  OR2_X1 U9841 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  INV_X1 U9842 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9361) );
  INV_X1 U9843 ( .A(n14174), .ZN(n12321) );
  INV_X1 U9844 ( .A(n12775), .ZN(n9159) );
  NAND2_X1 U9845 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  AND2_X1 U9846 ( .A1(n8142), .A2(n8141), .ZN(n8153) );
  NOR2_X1 U9847 ( .A1(n12588), .A2(n12893), .ZN(n8254) );
  INV_X1 U9848 ( .A(n11777), .ZN(n12698) );
  NAND2_X1 U9849 ( .A1(n12640), .A2(n12647), .ZN(n8256) );
  AND2_X1 U9850 ( .A1(n9129), .A2(n13199), .ZN(n9241) );
  INV_X1 U9851 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7745) );
  INV_X1 U9852 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8621) );
  NOR2_X1 U9853 ( .A1(n8824), .A2(n13235), .ZN(n8840) );
  AOI21_X1 U9854 ( .B1(n9733), .B2(n12069), .A(n9961), .ZN(n9962) );
  NAND2_X1 U9855 ( .A1(n8803), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8824) );
  OR2_X1 U9856 ( .A1(n8737), .A2(n8719), .ZN(n8761) );
  OR2_X1 U9857 ( .A1(n8528), .A2(n8527), .ZN(n8551) );
  AND2_X1 U9858 ( .A1(n14758), .A2(n11488), .ZN(n14759) );
  INV_X1 U9859 ( .A(n13495), .ZN(n12031) );
  NAND2_X1 U9860 ( .A1(n10620), .A2(n10768), .ZN(n10784) );
  OR2_X1 U9861 ( .A1(n12399), .A2(n12398), .ZN(n12400) );
  INV_X1 U9862 ( .A(n14578), .ZN(n11323) );
  INV_X1 U9863 ( .A(n9588), .ZN(n9589) );
  NAND2_X1 U9864 ( .A1(n9569), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9577) );
  AND2_X1 U9865 ( .A1(n14275), .A2(n13749), .ZN(n9708) );
  INV_X1 U9866 ( .A(n12324), .ZN(n14118) );
  OR2_X1 U9867 ( .A1(n9522), .A2(n9521), .ZN(n9533) );
  INV_X1 U9868 ( .A(n12171), .ZN(n12170) );
  NAND2_X1 U9869 ( .A1(n12098), .A2(n9679), .ZN(n10736) );
  OAI22_X1 U9870 ( .A1(n9095), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n9094), .B2(
        n9093), .ZN(n9101) );
  INV_X1 U9871 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12795) );
  NAND2_X1 U9872 ( .A1(n9160), .A2(n9159), .ZN(n9161) );
  INV_X1 U9873 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10959) );
  INV_X1 U9874 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12552) );
  OR2_X1 U9875 ( .A1(n7963), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7999) );
  AND2_X1 U9876 ( .A1(n10542), .A2(n10540), .ZN(n10556) );
  AOI21_X1 U9877 ( .B1(n12927), .B2(n15061), .A(n8254), .ZN(n8255) );
  AND2_X1 U9878 ( .A1(n12687), .A2(n12680), .ZN(n11587) );
  INV_X1 U9879 ( .A(n15071), .ZN(n15045) );
  INV_X1 U9880 ( .A(n12772), .ZN(n11803) );
  AND2_X1 U9881 ( .A1(n8309), .A2(n12619), .ZN(n13063) );
  INV_X1 U9882 ( .A(n8256), .ZN(n12593) );
  NAND2_X1 U9883 ( .A1(n8251), .A2(n12746), .ZN(n15050) );
  AND2_X1 U9884 ( .A1(n7772), .A2(n7771), .ZN(n8054) );
  INV_X1 U9885 ( .A(n8954), .ZN(n8956) );
  NOR2_X1 U9886 ( .A1(n8862), .A2(n8863), .ZN(n8882) );
  OR2_X1 U9887 ( .A1(n8622), .A2(n8621), .ZN(n8644) );
  AND2_X1 U9888 ( .A1(n8448), .A2(n8447), .ZN(n10505) );
  OR2_X1 U9889 ( .A1(n10581), .A2(n9018), .ZN(n9019) );
  AND2_X1 U9890 ( .A1(n8781), .A2(n8780), .ZN(n13548) );
  OR2_X1 U9891 ( .A1(n10401), .A2(n10400), .ZN(n10434) );
  AND2_X1 U9892 ( .A1(n8958), .A2(n8957), .ZN(n13407) );
  INV_X1 U9893 ( .A(n13485), .ZN(n13523) );
  AND2_X1 U9894 ( .A1(n9993), .A2(n8377), .ZN(n10143) );
  INV_X1 U9895 ( .A(n13315), .ZN(n11152) );
  NAND2_X1 U9896 ( .A1(n13562), .A2(n10713), .ZN(n14803) );
  INV_X1 U9897 ( .A(n14872), .ZN(n14847) );
  NOR2_X1 U9898 ( .A1(n10629), .A2(n10628), .ZN(n13520) );
  XNOR2_X1 U9899 ( .A(n8981), .B(n8980), .ZN(n10142) );
  OR2_X1 U9900 ( .A1(n8713), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8639) );
  INV_X1 U9901 ( .A(n14033), .ZN(n13749) );
  OR2_X1 U9902 ( .A1(n9545), .A2(n10051), .ZN(n9293) );
  AND2_X1 U9903 ( .A1(n11825), .A2(n11826), .ZN(n11823) );
  AND2_X1 U9904 ( .A1(n9548), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9558) );
  AND2_X1 U9905 ( .A1(n9541), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9548) );
  NAND2_X1 U9906 ( .A1(n9719), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9310) );
  INV_X1 U9907 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n13863) );
  INV_X1 U9908 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10122) );
  INV_X1 U9909 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10215) );
  INV_X1 U9910 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15351) );
  INV_X1 U9911 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13732) );
  INV_X1 U9912 ( .A(n14371), .ZN(n10237) );
  INV_X1 U9913 ( .A(n13845), .ZN(n14220) );
  NAND2_X1 U9914 ( .A1(n14622), .A2(n14143), .ZN(n10360) );
  INV_X1 U9915 ( .A(n10068), .ZN(n9676) );
  INV_X1 U9916 ( .A(n14611), .ZN(n14234) );
  INV_X1 U9917 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9279) );
  OAI22_X1 U9918 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n15210), .B1(n9102), .B2(
        n9101), .ZN(n9104) );
  NAND2_X1 U9919 ( .A1(n9245), .A2(n9243), .ZN(n9232) );
  INV_X1 U9920 ( .A(n12574), .ZN(n14441) );
  OR2_X1 U9921 ( .A1(n7841), .A2(n12894), .ZN(n12582) );
  AOI21_X1 U9922 ( .B1(n12970), .B2(n8222), .A(n8184), .ZN(n12978) );
  INV_X1 U9923 ( .A(n11053), .ZN(n14951) );
  INV_X1 U9924 ( .A(n14908), .ZN(n15023) );
  AND2_X1 U9925 ( .A1(n12941), .A2(n12940), .ZN(n13089) );
  AND2_X1 U9926 ( .A1(n13016), .A2(n13015), .ZN(n13115) );
  INV_X1 U9927 ( .A(n13063), .ZN(n15067) );
  INV_X1 U9928 ( .A(n11587), .ZN(n12604) );
  NAND2_X1 U9929 ( .A1(n10489), .A2(n15045), .ZN(n15072) );
  NAND2_X1 U9930 ( .A1(n12872), .A2(n10577), .ZN(n15071) );
  AND2_X1 U9931 ( .A1(n9247), .A2(n9246), .ZN(n10488) );
  NOR2_X1 U9932 ( .A1(n15130), .A2(n8321), .ZN(n8322) );
  NOR2_X1 U9933 ( .A1(n15071), .A2(n12761), .ZN(n15129) );
  INV_X1 U9934 ( .A(n15124), .ZN(n15105) );
  INV_X1 U9935 ( .A(SI_11_), .ZN(n15455) );
  AND2_X1 U9936 ( .A1(n10006), .A2(P3_U3151), .ZN(n14386) );
  INV_X1 U9937 ( .A(n11176), .ZN(n9988) );
  INV_X1 U9938 ( .A(n9931), .ZN(n9900) );
  NAND2_X1 U9939 ( .A1(n8576), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8376) );
  INV_X1 U9940 ( .A(n14744), .ZN(n14790) );
  OR2_X1 U9941 ( .A1(n10145), .A2(n10144), .ZN(n10169) );
  INV_X1 U9942 ( .A(n13571), .ZN(n14800) );
  INV_X1 U9943 ( .A(n13524), .ZN(n13538) );
  NAND2_X1 U9944 ( .A1(n8986), .A2(n8985), .ZN(n10642) );
  AND2_X1 U9945 ( .A1(n11185), .A2(n14827), .ZN(n14840) );
  NOR2_X1 U9946 ( .A1(n9735), .A2(n9988), .ZN(n14877) );
  AND2_X1 U9947 ( .A1(n9997), .A2(n10142), .ZN(n9017) );
  OR2_X1 U9948 ( .A1(n8973), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n8974) );
  AND2_X1 U9949 ( .A1(n8595), .A2(n8639), .ZN(n11487) );
  AND2_X1 U9950 ( .A1(n10006), .A2(P2_U3088), .ZN(n11668) );
  INV_X1 U9951 ( .A(n13832), .ZN(n13814) );
  AND2_X1 U9952 ( .A1(n10587), .A2(n10364), .ZN(n13834) );
  AND4_X1 U9953 ( .A1(n9489), .A2(n9488), .A3(n9487), .A4(n9486), .ZN(n14217)
         );
  INV_X1 U9954 ( .A(n14592), .ZN(n13984) );
  INV_X1 U9955 ( .A(n14588), .ZN(n14012) );
  AND2_X1 U9956 ( .A1(n13840), .A2(n14209), .ZN(n12053) );
  INV_X1 U9957 ( .A(n14014), .ZN(n14143) );
  OR2_X1 U9958 ( .A1(n10360), .A2(n10363), .ZN(n14637) );
  INV_X1 U9959 ( .A(n14637), .ZN(n14599) );
  INV_X1 U9960 ( .A(n14196), .ZN(n14626) );
  AND2_X1 U9961 ( .A1(n12346), .A2(n10352), .ZN(n10246) );
  INV_X1 U9962 ( .A(n14097), .ZN(n14288) );
  NAND2_X1 U9963 ( .A1(n12450), .A2(n9678), .ZN(n14404) );
  INV_X1 U9964 ( .A(n14702), .ZN(n14697) );
  INV_X1 U9965 ( .A(n14404), .ZN(n14707) );
  NOR2_X1 U9966 ( .A1(n10234), .A2(n10354), .ZN(n10247) );
  OR2_X1 U9967 ( .A1(n9660), .A2(n11976), .ZN(n10068) );
  AND2_X1 U9968 ( .A1(n9342), .A2(n9341), .ZN(n13917) );
  AND2_X1 U9969 ( .A1(n10542), .A2(n10541), .ZN(n14990) );
  OR2_X1 U9970 ( .A1(n9232), .A2(n12760), .ZN(n14446) );
  AND2_X1 U9971 ( .A1(n9231), .A2(n9230), .ZN(n14433) );
  INV_X1 U9972 ( .A(n14439), .ZN(n14427) );
  AND4_X1 U9973 ( .A1(n12582), .A2(n8250), .A3(n8249), .A4(n8248), .ZN(n12588)
         );
  INV_X1 U9974 ( .A(n13021), .ZN(n12768) );
  INV_X1 U9975 ( .A(n14990), .ZN(n15041) );
  INV_X1 U9976 ( .A(n15031), .ZN(n15010) );
  INV_X1 U9977 ( .A(n14474), .ZN(n15036) );
  AND2_X1 U9978 ( .A1(n13038), .A2(n13037), .ZN(n13120) );
  INV_X1 U9979 ( .A(n15077), .ZN(n13011) );
  NAND2_X1 U9980 ( .A1(n15077), .A2(n10856), .ZN(n13029) );
  INV_X1 U9981 ( .A(n15144), .ZN(n15141) );
  INV_X1 U9982 ( .A(n12920), .ZN(n13153) );
  AND3_X1 U9983 ( .A1(n15112), .A2(n15111), .A3(n15110), .ZN(n15137) );
  NAND2_X1 U9984 ( .A1(n8295), .A2(n10066), .ZN(n12085) );
  INV_X1 U9985 ( .A(SI_13_), .ZN(n10139) );
  AND2_X1 U9986 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  INV_X1 U9987 ( .A(n13302), .ZN(n11948) );
  INV_X1 U9988 ( .A(n13278), .ZN(n13304) );
  NAND2_X1 U9989 ( .A1(n10169), .A2(n10146), .ZN(n14795) );
  INV_X1 U9990 ( .A(n14797), .ZN(n13494) );
  INV_X1 U9991 ( .A(n13562), .ZN(n14809) );
  INV_X1 U9992 ( .A(n14806), .ZN(n13576) );
  OR2_X1 U9993 ( .A1(n10637), .A2(n10642), .ZN(n14888) );
  AND4_X1 U9994 ( .A1(n14854), .A2(n14853), .A3(n14852), .A4(n14851), .ZN(
        n14885) );
  OR2_X1 U9995 ( .A1(n10637), .A2(n10606), .ZN(n14878) );
  INV_X1 U9996 ( .A(n14818), .ZN(n14815) );
  NOR2_X1 U9997 ( .A1(n14810), .A2(n14815), .ZN(n14814) );
  INV_X1 U9998 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n15238) );
  INV_X1 U9999 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10389) );
  INV_X1 U10000 ( .A(n14513), .ZN(n14525) );
  AND2_X1 U10001 ( .A1(n10589), .A2(n12349), .ZN(n13832) );
  INV_X1 U10002 ( .A(n14128), .ZN(n14298) );
  INV_X1 U10003 ( .A(n12291), .ZN(n14021) );
  OAI21_X1 U10004 ( .B1(n14145), .B2(n9598), .A(n9553), .ZN(n14152) );
  INV_X1 U10005 ( .A(n12166), .ZN(n13848) );
  INV_X1 U10006 ( .A(n12114), .ZN(n13857) );
  OR2_X1 U10007 ( .A1(n14570), .A2(n10094), .ZN(n14588) );
  INV_X1 U10008 ( .A(n14568), .ZN(n14596) );
  OR2_X1 U10009 ( .A1(n14642), .A2(n14630), .ZN(n14616) );
  NAND2_X1 U10010 ( .A1(n9715), .A2(n14637), .ZN(n14226) );
  OR2_X1 U10011 ( .A1(n14642), .A2(n14404), .ZN(n14249) );
  INV_X1 U10012 ( .A(n14720), .ZN(n14718) );
  AND3_X2 U10013 ( .A1(n10247), .A2(n10353), .A3(n10246), .ZN(n14720) );
  AND3_X1 U10014 ( .A1(n14408), .A2(n14407), .A3(n14406), .ZN(n14410) );
  INV_X1 U10015 ( .A(n14710), .ZN(n14708) );
  AND2_X2 U10016 ( .A1(n10357), .A2(n10068), .ZN(n14669) );
  INV_X1 U10017 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11667) );
  INV_X1 U10018 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10572) );
  INV_X1 U10019 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10202) );
  INV_X1 U10020 ( .A(n10942), .ZN(P3_U3897) );
  AND2_X1 U10021 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10145), .ZN(P2_U3947) );
  AND2_X1 U10022 ( .A1(n10343), .A2(n10072), .ZN(P1_U4016) );
  NAND2_X1 U10023 ( .A1(n7698), .A2(n9731), .ZN(P1_U3356) );
  NOR2_X1 U10024 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n7708) );
  NAND4_X1 U10025 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n8108)
         );
  NAND3_X1 U10026 ( .A1(n7995), .A2(n15406), .A3(n7709), .ZN(n7710) );
  NOR2_X1 U10027 ( .A1(n7712), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U10028 ( .A1(n7833), .A2(n7279), .ZN(n7850) );
  NOR2_X1 U10029 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), 
        .ZN(n7718) );
  NOR2_X1 U10030 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n7717) );
  INV_X1 U10031 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7720) );
  MUX2_X1 U10032 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7722), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7723) );
  INV_X1 U10033 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U10034 ( .A1(n7885), .A2(n10564), .ZN(n7904) );
  NAND2_X1 U10035 ( .A1(n15291), .A2(n11733), .ZN(n7724) );
  NAND2_X1 U10036 ( .A1(n8025), .A2(n12795), .ZN(n8045) );
  INV_X1 U10037 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10038 ( .A1(n7725), .A2(n8218), .ZN(n8221) );
  INV_X1 U10039 ( .A(n8221), .ZN(n7727) );
  INV_X1 U10040 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10041 ( .A1(n7727), .A2(n7726), .ZN(n12894) );
  NAND2_X1 U10042 ( .A1(n8221), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7728) );
  NAND2_X1 U10043 ( .A1(n12894), .A2(n7728), .ZN(n12921) );
  NAND2_X1 U10044 ( .A1(n8222), .A2(n12921), .ZN(n7735) );
  NAND2_X1 U10045 ( .A1(n7842), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7734) );
  NAND2_X1 U10046 ( .A1(n12365), .A2(n13207), .ZN(n7856) );
  INV_X1 U10047 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13152) );
  OR2_X1 U10048 ( .A1(n8247), .A2(n13152), .ZN(n7733) );
  NAND2_X2 U10049 ( .A1(n7730), .A2(n13207), .ZN(n8117) );
  INV_X1 U10050 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n7731) );
  OR2_X1 U10051 ( .A1(n6561), .A2(n7731), .ZN(n7732) );
  NAND4_X1 U10052 ( .A1(n7735), .A2(n7734), .A3(n7733), .A4(n7732), .ZN(n12927) );
  XNOR2_X1 U10053 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7831) );
  INV_X1 U10054 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U10055 ( .A1(n8390), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7830) );
  INV_X1 U10056 ( .A(n7830), .ZN(n7736) );
  NAND2_X1 U10057 ( .A1(n7831), .A2(n7736), .ZN(n7738) );
  INV_X1 U10058 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10005) );
  NAND2_X1 U10059 ( .A1(n10005), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10060 ( .A1(n7738), .A2(n7737), .ZN(n7849) );
  NAND2_X1 U10061 ( .A1(n10053), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U10062 ( .A1(n7849), .A2(n7739), .ZN(n7741) );
  NAND2_X1 U10063 ( .A1(n10034), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10064 ( .A1(n7741), .A2(n7740), .ZN(n7862) );
  NAND2_X1 U10065 ( .A1(n10028), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7743) );
  INV_X1 U10066 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10067 ( .A1(n7894), .A2(n7893), .ZN(n7747) );
  NAND2_X1 U10068 ( .A1(n7745), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U10069 ( .A1(n10039), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U10070 ( .A1(n10047), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7748) );
  INV_X1 U10071 ( .A(n7911), .ZN(n7749) );
  NAND2_X1 U10072 ( .A1(n10058), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7752) );
  NAND2_X1 U10073 ( .A1(n10063), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7753) );
  XNOR2_X1 U10074 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7970) );
  NAND2_X1 U10075 ( .A1(n7971), .A2(n7970), .ZN(n7755) );
  NAND2_X1 U10076 ( .A1(n10078), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U10077 ( .A1(n10138), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U10078 ( .A1(n10202), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10079 ( .A1(n10204), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U10080 ( .A1(n7759), .A2(n7758), .ZN(n7993) );
  NAND2_X1 U10081 ( .A1(n15357), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U10082 ( .A1(n15428), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U10083 ( .A1(n7767), .A2(n7765), .ZN(n8020) );
  INV_X1 U10084 ( .A(n8020), .ZN(n7766) );
  NAND2_X1 U10085 ( .A1(n8021), .A2(n7766), .ZN(n7768) );
  NAND2_X1 U10086 ( .A1(n7768), .A2(n7767), .ZN(n8035) );
  NAND2_X1 U10087 ( .A1(n10385), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7770) );
  INV_X1 U10088 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10387) );
  NAND2_X1 U10089 ( .A1(n10387), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U10090 ( .A1(n15293), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10091 ( .A1(n10333), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U10092 ( .A1(n10390), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U10093 ( .A1(n10389), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U10094 ( .A1(n7775), .A2(n7773), .ZN(n8075) );
  INV_X1 U10095 ( .A(n8075), .ZN(n7774) );
  NAND2_X1 U10096 ( .A1(n10572), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7777) );
  NAND2_X1 U10097 ( .A1(n10573), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7776) );
  INV_X1 U10098 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U10099 ( .A1(n10853), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7779) );
  INV_X1 U10100 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U10101 ( .A1(n10855), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7778) );
  INV_X1 U10102 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U10103 ( .A1(n11174), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7781) );
  INV_X1 U10104 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U10105 ( .A1(n11177), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7780) );
  INV_X1 U10106 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n15421) );
  NAND2_X1 U10107 ( .A1(n15421), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7783) );
  INV_X1 U10108 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U10109 ( .A1(n11361), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7782) );
  AND2_X1 U10110 ( .A1(n7783), .A2(n7782), .ZN(n8135) );
  INV_X1 U10111 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U10112 ( .A1(n7784), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7786) );
  INV_X1 U10113 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12072) );
  NAND2_X1 U10114 ( .A1(n12072), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7785) );
  AND2_X1 U10115 ( .A1(n7786), .A2(n7785), .ZN(n8147) );
  XNOR2_X1 U10116 ( .A(n15238), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U10117 ( .A1(n15238), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10118 ( .A1(n7788), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7789) );
  INV_X1 U10119 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11740) );
  INV_X1 U10120 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U10121 ( .A1(n8896), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7792) );
  INV_X1 U10122 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U10123 ( .A1(n15247), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7791) );
  AND2_X1 U10124 ( .A1(n7792), .A2(n7791), .ZN(n8187) );
  INV_X1 U10125 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11974) );
  NAND2_X1 U10126 ( .A1(n11974), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7795) );
  INV_X1 U10127 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11972) );
  NAND2_X1 U10128 ( .A1(n11972), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U10129 ( .A1(n7795), .A2(n7793), .ZN(n8202) );
  INV_X1 U10130 ( .A(n8202), .ZN(n7794) );
  INV_X1 U10131 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14367) );
  NAND2_X1 U10132 ( .A1(n14367), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7798) );
  INV_X1 U10133 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12051) );
  NAND2_X1 U10134 ( .A1(n12051), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U10135 ( .A1(n7798), .A2(n7796), .ZN(n8212) );
  INV_X1 U10136 ( .A(n8212), .ZN(n7797) );
  NAND2_X1 U10137 ( .A1(n8213), .A2(n7797), .ZN(n7799) );
  NAND2_X1 U10138 ( .A1(n7799), .A2(n7798), .ZN(n7803) );
  INV_X1 U10139 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15279) );
  NAND2_X1 U10140 ( .A1(n15279), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8230) );
  INV_X1 U10141 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10142 ( .A1(n7800), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7801) );
  AND2_X1 U10143 ( .A1(n8230), .A2(n7801), .ZN(n7802) );
  NAND2_X1 U10144 ( .A1(n7803), .A2(n7802), .ZN(n8231) );
  OR2_X1 U10145 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  NAND2_X1 U10146 ( .A1(n8231), .A2(n7804), .ZN(n12364) );
  NAND2_X1 U10147 ( .A1(n8215), .A2(SI_28_), .ZN(n7816) );
  INV_X1 U10148 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n7818) );
  OR2_X1 U10149 ( .A1(n7841), .A2(n7818), .ZN(n7822) );
  INV_X1 U10150 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10552) );
  OR2_X1 U10151 ( .A1(n8117), .A2(n10552), .ZN(n7821) );
  INV_X1 U10152 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n7819) );
  OR2_X1 U10153 ( .A1(n7856), .A2(n7819), .ZN(n7820) );
  INV_X1 U10154 ( .A(SI_0_), .ZN(n10019) );
  INV_X1 U10155 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U10156 ( .A1(n9302), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10157 ( .A1(n7830), .A2(n7823), .ZN(n10018) );
  NAND2_X1 U10158 ( .A1(n8214), .A2(n10018), .ZN(n7824) );
  NAND2_X1 U10159 ( .A1(n7842), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7829) );
  INV_X1 U10160 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10544) );
  OR2_X1 U10161 ( .A1(n6561), .A2(n10544), .ZN(n7828) );
  INV_X1 U10162 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15073) );
  OR2_X1 U10163 ( .A1(n7841), .A2(n15073), .ZN(n7827) );
  INV_X1 U10164 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7825) );
  OR2_X1 U10165 ( .A1(n7856), .A2(n7825), .ZN(n7826) );
  XNOR2_X1 U10166 ( .A(n7831), .B(n7830), .ZN(n10007) );
  NAND2_X1 U10167 ( .A1(n8215), .A2(SI_1_), .ZN(n7837) );
  NAND2_X1 U10168 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n7832) );
  INV_X1 U10169 ( .A(n7833), .ZN(n7834) );
  OAI211_X1 U10170 ( .C1(n7847), .C2(n10007), .A(n7837), .B(n7702), .ZN(n9133)
         );
  NAND2_X1 U10171 ( .A1(n12782), .A2(n15059), .ZN(n12638) );
  NAND2_X1 U10172 ( .A1(n7838), .A2(n9133), .ZN(n12634) );
  NAND2_X1 U10173 ( .A1(n12638), .A2(n12634), .ZN(n15066) );
  NAND2_X1 U10174 ( .A1(n15065), .A2(n15066), .ZN(n7840) );
  NAND2_X1 U10175 ( .A1(n7838), .A2(n15059), .ZN(n7839) );
  NAND2_X1 U10176 ( .A1(n7840), .A2(n7839), .ZN(n15048) );
  INV_X1 U10177 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15046) );
  OR2_X1 U10178 ( .A1(n7841), .A2(n15046), .ZN(n7846) );
  NAND2_X1 U10179 ( .A1(n7842), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7845) );
  INV_X1 U10180 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10669) );
  INV_X1 U10181 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7843) );
  INV_X2 U10182 ( .A(n7847), .ZN(n8214) );
  XNOR2_X1 U10183 ( .A(n10034), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n7848) );
  XNOR2_X1 U10184 ( .A(n7849), .B(n7848), .ZN(n10017) );
  NAND2_X1 U10185 ( .A1(n8214), .A2(n10017), .ZN(n7852) );
  NAND2_X1 U10186 ( .A1(n8113), .A2(n6564), .ZN(n7851) );
  INV_X1 U10187 ( .A(n15043), .ZN(n10337) );
  NAND2_X1 U10188 ( .A1(n12355), .A2(n10337), .ZN(n12626) );
  NAND2_X1 U10189 ( .A1(n15063), .A2(n15043), .ZN(n12635) );
  NAND2_X1 U10190 ( .A1(n15048), .A2(n15047), .ZN(n7854) );
  NAND2_X1 U10191 ( .A1(n12355), .A2(n15043), .ZN(n7853) );
  NAND2_X1 U10192 ( .A1(n7854), .A2(n7853), .ZN(n10868) );
  INV_X1 U10193 ( .A(n10868), .ZN(n7867) );
  OR2_X1 U10194 ( .A1(n7841), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n7860) );
  INV_X2 U10195 ( .A(n12584), .ZN(n8246) );
  NAND2_X1 U10196 ( .A1(n8246), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7859) );
  INV_X1 U10197 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11037) );
  OR2_X1 U10198 ( .A1(n8117), .A2(n11037), .ZN(n7858) );
  INV_X1 U10199 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7855) );
  OR2_X1 U10200 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  NAND4_X1 U10201 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n12781) );
  INV_X1 U10202 ( .A(n12781), .ZN(n15051) );
  XNOR2_X1 U10203 ( .A(n10033), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n7861) );
  XNOR2_X1 U10204 ( .A(n7862), .B(n7861), .ZN(n10015) );
  NAND2_X1 U10205 ( .A1(n8214), .A2(n10015), .ZN(n7866) );
  NAND2_X1 U10206 ( .A1(n7850), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7863) );
  MUX2_X1 U10207 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7863), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n7864) );
  NAND2_X1 U10208 ( .A1(n7864), .A2(n7877), .ZN(n11039) );
  NAND2_X1 U10209 ( .A1(n8113), .A2(n11039), .ZN(n7865) );
  INV_X1 U10210 ( .A(n15089), .ZN(n10874) );
  NAND2_X1 U10211 ( .A1(n15051), .A2(n10874), .ZN(n12640) );
  NAND2_X1 U10212 ( .A1(n12781), .A2(n15089), .ZN(n12647) );
  NAND2_X1 U10213 ( .A1(n12781), .A2(n10874), .ZN(n7868) );
  AND2_X1 U10214 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7869) );
  NOR2_X1 U10215 ( .A1(n7885), .A2(n7869), .ZN(n10863) );
  OR2_X1 U10216 ( .A1(n7841), .A2(n10863), .ZN(n7874) );
  NAND2_X1 U10217 ( .A1(n8246), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7873) );
  INV_X1 U10218 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n7870) );
  OR2_X1 U10219 ( .A1(n8247), .A2(n7870), .ZN(n7872) );
  INV_X1 U10220 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11044) );
  OR2_X1 U10221 ( .A1(n8117), .A2(n11044), .ZN(n7871) );
  NAND4_X1 U10222 ( .A1(n7874), .A2(n7873), .A3(n7872), .A4(n7871), .ZN(n12780) );
  XNOR2_X1 U10223 ( .A(n7876), .B(n7875), .ZN(n10010) );
  NAND2_X1 U10224 ( .A1(n8214), .A2(n10010), .ZN(n7883) );
  INV_X1 U10225 ( .A(n7897), .ZN(n7881) );
  NAND2_X1 U10226 ( .A1(n7877), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7879) );
  MUX2_X1 U10227 ( .A(n7879), .B(P3_IR_REG_31__SCAN_IN), .S(n7878), .Z(n7880)
         );
  NAND2_X1 U10228 ( .A1(n7881), .A2(n7880), .ZN(n11046) );
  NAND2_X1 U10229 ( .A1(n8113), .A2(n11046), .ZN(n7882) );
  OAI211_X1 U10230 ( .C1(n12585), .C2(SI_4_), .A(n7883), .B(n7882), .ZN(n9142)
         );
  INV_X1 U10231 ( .A(n9142), .ZN(n15096) );
  NAND2_X1 U10232 ( .A1(n9144), .A2(n15096), .ZN(n12648) );
  NAND2_X1 U10233 ( .A1(n12780), .A2(n9142), .ZN(n12651) );
  NAND2_X1 U10234 ( .A1(n12648), .A2(n12651), .ZN(n10859) );
  NAND2_X1 U10235 ( .A1(n12780), .A2(n15096), .ZN(n7884) );
  OR2_X1 U10236 ( .A1(n7885), .A2(n10564), .ZN(n7886) );
  NAND2_X1 U10237 ( .A1(n7904), .A2(n7886), .ZN(n10697) );
  NAND2_X1 U10238 ( .A1(n8222), .A2(n10697), .ZN(n7892) );
  NAND2_X1 U10239 ( .A1(n8246), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7891) );
  INV_X1 U10240 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n7888) );
  OR2_X1 U10241 ( .A1(n8247), .A2(n7888), .ZN(n7890) );
  INV_X1 U10242 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11051) );
  OR2_X1 U10243 ( .A1(n8117), .A2(n11051), .ZN(n7889) );
  NAND4_X1 U10244 ( .A1(n7892), .A2(n7891), .A3(n7890), .A4(n7889), .ZN(n12779) );
  INV_X1 U10245 ( .A(n12779), .ZN(n9148) );
  XNOR2_X1 U10246 ( .A(n7894), .B(n7893), .ZN(n10012) );
  NAND2_X1 U10247 ( .A1(n8214), .A2(n10012), .ZN(n7901) );
  NOR2_X1 U10248 ( .A1(n7897), .A2(n8285), .ZN(n7895) );
  MUX2_X1 U10249 ( .A(n8285), .B(n7895), .S(P3_IR_REG_5__SCAN_IN), .Z(n7899)
         );
  NAND2_X1 U10250 ( .A1(n7897), .A2(n7896), .ZN(n7927) );
  INV_X1 U10251 ( .A(n7927), .ZN(n7898) );
  NAND2_X1 U10252 ( .A1(n8113), .A2(n11053), .ZN(n7900) );
  OAI211_X1 U10253 ( .C1(n12585), .C2(SI_5_), .A(n7901), .B(n7900), .ZN(n15097) );
  INV_X1 U10254 ( .A(n15097), .ZN(n10698) );
  NAND2_X1 U10255 ( .A1(n9148), .A2(n10698), .ZN(n12654) );
  NAND2_X1 U10256 ( .A1(n12779), .A2(n15097), .ZN(n12649) );
  NAND2_X1 U10257 ( .A1(n9148), .A2(n15097), .ZN(n7903) );
  NAND2_X1 U10258 ( .A1(n7904), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U10259 ( .A1(n7918), .A2(n7905), .ZN(n10996) );
  NAND2_X1 U10260 ( .A1(n8222), .A2(n10996), .ZN(n7910) );
  NAND2_X1 U10261 ( .A1(n8246), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7909) );
  INV_X1 U10262 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n7906) );
  OR2_X1 U10263 ( .A1(n8247), .A2(n7906), .ZN(n7908) );
  INV_X1 U10264 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11058) );
  OR2_X1 U10265 ( .A1(n8117), .A2(n11058), .ZN(n7907) );
  NAND4_X1 U10266 ( .A1(n7910), .A2(n7909), .A3(n7908), .A4(n7907), .ZN(n12778) );
  INV_X1 U10267 ( .A(n12778), .ZN(n7916) );
  XNOR2_X1 U10268 ( .A(n7912), .B(n7911), .ZN(n10014) );
  NAND2_X1 U10269 ( .A1(n8215), .A2(SI_6_), .ZN(n7915) );
  NAND2_X1 U10270 ( .A1(n7927), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7913) );
  XNOR2_X1 U10271 ( .A(n7913), .B(P3_IR_REG_6__SCAN_IN), .ZN(n14972) );
  NAND2_X1 U10272 ( .A1(n8113), .A2(n14972), .ZN(n7914) );
  OAI211_X1 U10273 ( .C1(n8191), .C2(n10014), .A(n7915), .B(n7914), .ZN(n15104) );
  NAND2_X1 U10274 ( .A1(n7916), .A2(n15104), .ZN(n12660) );
  INV_X1 U10275 ( .A(n15104), .ZN(n10991) );
  NAND2_X1 U10276 ( .A1(n12778), .A2(n10991), .ZN(n12656) );
  NAND2_X1 U10277 ( .A1(n12660), .A2(n12656), .ZN(n10896) );
  NAND2_X1 U10278 ( .A1(n10897), .A2(n10896), .ZN(n10895) );
  NAND2_X1 U10279 ( .A1(n12778), .A2(n15104), .ZN(n7917) );
  AND2_X1 U10280 ( .A1(n7918), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7919) );
  NOR2_X1 U10281 ( .A1(n7934), .A2(n7919), .ZN(n11118) );
  OR2_X1 U10282 ( .A1(n7841), .A2(n11118), .ZN(n7924) );
  NAND2_X1 U10283 ( .A1(n8246), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7923) );
  INV_X1 U10284 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n7920) );
  OR2_X1 U10285 ( .A1(n8247), .A2(n7920), .ZN(n7922) );
  INV_X1 U10286 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11117) );
  OR2_X1 U10287 ( .A1(n8117), .A2(n11117), .ZN(n7921) );
  NAND4_X1 U10288 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), .ZN(n12777) );
  XNOR2_X1 U10289 ( .A(n7926), .B(n7925), .ZN(n10022) );
  NAND2_X1 U10290 ( .A1(n8214), .A2(n10022), .ZN(n7932) );
  INV_X1 U10291 ( .A(SI_7_), .ZN(n10021) );
  NAND2_X1 U10292 ( .A1(n8215), .A2(n10021), .ZN(n7931) );
  OAI21_X1 U10293 ( .B1(n7927), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7929) );
  INV_X1 U10294 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7928) );
  XNOR2_X1 U10295 ( .A(n7929), .B(n7928), .ZN(n14986) );
  NAND2_X1 U10296 ( .A1(n8113), .A2(n14986), .ZN(n7930) );
  XNOR2_X1 U10297 ( .A(n12777), .B(n12661), .ZN(n12659) );
  NAND2_X1 U10298 ( .A1(n12777), .A2(n12661), .ZN(n7933) );
  NOR2_X1 U10299 ( .A1(n7934), .A2(n10959), .ZN(n7935) );
  OR2_X1 U10300 ( .A1(n7948), .A2(n7935), .ZN(n10953) );
  NAND2_X1 U10301 ( .A1(n8222), .A2(n10953), .ZN(n7940) );
  NAND2_X1 U10302 ( .A1(n8246), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7939) );
  INV_X1 U10303 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n7936) );
  OR2_X1 U10304 ( .A1(n8247), .A2(n7936), .ZN(n7938) );
  INV_X1 U10305 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11070) );
  OR2_X1 U10306 ( .A1(n8117), .A2(n11070), .ZN(n7937) );
  NAND4_X1 U10307 ( .A1(n7940), .A2(n7939), .A3(n7938), .A4(n7937), .ZN(n12776) );
  INV_X1 U10308 ( .A(n12776), .ZN(n11197) );
  XNOR2_X1 U10309 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7941) );
  XNOR2_X1 U10310 ( .A(n7942), .B(n7941), .ZN(n10024) );
  NAND2_X1 U10311 ( .A1(n8215), .A2(SI_8_), .ZN(n7946) );
  NAND2_X1 U10312 ( .A1(n7943), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7944) );
  XNOR2_X1 U10313 ( .A(n7944), .B(P3_IR_REG_8__SCAN_IN), .ZN(n15002) );
  NAND2_X1 U10314 ( .A1(n8113), .A2(n15002), .ZN(n7945) );
  OAI211_X1 U10315 ( .C1(n8191), .C2(n10024), .A(n7946), .B(n7945), .ZN(n10961) );
  NAND2_X1 U10316 ( .A1(n11197), .A2(n10961), .ZN(n12666) );
  INV_X1 U10317 ( .A(n10961), .ZN(n15113) );
  NAND2_X1 U10318 ( .A1(n12776), .A2(n15113), .ZN(n12667) );
  OR2_X1 U10319 ( .A1(n7948), .A2(n15369), .ZN(n7949) );
  NAND2_X1 U10320 ( .A1(n7963), .A2(n7949), .ZN(n11287) );
  NAND2_X1 U10321 ( .A1(n8222), .A2(n11287), .ZN(n7954) );
  NAND2_X1 U10322 ( .A1(n7842), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7953) );
  INV_X1 U10323 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11077) );
  OR2_X1 U10324 ( .A1(n8117), .A2(n11077), .ZN(n7952) );
  INV_X1 U10325 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n7950) );
  OR2_X1 U10326 ( .A1(n8247), .A2(n7950), .ZN(n7951) );
  NAND4_X1 U10327 ( .A1(n7954), .A2(n7953), .A3(n7952), .A4(n7951), .ZN(n12775) );
  XNOR2_X1 U10328 ( .A(n10065), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n7955) );
  XNOR2_X1 U10329 ( .A(n7956), .B(n7955), .ZN(n14381) );
  NAND2_X1 U10330 ( .A1(n8214), .A2(n14381), .ZN(n7960) );
  OR2_X1 U10331 ( .A1(n7957), .A2(n8285), .ZN(n7958) );
  XNOR2_X1 U10332 ( .A(n7958), .B(n7972), .ZN(n14384) );
  NAND2_X1 U10333 ( .A1(n8113), .A2(n14384), .ZN(n7959) );
  OAI211_X1 U10334 ( .C1(n12585), .C2(SI_9_), .A(n7960), .B(n7959), .ZN(n15120) );
  XNOR2_X1 U10335 ( .A(n12775), .B(n15120), .ZN(n12598) );
  NAND2_X1 U10336 ( .A1(n11197), .A2(n15113), .ZN(n11280) );
  AND2_X1 U10337 ( .A1(n12598), .A2(n11280), .ZN(n7961) );
  INV_X1 U10338 ( .A(n15120), .ZN(n11288) );
  NAND2_X1 U10339 ( .A1(n12775), .A2(n11288), .ZN(n7962) );
  NAND2_X1 U10340 ( .A1(n7963), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10341 ( .A1(n7999), .A2(n7964), .ZN(n11531) );
  NAND2_X1 U10342 ( .A1(n8222), .A2(n11531), .ZN(n7969) );
  NAND2_X1 U10343 ( .A1(n8246), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7968) );
  INV_X1 U10344 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n7965) );
  OR2_X1 U10345 ( .A1(n8247), .A2(n7965), .ZN(n7967) );
  INV_X1 U10346 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11082) );
  OR2_X1 U10347 ( .A1(n8117), .A2(n11082), .ZN(n7966) );
  NAND4_X1 U10348 ( .A1(n7969), .A2(n7968), .A3(n7967), .A4(n7966), .ZN(n12774) );
  INV_X1 U10349 ( .A(n12774), .ZN(n11448) );
  XNOR2_X1 U10350 ( .A(n7971), .B(n7970), .ZN(n10037) );
  NAND2_X1 U10351 ( .A1(n10037), .A2(n8214), .ZN(n7980) );
  INV_X1 U10352 ( .A(SI_10_), .ZN(n15294) );
  AND2_X1 U10353 ( .A1(n7957), .A2(n7972), .ZN(n7973) );
  NOR2_X1 U10354 ( .A1(n7973), .A2(n8285), .ZN(n7974) );
  MUX2_X1 U10355 ( .A(n8285), .B(n7974), .S(P3_IR_REG_10__SCAN_IN), .Z(n7975)
         );
  INV_X1 U10356 ( .A(n7975), .ZN(n7978) );
  INV_X1 U10357 ( .A(n8111), .ZN(n7977) );
  AOI22_X1 U10358 ( .A1(n8215), .A2(n15294), .B1(n8113), .B2(n11462), .ZN(
        n7979) );
  NAND2_X1 U10359 ( .A1(n11448), .A2(n11353), .ZN(n12674) );
  INV_X1 U10360 ( .A(n11353), .ZN(n15125) );
  NAND2_X1 U10361 ( .A1(n15125), .A2(n12774), .ZN(n12675) );
  NAND2_X1 U10362 ( .A1(n12674), .A2(n12675), .ZN(n11348) );
  XNOR2_X1 U10363 ( .A(n7999), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n11636) );
  NAND2_X1 U10364 ( .A1(n8222), .A2(n11636), .ZN(n7986) );
  NAND2_X1 U10365 ( .A1(n8246), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7985) );
  INV_X1 U10366 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n7981) );
  OR2_X1 U10367 ( .A1(n8247), .A2(n7981), .ZN(n7984) );
  INV_X1 U10368 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7982) );
  OR2_X1 U10369 ( .A1(n6561), .A2(n7982), .ZN(n7983) );
  NAND4_X1 U10370 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n12773) );
  XNOR2_X1 U10371 ( .A(n10138), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n7987) );
  XNOR2_X1 U10372 ( .A(n7988), .B(n7987), .ZN(n15453) );
  NAND2_X1 U10373 ( .A1(n15453), .A2(n8214), .ZN(n7991) );
  OR2_X1 U10374 ( .A1(n8111), .A2(n8285), .ZN(n7989) );
  XNOR2_X1 U10375 ( .A(n7989), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U10376 ( .A1(n8215), .A2(SI_11_), .B1(n8113), .B2(n11652), .ZN(
        n7990) );
  NAND2_X1 U10377 ( .A1(n7991), .A2(n7990), .ZN(n11451) );
  XNOR2_X1 U10378 ( .A(n11631), .B(n11451), .ZN(n12676) );
  NAND2_X1 U10379 ( .A1(n11451), .A2(n12773), .ZN(n7992) );
  XNOR2_X1 U10380 ( .A(n7994), .B(n7993), .ZN(n14385) );
  NAND2_X1 U10381 ( .A1(n14385), .A2(n8214), .ZN(n7998) );
  NAND2_X1 U10382 ( .A1(n8111), .A2(n15406), .ZN(n8009) );
  NAND2_X1 U10383 ( .A1(n8009), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7996) );
  XNOR2_X1 U10384 ( .A(n7996), .B(n7995), .ZN(n14390) );
  AOI22_X1 U10385 ( .A1(n8215), .A2(n8614), .B1(n8113), .B2(n14390), .ZN(n7997) );
  NAND2_X1 U10386 ( .A1(n7998), .A2(n7997), .ZN(n14492) );
  OAI21_X1 U10387 ( .B1(n7999), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10388 ( .A1(n8000), .A2(n8012), .ZN(n11591) );
  NAND2_X1 U10389 ( .A1(n8222), .A2(n11591), .ZN(n8005) );
  NAND2_X1 U10390 ( .A1(n8246), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8004) );
  INV_X1 U10391 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8001) );
  OR2_X1 U10392 ( .A1(n8247), .A2(n8001), .ZN(n8003) );
  INV_X1 U10393 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11592) );
  OR2_X1 U10394 ( .A1(n6561), .A2(n11592), .ZN(n8002) );
  NAND4_X1 U10395 ( .A1(n8005), .A2(n8004), .A3(n8003), .A4(n8002), .ZN(n12772) );
  NAND2_X1 U10396 ( .A1(n14492), .A2(n11803), .ZN(n8006) );
  OR2_X1 U10397 ( .A1(n14492), .A2(n11803), .ZN(n8007) );
  XNOR2_X1 U10398 ( .A(n8008), .B(n10245), .ZN(n10140) );
  NAND2_X1 U10399 ( .A1(n6571), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8010) );
  XNOR2_X1 U10400 ( .A(n8010), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12801) );
  AND2_X1 U10401 ( .A1(n8012), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8013) );
  NOR2_X1 U10402 ( .A1(n8025), .A2(n8013), .ZN(n11804) );
  OR2_X1 U10403 ( .A1(n7841), .A2(n11804), .ZN(n8018) );
  NAND2_X1 U10404 ( .A1(n8246), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8017) );
  INV_X1 U10405 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11805) );
  OR2_X1 U10406 ( .A1(n6561), .A2(n11805), .ZN(n8016) );
  INV_X1 U10407 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n8014) );
  OR2_X1 U10408 ( .A1(n8247), .A2(n8014), .ZN(n8015) );
  NAND4_X1 U10409 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n12771) );
  INV_X1 U10410 ( .A(n12771), .ZN(n14419) );
  OR2_X1 U10411 ( .A1(n14490), .A2(n14419), .ZN(n12691) );
  NAND2_X1 U10412 ( .A1(n14490), .A2(n14419), .ZN(n12688) );
  XNOR2_X1 U10413 ( .A(n8021), .B(n8020), .ZN(n10231) );
  NAND2_X1 U10414 ( .A1(n10231), .A2(n8214), .ZN(n8024) );
  NOR2_X1 U10415 ( .A1(n6571), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8039) );
  OR2_X1 U10416 ( .A1(n8039), .A2(n8285), .ZN(n8022) );
  XNOR2_X1 U10417 ( .A(n8022), .B(n8038), .ZN(n12787) );
  INV_X1 U10418 ( .A(n12787), .ZN(n12799) );
  AOI22_X1 U10419 ( .A1(n8215), .A2(SI_14_), .B1(n8113), .B2(n12799), .ZN(
        n8023) );
  OR2_X1 U10420 ( .A1(n8025), .A2(n12795), .ZN(n8026) );
  AND2_X1 U10421 ( .A1(n8026), .A2(n8045), .ZN(n14434) );
  OR2_X1 U10422 ( .A1(n7841), .A2(n14434), .ZN(n8031) );
  NAND2_X1 U10423 ( .A1(n8246), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8030) );
  INV_X1 U10424 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11750) );
  OR2_X1 U10425 ( .A1(n8117), .A2(n11750), .ZN(n8029) );
  INV_X1 U10426 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n8027) );
  OR2_X1 U10427 ( .A1(n8247), .A2(n8027), .ZN(n8028) );
  NAND4_X1 U10428 ( .A1(n8031), .A2(n8030), .A3(n8029), .A4(n8028), .ZN(n12770) );
  INV_X1 U10429 ( .A(n12770), .ZN(n12079) );
  OR2_X1 U10430 ( .A1(n14481), .A2(n12079), .ZN(n12689) );
  NAND2_X1 U10431 ( .A1(n14481), .A2(n12079), .ZN(n12694) );
  NAND2_X1 U10432 ( .A1(n12689), .A2(n12694), .ZN(n12592) );
  OR2_X1 U10433 ( .A1(n14490), .A2(n12771), .ZN(n11746) );
  AND2_X1 U10434 ( .A1(n12592), .A2(n11746), .ZN(n8032) );
  NAND2_X1 U10435 ( .A1(n11800), .A2(n8032), .ZN(n11745) );
  NAND2_X1 U10436 ( .A1(n14481), .A2(n12770), .ZN(n8033) );
  NAND2_X1 U10437 ( .A1(n11745), .A2(n8033), .ZN(n11773) );
  INV_X1 U10438 ( .A(n11773), .ZN(n8052) );
  OR2_X1 U10439 ( .A1(n8035), .A2(n8034), .ZN(n8036) );
  NAND2_X1 U10440 ( .A1(n8037), .A2(n8036), .ZN(n10251) );
  NAND2_X1 U10441 ( .A1(n8039), .A2(n8038), .ZN(n8041) );
  NAND2_X1 U10442 ( .A1(n8041), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8040) );
  MUX2_X1 U10443 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8040), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n8042) );
  AOI22_X1 U10444 ( .A1(n8215), .A2(SI_15_), .B1(n8113), .B2(n12853), .ZN(
        n8043) );
  NAND2_X1 U10445 ( .A1(n8045), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10446 ( .A1(n8066), .A2(n8046), .ZN(n12081) );
  NAND2_X1 U10447 ( .A1(n8222), .A2(n12081), .ZN(n8051) );
  NAND2_X1 U10448 ( .A1(n7842), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8050) );
  INV_X1 U10449 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n8047) );
  OR2_X1 U10450 ( .A1(n8247), .A2(n8047), .ZN(n8049) );
  INV_X1 U10451 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12825) );
  OR2_X1 U10452 ( .A1(n6561), .A2(n12825), .ZN(n8048) );
  NAND4_X1 U10453 ( .A1(n8051), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(n14415) );
  OR2_X1 U10454 ( .A1(n13137), .A2(n14415), .ZN(n8053) );
  OR2_X1 U10455 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  NAND2_X1 U10456 ( .A1(n8057), .A2(n8056), .ZN(n10295) );
  NAND2_X1 U10457 ( .A1(n8059), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8058) );
  MUX2_X1 U10458 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8058), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n8062) );
  INV_X1 U10459 ( .A(n8059), .ZN(n8061) );
  INV_X1 U10460 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10461 ( .A1(n8061), .A2(n8060), .ZN(n8092) );
  NAND2_X1 U10462 ( .A1(n8062), .A2(n8092), .ZN(n12845) );
  INV_X1 U10463 ( .A(n8063), .ZN(n8064) );
  INV_X1 U10464 ( .A(n8081), .ZN(n8068) );
  NAND2_X1 U10465 ( .A1(n8066), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10466 ( .A1(n8068), .A2(n8067), .ZN(n14443) );
  NAND2_X1 U10467 ( .A1(n8222), .A2(n14443), .ZN(n8072) );
  NAND2_X1 U10468 ( .A1(n8246), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8071) );
  INV_X1 U10469 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13194) );
  OR2_X1 U10470 ( .A1(n8247), .A2(n13194), .ZN(n8070) );
  INV_X1 U10471 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12855) );
  OR2_X1 U10472 ( .A1(n8117), .A2(n12855), .ZN(n8069) );
  NAND4_X1 U10473 ( .A1(n8072), .A2(n8071), .A3(n8070), .A4(n8069), .ZN(n12769) );
  NAND2_X1 U10474 ( .A1(n14442), .A2(n12769), .ZN(n8073) );
  XNOR2_X1 U10475 ( .A(n8076), .B(n8075), .ZN(n10381) );
  NAND2_X1 U10476 ( .A1(n10381), .A2(n8214), .ZN(n8079) );
  NAND2_X1 U10477 ( .A1(n8092), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8077) );
  XNOR2_X1 U10478 ( .A(n8077), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U10479 ( .A1(n8113), .A2(n14466), .B1(n8215), .B2(SI_17_), .ZN(
        n8078) );
  NAND2_X1 U10480 ( .A1(n8079), .A2(n8078), .ZN(n12521) );
  NOR2_X1 U10481 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  OR2_X1 U10482 ( .A1(n8096), .A2(n8082), .ZN(n13068) );
  NAND2_X1 U10483 ( .A1(n8222), .A2(n13068), .ZN(n8086) );
  NAND2_X1 U10484 ( .A1(n8246), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8085) );
  INV_X1 U10485 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13190) );
  OR2_X1 U10486 ( .A1(n8247), .A2(n13190), .ZN(n8084) );
  INV_X1 U10487 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14476) );
  OR2_X1 U10488 ( .A1(n8117), .A2(n14476), .ZN(n8083) );
  NAND4_X1 U10489 ( .A1(n8086), .A2(n8085), .A3(n8084), .A4(n8083), .ZN(n13050) );
  INV_X1 U10490 ( .A(n13050), .ZN(n12562) );
  OR2_X1 U10491 ( .A1(n12521), .A2(n12562), .ZN(n12706) );
  NAND2_X1 U10492 ( .A1(n12521), .A2(n12562), .ZN(n12705) );
  NAND2_X1 U10493 ( .A1(n12706), .A2(n12705), .ZN(n13061) );
  AND2_X1 U10494 ( .A1(n12521), .A2(n13050), .ZN(n8087) );
  OR2_X1 U10495 ( .A1(n8089), .A2(n8088), .ZN(n8090) );
  NAND2_X1 U10496 ( .A1(n8091), .A2(n8090), .ZN(n10408) );
  OAI21_X1 U10497 ( .B1(n8092), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8093) );
  XNOR2_X1 U10498 ( .A(n8093), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12884) );
  AOI22_X1 U10499 ( .A1(n12884), .A2(n8113), .B1(SI_18_), .B2(n8215), .ZN(
        n8094) );
  OR2_X1 U10500 ( .A1(n8096), .A2(n12559), .ZN(n8097) );
  NAND2_X1 U10501 ( .A1(n8116), .A2(n8097), .ZN(n13057) );
  NAND2_X1 U10502 ( .A1(n8222), .A2(n13057), .ZN(n8102) );
  NAND2_X1 U10503 ( .A1(n8246), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8101) );
  INV_X1 U10504 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8098) );
  OR2_X1 U10505 ( .A1(n6561), .A2(n8098), .ZN(n8100) );
  INV_X1 U10506 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13186) );
  OR2_X1 U10507 ( .A1(n8247), .A2(n13186), .ZN(n8099) );
  NAND4_X1 U10508 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n13035) );
  NAND2_X1 U10509 ( .A1(n13056), .A2(n13065), .ZN(n12712) );
  NAND2_X1 U10510 ( .A1(n13039), .A2(n12712), .ZN(n13055) );
  OR2_X1 U10511 ( .A1(n13056), .A2(n13035), .ZN(n8103) );
  OR2_X1 U10512 ( .A1(n8105), .A2(n8104), .ZN(n8106) );
  NAND2_X1 U10513 ( .A1(n8107), .A2(n8106), .ZN(n10529) );
  NAND2_X1 U10514 ( .A1(n10529), .A2(n8214), .ZN(n8115) );
  NAND2_X1 U10515 ( .A1(n8111), .A2(n8110), .ZN(n8242) );
  AOI22_X1 U10516 ( .A1(n8215), .A2(n10530), .B1(n8113), .B2(n12883), .ZN(
        n8114) );
  XNOR2_X1 U10517 ( .A(n8116), .B(P3_REG3_REG_19__SCAN_IN), .ZN(n13043) );
  NAND2_X1 U10518 ( .A1(n13043), .A2(n8222), .ZN(n8121) );
  INV_X1 U10519 ( .A(n8117), .ZN(n12580) );
  NAND2_X1 U10520 ( .A1(n12580), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10521 ( .A1(n8246), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10522 ( .A1(n7887), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8118) );
  NAND4_X1 U10523 ( .A1(n8121), .A2(n8120), .A3(n8119), .A4(n8118), .ZN(n13049) );
  NAND2_X1 U10524 ( .A1(n13184), .A2(n13049), .ZN(n12719) );
  INV_X1 U10525 ( .A(n13049), .ZN(n13020) );
  OR2_X1 U10526 ( .A1(n13184), .A2(n13020), .ZN(n8123) );
  NAND2_X1 U10527 ( .A1(n13031), .A2(n8123), .ZN(n13018) );
  OR2_X1 U10528 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  NAND2_X1 U10529 ( .A1(n8127), .A2(n8126), .ZN(n10575) );
  NAND2_X1 U10530 ( .A1(n8215), .A2(SI_20_), .ZN(n8128) );
  INV_X1 U10531 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13178) );
  AND2_X1 U10532 ( .A1(n8130), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8131) );
  OR2_X1 U10533 ( .A1(n8131), .A2(n8142), .ZN(n13022) );
  NAND2_X1 U10534 ( .A1(n13022), .A2(n8222), .ZN(n8133) );
  AOI22_X1 U10535 ( .A1(n12580), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n7842), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n8132) );
  OAI211_X1 U10536 ( .C1(n8247), .C2(n13178), .A(n8133), .B(n8132), .ZN(n13036) );
  INV_X1 U10537 ( .A(n13036), .ZN(n13003) );
  NAND2_X1 U10538 ( .A1(n13113), .A2(n13003), .ZN(n12723) );
  NAND2_X1 U10539 ( .A1(n12722), .A2(n12723), .ZN(n13017) );
  NAND2_X1 U10540 ( .A1(n13113), .A2(n13036), .ZN(n8134) );
  OR2_X1 U10541 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  NAND2_X1 U10542 ( .A1(n8138), .A2(n8137), .ZN(n10825) );
  NAND2_X1 U10543 ( .A1(n8215), .A2(SI_21_), .ZN(n8139) );
  NOR2_X1 U10544 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  OR2_X1 U10545 ( .A1(n8153), .A2(n8143), .ZN(n13007) );
  NAND2_X1 U10546 ( .A1(n13007), .A2(n8222), .ZN(n8146) );
  AOI22_X1 U10547 ( .A1(n12580), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n7842), 
        .B2(P3_REG1_REG_21__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10548 ( .A1(n7887), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8144) );
  AND2_X1 U10549 ( .A1(n13006), .A2(n12768), .ZN(n12590) );
  OR2_X1 U10550 ( .A1(n13006), .A2(n12768), .ZN(n12589) );
  OR2_X1 U10551 ( .A1(n8148), .A2(n8147), .ZN(n8149) );
  NAND2_X1 U10552 ( .A1(n8150), .A2(n8149), .ZN(n10851) );
  NAND2_X1 U10553 ( .A1(n8215), .A2(SI_22_), .ZN(n8151) );
  OR2_X1 U10554 ( .A1(n8153), .A2(n12552), .ZN(n8154) );
  NAND2_X1 U10555 ( .A1(n8166), .A2(n8154), .ZN(n12995) );
  NAND2_X1 U10556 ( .A1(n12995), .A2(n8222), .ZN(n8160) );
  INV_X1 U10557 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10558 ( .A1(n8246), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U10559 ( .A1(n7887), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8155) );
  OAI211_X1 U10560 ( .C1(n6561), .C2(n8157), .A(n8156), .B(n8155), .ZN(n8158)
         );
  INV_X1 U10561 ( .A(n8158), .ZN(n8159) );
  NAND2_X1 U10562 ( .A1(n8160), .A2(n8159), .ZN(n12551) );
  NOR2_X1 U10563 ( .A1(n9197), .A2(n12551), .ZN(n8161) );
  XNOR2_X1 U10564 ( .A(n8163), .B(n8162), .ZN(n10964) );
  NAND2_X1 U10565 ( .A1(n10964), .A2(n8214), .ZN(n8165) );
  NAND2_X1 U10566 ( .A1(n8215), .A2(SI_23_), .ZN(n8164) );
  NAND2_X1 U10567 ( .A1(n8166), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10568 ( .A1(n8179), .A2(n8167), .ZN(n12982) );
  NAND2_X1 U10569 ( .A1(n12982), .A2(n8222), .ZN(n8172) );
  INV_X1 U10570 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n15364) );
  NAND2_X1 U10571 ( .A1(n8246), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10572 ( .A1(n12580), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8168) );
  OAI211_X1 U10573 ( .C1(n8247), .C2(n15364), .A(n8169), .B(n8168), .ZN(n8170)
         );
  INV_X1 U10574 ( .A(n8170), .ZN(n8171) );
  INV_X1 U10575 ( .A(n12731), .ZN(n8173) );
  NAND2_X1 U10576 ( .A1(n12986), .A2(n8173), .ZN(n8174) );
  NAND2_X1 U10577 ( .A1(n12986), .A2(n12731), .ZN(n8175) );
  XNOR2_X1 U10578 ( .A(n8176), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11384) );
  NAND2_X1 U10579 ( .A1(n11384), .A2(n8214), .ZN(n8178) );
  NAND2_X1 U10580 ( .A1(n8215), .A2(SI_24_), .ZN(n8177) );
  NAND2_X1 U10581 ( .A1(n8179), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10582 ( .A1(n8194), .A2(n8180), .ZN(n12970) );
  INV_X1 U10583 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10584 ( .A1(n7887), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10585 ( .A1(n8246), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8181) );
  OAI211_X1 U10586 ( .C1(n6561), .C2(n8183), .A(n8182), .B(n8181), .ZN(n8184)
         );
  INV_X1 U10587 ( .A(n12978), .ZN(n12767) );
  OR2_X1 U10588 ( .A1(n12531), .A2(n12767), .ZN(n8185) );
  NAND2_X1 U10589 ( .A1(n8186), .A2(n8185), .ZN(n12953) );
  OR2_X1 U10590 ( .A1(n8188), .A2(n8187), .ZN(n8189) );
  NAND2_X1 U10591 ( .A1(n8190), .A2(n8189), .ZN(n11423) );
  NAND2_X1 U10592 ( .A1(n8215), .A2(SI_25_), .ZN(n8192) );
  NAND2_X1 U10593 ( .A1(n8194), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10594 ( .A1(n8195), .A2(n6599), .ZN(n12961) );
  INV_X1 U10595 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10596 ( .A1(n7887), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10597 ( .A1(n7842), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U10598 ( .C1(n8117), .C2(n8198), .A(n8197), .B(n8196), .ZN(n8199)
         );
  AOI21_X1 U10599 ( .B1(n12961), .B2(n8222), .A(n8199), .ZN(n9210) );
  OR2_X1 U10600 ( .A1(n12960), .A2(n9210), .ZN(n12739) );
  NAND2_X1 U10601 ( .A1(n12960), .A2(n9210), .ZN(n12938) );
  INV_X1 U10602 ( .A(n9210), .ZN(n12766) );
  NAND2_X1 U10603 ( .A1(n12960), .A2(n12766), .ZN(n8201) );
  XNOR2_X1 U10604 ( .A(n8203), .B(n8202), .ZN(n11625) );
  NAND2_X1 U10605 ( .A1(n11625), .A2(n8214), .ZN(n8205) );
  NAND2_X1 U10606 ( .A1(n8215), .A2(SI_26_), .ZN(n8204) );
  AOI21_X1 U10607 ( .B1(P3_REG3_REG_26__SCAN_IN), .B2(n6599), .A(n8218), .ZN(
        n12946) );
  NAND2_X1 U10608 ( .A1(n7842), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8208) );
  INV_X1 U10609 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12947) );
  OR2_X1 U10610 ( .A1(n8117), .A2(n12947), .ZN(n8207) );
  INV_X1 U10611 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n15254) );
  OR2_X1 U10612 ( .A1(n8247), .A2(n15254), .ZN(n8206) );
  OR2_X1 U10613 ( .A1(n12949), .A2(n12928), .ZN(n8211) );
  AND2_X1 U10614 ( .A1(n12949), .A2(n12928), .ZN(n8210) );
  XNOR2_X1 U10615 ( .A(n8213), .B(n8212), .ZN(n11713) );
  NAND2_X1 U10616 ( .A1(n11713), .A2(n8214), .ZN(n8217) );
  NAND2_X1 U10617 ( .A1(n8215), .A2(SI_27_), .ZN(n8216) );
  INV_X1 U10618 ( .A(n8218), .ZN(n8219) );
  NAND2_X1 U10619 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8219), .ZN(n8220) );
  NAND2_X1 U10620 ( .A1(n8221), .A2(n8220), .ZN(n12930) );
  NAND2_X1 U10621 ( .A1(n8222), .A2(n12930), .ZN(n8227) );
  NAND2_X1 U10622 ( .A1(n7842), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8226) );
  INV_X1 U10623 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12932) );
  OR2_X1 U10624 ( .A1(n8117), .A2(n12932), .ZN(n8225) );
  INV_X1 U10625 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8223) );
  OR2_X1 U10626 ( .A1(n8247), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U10627 ( .A1(n13084), .A2(n8228), .ZN(n12917) );
  NAND2_X1 U10628 ( .A1(n12920), .A2(n8245), .ZN(n8273) );
  NAND2_X1 U10629 ( .A1(n12621), .A2(n8273), .ZN(n12475) );
  NOR2_X1 U10630 ( .A1(n12909), .A2(n12918), .ZN(n12912) );
  AOI21_X1 U10631 ( .B1(n12927), .B2(n12920), .A(n12912), .ZN(n8229) );
  INV_X1 U10632 ( .A(n8229), .ZN(n8238) );
  NAND2_X1 U10633 ( .A1(n8231), .A2(n8230), .ZN(n12367) );
  INV_X1 U10634 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13695) );
  XNOR2_X1 U10635 ( .A(n13695), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n8232) );
  XNOR2_X1 U10636 ( .A(n12367), .B(n8232), .ZN(n13205) );
  NAND2_X1 U10637 ( .A1(n13205), .A2(n8214), .ZN(n8234) );
  NAND2_X1 U10638 ( .A1(n8215), .A2(SI_29_), .ZN(n8233) );
  NAND2_X1 U10639 ( .A1(n7842), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8237) );
  INV_X1 U10640 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12902) );
  OR2_X1 U10641 ( .A1(n6561), .A2(n12902), .ZN(n8236) );
  INV_X1 U10642 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8321) );
  OR2_X1 U10643 ( .A1(n8247), .A2(n8321), .ZN(n8235) );
  NAND2_X1 U10644 ( .A1(n12905), .A2(n12765), .ZN(n12614) );
  NAND2_X1 U10645 ( .A1(n12612), .A2(n12614), .ZN(n12611) );
  NAND2_X1 U10646 ( .A1(n6679), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10647 ( .A1(n12872), .A2(n12761), .ZN(n8309) );
  NAND2_X1 U10648 ( .A1(n8240), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10649 ( .A1(n8242), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10650 ( .A1(n12630), .A2(n9250), .ZN(n12619) );
  INV_X1 U10651 ( .A(n12759), .ZN(n10534) );
  INV_X1 U10652 ( .A(n6973), .ZN(n12805) );
  NAND2_X1 U10653 ( .A1(n10534), .A2(n12805), .ZN(n10554) );
  NAND2_X1 U10654 ( .A1(n8246), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8250) );
  OR2_X1 U10655 ( .A1(n8247), .A2(n13150), .ZN(n8249) );
  INV_X1 U10656 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n12899) );
  OR2_X1 U10657 ( .A1(n6561), .A2(n12899), .ZN(n8248) );
  INV_X1 U10658 ( .A(P3_B_REG_SCAN_IN), .ZN(n8252) );
  NOR2_X1 U10659 ( .A1(n12759), .A2(n8252), .ZN(n8253) );
  OR2_X1 U10660 ( .A1(n15050), .A2(n8253), .ZN(n12893) );
  NAND2_X1 U10661 ( .A1(n10867), .A2(n12593), .ZN(n8257) );
  NAND2_X1 U10662 ( .A1(n8257), .A2(n12640), .ZN(n10857) );
  INV_X1 U10663 ( .A(n10859), .ZN(n12645) );
  NAND2_X1 U10664 ( .A1(n10857), .A2(n12645), .ZN(n8258) );
  INV_X1 U10665 ( .A(n10896), .ZN(n12594) );
  NAND2_X1 U10666 ( .A1(n8259), .A2(n12660), .ZN(n11112) );
  NAND2_X1 U10667 ( .A1(n11112), .A2(n12659), .ZN(n8261) );
  INV_X1 U10668 ( .A(n12777), .ZN(n8260) );
  NAND2_X1 U10669 ( .A1(n8260), .A2(n12661), .ZN(n12662) );
  NOR2_X1 U10670 ( .A1(n12775), .A2(n15120), .ZN(n8262) );
  NAND2_X1 U10671 ( .A1(n12775), .A2(n15120), .ZN(n8263) );
  INV_X1 U10672 ( .A(n12675), .ZN(n8264) );
  NAND2_X1 U10673 ( .A1(n11631), .A2(n11451), .ZN(n12679) );
  OR2_X1 U10674 ( .A1(n14492), .A2(n12772), .ZN(n12687) );
  NAND2_X1 U10675 ( .A1(n14492), .A2(n12772), .ZN(n12680) );
  NAND2_X1 U10676 ( .A1(n11588), .A2(n11587), .ZN(n8265) );
  INV_X1 U10677 ( .A(n12688), .ZN(n8266) );
  INV_X1 U10678 ( .A(n14415), .ZN(n8267) );
  OR2_X1 U10679 ( .A1(n13137), .A2(n8267), .ZN(n12696) );
  NAND2_X1 U10680 ( .A1(n13137), .A2(n8267), .ZN(n12700) );
  NAND2_X1 U10681 ( .A1(n12696), .A2(n12700), .ZN(n11777) );
  INV_X1 U10682 ( .A(n12769), .ZN(n13066) );
  OR2_X1 U10683 ( .A1(n14442), .A2(n13066), .ZN(n12702) );
  NAND2_X1 U10684 ( .A1(n14442), .A2(n13066), .ZN(n12701) );
  INV_X1 U10685 ( .A(n13039), .ZN(n12708) );
  NOR2_X1 U10686 ( .A1(n8122), .A2(n12708), .ZN(n8269) );
  INV_X1 U10687 ( .A(n13013), .ZN(n12714) );
  NOR2_X1 U10688 ( .A1(n13017), .A2(n12714), .ZN(n8270) );
  NAND2_X1 U10689 ( .A1(n13015), .A2(n12722), .ZN(n13004) );
  NOR2_X1 U10690 ( .A1(n13006), .A2(n13021), .ZN(n12725) );
  NAND2_X1 U10691 ( .A1(n13006), .A2(n13021), .ZN(n12727) );
  AND2_X1 U10692 ( .A1(n9197), .A2(n13002), .ZN(n12624) );
  OR2_X1 U10693 ( .A1(n12531), .A2(n12978), .ZN(n12735) );
  NAND2_X1 U10694 ( .A1(n12531), .A2(n12978), .ZN(n12734) );
  NAND2_X1 U10695 ( .A1(n12735), .A2(n12734), .ZN(n12968) );
  NAND2_X1 U10696 ( .A1(n12969), .A2(n12734), .ZN(n12959) );
  INV_X1 U10697 ( .A(n12928), .ZN(n9234) );
  NAND2_X1 U10698 ( .A1(n12949), .A2(n9234), .ZN(n12744) );
  NAND2_X1 U10699 ( .A1(n12743), .A2(n12744), .ZN(n12942) );
  INV_X1 U10700 ( .A(n12938), .ZN(n8271) );
  NOR2_X1 U10701 ( .A1(n12942), .A2(n8271), .ZN(n8272) );
  NAND2_X1 U10702 ( .A1(n8273), .A2(n12917), .ZN(n12622) );
  XNOR2_X1 U10703 ( .A(n12613), .B(n12611), .ZN(n12900) );
  NAND2_X1 U10704 ( .A1(n10827), .A2(n10577), .ZN(n8274) );
  XNOR2_X1 U10705 ( .A(n12761), .B(n8274), .ZN(n8276) );
  NAND2_X1 U10706 ( .A1(n12883), .A2(n10827), .ZN(n8275) );
  NAND2_X1 U10707 ( .A1(n8276), .A2(n8275), .ZN(n9225) );
  INV_X1 U10708 ( .A(n9251), .ZN(n12756) );
  INV_X1 U10709 ( .A(n12761), .ZN(n8277) );
  AND2_X1 U10710 ( .A1(n12756), .A2(n15124), .ZN(n8278) );
  NAND2_X1 U10711 ( .A1(n9225), .A2(n8278), .ZN(n8279) );
  NAND3_X1 U10712 ( .A1(n12761), .A2(n9250), .A3(n12883), .ZN(n9248) );
  NAND2_X1 U10713 ( .A1(n8279), .A2(n9248), .ZN(n15118) );
  INV_X1 U10714 ( .A(n8286), .ZN(n8290) );
  NAND2_X1 U10715 ( .A1(n8317), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8283) );
  MUX2_X1 U10716 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8283), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8284) );
  XNOR2_X1 U10717 ( .A(n8294), .B(P3_B_REG_SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10718 ( .A1(n8289), .A2(n11422), .ZN(n8292) );
  OR2_X1 U10719 ( .A1(n8295), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10720 ( .A1(n11628), .A2(n11422), .ZN(n8296) );
  INV_X1 U10721 ( .A(n10485), .ZN(n13199) );
  NOR2_X1 U10722 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .ZN(
        n8301) );
  NOR4_X1 U10723 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8300) );
  NOR4_X1 U10724 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8299) );
  NOR4_X1 U10725 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8298) );
  NAND4_X1 U10726 ( .A1(n8301), .A2(n8300), .A3(n8299), .A4(n8298), .ZN(n8307)
         );
  NOR4_X1 U10727 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8305) );
  NOR4_X1 U10728 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8304) );
  NOR4_X1 U10729 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8303) );
  NOR4_X1 U10730 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8302) );
  NAND4_X1 U10731 ( .A1(n8305), .A2(n8304), .A3(n8303), .A4(n8302), .ZN(n8306)
         );
  NOR2_X1 U10732 ( .A1(n8307), .A2(n8306), .ZN(n8308) );
  OR2_X1 U10733 ( .A1(n8295), .A2(n8308), .ZN(n9243) );
  NAND2_X1 U10734 ( .A1(n9241), .A2(n9243), .ZN(n9226) );
  NAND2_X1 U10735 ( .A1(n10827), .A2(n9250), .ZN(n9128) );
  NOR2_X1 U10736 ( .A1(n8309), .A2(n9128), .ZN(n9224) );
  NOR2_X1 U10737 ( .A1(n9224), .A2(n10286), .ZN(n8312) );
  INV_X1 U10738 ( .A(n9225), .ZN(n8311) );
  OAI22_X1 U10739 ( .A1(n9226), .A2(n8312), .B1(n9232), .B2(n8311), .ZN(n8318)
         );
  INV_X1 U10740 ( .A(n11422), .ZN(n8313) );
  NAND2_X1 U10741 ( .A1(n8313), .A2(n6781), .ZN(n8314) );
  NAND2_X1 U10742 ( .A1(n6738), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8315) );
  MUX2_X1 U10743 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8315), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8316) );
  INV_X1 U10744 ( .A(n13200), .ZN(n10066) );
  INV_X1 U10745 ( .A(n12905), .ZN(n9260) );
  NOR2_X1 U10746 ( .A1(n8320), .A2(n8322), .ZN(n8323) );
  NAND2_X1 U10747 ( .A1(n8324), .A2(n8323), .ZN(P3_U3456) );
  NAND4_X1 U10748 ( .A1(n8329), .A2(n15399), .A3(n8328), .A4(n8327), .ZN(n8712) );
  NAND4_X1 U10749 ( .A1(n8331), .A2(n8330), .A3(n8592), .A4(n15400), .ZN(n8332) );
  NOR2_X1 U10750 ( .A1(n8712), .A2(n8332), .ZN(n8333) );
  INV_X1 U10751 ( .A(n8971), .ZN(n8335) );
  INV_X1 U10752 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10753 ( .A1(n8335), .A2(n8334), .ZN(n8337) );
  INV_X1 U10754 ( .A(n8967), .ZN(n8979) );
  OAI21_X1 U10755 ( .B1(P2_IR_REG_21__SCAN_IN), .B2(P2_IR_REG_20__SCAN_IN), 
        .A(P2_IR_REG_22__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10756 ( .A1(n8338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8339) );
  OAI21_X1 U10757 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n8340), .A(n8339), .ZN(
        n8343) );
  OR2_X1 U10758 ( .A1(n8341), .A2(n8340), .ZN(n8342) );
  INV_X1 U10759 ( .A(n8352), .ZN(n8344) );
  NAND2_X2 U10760 ( .A1(n9732), .A2(n11185), .ZN(n8410) );
  NOR2_X1 U10761 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8347) );
  NOR2_X1 U10762 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8346) );
  NAND3_X1 U10763 ( .A1(n8349), .A2(n8354), .A3(n8348), .ZN(n8350) );
  AND2_X1 U10764 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n8359) );
  INV_X1 U10765 ( .A(n8970), .ZN(n8357) );
  AND2_X1 U10766 ( .A1(n8354), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n8356) );
  INV_X1 U10767 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8568) );
  XNOR2_X1 U10768 ( .A(n8568), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8355) );
  AOI21_X1 U10769 ( .B1(n8357), .B2(n8356), .A(n8355), .ZN(n8358) );
  INV_X1 U10770 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10052) );
  OAI21_X1 U10771 ( .B1(n8417), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n8360), .ZN(
        n8396) );
  AND2_X1 U10772 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8361) );
  NAND2_X1 U10773 ( .A1(n6566), .A2(n8361), .ZN(n9304) );
  AND2_X1 U10774 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10775 ( .A1(n8417), .A2(n8362), .ZN(n8392) );
  XNOR2_X1 U10776 ( .A(n8398), .B(n8397), .ZN(n10051) );
  NAND2_X1 U10777 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8364) );
  MUX2_X1 U10778 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8364), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8367) );
  INV_X1 U10779 ( .A(n8365), .ZN(n8366) );
  NAND2_X1 U10780 ( .A1(n8367), .A2(n8366), .ZN(n10331) );
  INV_X1 U10781 ( .A(n10331), .ZN(n10170) );
  NAND2_X1 U10782 ( .A1(n8380), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10783 ( .A1(n8386), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10784 ( .A1(n13325), .A2(n6569), .ZN(n8379) );
  NAND2_X1 U10785 ( .A1(n8378), .A2(n8379), .ZN(n8395) );
  NAND2_X1 U10786 ( .A1(n8576), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8389) );
  INV_X1 U10787 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8381) );
  NOR2_X1 U10788 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  NOR2_X1 U10789 ( .A1(n8385), .A2(n8384), .ZN(n8388) );
  NAND2_X1 U10790 ( .A1(n8386), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8387) );
  NAND3_X1 U10791 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n9734) );
  NAND2_X1 U10792 ( .A1(n10006), .A2(SI_0_), .ZN(n8391) );
  NAND2_X1 U10793 ( .A1(n8391), .A2(n8390), .ZN(n8393) );
  NAND2_X1 U10794 ( .A1(n8393), .A2(n8392), .ZN(n13701) );
  INV_X1 U10795 ( .A(n8811), .ZN(n13525) );
  OAI22_X1 U10796 ( .A1(n10607), .A2(n13525), .B1(n8410), .B2(n10807), .ZN(
        n10731) );
  NAND2_X1 U10797 ( .A1(n10728), .A2(n8395), .ZN(n10579) );
  INV_X1 U10798 ( .A(SI_1_), .ZN(n10008) );
  MUX2_X1 U10799 ( .A(n10053), .B(n10034), .S(n8417), .Z(n8414) );
  XNOR2_X1 U10800 ( .A(n8414), .B(SI_2_), .ZN(n8412) );
  XNOR2_X1 U10801 ( .A(n8411), .B(n8412), .ZN(n9312) );
  OR2_X1 U10802 ( .A1(n8365), .A2(n8568), .ZN(n8399) );
  XNOR2_X1 U10803 ( .A(n8399), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U10804 ( .A1(n10141), .A2(n10222), .ZN(n8400) );
  XNOR2_X1 U10805 ( .A(n8410), .B(n10776), .ZN(n8407) );
  NAND2_X1 U10806 ( .A1(n8380), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U10807 ( .A1(n8576), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U10808 ( .A1(n9931), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10809 ( .A1(n8386), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8402) );
  INV_X1 U10810 ( .A(n8811), .ZN(n11860) );
  NAND2_X1 U10811 ( .A1(n13323), .A2(n8811), .ZN(n8406) );
  NAND2_X1 U10812 ( .A1(n8407), .A2(n8406), .ZN(n8409) );
  OR2_X1 U10813 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  AND2_X1 U10814 ( .A1(n8409), .A2(n8408), .ZN(n10580) );
  NAND2_X1 U10815 ( .A1(n10579), .A2(n10580), .ZN(n10578) );
  INV_X1 U10816 ( .A(n8414), .ZN(n8415) );
  NAND2_X1 U10817 ( .A1(n8415), .A2(SI_2_), .ZN(n8416) );
  MUX2_X1 U10818 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8417), .Z(n8432) );
  XNOR2_X1 U10819 ( .A(n8431), .B(n8429), .ZN(n10026) );
  NAND2_X1 U10820 ( .A1(n10026), .A2(n8434), .ZN(n8421) );
  NAND2_X1 U10821 ( .A1(n8418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8419) );
  XNOR2_X1 U10822 ( .A(n8419), .B(P2_IR_REG_3__SCAN_IN), .ZN(n13335) );
  AOI22_X1 U10823 ( .A1(n9926), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10141), 
        .B2(n13335), .ZN(n8420) );
  XNOR2_X1 U10824 ( .A(n8410), .B(n14837), .ZN(n8428) );
  INV_X2 U10825 ( .A(n8422), .ZN(n9020) );
  INV_X1 U10826 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10827 ( .A1(n8526), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U10828 ( .A1(n6565), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10829 ( .A1(n9931), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8424) );
  AND2_X1 U10830 ( .A1(n13322), .A2(n8811), .ZN(n8427) );
  XNOR2_X1 U10831 ( .A(n8428), .B(n8427), .ZN(n10657) );
  NAND2_X1 U10832 ( .A1(n8432), .A2(SI_3_), .ZN(n8433) );
  XNOR2_X1 U10833 ( .A(n8452), .B(SI_4_), .ZN(n8449) );
  XNOR2_X1 U10834 ( .A(n8451), .B(n8449), .ZN(n10035) );
  CLKBUF_X3 U10835 ( .A(n8434), .Z(n9894) );
  NAND2_X1 U10836 ( .A1(n10035), .A2(n9894), .ZN(n8438) );
  NAND2_X1 U10837 ( .A1(n8435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8436) );
  XNOR2_X1 U10838 ( .A(n8436), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U10839 ( .A1(n9926), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10141), 
        .B2(n10174), .ZN(n8437) );
  NAND2_X1 U10840 ( .A1(n8438), .A2(n8437), .ZN(n14848) );
  XNOR2_X1 U10841 ( .A(n14848), .B(n8964), .ZN(n8443) );
  NAND2_X1 U10842 ( .A1(n9931), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10843 ( .A1(n8526), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8441) );
  INV_X1 U10844 ( .A(n8460), .ZN(n8461) );
  OAI21_X1 U10845 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8461), .ZN(n10761) );
  INV_X1 U10846 ( .A(n10761), .ZN(n10513) );
  NAND2_X1 U10847 ( .A1(n9020), .A2(n10513), .ZN(n8440) );
  NAND2_X1 U10848 ( .A1(n6565), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8439) );
  NAND4_X1 U10849 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n13321) );
  NAND2_X1 U10850 ( .A1(n13321), .A2(n8811), .ZN(n8444) );
  NAND2_X1 U10851 ( .A1(n8443), .A2(n8444), .ZN(n8448) );
  INV_X1 U10852 ( .A(n8443), .ZN(n8446) );
  INV_X1 U10853 ( .A(n8444), .ZN(n8445) );
  NAND2_X1 U10854 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  INV_X1 U10855 ( .A(n8449), .ZN(n8450) );
  NAND2_X1 U10856 ( .A1(n8451), .A2(n8450), .ZN(n8454) );
  NAND2_X1 U10857 ( .A1(n8452), .A2(SI_4_), .ZN(n8453) );
  MUX2_X1 U10858 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10025), .Z(n8477) );
  XNOR2_X1 U10859 ( .A(n8477), .B(SI_5_), .ZN(n8474) );
  XNOR2_X1 U10860 ( .A(n8476), .B(n8474), .ZN(n10029) );
  NAND2_X1 U10861 ( .A1(n10029), .A2(n9894), .ZN(n8459) );
  INV_X1 U10862 ( .A(n8435), .ZN(n8456) );
  NAND2_X1 U10863 ( .A1(n8456), .A2(n8455), .ZN(n8479) );
  NAND2_X1 U10864 ( .A1(n8479), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8457) );
  XNOR2_X1 U10865 ( .A(n8457), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U10866 ( .A1(n9926), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10141), 
        .B2(n10187), .ZN(n8458) );
  NAND2_X1 U10867 ( .A1(n8459), .A2(n8458), .ZN(n10919) );
  XNOR2_X1 U10868 ( .A(n10919), .B(n8964), .ZN(n8468) );
  NAND2_X1 U10869 ( .A1(n9931), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10870 ( .A1(n8526), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10871 ( .A1(n8460), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8486) );
  INV_X1 U10872 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n15220) );
  NAND2_X1 U10873 ( .A1(n8461), .A2(n15220), .ZN(n8462) );
  AND2_X1 U10874 ( .A1(n8486), .A2(n8462), .ZN(n10918) );
  NAND2_X1 U10875 ( .A1(n9020), .A2(n10918), .ZN(n8465) );
  NAND2_X1 U10876 ( .A1(n6565), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8464) );
  NAND4_X1 U10877 ( .A1(n8467), .A2(n8466), .A3(n8465), .A4(n8464), .ZN(n13320) );
  NAND2_X1 U10878 ( .A1(n13320), .A2(n8811), .ZN(n8469) );
  NAND2_X1 U10879 ( .A1(n8468), .A2(n8469), .ZN(n8473) );
  INV_X1 U10880 ( .A(n8468), .ZN(n8471) );
  INV_X1 U10881 ( .A(n8469), .ZN(n8470) );
  NAND2_X1 U10882 ( .A1(n8471), .A2(n8470), .ZN(n8472) );
  AND2_X1 U10883 ( .A1(n8473), .A2(n8472), .ZN(n10498) );
  NAND2_X1 U10884 ( .A1(n10497), .A2(n10498), .ZN(n10496) );
  INV_X1 U10885 ( .A(n8474), .ZN(n8475) );
  NAND2_X1 U10886 ( .A1(n8477), .A2(SI_5_), .ZN(n8478) );
  MUX2_X1 U10887 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10006), .Z(n8500) );
  XNOR2_X1 U10888 ( .A(n8500), .B(SI_6_), .ZN(n8497) );
  XNOR2_X1 U10889 ( .A(n8499), .B(n8497), .ZN(n10038) );
  NAND2_X1 U10890 ( .A1(n10038), .A2(n9894), .ZN(n8484) );
  INV_X1 U10891 ( .A(n8479), .ZN(n8481) );
  INV_X1 U10892 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U10893 ( .A1(n8481), .A2(n8480), .ZN(n8502) );
  NAND2_X1 U10894 ( .A1(n8502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8482) );
  XNOR2_X1 U10895 ( .A(n8482), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U10896 ( .A1(n9926), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10141), 
        .B2(n10176), .ZN(n8483) );
  NAND2_X1 U10897 ( .A1(n8484), .A2(n8483), .ZN(n10835) );
  XNOR2_X1 U10898 ( .A(n10835), .B(n8964), .ZN(n8492) );
  NAND2_X1 U10899 ( .A1(n8526), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U10900 ( .A1(n6565), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8490) );
  NOR2_X1 U10901 ( .A1(n8486), .A2(n8485), .ZN(n8506) );
  INV_X1 U10902 ( .A(n8506), .ZN(n8508) );
  NAND2_X1 U10903 ( .A1(n8486), .A2(n8485), .ZN(n8487) );
  AND2_X1 U10904 ( .A1(n8508), .A2(n8487), .ZN(n10466) );
  NAND2_X1 U10905 ( .A1(n9020), .A2(n10466), .ZN(n8489) );
  NAND2_X1 U10906 ( .A1(n9931), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8488) );
  NAND4_X1 U10907 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(n13319) );
  NAND2_X1 U10908 ( .A1(n13319), .A2(n8811), .ZN(n8493) );
  XNOR2_X1 U10909 ( .A(n8492), .B(n8493), .ZN(n10464) );
  INV_X1 U10910 ( .A(n8492), .ZN(n8495) );
  INV_X1 U10911 ( .A(n8493), .ZN(n8494) );
  NAND2_X1 U10912 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  INV_X1 U10913 ( .A(n8497), .ZN(n8498) );
  NAND2_X1 U10914 ( .A1(n8500), .A2(SI_6_), .ZN(n8501) );
  MUX2_X1 U10915 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10006), .Z(n8521) );
  XNOR2_X1 U10916 ( .A(n8521), .B(SI_7_), .ZN(n8518) );
  XNOR2_X1 U10917 ( .A(n8520), .B(n8518), .ZN(n10044) );
  NAND2_X1 U10918 ( .A1(n10044), .A2(n9894), .ZN(n8505) );
  NAND2_X1 U10919 ( .A1(n8522), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8503) );
  XNOR2_X1 U10920 ( .A(n8503), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U10921 ( .A1(n9926), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10141), 
        .B2(n10274), .ZN(n8504) );
  NAND2_X1 U10922 ( .A1(n8505), .A2(n8504), .ZN(n14796) );
  XNOR2_X1 U10923 ( .A(n14796), .B(n8410), .ZN(n8516) );
  NAND2_X1 U10924 ( .A1(n8506), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8528) );
  INV_X1 U10925 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10926 ( .A1(n8508), .A2(n8507), .ZN(n8509) );
  AND2_X1 U10927 ( .A1(n8528), .A2(n8509), .ZN(n14799) );
  NAND2_X1 U10928 ( .A1(n9020), .A2(n14799), .ZN(n8513) );
  NAND2_X1 U10929 ( .A1(n8526), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10930 ( .A1(n6565), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U10931 ( .A1(n9931), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8510) );
  NAND4_X1 U10932 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), .ZN(n13318) );
  NAND2_X1 U10933 ( .A1(n13318), .A2(n8811), .ZN(n8514) );
  XNOR2_X1 U10934 ( .A(n8516), .B(n8514), .ZN(n10909) );
  INV_X1 U10935 ( .A(n8514), .ZN(n8515) );
  AND2_X1 U10936 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  INV_X1 U10937 ( .A(n8518), .ZN(n8519) );
  MUX2_X1 U10938 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10006), .Z(n8543) );
  XNOR2_X1 U10939 ( .A(n8543), .B(SI_8_), .ZN(n8540) );
  XNOR2_X1 U10940 ( .A(n8542), .B(n8540), .ZN(n10057) );
  NAND2_X1 U10941 ( .A1(n10057), .A2(n9894), .ZN(n8525) );
  OAI21_X1 U10942 ( .B1(n8522), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8523) );
  XNOR2_X1 U10943 ( .A(n8523), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U10944 ( .A1(n9926), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10141), 
        .B2(n10276), .ZN(n8524) );
  NAND2_X1 U10945 ( .A1(n8525), .A2(n8524), .ZN(n11141) );
  XNOR2_X1 U10946 ( .A(n11141), .B(n8964), .ZN(n8534) );
  NAND2_X1 U10947 ( .A1(n8526), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10948 ( .A1(n6565), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8532) );
  INV_X1 U10949 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10950 ( .A1(n8528), .A2(n8527), .ZN(n8529) );
  AND2_X1 U10951 ( .A1(n8551), .A2(n8529), .ZN(n10984) );
  NAND2_X1 U10952 ( .A1(n9020), .A2(n10984), .ZN(n8531) );
  NAND2_X1 U10953 ( .A1(n9931), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8530) );
  NAND4_X1 U10954 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n13317) );
  NAND2_X1 U10955 ( .A1(n13317), .A2(n8811), .ZN(n8535) );
  NAND2_X1 U10956 ( .A1(n8534), .A2(n8535), .ZN(n8539) );
  INV_X1 U10957 ( .A(n8534), .ZN(n8537) );
  INV_X1 U10958 ( .A(n8535), .ZN(n8536) );
  NAND2_X1 U10959 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  AND2_X1 U10960 ( .A1(n8539), .A2(n8538), .ZN(n10879) );
  INV_X1 U10961 ( .A(n8540), .ZN(n8541) );
  NAND2_X1 U10962 ( .A1(n8542), .A2(n8541), .ZN(n8545) );
  NAND2_X1 U10963 ( .A1(n8543), .A2(SI_8_), .ZN(n8544) );
  MUX2_X1 U10964 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10006), .Z(n8566) );
  XNOR2_X1 U10965 ( .A(n8566), .B(SI_9_), .ZN(n8563) );
  XNOR2_X1 U10966 ( .A(n8565), .B(n8563), .ZN(n10061) );
  NAND2_X1 U10967 ( .A1(n10061), .A2(n9894), .ZN(n8549) );
  OR2_X1 U10968 ( .A1(n8546), .A2(n8568), .ZN(n8547) );
  XNOR2_X1 U10969 ( .A(n8547), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U10970 ( .A1(n9926), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10141), 
        .B2(n10396), .ZN(n8548) );
  NAND2_X1 U10971 ( .A1(n8549), .A2(n8548), .ZN(n11334) );
  XNOR2_X1 U10972 ( .A(n11334), .B(n8964), .ZN(n8557) );
  NAND2_X1 U10973 ( .A1(n9931), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U10974 ( .A1(n8526), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8555) );
  INV_X1 U10975 ( .A(n8572), .ZN(n8574) );
  NAND2_X1 U10976 ( .A1(n8551), .A2(n8550), .ZN(n8552) );
  AND2_X1 U10977 ( .A1(n8574), .A2(n8552), .ZN(n11333) );
  NAND2_X1 U10978 ( .A1(n9020), .A2(n11333), .ZN(n8554) );
  NAND2_X1 U10979 ( .A1(n6565), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8553) );
  NAND4_X1 U10980 ( .A1(n8556), .A2(n8555), .A3(n8554), .A4(n8553), .ZN(n13316) );
  NAND2_X1 U10981 ( .A1(n13316), .A2(n8811), .ZN(n8558) );
  NAND2_X1 U10982 ( .A1(n8557), .A2(n8558), .ZN(n8562) );
  INV_X1 U10983 ( .A(n8557), .ZN(n8560) );
  INV_X1 U10984 ( .A(n8558), .ZN(n8559) );
  NAND2_X1 U10985 ( .A1(n8560), .A2(n8559), .ZN(n8561) );
  AND2_X1 U10986 ( .A1(n8562), .A2(n8561), .ZN(n10945) );
  INV_X1 U10987 ( .A(n8563), .ZN(n8564) );
  NAND2_X1 U10988 ( .A1(n8566), .A2(SI_9_), .ZN(n8567) );
  MUX2_X1 U10989 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10006), .Z(n8588) );
  XNOR2_X1 U10990 ( .A(n8588), .B(SI_10_), .ZN(n8585) );
  XNOR2_X1 U10991 ( .A(n8587), .B(n8585), .ZN(n10077) );
  NAND2_X1 U10992 ( .A1(n10077), .A2(n9894), .ZN(n8571) );
  AND2_X1 U10993 ( .A1(n8546), .A2(n15400), .ZN(n8593) );
  OR2_X1 U10994 ( .A1(n8593), .A2(n8568), .ZN(n8569) );
  XNOR2_X1 U10995 ( .A(n8569), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U10996 ( .A1(n9926), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10141), 
        .B2(n10428), .ZN(n8570) );
  XNOR2_X1 U10997 ( .A(n11190), .B(n8964), .ZN(n8581) );
  NAND2_X1 U10998 ( .A1(n9931), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U10999 ( .A1(n8526), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8579) );
  INV_X1 U11000 ( .A(n8599), .ZN(n8600) );
  INV_X1 U11001 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11002 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  AND2_X1 U11003 ( .A1(n8600), .A2(n8575), .ZN(n11000) );
  NAND2_X1 U11004 ( .A1(n9020), .A2(n11000), .ZN(n8578) );
  NAND2_X1 U11005 ( .A1(n6565), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8577) );
  NAND4_X1 U11006 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(n13315) );
  NAND2_X1 U11007 ( .A1(n13315), .A2(n8811), .ZN(n8582) );
  XNOR2_X1 U11008 ( .A(n8581), .B(n8582), .ZN(n10998) );
  INV_X1 U11009 ( .A(n8581), .ZN(n8584) );
  INV_X1 U11010 ( .A(n8582), .ZN(n8583) );
  INV_X1 U11011 ( .A(n8585), .ZN(n8586) );
  INV_X1 U11012 ( .A(n8589), .ZN(n8590) );
  NAND2_X1 U11013 ( .A1(n8590), .A2(SI_11_), .ZN(n8591) );
  XNOR2_X1 U11014 ( .A(n8613), .B(n8612), .ZN(n10135) );
  NAND2_X1 U11015 ( .A1(n10135), .A2(n9894), .ZN(n8597) );
  NAND2_X1 U11016 ( .A1(n8593), .A2(n8592), .ZN(n8713) );
  NAND2_X1 U11017 ( .A1(n8713), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8594) );
  MUX2_X1 U11018 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8594), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n8595) );
  AOI22_X1 U11019 ( .A1(n9926), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10141), 
        .B2(n11487), .ZN(n8596) );
  XNOR2_X1 U11020 ( .A(n11389), .B(n8964), .ZN(n8606) );
  NAND2_X1 U11021 ( .A1(n9931), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U11022 ( .A1(n8526), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11023 ( .A1(n8599), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8622) );
  INV_X1 U11024 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n15250) );
  NAND2_X1 U11025 ( .A1(n8600), .A2(n15250), .ZN(n8601) );
  AND2_X1 U11026 ( .A1(n8622), .A2(n8601), .ZN(n11366) );
  NAND2_X1 U11027 ( .A1(n9020), .A2(n11366), .ZN(n8603) );
  NAND2_X1 U11028 ( .A1(n6565), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8602) );
  NAND4_X1 U11029 ( .A1(n8605), .A2(n8604), .A3(n8603), .A4(n8602), .ZN(n13314) );
  NAND2_X1 U11030 ( .A1(n13314), .A2(n8811), .ZN(n8607) );
  NAND2_X1 U11031 ( .A1(n8606), .A2(n8607), .ZN(n8611) );
  INV_X1 U11032 ( .A(n8606), .ZN(n8609) );
  INV_X1 U11033 ( .A(n8607), .ZN(n8608) );
  NAND2_X1 U11034 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U11035 ( .A1(n8611), .A2(n8610), .ZN(n11364) );
  MUX2_X1 U11036 ( .A(n10202), .B(n10204), .S(n10006), .Z(n8615) );
  NAND2_X1 U11037 ( .A1(n8615), .A2(n8614), .ZN(n8635) );
  INV_X1 U11038 ( .A(n8615), .ZN(n8616) );
  NAND2_X1 U11039 ( .A1(n8616), .A2(SI_12_), .ZN(n8617) );
  NAND2_X1 U11040 ( .A1(n10201), .A2(n9894), .ZN(n8620) );
  NAND2_X1 U11041 ( .A1(n8639), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8618) );
  XNOR2_X1 U11042 ( .A(n8618), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U11043 ( .A1(n9926), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10141), 
        .B2(n11486), .ZN(n8619) );
  XNOR2_X1 U11044 ( .A(n13667), .B(n8964), .ZN(n8628) );
  NAND2_X1 U11045 ( .A1(n8526), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11046 ( .A1(n9931), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11047 ( .A1(n8622), .A2(n8621), .ZN(n8623) );
  AND2_X1 U11048 ( .A1(n8644), .A2(n8623), .ZN(n11417) );
  NAND2_X1 U11049 ( .A1(n9020), .A2(n11417), .ZN(n8625) );
  NAND2_X1 U11050 ( .A1(n6565), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8624) );
  NAND4_X1 U11051 ( .A1(n8627), .A2(n8626), .A3(n8625), .A4(n8624), .ZN(n13313) );
  NAND2_X1 U11052 ( .A1(n13313), .A2(n8811), .ZN(n8629) );
  NAND2_X1 U11053 ( .A1(n8628), .A2(n8629), .ZN(n8633) );
  INV_X1 U11054 ( .A(n8628), .ZN(n8631) );
  INV_X1 U11055 ( .A(n8629), .ZN(n8630) );
  NAND2_X1 U11056 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  AND2_X1 U11057 ( .A1(n8633), .A2(n8632), .ZN(n11413) );
  MUX2_X1 U11058 ( .A(n10243), .B(n10245), .S(n10006), .Z(n8636) );
  INV_X1 U11059 ( .A(n8636), .ZN(n8637) );
  NAND2_X1 U11060 ( .A1(n8637), .A2(SI_13_), .ZN(n8638) );
  XNOR2_X1 U11061 ( .A(n8655), .B(n7700), .ZN(n10242) );
  NAND2_X1 U11062 ( .A1(n10242), .A2(n9894), .ZN(n8642) );
  NOR2_X1 U11063 ( .A1(n8639), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8657) );
  OR2_X1 U11064 ( .A1(n8657), .A2(n8568), .ZN(n8640) );
  XNOR2_X1 U11065 ( .A(n8640), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U11066 ( .A1(n11478), .A2(n10141), .B1(n9926), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n8641) );
  XNOR2_X1 U11067 ( .A(n11692), .B(n8964), .ZN(n8650) );
  NAND2_X1 U11068 ( .A1(n8526), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U11069 ( .A1(n6565), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8648) );
  INV_X1 U11070 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11071 ( .A1(n8644), .A2(n8643), .ZN(n8645) );
  AND2_X1 U11072 ( .A1(n8665), .A2(n8645), .ZN(n11439) );
  NAND2_X1 U11073 ( .A1(n9020), .A2(n11439), .ZN(n8647) );
  NAND2_X1 U11074 ( .A1(n9931), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8646) );
  NAND4_X1 U11075 ( .A1(n8649), .A2(n8648), .A3(n8647), .A4(n8646), .ZN(n13312) );
  NAND2_X1 U11076 ( .A1(n13312), .A2(n8811), .ZN(n8651) );
  XNOR2_X1 U11077 ( .A(n8650), .B(n8651), .ZN(n11437) );
  INV_X1 U11078 ( .A(n8650), .ZN(n8653) );
  INV_X1 U11079 ( .A(n8651), .ZN(n8652) );
  NAND2_X1 U11080 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  XNOR2_X1 U11081 ( .A(n8700), .B(SI_14_), .ZN(n8675) );
  MUX2_X1 U11082 ( .A(n15357), .B(n15428), .S(n10006), .Z(n8697) );
  XNOR2_X1 U11083 ( .A(n8675), .B(n8697), .ZN(n10368) );
  NAND2_X1 U11084 ( .A1(n10368), .A2(n9894), .ZN(n8661) );
  NAND2_X1 U11085 ( .A1(n8657), .A2(n15399), .ZN(n8680) );
  NAND2_X1 U11086 ( .A1(n8680), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8658) );
  XNOR2_X1 U11087 ( .A(n8658), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11482) );
  NOR2_X1 U11088 ( .A1(n6559), .A2(n15428), .ZN(n8659) );
  AOI21_X1 U11089 ( .B1(n11482), .B2(n10141), .A(n8659), .ZN(n8660) );
  XNOR2_X1 U11090 ( .A(n13661), .B(n8964), .ZN(n8670) );
  INV_X1 U11091 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11092 ( .A1(n9931), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U11093 ( .A1(n8526), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8662) );
  AND2_X1 U11094 ( .A1(n8663), .A2(n8662), .ZN(n8668) );
  INV_X1 U11095 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8664) );
  INV_X1 U11096 ( .A(n8686), .ZN(n8688) );
  NAND2_X1 U11097 ( .A1(n8665), .A2(n8664), .ZN(n8666) );
  NAND2_X1 U11098 ( .A1(n8688), .A2(n8666), .ZN(n11722) );
  OR2_X1 U11099 ( .A1(n11722), .A2(n8422), .ZN(n8667) );
  OAI211_X1 U11100 ( .C1(n8463), .C2(n8669), .A(n8668), .B(n8667), .ZN(n13311)
         );
  NAND2_X1 U11101 ( .A1(n13311), .A2(n6569), .ZN(n8671) );
  NAND2_X1 U11102 ( .A1(n8670), .A2(n8671), .ZN(n8685) );
  INV_X1 U11103 ( .A(n8670), .ZN(n8673) );
  INV_X1 U11104 ( .A(n8671), .ZN(n8672) );
  NAND2_X1 U11105 ( .A1(n8673), .A2(n8672), .ZN(n8684) );
  AND2_X1 U11106 ( .A1(n8685), .A2(n8684), .ZN(n11706) );
  INV_X1 U11107 ( .A(n8697), .ZN(n8701) );
  NOR2_X1 U11108 ( .A1(n8700), .A2(n10232), .ZN(n8674) );
  AOI21_X1 U11109 ( .B1(n8675), .B2(n8701), .A(n8674), .ZN(n8679) );
  MUX2_X1 U11110 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10006), .Z(n8676) );
  NAND2_X1 U11111 ( .A1(n8676), .A2(SI_15_), .ZN(n8704) );
  INV_X1 U11112 ( .A(n8676), .ZN(n8677) );
  NAND2_X1 U11113 ( .A1(n8677), .A2(n10250), .ZN(n8702) );
  AND2_X1 U11114 ( .A1(n8704), .A2(n8702), .ZN(n8678) );
  XNOR2_X1 U11115 ( .A(n8679), .B(n8678), .ZN(n10384) );
  NAND2_X1 U11116 ( .A1(n10384), .A2(n9894), .ZN(n8683) );
  OAI21_X1 U11117 ( .B1(n8680), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8681) );
  XNOR2_X1 U11118 ( .A(n8681), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U11119 ( .A1(n11616), .A2(n10141), .B1(n9926), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8682) );
  XNOR2_X1 U11120 ( .A(n13656), .B(n6567), .ZN(n11755) );
  INV_X1 U11121 ( .A(n11755), .ZN(n8694) );
  NAND3_X1 U11122 ( .A1(n11707), .A2(n8694), .A3(n8684), .ZN(n8696) );
  INV_X1 U11123 ( .A(n8685), .ZN(n8693) );
  INV_X1 U11124 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8692) );
  INV_X1 U11125 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11126 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U11127 ( .A1(n8737), .A2(n8689), .ZN(n11759) );
  OR2_X1 U11128 ( .A1(n11759), .A2(n8422), .ZN(n8691) );
  AOI22_X1 U11129 ( .A1(n8526), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n6565), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n8690) );
  OAI211_X1 U11130 ( .C1(n9900), .C2(n8692), .A(n8691), .B(n8690), .ZN(n13310)
         );
  NAND2_X1 U11131 ( .A1(n13310), .A2(n6569), .ZN(n11754) );
  AOI21_X1 U11132 ( .B1(n8694), .B2(n8693), .A(n11754), .ZN(n8695) );
  OAI21_X1 U11133 ( .B1(n10232), .B2(n8697), .A(n8704), .ZN(n8698) );
  INV_X1 U11134 ( .A(n8698), .ZN(n8699) );
  NOR2_X1 U11135 ( .A1(n8701), .A2(SI_14_), .ZN(n8705) );
  INV_X1 U11136 ( .A(n8702), .ZN(n8703) );
  AOI21_X1 U11137 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8706) );
  MUX2_X1 U11138 ( .A(n15293), .B(n10333), .S(n10006), .Z(n8707) );
  INV_X1 U11139 ( .A(n8707), .ZN(n8708) );
  NAND2_X1 U11140 ( .A1(n8708), .A2(SI_16_), .ZN(n8709) );
  MUX2_X1 U11141 ( .A(n10390), .B(n10389), .S(n10006), .Z(n8750) );
  XNOR2_X1 U11142 ( .A(n8750), .B(SI_17_), .ZN(n8711) );
  XNOR2_X1 U11143 ( .A(n8751), .B(n8711), .ZN(n10388) );
  NAND2_X1 U11144 ( .A1(n10388), .A2(n9894), .ZN(n8716) );
  OR2_X1 U11145 ( .A1(n8713), .A2(n8712), .ZN(n8733) );
  NAND2_X1 U11146 ( .A1(n8757), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8714) );
  XNOR2_X1 U11147 ( .A(n8714), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U11148 ( .A1(n9926), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n13344), 
        .B2(n10141), .ZN(n8715) );
  XNOR2_X1 U11149 ( .A(n13651), .B(n8964), .ZN(n8726) );
  INV_X1 U11150 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8718) );
  INV_X1 U11151 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8717) );
  OAI21_X1 U11152 ( .B1(n8737), .B2(n8718), .A(n8717), .ZN(n8720) );
  NAND2_X1 U11153 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n8719) );
  AND2_X1 U11154 ( .A1(n8720), .A2(n8761), .ZN(n13249) );
  NAND2_X1 U11155 ( .A1(n13249), .A2(n9020), .ZN(n8725) );
  INV_X1 U11156 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13354) );
  NAND2_X1 U11157 ( .A1(n8526), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11158 ( .A1(n6565), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8721) );
  OAI211_X1 U11159 ( .C1(n13354), .C2(n9900), .A(n8722), .B(n8721), .ZN(n8723)
         );
  INV_X1 U11160 ( .A(n8723), .ZN(n8724) );
  NAND2_X1 U11161 ( .A1(n8725), .A2(n8724), .ZN(n13308) );
  NAND2_X1 U11162 ( .A1(n13308), .A2(n8811), .ZN(n8727) );
  NAND2_X1 U11163 ( .A1(n8726), .A2(n8727), .ZN(n8749) );
  INV_X1 U11164 ( .A(n8726), .ZN(n8729) );
  INV_X1 U11165 ( .A(n8727), .ZN(n8728) );
  NAND2_X1 U11166 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U11167 ( .A1(n8749), .A2(n8730), .ZN(n13255) );
  XNOR2_X1 U11168 ( .A(n8731), .B(n8732), .ZN(n10332) );
  NAND2_X1 U11169 ( .A1(n10332), .A2(n9894), .ZN(n8736) );
  NAND2_X1 U11170 ( .A1(n8733), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8734) );
  XNOR2_X1 U11171 ( .A(n8734), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U11172 ( .A1(n9926), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10141), 
        .B2(n11611), .ZN(n8735) );
  XNOR2_X1 U11173 ( .A(n11884), .B(n8410), .ZN(n8745) );
  XNOR2_X1 U11174 ( .A(n8737), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U11175 ( .A1(n11945), .A2(n9020), .ZN(n8743) );
  INV_X1 U11176 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11177 ( .A1(n6565), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11178 ( .A1(n9931), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8738) );
  OAI211_X1 U11179 ( .C1(n8598), .C2(n8740), .A(n8739), .B(n8738), .ZN(n8741)
         );
  INV_X1 U11180 ( .A(n8741), .ZN(n8742) );
  NAND2_X1 U11181 ( .A1(n8743), .A2(n8742), .ZN(n13309) );
  AND2_X1 U11182 ( .A1(n13309), .A2(n8811), .ZN(n8746) );
  AND2_X1 U11183 ( .A1(n8745), .A2(n8746), .ZN(n11935) );
  NOR2_X1 U11184 ( .A1(n13255), .A2(n11935), .ZN(n8744) );
  INV_X1 U11185 ( .A(n8745), .ZN(n8748) );
  INV_X1 U11186 ( .A(n8746), .ZN(n8747) );
  NAND2_X1 U11187 ( .A1(n8748), .A2(n8747), .ZN(n13254) );
  MUX2_X1 U11188 ( .A(n10572), .B(n10573), .S(n10025), .Z(n8754) );
  NAND2_X1 U11189 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  NAND2_X1 U11190 ( .A1(n8774), .A2(n8756), .ZN(n10574) );
  OR2_X1 U11191 ( .A1(n10574), .A2(n8821), .ZN(n8760) );
  OAI21_X1 U11192 ( .B1(n8757), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8758) );
  XNOR2_X1 U11193 ( .A(n8758), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U11194 ( .A1(n13364), .A2(n10141), .B1(n9926), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8759) );
  XNOR2_X1 U11195 ( .A(n13645), .B(n8964), .ZN(n8768) );
  INV_X1 U11196 ( .A(n8777), .ZN(n8779) );
  NAND2_X1 U11197 ( .A1(n8761), .A2(n15363), .ZN(n8762) );
  NAND2_X1 U11198 ( .A1(n8779), .A2(n8762), .ZN(n13572) );
  OR2_X1 U11199 ( .A1(n13572), .A2(n8422), .ZN(n8767) );
  INV_X1 U11200 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n15432) );
  NAND2_X1 U11201 ( .A1(n8526), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11202 ( .A1(n9931), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8763) );
  OAI211_X1 U11203 ( .C1(n8463), .C2(n15432), .A(n8764), .B(n8763), .ZN(n8765)
         );
  INV_X1 U11204 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U11205 ( .A1(n8767), .A2(n8766), .ZN(n13541) );
  NAND2_X1 U11206 ( .A1(n13541), .A2(n6569), .ZN(n8769) );
  XNOR2_X1 U11207 ( .A(n8768), .B(n8769), .ZN(n11965) );
  INV_X1 U11208 ( .A(n8768), .ZN(n8771) );
  INV_X1 U11209 ( .A(n8769), .ZN(n8770) );
  NAND2_X1 U11210 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  MUX2_X1 U11211 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10006), .Z(n8795) );
  XNOR2_X1 U11212 ( .A(n8795), .B(SI_19_), .ZN(n8794) );
  XNOR2_X1 U11213 ( .A(n8793), .B(n8794), .ZN(n10852) );
  NAND2_X1 U11214 ( .A1(n10852), .A2(n9894), .ZN(n8776) );
  AOI22_X1 U11215 ( .A1(n9926), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10141), 
        .B2(n10646), .ZN(n8775) );
  XNOR2_X1 U11216 ( .A(n13640), .B(n8964), .ZN(n8788) );
  INV_X1 U11217 ( .A(n8803), .ZN(n8781) );
  INV_X1 U11218 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11219 ( .A1(n8779), .A2(n8778), .ZN(n8780) );
  NAND2_X1 U11220 ( .A1(n13548), .A2(n9020), .ZN(n8787) );
  INV_X1 U11221 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11222 ( .A1(n6565), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U11223 ( .A1(n8526), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8782) );
  OAI211_X1 U11224 ( .C1(n9900), .C2(n8784), .A(n8783), .B(n8782), .ZN(n8785)
         );
  INV_X1 U11225 ( .A(n8785), .ZN(n8786) );
  NAND2_X1 U11226 ( .A1(n8787), .A2(n8786), .ZN(n13307) );
  NAND2_X1 U11227 ( .A1(n13307), .A2(n6569), .ZN(n8789) );
  NAND2_X1 U11228 ( .A1(n8788), .A2(n8789), .ZN(n13225) );
  INV_X1 U11229 ( .A(n8788), .ZN(n8791) );
  INV_X1 U11230 ( .A(n8789), .ZN(n8790) );
  NAND2_X1 U11231 ( .A1(n8791), .A2(n8790), .ZN(n13224) );
  INV_X1 U11232 ( .A(n8795), .ZN(n8796) );
  MUX2_X1 U11233 ( .A(n11174), .B(n11177), .S(n10006), .Z(n8799) );
  NAND2_X1 U11234 ( .A1(n8798), .A2(n8799), .ZN(n8800) );
  NAND2_X1 U11235 ( .A1(n8815), .A2(n8800), .ZN(n11175) );
  OR2_X1 U11236 ( .A1(n11175), .A2(n8821), .ZN(n8802) );
  NAND2_X1 U11237 ( .A1(n9926), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8801) );
  XNOR2_X1 U11238 ( .A(n13635), .B(n8964), .ZN(n8813) );
  OR2_X1 U11239 ( .A1(n8803), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8804) );
  AND2_X1 U11240 ( .A1(n8824), .A2(n8804), .ZN(n13528) );
  NAND2_X1 U11241 ( .A1(n13528), .A2(n9020), .ZN(n8810) );
  INV_X1 U11242 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U11243 ( .A1(n9931), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U11244 ( .A1(n6565), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8805) );
  OAI211_X1 U11245 ( .C1(n8598), .C2(n8807), .A(n8806), .B(n8805), .ZN(n8808)
         );
  INV_X1 U11246 ( .A(n8808), .ZN(n8809) );
  NAND2_X1 U11247 ( .A1(n8810), .A2(n8809), .ZN(n13539) );
  NAND2_X1 U11248 ( .A1(n13539), .A2(n6569), .ZN(n8812) );
  XNOR2_X1 U11249 ( .A(n8813), .B(n8812), .ZN(n13271) );
  MUX2_X1 U11250 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10025), .Z(n8816) );
  NAND2_X1 U11251 ( .A1(n8816), .A2(SI_21_), .ZN(n8851) );
  OAI21_X1 U11252 ( .B1(SI_21_), .B2(n8816), .A(n8851), .ZN(n8817) );
  INV_X1 U11253 ( .A(n8817), .ZN(n8818) );
  OR2_X1 U11254 ( .A1(n8819), .A2(n8818), .ZN(n8820) );
  NAND2_X1 U11255 ( .A1(n8852), .A2(n8820), .ZN(n11359) );
  OR2_X1 U11256 ( .A1(n11359), .A2(n8821), .ZN(n8823) );
  NAND2_X1 U11257 ( .A1(n9926), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8822) );
  XNOR2_X1 U11258 ( .A(n13629), .B(n8410), .ZN(n8835) );
  INV_X1 U11259 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13235) );
  NAND2_X1 U11260 ( .A1(n8824), .A2(n13235), .ZN(n8826) );
  INV_X1 U11261 ( .A(n8840), .ZN(n8825) );
  NAND2_X1 U11262 ( .A1(n8826), .A2(n8825), .ZN(n13505) );
  OR2_X1 U11263 ( .A1(n13505), .A2(n8422), .ZN(n8832) );
  INV_X1 U11264 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11265 ( .A1(n6565), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U11266 ( .A1(n8526), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8827) );
  OAI211_X1 U11267 ( .C1(n9900), .C2(n8829), .A(n8828), .B(n8827), .ZN(n8830)
         );
  INV_X1 U11268 ( .A(n8830), .ZN(n8831) );
  NAND2_X1 U11269 ( .A1(n8832), .A2(n8831), .ZN(n13485) );
  NAND2_X1 U11270 ( .A1(n13485), .A2(n6569), .ZN(n8833) );
  XNOR2_X1 U11271 ( .A(n8835), .B(n8833), .ZN(n13233) );
  INV_X1 U11272 ( .A(n8833), .ZN(n8834) );
  NAND2_X1 U11273 ( .A1(n8835), .A2(n8834), .ZN(n8836) );
  NAND2_X1 U11274 ( .A1(n8852), .A2(n8851), .ZN(n8837) );
  MUX2_X1 U11275 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10006), .Z(n8853) );
  XNOR2_X1 U11276 ( .A(n9556), .B(n8853), .ZN(n12068) );
  NAND2_X1 U11277 ( .A1(n12068), .A2(n9894), .ZN(n8839) );
  NAND2_X1 U11278 ( .A1(n9926), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8838) );
  XNOR2_X1 U11279 ( .A(n13621), .B(n8964), .ZN(n8846) );
  NAND2_X1 U11280 ( .A1(n9931), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11281 ( .A1(n8380), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8844) );
  NAND2_X1 U11282 ( .A1(n8840), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8862) );
  OAI21_X1 U11283 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n8840), .A(n8862), .ZN(
        n8841) );
  INV_X1 U11284 ( .A(n8841), .ZN(n13491) );
  NAND2_X1 U11285 ( .A1(n9020), .A2(n13491), .ZN(n8843) );
  NAND2_X1 U11286 ( .A1(n6565), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8842) );
  NAND4_X1 U11287 ( .A1(n8845), .A2(n8844), .A3(n8843), .A4(n8842), .ZN(n13502) );
  AND2_X1 U11288 ( .A1(n13502), .A2(n6569), .ZN(n13280) );
  INV_X1 U11289 ( .A(n8846), .ZN(n8847) );
  NAND2_X1 U11290 ( .A1(n8848), .A2(n8847), .ZN(n8849) );
  NAND2_X1 U11291 ( .A1(n8853), .A2(SI_22_), .ZN(n8850) );
  INV_X1 U11292 ( .A(n8853), .ZN(n8855) );
  INV_X1 U11293 ( .A(SI_22_), .ZN(n8854) );
  NAND2_X1 U11294 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  MUX2_X1 U11295 ( .A(n11667), .B(n15238), .S(n10006), .Z(n8857) );
  NAND2_X1 U11296 ( .A1(n8873), .A2(n8874), .ZN(n8859) );
  NAND2_X1 U11297 ( .A1(n11669), .A2(n9894), .ZN(n8861) );
  NAND2_X1 U11298 ( .A1(n9926), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8860) );
  XNOR2_X1 U11299 ( .A(n13614), .B(n8964), .ZN(n8868) );
  NAND2_X1 U11300 ( .A1(n9931), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U11301 ( .A1(n8380), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8866) );
  INV_X1 U11302 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8863) );
  AOI21_X1 U11303 ( .B1(n8863), .B2(n8862), .A(n8882), .ZN(n13473) );
  NAND2_X1 U11304 ( .A1(n9020), .A2(n13473), .ZN(n8865) );
  NAND2_X1 U11305 ( .A1(n6565), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8864) );
  NAND4_X1 U11306 ( .A1(n8867), .A2(n8866), .A3(n8865), .A4(n8864), .ZN(n13484) );
  AND2_X1 U11307 ( .A1(n13484), .A2(n6569), .ZN(n13218) );
  INV_X1 U11308 ( .A(n8868), .ZN(n8869) );
  INV_X1 U11309 ( .A(SI_23_), .ZN(n8872) );
  MUX2_X1 U11310 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10006), .Z(n8875) );
  NAND2_X1 U11311 ( .A1(n8875), .A2(SI_24_), .ZN(n8895) );
  OAI21_X1 U11312 ( .B1(SI_24_), .B2(n8875), .A(n8895), .ZN(n8877) );
  NAND2_X1 U11313 ( .A1(n8878), .A2(n8877), .ZN(n8879) );
  AND2_X1 U11314 ( .A1(n8894), .A2(n8879), .ZN(n11715) );
  NAND2_X1 U11315 ( .A1(n11715), .A2(n9894), .ZN(n8881) );
  NAND2_X1 U11316 ( .A1(n9926), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8880) );
  XNOR2_X1 U11317 ( .A(n13607), .B(n8410), .ZN(n8888) );
  NAND2_X1 U11318 ( .A1(n9931), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U11319 ( .A1(n8380), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U11320 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n8882), .ZN(n8900) );
  OAI21_X1 U11321 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8882), .A(n8900), .ZN(
        n8883) );
  INV_X1 U11322 ( .A(n8883), .ZN(n13463) );
  NAND2_X1 U11323 ( .A1(n9020), .A2(n13463), .ZN(n8885) );
  NAND2_X1 U11324 ( .A1(n6565), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8884) );
  NAND4_X1 U11325 ( .A1(n8887), .A2(n8886), .A3(n8885), .A4(n8884), .ZN(n13471) );
  AND2_X1 U11326 ( .A1(n13471), .A2(n6569), .ZN(n8889) );
  NAND2_X1 U11327 ( .A1(n8888), .A2(n8889), .ZN(n8893) );
  INV_X1 U11328 ( .A(n8888), .ZN(n8891) );
  INV_X1 U11329 ( .A(n8889), .ZN(n8890) );
  NAND2_X1 U11330 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  AND2_X1 U11331 ( .A1(n8893), .A2(n8892), .ZN(n13263) );
  MUX2_X1 U11332 ( .A(n8896), .B(n15247), .S(n10006), .Z(n8912) );
  NAND2_X1 U11333 ( .A1(n11895), .A2(n9894), .ZN(n8898) );
  NAND2_X1 U11334 ( .A1(n9926), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8897) );
  XNOR2_X1 U11335 ( .A(n13603), .B(n8410), .ZN(n8906) );
  NAND2_X1 U11336 ( .A1(n9931), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U11337 ( .A1(n8526), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8904) );
  INV_X1 U11338 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8901) );
  INV_X1 U11339 ( .A(n8900), .ZN(n8899) );
  NAND2_X1 U11340 ( .A1(n8899), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8917) );
  INV_X1 U11341 ( .A(n8917), .ZN(n8918) );
  AOI21_X1 U11342 ( .B1(n8901), .B2(n8900), .A(n8918), .ZN(n13442) );
  NAND2_X1 U11343 ( .A1(n9020), .A2(n13442), .ZN(n8903) );
  NAND2_X1 U11344 ( .A1(n6565), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8902) );
  NAND4_X1 U11345 ( .A1(n8905), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(n13456) );
  AND2_X1 U11346 ( .A1(n13456), .A2(n6569), .ZN(n8907) );
  NAND2_X1 U11347 ( .A1(n8906), .A2(n8907), .ZN(n8911) );
  INV_X1 U11348 ( .A(n8906), .ZN(n8909) );
  INV_X1 U11349 ( .A(n8907), .ZN(n8908) );
  NAND2_X1 U11350 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  AND2_X1 U11351 ( .A1(n8911), .A2(n8910), .ZN(n13243) );
  INV_X1 U11352 ( .A(SI_25_), .ZN(n11421) );
  NAND2_X1 U11353 ( .A1(n8912), .A2(n11421), .ZN(n8913) );
  MUX2_X1 U11354 ( .A(n11974), .B(n11972), .S(n10006), .Z(n8929) );
  XNOR2_X1 U11355 ( .A(n8929), .B(SI_26_), .ZN(n8914) );
  XNOR2_X1 U11356 ( .A(n8928), .B(n8914), .ZN(n11971) );
  NAND2_X1 U11357 ( .A1(n11971), .A2(n9894), .ZN(n8916) );
  NAND2_X1 U11358 ( .A1(n9926), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8915) );
  XNOR2_X1 U11359 ( .A(n13598), .B(n8964), .ZN(n8925) );
  NAND2_X1 U11360 ( .A1(n9931), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U11361 ( .A1(n8380), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8922) );
  INV_X1 U11362 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13293) );
  NAND2_X1 U11363 ( .A1(n13293), .A2(n8917), .ZN(n8919) );
  NAND2_X1 U11364 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8918), .ZN(n8941) );
  AND2_X1 U11365 ( .A1(n8919), .A2(n8941), .ZN(n13434) );
  NAND2_X1 U11366 ( .A1(n9020), .A2(n13434), .ZN(n8921) );
  NAND2_X1 U11367 ( .A1(n6565), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8920) );
  NAND4_X1 U11368 ( .A1(n8923), .A2(n8922), .A3(n8921), .A4(n8920), .ZN(n13448) );
  NAND2_X1 U11369 ( .A1(n13448), .A2(n6569), .ZN(n8924) );
  XNOR2_X1 U11370 ( .A(n8925), .B(n8924), .ZN(n13292) );
  NAND2_X1 U11371 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  INV_X1 U11372 ( .A(n8928), .ZN(n8927) );
  INV_X1 U11373 ( .A(SI_26_), .ZN(n11626) );
  NAND2_X1 U11374 ( .A1(n8928), .A2(n11626), .ZN(n8931) );
  INV_X1 U11375 ( .A(n8929), .ZN(n8930) );
  NAND2_X1 U11376 ( .A1(n8931), .A2(n8930), .ZN(n8932) );
  MUX2_X1 U11377 ( .A(n14367), .B(n12051), .S(n10006), .Z(n9003) );
  XNOR2_X1 U11378 ( .A(n9003), .B(SI_27_), .ZN(n8934) );
  NAND2_X1 U11379 ( .A1(n12049), .A2(n9894), .ZN(n8938) );
  NAND2_X1 U11380 ( .A1(n9926), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8937) );
  XNOR2_X1 U11381 ( .A(n13591), .B(n6567), .ZN(n8947) );
  NAND2_X1 U11382 ( .A1(n9931), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U11383 ( .A1(n8380), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8945) );
  INV_X1 U11384 ( .A(n8941), .ZN(n8939) );
  INV_X1 U11385 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U11386 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  NAND2_X1 U11387 ( .A1(n9020), .A2(n13419), .ZN(n8944) );
  NAND2_X1 U11388 ( .A1(n6565), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8943) );
  NAND4_X1 U11389 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n13428) );
  AND2_X1 U11390 ( .A1(n13428), .A2(n6569), .ZN(n8948) );
  NAND2_X1 U11391 ( .A1(n8947), .A2(n8948), .ZN(n8953) );
  INV_X1 U11392 ( .A(n8947), .ZN(n8950) );
  INV_X1 U11393 ( .A(n8948), .ZN(n8949) );
  NAND2_X1 U11394 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  NAND2_X1 U11395 ( .A1(n8953), .A2(n8951), .ZN(n13209) );
  INV_X1 U11396 ( .A(n13209), .ZN(n8952) );
  NAND2_X1 U11397 ( .A1(n9931), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11398 ( .A1(n8380), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8961) );
  INV_X1 U11399 ( .A(n12041), .ZN(n8958) );
  INV_X1 U11400 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11401 ( .A1(n8956), .A2(n8955), .ZN(n8957) );
  NAND2_X1 U11402 ( .A1(n9020), .A2(n13407), .ZN(n8960) );
  NAND2_X1 U11403 ( .A1(n6565), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8959) );
  NAND4_X1 U11404 ( .A1(n8962), .A2(n8961), .A3(n8960), .A4(n8959), .ZN(n13414) );
  NAND2_X1 U11405 ( .A1(n13414), .A2(n8811), .ZN(n8963) );
  XNOR2_X1 U11406 ( .A(n8964), .B(n8963), .ZN(n8965) );
  XNOR2_X1 U11407 ( .A(n8966), .B(n8965), .ZN(n9010) );
  NAND2_X1 U11408 ( .A1(n8967), .A2(n8980), .ZN(n8976) );
  OAI21_X1 U11409 ( .B1(n8976), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U11410 ( .A1(n8973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8972) );
  MUX2_X1 U11411 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8972), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8975) );
  NAND2_X1 U11412 ( .A1(n8976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11413 ( .A1(n8979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8981) );
  INV_X1 U11414 ( .A(P2_B_REG_SCAN_IN), .ZN(n15383) );
  XOR2_X1 U11415 ( .A(n11742), .B(n15383), .Z(n8982) );
  NAND2_X1 U11416 ( .A1(n11924), .A2(n8982), .ZN(n8984) );
  INV_X1 U11417 ( .A(n11973), .ZN(n8983) );
  INV_X1 U11418 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U11419 ( .A1(n14810), .A2(n14812), .ZN(n8986) );
  AND2_X1 U11420 ( .A1(n11742), .A2(n11973), .ZN(n14813) );
  INV_X1 U11421 ( .A(n14813), .ZN(n8985) );
  NOR4_X1 U11422 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8995) );
  INV_X1 U11423 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15397) );
  INV_X1 U11424 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15341) );
  INV_X1 U11425 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15371) );
  INV_X1 U11426 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15304) );
  NAND4_X1 U11427 ( .A1(n15397), .A2(n15341), .A3(n15371), .A4(n15304), .ZN(
        n8992) );
  NOR4_X1 U11428 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8990) );
  NOR4_X1 U11429 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8989) );
  NOR4_X1 U11430 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8988) );
  NOR4_X1 U11431 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8987) );
  NAND4_X1 U11432 ( .A1(n8990), .A2(n8989), .A3(n8988), .A4(n8987), .ZN(n8991)
         );
  NOR4_X1 U11433 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8992), .A4(n8991), .ZN(n8994) );
  NOR4_X1 U11434 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8993) );
  NAND3_X1 U11435 ( .A1(n8995), .A2(n8994), .A3(n8993), .ZN(n8996) );
  NAND2_X1 U11436 ( .A1(n8996), .A2(n14810), .ZN(n10605) );
  INV_X1 U11437 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14816) );
  NAND2_X1 U11438 ( .A1(n14810), .A2(n14816), .ZN(n8998) );
  NAND2_X1 U11439 ( .A1(n11924), .A2(n11973), .ZN(n8997) );
  NAND2_X1 U11440 ( .A1(n8998), .A2(n8997), .ZN(n14817) );
  INV_X1 U11441 ( .A(n14817), .ZN(n8999) );
  AND2_X1 U11442 ( .A1(n10605), .A2(n8999), .ZN(n10641) );
  INV_X1 U11443 ( .A(n10641), .ZN(n9000) );
  OR2_X1 U11444 ( .A1(n10642), .A2(n9000), .ZN(n9015) );
  OR2_X1 U11445 ( .A1(n14815), .A2(n9015), .ZN(n9011) );
  NAND2_X1 U11446 ( .A1(n11176), .A2(n13373), .ZN(n9990) );
  NAND2_X1 U11447 ( .A1(n10647), .A2(n9990), .ZN(n14872) );
  INV_X1 U11448 ( .A(n10143), .ZN(n9001) );
  NAND2_X1 U11449 ( .A1(n14872), .A2(n9001), .ZN(n9002) );
  INV_X1 U11450 ( .A(n9003), .ZN(n9004) );
  NAND2_X1 U11451 ( .A1(n9004), .A2(SI_27_), .ZN(n9005) );
  MUX2_X1 U11452 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10025), .Z(n9624) );
  XNOR2_X1 U11453 ( .A(n9624), .B(SI_28_), .ZN(n9627) );
  NAND2_X1 U11454 ( .A1(n12048), .A2(n9894), .ZN(n9008) );
  NAND2_X1 U11455 ( .A1(n9926), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11456 ( .A1(n10647), .A2(n9988), .ZN(n10712) );
  INV_X1 U11457 ( .A(n9993), .ZN(n12069) );
  NAND2_X1 U11458 ( .A1(n12069), .A2(n10646), .ZN(n9735) );
  INV_X1 U11459 ( .A(n8377), .ZN(n11360) );
  INV_X1 U11460 ( .A(n9012), .ZN(n9013) );
  AND2_X2 U11461 ( .A1(n10143), .A2(n9013), .ZN(n13540) );
  NOR2_X2 U11462 ( .A1(n13252), .A2(n13522), .ZN(n13282) );
  INV_X1 U11463 ( .A(n10603), .ZN(n9014) );
  NAND2_X1 U11464 ( .A1(n9015), .A2(n9014), .ZN(n9016) );
  AND2_X1 U11465 ( .A1(n9990), .A2(n8377), .ZN(n9929) );
  NAND2_X1 U11466 ( .A1(n9929), .A2(n9993), .ZN(n10640) );
  NAND2_X1 U11467 ( .A1(n9016), .A2(n10640), .ZN(n10581) );
  INV_X1 U11468 ( .A(n9017), .ZN(n9018) );
  AOI22_X1 U11469 ( .A1(n13282), .A2(n13428), .B1(n13283), .B2(n13407), .ZN(
        n9026) );
  NAND2_X1 U11470 ( .A1(n10143), .A2(n9012), .ZN(n13524) );
  NAND2_X1 U11471 ( .A1(n9931), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U11472 ( .A1(n8380), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11473 ( .A1(n9020), .A2(n12041), .ZN(n9022) );
  NAND2_X1 U11474 ( .A1(n6565), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9021) );
  NAND4_X1 U11475 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(n13392) );
  AOI22_X1 U11476 ( .A1(n13284), .A2(n13392), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9025) );
  INV_X1 U11477 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15321) );
  INV_X1 U11478 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14768) );
  INV_X1 U11479 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14544) );
  XNOR2_X1 U11480 ( .A(n9028), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n9041) );
  NOR2_X1 U11481 ( .A1(n9031), .A2(n14954), .ZN(n9032) );
  INV_X1 U11482 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9033) );
  NOR2_X1 U11483 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n9033), .ZN(n9034) );
  NOR2_X1 U11484 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9035), .ZN(n9037) );
  XNOR2_X1 U11485 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9035), .ZN(n9064) );
  INV_X1 U11486 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13940) );
  XOR2_X1 U11487 ( .A(n15016), .B(n10122), .Z(n9069) );
  XOR2_X1 U11488 ( .A(n9070), .B(n9069), .Z(n9068) );
  NAND2_X1 U11489 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9039), .ZN(n9054) );
  XNOR2_X1 U11490 ( .A(n9040), .B(n9041), .ZN(n9048) );
  INV_X1 U11491 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15309) );
  XNOR2_X1 U11492 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n9042) );
  XOR2_X1 U11493 ( .A(n9043), .B(n9042), .Z(n9044) );
  OR2_X1 U11494 ( .A1(n15309), .A2(n9044), .ZN(n9046) );
  AOI21_X1 U11495 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14899), .A(n9043), .ZN(
        n15465) );
  INV_X1 U11496 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15464) );
  NOR2_X1 U11497 ( .A1(n15465), .A2(n15464), .ZN(n15473) );
  NAND2_X1 U11498 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  NOR2_X1 U11499 ( .A1(n9048), .A2(n9047), .ZN(n14378) );
  NOR2_X1 U11500 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n14377), .ZN(n9049) );
  XNOR2_X1 U11501 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9050), .ZN(n15470) );
  INV_X1 U11502 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9051) );
  NAND2_X1 U11503 ( .A1(n15469), .A2(n15470), .ZN(n15468) );
  NAND2_X1 U11504 ( .A1(n15462), .A2(n15461), .ZN(n9053) );
  NAND2_X1 U11505 ( .A1(n9054), .A2(n9053), .ZN(n9057) );
  XNOR2_X1 U11506 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9055), .ZN(n9056) );
  NOR2_X1 U11507 ( .A1(n9057), .A2(n9056), .ZN(n9059) );
  XNOR2_X1 U11508 ( .A(n9057), .B(n9056), .ZN(n15463) );
  NOR2_X1 U11509 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15463), .ZN(n9058) );
  NAND2_X1 U11510 ( .A1(n9060), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9063) );
  XNOR2_X1 U11511 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n9062) );
  XOR2_X1 U11512 ( .A(n9062), .B(n9061), .Z(n14391) );
  NAND2_X1 U11513 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9065), .ZN(n9066) );
  XNOR2_X1 U11514 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9064), .ZN(n15467) );
  XNOR2_X1 U11515 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9073) );
  XNOR2_X1 U11516 ( .A(n9073), .B(n9072), .ZN(n14395) );
  NAND2_X1 U11517 ( .A1(n10215), .A2(n9074), .ZN(n9080) );
  NAND2_X1 U11518 ( .A1(n9078), .A2(n9080), .ZN(n9075) );
  XNOR2_X1 U11519 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n9075), .ZN(n9077) );
  XNOR2_X1 U11520 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .ZN(n9081) );
  NAND2_X1 U11521 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n9078), .ZN(n9079) );
  XNOR2_X1 U11522 ( .A(n9081), .B(n9084), .ZN(n14543) );
  NAND2_X1 U11523 ( .A1(n14542), .A2(n14543), .ZN(n9082) );
  NOR2_X1 U11524 ( .A1(n14542), .A2(n14543), .ZN(n14541) );
  INV_X1 U11525 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15266) );
  NAND2_X1 U11526 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n15266), .ZN(n9083) );
  XOR2_X1 U11527 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n9085) );
  XNOR2_X1 U11528 ( .A(n9088), .B(n9085), .ZN(n14548) );
  NAND2_X1 U11529 ( .A1(n14547), .A2(n14548), .ZN(n9086) );
  XNOR2_X1 U11530 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9089) );
  AND2_X1 U11531 ( .A1(n15353), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n9087) );
  XOR2_X1 U11532 ( .A(n9089), .B(n9092), .Z(n9090) );
  INV_X1 U11533 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9095) );
  INV_X1 U11534 ( .A(n9092), .ZN(n9094) );
  AND2_X1 U11535 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n9095), .ZN(n9093) );
  XOR2_X1 U11536 ( .A(P1_ADDR_REG_14__SCAN_IN), .B(P3_ADDR_REG_14__SCAN_IN), 
        .Z(n9096) );
  XOR2_X1 U11537 ( .A(n9101), .B(n9096), .Z(n9097) );
  NOR2_X1 U11538 ( .A1(n9098), .A2(n9097), .ZN(n14554) );
  INV_X1 U11539 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14582) );
  NOR2_X1 U11540 ( .A1(n14582), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n9105) );
  AOI21_X1 U11541 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n14582), .A(n9105), .ZN(
        n9103) );
  INV_X1 U11542 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15210) );
  INV_X1 U11543 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9100) );
  NOR2_X1 U11544 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n9100), .ZN(n9102) );
  XOR2_X1 U11545 ( .A(n9103), .B(n9104), .Z(n14557) );
  XNOR2_X1 U11546 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9106) );
  INV_X1 U11547 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15281) );
  OAI22_X1 U11548 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15281), .B1(n9105), 
        .B2(n9104), .ZN(n9111) );
  XOR2_X1 U11549 ( .A(n9106), .B(n9111), .Z(n9107) );
  INV_X1 U11550 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9110) );
  AND2_X1 U11551 ( .A1(n9110), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n9112) );
  OAI22_X1 U11552 ( .A1(n9112), .A2(n9111), .B1(P3_ADDR_REG_16__SCAN_IN), .B2(
        n9110), .ZN(n9116) );
  XOR2_X1 U11553 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9116), .Z(n9117) );
  XNOR2_X1 U11554 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n9117), .ZN(n9114) );
  NOR2_X1 U11555 ( .A1(n9113), .A2(n9114), .ZN(n14412) );
  NOR2_X1 U11556 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n14411), .ZN(n9115) );
  NOR2_X1 U11557 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n9116), .ZN(n9119) );
  AND2_X1 U11558 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9117), .ZN(n9118) );
  NOR2_X1 U11559 ( .A1(n9119), .A2(n9118), .ZN(n9123) );
  XOR2_X1 U11560 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n9122) );
  XNOR2_X1 U11561 ( .A(n9123), .B(n9122), .ZN(n9120) );
  INV_X1 U11562 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14597) );
  NOR2_X1 U11563 ( .A1(n9123), .A2(n9122), .ZN(n9124) );
  AOI21_X1 U11564 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14597), .A(n9124), .ZN(
        n9126) );
  XNOR2_X1 U11565 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9125) );
  XNOR2_X1 U11566 ( .A(n9126), .B(n9125), .ZN(n9127) );
  INV_X1 U11567 ( .A(n9128), .ZN(n12758) );
  NAND2_X1 U11568 ( .A1(n12630), .A2(n10577), .ZN(n9130) );
  INV_X2 U11569 ( .A(n9139), .ZN(n12352) );
  XNOR2_X1 U11570 ( .A(n13084), .B(n12352), .ZN(n12482) );
  NOR2_X1 U11571 ( .A1(n12482), .A2(n12913), .ZN(n12477) );
  AOI21_X1 U11572 ( .B1(n12482), .B2(n12913), .A(n12477), .ZN(n9218) );
  XNOR2_X1 U11573 ( .A(n6568), .B(n15089), .ZN(n9141) );
  NAND2_X1 U11574 ( .A1(n12352), .A2(n15065), .ZN(n9136) );
  NAND2_X1 U11575 ( .A1(n12782), .A2(n9133), .ZN(n9135) );
  NAND2_X1 U11576 ( .A1(n9138), .A2(n7838), .ZN(n9134) );
  OAI21_X1 U11577 ( .B1(n9139), .B2(n9135), .A(n9134), .ZN(n12351) );
  XNOR2_X1 U11578 ( .A(n9139), .B(n15043), .ZN(n9140) );
  XNOR2_X1 U11579 ( .A(n9140), .B(n15063), .ZN(n10336) );
  XNOR2_X1 U11580 ( .A(n9141), .B(n12781), .ZN(n10001) );
  XNOR2_X1 U11581 ( .A(n12474), .B(n9142), .ZN(n9143) );
  XOR2_X1 U11582 ( .A(n12780), .B(n9143), .Z(n10476) );
  NAND2_X1 U11583 ( .A1(n10475), .A2(n10476), .ZN(n10474) );
  INV_X1 U11584 ( .A(n9143), .ZN(n9145) );
  XNOR2_X1 U11585 ( .A(n12474), .B(n15097), .ZN(n9147) );
  XOR2_X1 U11586 ( .A(n12779), .B(n9147), .Z(n10562) );
  INV_X1 U11587 ( .A(n9147), .ZN(n9149) );
  NAND2_X1 U11588 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  INV_X4 U11589 ( .A(n12352), .ZN(n12474) );
  XNOR2_X1 U11590 ( .A(n12474), .B(n15104), .ZN(n9151) );
  XOR2_X1 U11591 ( .A(n12778), .B(n9151), .Z(n10993) );
  INV_X1 U11592 ( .A(n9151), .ZN(n9152) );
  XNOR2_X1 U11593 ( .A(n12474), .B(n12659), .ZN(n10887) );
  INV_X1 U11594 ( .A(n10887), .ZN(n9153) );
  NAND2_X1 U11595 ( .A1(n9153), .A2(n12777), .ZN(n9154) );
  NAND2_X1 U11596 ( .A1(n10886), .A2(n9154), .ZN(n10956) );
  XNOR2_X1 U11597 ( .A(n12474), .B(n10961), .ZN(n9155) );
  XNOR2_X1 U11598 ( .A(n9155), .B(n12776), .ZN(n10955) );
  NAND2_X1 U11599 ( .A1(n10956), .A2(n10955), .ZN(n10954) );
  INV_X1 U11600 ( .A(n9155), .ZN(n9156) );
  NAND2_X1 U11601 ( .A1(n9156), .A2(n12776), .ZN(n9157) );
  XNOR2_X1 U11602 ( .A(n12474), .B(n15120), .ZN(n9158) );
  XNOR2_X1 U11603 ( .A(n9158), .B(n12775), .ZN(n11196) );
  INV_X1 U11604 ( .A(n9158), .ZN(n9160) );
  XNOR2_X1 U11605 ( .A(n12474), .B(n11353), .ZN(n9162) );
  XOR2_X1 U11606 ( .A(n12774), .B(n9162), .Z(n11530) );
  INV_X1 U11607 ( .A(n9162), .ZN(n9163) );
  XOR2_X1 U11608 ( .A(n11451), .B(n12474), .Z(n9164) );
  OR2_X2 U11609 ( .A1(n9165), .A2(n9164), .ZN(n11630) );
  NAND2_X1 U11610 ( .A1(n9165), .A2(n9164), .ZN(n11629) );
  INV_X1 U11611 ( .A(n11629), .ZN(n9166) );
  XNOR2_X1 U11612 ( .A(n12474), .B(n14492), .ZN(n9169) );
  XOR2_X1 U11613 ( .A(n12772), .B(n9169), .Z(n11731) );
  XNOR2_X1 U11614 ( .A(n14481), .B(n12474), .ZN(n9174) );
  XOR2_X1 U11615 ( .A(n12770), .B(n9174), .Z(n14425) );
  INV_X1 U11616 ( .A(n14425), .ZN(n9167) );
  XOR2_X1 U11617 ( .A(n12474), .B(n14490), .Z(n11766) );
  NAND2_X1 U11618 ( .A1(n11766), .A2(n12771), .ZN(n14423) );
  AND2_X1 U11619 ( .A1(n9167), .A2(n14423), .ZN(n14422) );
  AND2_X1 U11620 ( .A1(n11731), .A2(n14422), .ZN(n9168) );
  INV_X1 U11621 ( .A(n14422), .ZN(n9173) );
  NOR2_X1 U11622 ( .A1(n11766), .A2(n12771), .ZN(n14420) );
  INV_X1 U11623 ( .A(n14420), .ZN(n9171) );
  INV_X1 U11624 ( .A(n9169), .ZN(n9170) );
  NAND2_X1 U11625 ( .A1(n9170), .A2(n11803), .ZN(n11764) );
  AND2_X1 U11626 ( .A1(n9171), .A2(n11764), .ZN(n9172) );
  INV_X1 U11627 ( .A(n9174), .ZN(n9175) );
  XNOR2_X1 U11628 ( .A(n13137), .B(n12474), .ZN(n9179) );
  XOR2_X1 U11629 ( .A(n14415), .B(n9179), .Z(n12075) );
  INV_X1 U11630 ( .A(n12075), .ZN(n9178) );
  INV_X1 U11631 ( .A(n9179), .ZN(n9180) );
  NAND2_X1 U11632 ( .A1(n9180), .A2(n14415), .ZN(n9181) );
  XNOR2_X1 U11633 ( .A(n14442), .B(n12474), .ZN(n9182) );
  XOR2_X1 U11634 ( .A(n12769), .B(n9182), .Z(n14435) );
  XNOR2_X1 U11635 ( .A(n12521), .B(n12474), .ZN(n9184) );
  XOR2_X1 U11636 ( .A(n13050), .B(n9184), .Z(n12522) );
  XNOR2_X1 U11637 ( .A(n13056), .B(n12474), .ZN(n9185) );
  XNOR2_X1 U11638 ( .A(n9185), .B(n13035), .ZN(n12557) );
  INV_X1 U11639 ( .A(n9185), .ZN(n9186) );
  NAND2_X1 U11640 ( .A1(n9186), .A2(n13035), .ZN(n9187) );
  XNOR2_X1 U11641 ( .A(n13184), .B(n12474), .ZN(n9189) );
  XOR2_X1 U11642 ( .A(n13049), .B(n9189), .Z(n12494) );
  NAND2_X1 U11643 ( .A1(n12495), .A2(n12494), .ZN(n9191) );
  NAND2_X1 U11644 ( .A1(n9189), .A2(n13049), .ZN(n9190) );
  XNOR2_X1 U11645 ( .A(n13113), .B(n12474), .ZN(n9192) );
  XNOR2_X1 U11646 ( .A(n9192), .B(n13036), .ZN(n12541) );
  INV_X1 U11647 ( .A(n9192), .ZN(n9193) );
  NAND2_X1 U11648 ( .A1(n9193), .A2(n13036), .ZN(n9194) );
  XNOR2_X1 U11649 ( .A(n13006), .B(n6568), .ZN(n9195) );
  NAND2_X1 U11650 ( .A1(n9195), .A2(n13021), .ZN(n9196) );
  OAI21_X1 U11651 ( .B1(n9195), .B2(n13021), .A(n9196), .ZN(n12502) );
  XNOR2_X1 U11652 ( .A(n9197), .B(n12474), .ZN(n9198) );
  NAND2_X1 U11653 ( .A1(n9199), .A2(n9198), .ZN(n9200) );
  NAND2_X1 U11654 ( .A1(n12548), .A2(n9200), .ZN(n9201) );
  XNOR2_X1 U11655 ( .A(n12986), .B(n12474), .ZN(n9202) );
  INV_X1 U11656 ( .A(n9201), .ZN(n9204) );
  INV_X1 U11657 ( .A(n9202), .ZN(n9203) );
  XNOR2_X1 U11658 ( .A(n12531), .B(n6568), .ZN(n9206) );
  NAND2_X1 U11659 ( .A1(n9206), .A2(n12978), .ZN(n12516) );
  INV_X1 U11660 ( .A(n9206), .ZN(n9207) );
  NAND2_X1 U11661 ( .A1(n9207), .A2(n12767), .ZN(n9208) );
  AND2_X1 U11662 ( .A1(n12516), .A2(n9208), .ZN(n12533) );
  NAND2_X1 U11663 ( .A1(n12513), .A2(n12516), .ZN(n9214) );
  XNOR2_X1 U11664 ( .A(n12960), .B(n12474), .ZN(n9211) );
  NAND2_X1 U11665 ( .A1(n9211), .A2(n9210), .ZN(n9215) );
  INV_X1 U11666 ( .A(n9211), .ZN(n9212) );
  NAND2_X1 U11667 ( .A1(n9212), .A2(n12766), .ZN(n9213) );
  AND2_X1 U11668 ( .A1(n9215), .A2(n9213), .ZN(n12514) );
  XNOR2_X1 U11669 ( .A(n12949), .B(n12352), .ZN(n9216) );
  NOR2_X1 U11670 ( .A1(n9216), .A2(n12928), .ZN(n9217) );
  AOI21_X1 U11671 ( .B1(n9216), .B2(n12928), .A(n9217), .ZN(n12568) );
  NAND2_X1 U11672 ( .A1(n9225), .A2(n15124), .ZN(n9220) );
  INV_X1 U11673 ( .A(n9224), .ZN(n9219) );
  OAI22_X1 U11674 ( .A1(n9226), .A2(n9220), .B1(n9232), .B2(n9219), .ZN(n9221)
         );
  INV_X1 U11675 ( .A(n13084), .ZN(n9237) );
  NAND2_X1 U11676 ( .A1(n9226), .A2(n15071), .ZN(n9222) );
  INV_X1 U11677 ( .A(n9242), .ZN(n10532) );
  NAND2_X1 U11678 ( .A1(n12746), .A2(n9251), .ZN(n10487) );
  NAND3_X1 U11679 ( .A1(n9998), .A2(n10533), .A3(n10487), .ZN(n9223) );
  AOI21_X1 U11680 ( .B1(n9232), .B2(n9224), .A(n9223), .ZN(n9228) );
  NAND2_X1 U11681 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  NAND2_X1 U11682 ( .A1(n9228), .A2(n9227), .ZN(n9229) );
  NAND2_X1 U11683 ( .A1(n9229), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9231) );
  NAND3_X1 U11684 ( .A1(n9232), .A2(n9242), .A3(n10286), .ZN(n9230) );
  NAND2_X1 U11685 ( .A1(n9242), .A2(n12756), .ZN(n12760) );
  INV_X1 U11686 ( .A(n14446), .ZN(n12510) );
  NAND2_X1 U11687 ( .A1(n12510), .A2(n15061), .ZN(n14418) );
  NOR2_X2 U11688 ( .A1(n14446), .A2(n15050), .ZN(n14416) );
  AOI22_X1 U11689 ( .A1(n14416), .A2(n12927), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9233) );
  OAI21_X1 U11690 ( .B1(n9234), .B2(n14418), .A(n9233), .ZN(n9235) );
  AOI21_X1 U11691 ( .B1(n12930), .B2(n14444), .A(n9235), .ZN(n9236) );
  OAI21_X1 U11692 ( .B1(n9237), .B2(n12574), .A(n9236), .ZN(n9238) );
  INV_X1 U11693 ( .A(n9238), .ZN(n9239) );
  NAND2_X1 U11694 ( .A1(n9240), .A2(n9239), .ZN(P3_U3154) );
  INV_X1 U11695 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9259) );
  INV_X1 U11696 ( .A(n9241), .ZN(n9247) );
  NAND2_X1 U11697 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  NOR2_X1 U11698 ( .A1(n9245), .A2(n9244), .ZN(n9246) );
  NAND2_X1 U11699 ( .A1(n12750), .A2(n9248), .ZN(n10484) );
  AND2_X1 U11700 ( .A1(n10484), .A2(n10487), .ZN(n9256) );
  NAND2_X1 U11701 ( .A1(n12761), .A2(n12883), .ZN(n9249) );
  OAI21_X1 U11702 ( .B1(n15124), .B2(n9250), .A(n9249), .ZN(n9252) );
  NAND2_X1 U11703 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  NAND2_X1 U11704 ( .A1(n9253), .A2(n12750), .ZN(n9254) );
  NAND2_X1 U11705 ( .A1(n10485), .A2(n9254), .ZN(n9255) );
  OAI21_X1 U11706 ( .B1(n10485), .B2(n9256), .A(n9255), .ZN(n9257) );
  INV_X1 U11707 ( .A(n9257), .ZN(n9258) );
  NAND2_X1 U11708 ( .A1(n15144), .A2(n15105), .ZN(n13136) );
  NAND2_X1 U11709 ( .A1(n9261), .A2(n7697), .ZN(P3_U3488) );
  NOR2_X2 U11710 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9264) );
  NOR2_X1 U11711 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9272) );
  NOR2_X1 U11712 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n9271) );
  NAND4_X1 U11713 ( .A1(n9272), .A2(n9271), .A3(n9270), .A4(n9269), .ZN(n9645)
         );
  NOR2_X1 U11714 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9275) );
  NAND4_X1 U11715 ( .A1(n9275), .A2(n9657), .A3(n9274), .A4(n9273), .ZN(n9276)
         );
  INV_X1 U11716 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10084) );
  AND2_X4 U11717 ( .A1(n14364), .A2(n9282), .ZN(n9719) );
  INV_X1 U11718 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10096) );
  OR2_X1 U11719 ( .A1(n12266), .A2(n10096), .ZN(n9286) );
  INV_X1 U11720 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13862) );
  OR2_X1 U11721 ( .A1(n9598), .A2(n13862), .ZN(n9285) );
  NAND2_X1 U11722 ( .A1(n9289), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9291) );
  INV_X4 U11723 ( .A(n9305), .ZN(n9530) );
  NAND2_X1 U11724 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14566), .ZN(n9292) );
  XNOR2_X1 U11725 ( .A(n9292), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13865) );
  NAND2_X1 U11726 ( .A1(n9530), .A2(n13865), .ZN(n9295) );
  NAND2_X1 U11727 ( .A1(n12283), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11728 ( .A1(n9719), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9301) );
  INV_X1 U11729 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n14636) );
  OR2_X1 U11730 ( .A1(n9598), .A2(n14636), .ZN(n9300) );
  INV_X1 U11731 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9296) );
  INV_X1 U11732 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9297) );
  OR2_X1 U11733 ( .A1(n12266), .A2(n9297), .ZN(n9298) );
  OAI21_X1 U11734 ( .B1(n10006), .B2(n10019), .A(n9302), .ZN(n9303) );
  AND2_X1 U11735 ( .A1(n9304), .A2(n9303), .ZN(n14373) );
  MUX2_X1 U11736 ( .A(n14566), .B(n14373), .S(n9305), .Z(n14632) );
  NAND2_X1 U11737 ( .A1(n10342), .A2(n14632), .ZN(n10737) );
  NAND2_X1 U11738 ( .A1(n10736), .A2(n10737), .ZN(n9307) );
  INV_X1 U11739 ( .A(n12101), .ZN(n9306) );
  INV_X1 U11740 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9308) );
  INV_X1 U11741 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10703) );
  OR2_X1 U11742 ( .A1(n9598), .A2(n10703), .ZN(n9311) );
  INV_X1 U11743 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10095) );
  OR2_X1 U11744 ( .A1(n12266), .A2(n10095), .ZN(n9309) );
  AND4_X2 U11745 ( .A1(n7695), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(n9318)
         );
  INV_X1 U11746 ( .A(n9312), .ZN(n10054) );
  NAND2_X1 U11747 ( .A1(n12283), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9317) );
  NOR2_X1 U11748 ( .A1(n9313), .A2(n9287), .ZN(n9314) );
  MUX2_X1 U11749 ( .A(n9287), .B(n9314), .S(P1_IR_REG_2__SCAN_IN), .Z(n9316)
         );
  NOR2_X1 U11750 ( .A1(n9316), .A2(n6963), .ZN(n13890) );
  NAND2_X1 U11751 ( .A1(n9318), .A2(n10441), .ZN(n9319) );
  NAND2_X1 U11752 ( .A1(n9719), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9323) );
  INV_X1 U11753 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10089) );
  OR2_X1 U11754 ( .A1(n12264), .A2(n10089), .ZN(n9322) );
  INV_X1 U11755 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10819) );
  OR2_X1 U11756 ( .A1(n12266), .A2(n10819), .ZN(n9321) );
  OR2_X1 U11757 ( .A1(n9598), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9320) );
  INV_X1 U11758 ( .A(n12283), .ZN(n9449) );
  NAND2_X1 U11759 ( .A1(n9433), .A2(n10026), .ZN(n9326) );
  NAND2_X1 U11760 ( .A1(n9315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9324) );
  XNOR2_X1 U11761 ( .A(n9324), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13902) );
  NAND2_X1 U11762 ( .A1(n9530), .A2(n13902), .ZN(n9325) );
  NAND2_X1 U11763 ( .A1(n10596), .A2(n10822), .ZN(n12110) );
  INV_X1 U11764 ( .A(n10596), .ZN(n13858) );
  NAND2_X1 U11765 ( .A1(n13858), .A2(n7439), .ZN(n12111) );
  AND2_X2 U11766 ( .A1(n12110), .A2(n12111), .ZN(n12302) );
  INV_X1 U11767 ( .A(n12302), .ZN(n9327) );
  NAND2_X1 U11768 ( .A1(n10596), .A2(n7439), .ZN(n9328) );
  NAND2_X1 U11769 ( .A1(n9719), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9338) );
  INV_X1 U11770 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9330) );
  OR2_X1 U11771 ( .A1(n12264), .A2(n9330), .ZN(n9337) );
  INV_X1 U11772 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10100) );
  OR2_X1 U11773 ( .A1(n12266), .A2(n10100), .ZN(n9336) );
  AND2_X1 U11774 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9346) );
  INV_X1 U11775 ( .A(n9346), .ZN(n9334) );
  INV_X1 U11776 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9332) );
  INV_X1 U11777 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U11778 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  NAND2_X1 U11779 ( .A1(n9334), .A2(n9333), .ZN(n14613) );
  OR2_X1 U11780 ( .A1(n9598), .A2(n14613), .ZN(n9335) );
  NAND2_X1 U11781 ( .A1(n10035), .A2(n12259), .ZN(n9345) );
  NAND2_X1 U11782 ( .A1(n9340), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9339) );
  MUX2_X1 U11783 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9339), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9342) );
  NOR2_X1 U11784 ( .A1(n9340), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9357) );
  INV_X1 U11785 ( .A(n9357), .ZN(n9341) );
  NAND2_X1 U11786 ( .A1(n9530), .A2(n13917), .ZN(n9344) );
  NAND2_X1 U11787 ( .A1(n12283), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9343) );
  AND3_X2 U11788 ( .A1(n9345), .A2(n9344), .A3(n9343), .ZN(n14684) );
  OR2_X1 U11789 ( .A1(n13857), .A2(n12115), .ZN(n12300) );
  NAND2_X1 U11790 ( .A1(n13857), .A2(n12115), .ZN(n12299) );
  NAND2_X1 U11791 ( .A1(n9346), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9362) );
  OAI21_X1 U11792 ( .B1(n9346), .B2(P1_REG3_REG_5__SCAN_IN), .A(n9362), .ZN(
        n11989) );
  OR2_X1 U11793 ( .A1(n9598), .A2(n11989), .ZN(n9350) );
  NAND2_X1 U11794 ( .A1(n9631), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U11795 ( .A1(n9719), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11796 ( .A1(n9718), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U11797 ( .A1(n10029), .A2(n12259), .ZN(n9353) );
  OR2_X1 U11798 ( .A1(n9357), .A2(n9287), .ZN(n9351) );
  XNOR2_X1 U11799 ( .A(n9351), .B(P1_IR_REG_5__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U11800 ( .A1(n12283), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9530), 
        .B2(n13927), .ZN(n9352) );
  NAND2_X1 U11801 ( .A1(n9353), .A2(n9352), .ZN(n14692) );
  INV_X1 U11802 ( .A(n14692), .ZN(n11995) );
  NAND2_X1 U11803 ( .A1(n11204), .A2(n11995), .ZN(n9355) );
  NAND2_X1 U11804 ( .A1(n13856), .A2(n14692), .ZN(n9354) );
  AND2_X1 U11805 ( .A1(n9355), .A2(n9354), .ZN(n12304) );
  INV_X1 U11806 ( .A(n12304), .ZN(n11977) );
  NAND2_X1 U11807 ( .A1(n10038), .A2(n12259), .ZN(n9360) );
  INV_X1 U11808 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U11809 ( .A1(n9357), .A2(n9356), .ZN(n9370) );
  NAND2_X1 U11810 ( .A1(n9370), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9358) );
  XNOR2_X1 U11811 ( .A(n9358), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U11812 ( .A1(n12283), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9530), 
        .B2(n10105), .ZN(n9359) );
  NAND2_X1 U11813 ( .A1(n9360), .A2(n9359), .ZN(n14696) );
  NAND2_X1 U11814 ( .A1(n9631), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U11815 ( .A1(n9719), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9366) );
  NOR2_X1 U11816 ( .A1(n9362), .A2(n9361), .ZN(n9373) );
  AND2_X1 U11817 ( .A1(n9362), .A2(n9361), .ZN(n9363) );
  NOR2_X1 U11818 ( .A1(n9373), .A2(n9363), .ZN(n11098) );
  NAND2_X1 U11819 ( .A1(n9633), .A2(n11098), .ZN(n9365) );
  NAND2_X1 U11820 ( .A1(n9718), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9364) );
  NAND4_X1 U11821 ( .A1(n9367), .A2(n9366), .A3(n9365), .A4(n9364), .ZN(n13855) );
  OR2_X1 U11822 ( .A1(n14696), .A2(n13855), .ZN(n9369) );
  NAND2_X1 U11823 ( .A1(n14696), .A2(n13855), .ZN(n9368) );
  NAND2_X1 U11824 ( .A1(n9369), .A2(n9368), .ZN(n12306) );
  INV_X1 U11825 ( .A(n12306), .ZN(n11101) );
  NAND2_X1 U11826 ( .A1(n11100), .A2(n11101), .ZN(n11099) );
  NAND2_X1 U11827 ( .A1(n11099), .A2(n9369), .ZN(n11164) );
  NAND2_X1 U11828 ( .A1(n10044), .A2(n12259), .ZN(n9372) );
  NAND2_X1 U11829 ( .A1(n9409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9380) );
  XNOR2_X1 U11830 ( .A(n9380), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13950) );
  AOI22_X1 U11831 ( .A1(n12283), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9530), 
        .B2(n13950), .ZN(n9371) );
  NAND2_X1 U11832 ( .A1(n9372), .A2(n9371), .ZN(n12129) );
  NAND2_X1 U11833 ( .A1(n9373), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9398) );
  OR2_X1 U11834 ( .A1(n9373), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U11835 ( .A1(n9398), .A2(n9374), .ZN(n11572) );
  OR2_X1 U11836 ( .A1(n9598), .A2(n11572), .ZN(n9378) );
  NAND2_X1 U11837 ( .A1(n9631), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9377) );
  NAND2_X1 U11838 ( .A1(n9719), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11839 ( .A1(n9718), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9375) );
  NAND4_X1 U11840 ( .A1(n9378), .A2(n9377), .A3(n9376), .A4(n9375), .ZN(n13854) );
  XNOR2_X1 U11841 ( .A(n12129), .B(n13854), .ZN(n12307) );
  INV_X1 U11842 ( .A(n12307), .ZN(n11165) );
  OR2_X1 U11843 ( .A1(n12129), .A2(n13854), .ZN(n9379) );
  NAND2_X1 U11844 ( .A1(n11163), .A2(n9379), .ZN(n11131) );
  NAND2_X1 U11845 ( .A1(n10057), .A2(n12259), .ZN(n9383) );
  INV_X1 U11846 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n15337) );
  NAND2_X1 U11847 ( .A1(n9380), .A2(n15337), .ZN(n9381) );
  NAND2_X1 U11848 ( .A1(n9381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9390) );
  XNOR2_X1 U11849 ( .A(n9390), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U11850 ( .A1(n12283), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9530), 
        .B2(n10211), .ZN(n9382) );
  NAND2_X1 U11851 ( .A1(n9383), .A2(n9382), .ZN(n12132) );
  NAND2_X1 U11852 ( .A1(n9631), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U11853 ( .A1(n9719), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9386) );
  XNOR2_X1 U11854 ( .A(n9398), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U11855 ( .A1(n9633), .A2(n11584), .ZN(n9385) );
  NAND2_X1 U11856 ( .A1(n9718), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9384) );
  NAND4_X1 U11857 ( .A1(n9387), .A2(n9386), .A3(n9385), .A4(n9384), .ZN(n13853) );
  OR2_X1 U11858 ( .A1(n12132), .A2(n13853), .ZN(n9389) );
  NAND2_X1 U11859 ( .A1(n12132), .A2(n13853), .ZN(n9388) );
  NAND2_X1 U11860 ( .A1(n9389), .A2(n9388), .ZN(n12309) );
  NAND2_X1 U11861 ( .A1(n11131), .A2(n11130), .ZN(n11129) );
  NAND2_X1 U11862 ( .A1(n11129), .A2(n9389), .ZN(n11268) );
  NAND2_X1 U11863 ( .A1(n10061), .A2(n12259), .ZN(n9394) );
  NAND2_X1 U11864 ( .A1(n9390), .A2(n9406), .ZN(n9391) );
  NAND2_X1 U11865 ( .A1(n9391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9392) );
  XNOR2_X1 U11866 ( .A(n9392), .B(P1_IR_REG_9__SCAN_IN), .ZN(n13968) );
  AOI22_X1 U11867 ( .A1(n12283), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9530), 
        .B2(n13968), .ZN(n9393) );
  NAND2_X1 U11868 ( .A1(n9394), .A2(n9393), .ZN(n12141) );
  INV_X1 U11869 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9396) );
  INV_X1 U11870 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9395) );
  OAI21_X1 U11871 ( .B1(n9398), .B2(n9396), .A(n9395), .ZN(n9399) );
  NAND2_X1 U11872 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n9397) );
  NAND2_X1 U11873 ( .A1(n9399), .A2(n9416), .ZN(n11565) );
  OR2_X1 U11874 ( .A1(n9598), .A2(n11565), .ZN(n9403) );
  NAND2_X1 U11875 ( .A1(n9631), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9402) );
  NAND2_X1 U11876 ( .A1(n9719), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11877 ( .A1(n9718), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9400) );
  NAND4_X1 U11878 ( .A1(n9403), .A2(n9402), .A3(n9401), .A4(n9400), .ZN(n13852) );
  INV_X1 U11879 ( .A(n13852), .ZN(n11555) );
  XNOR2_X1 U11880 ( .A(n12141), .B(n11555), .ZN(n12311) );
  NAND2_X1 U11881 ( .A1(n11268), .A2(n12311), .ZN(n11267) );
  OR2_X1 U11882 ( .A1(n12141), .A2(n13852), .ZN(n9404) );
  NAND2_X1 U11883 ( .A1(n10077), .A2(n12259), .ZN(n9415) );
  INV_X1 U11884 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9405) );
  NAND3_X1 U11885 ( .A1(n15337), .A2(n9406), .A3(n9405), .ZN(n9408) );
  NOR2_X1 U11886 ( .A1(n9409), .A2(n9408), .ZN(n9412) );
  OR2_X1 U11887 ( .A1(n9412), .A2(n9287), .ZN(n9410) );
  MUX2_X1 U11888 ( .A(n9410), .B(P1_IR_REG_31__SCAN_IN), .S(n9411), .Z(n9413)
         );
  NAND2_X1 U11889 ( .A1(n9412), .A2(n9411), .ZN(n9434) );
  NAND2_X1 U11890 ( .A1(n9413), .A2(n9434), .ZN(n10297) );
  INV_X1 U11891 ( .A(n10297), .ZN(n10302) );
  AOI22_X1 U11892 ( .A1(n12283), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9530), 
        .B2(n10302), .ZN(n9414) );
  NAND2_X1 U11893 ( .A1(n9415), .A2(n9414), .ZN(n12150) );
  AND2_X1 U11894 ( .A1(n9416), .A2(n15303), .ZN(n9417) );
  NOR2_X1 U11895 ( .A1(n9424), .A2(n9417), .ZN(n14600) );
  NAND2_X1 U11896 ( .A1(n9633), .A2(n14600), .ZN(n9421) );
  NAND2_X1 U11897 ( .A1(n9631), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U11898 ( .A1(n9719), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U11899 ( .A1(n9718), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9418) );
  NAND4_X1 U11900 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(n13851) );
  XNOR2_X1 U11901 ( .A(n12150), .B(n13851), .ZN(n12312) );
  INV_X1 U11902 ( .A(n12312), .ZN(n11397) );
  OR2_X1 U11903 ( .A1(n12150), .A2(n13851), .ZN(n9422) );
  NAND2_X1 U11904 ( .A1(n9719), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9429) );
  INV_X1 U11905 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11379) );
  OR2_X1 U11906 ( .A1(n12266), .A2(n11379), .ZN(n9428) );
  INV_X1 U11907 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9423) );
  OR2_X1 U11908 ( .A1(n12264), .A2(n9423), .ZN(n9427) );
  NOR2_X1 U11909 ( .A1(n9424), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9425) );
  OR2_X1 U11910 ( .A1(n9438), .A2(n9425), .ZN(n11843) );
  OR2_X1 U11911 ( .A1(n9598), .A2(n11843), .ZN(n9426) );
  NAND2_X1 U11912 ( .A1(n10135), .A2(n12259), .ZN(n9432) );
  NAND2_X1 U11913 ( .A1(n9434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9430) );
  XNOR2_X1 U11914 ( .A(n9430), .B(P1_IR_REG_11__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U11915 ( .A1(n12283), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9530), 
        .B2(n13985), .ZN(n9431) );
  NAND2_X1 U11916 ( .A1(n10201), .A2(n12259), .ZN(n9437) );
  NAND2_X1 U11917 ( .A1(n9435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9447) );
  XNOR2_X1 U11918 ( .A(n9447), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U11919 ( .A1(n12283), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9530), 
        .B2(n10449), .ZN(n9436) );
  OR2_X1 U11920 ( .A1(n9438), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U11921 ( .A1(n9454), .A2(n9439), .ZN(n11829) );
  OR2_X1 U11922 ( .A1(n9598), .A2(n11829), .ZN(n9443) );
  NAND2_X1 U11923 ( .A1(n9718), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U11924 ( .A1(n9631), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U11925 ( .A1(n9719), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9440) );
  NAND4_X1 U11926 ( .A1(n9443), .A2(n9442), .A3(n9441), .A4(n9440), .ZN(n13849) );
  XNOR2_X1 U11927 ( .A(n14401), .B(n13849), .ZN(n12315) );
  INV_X1 U11928 ( .A(n12315), .ZN(n11600) );
  NOR2_X1 U11929 ( .A1(n14401), .A2(n13849), .ZN(n12155) );
  INV_X1 U11930 ( .A(n12155), .ZN(n9444) );
  NAND2_X1 U11931 ( .A1(n9445), .A2(n9444), .ZN(n11785) );
  NAND2_X1 U11932 ( .A1(n10242), .A2(n12259), .ZN(n9452) );
  NAND2_X1 U11933 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  NAND2_X1 U11934 ( .A1(n9448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9462) );
  INV_X1 U11935 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9461) );
  XNOR2_X1 U11936 ( .A(n9462), .B(n9461), .ZN(n10521) );
  OAI22_X1 U11937 ( .A1(n10521), .A2(n9305), .B1(n9449), .B2(n10243), .ZN(
        n9450) );
  INV_X1 U11938 ( .A(n9450), .ZN(n9451) );
  NAND2_X1 U11939 ( .A1(n9719), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9459) );
  INV_X1 U11940 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10457) );
  OR2_X1 U11941 ( .A1(n12264), .A2(n10457), .ZN(n9458) );
  INV_X1 U11942 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U11943 ( .A1(n9454), .A2(n9453), .ZN(n9455) );
  NAND2_X1 U11944 ( .A1(n9468), .A2(n9455), .ZN(n11961) );
  OR2_X1 U11945 ( .A1(n9598), .A2(n11961), .ZN(n9457) );
  INV_X1 U11946 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10452) );
  OR2_X1 U11947 ( .A1(n12266), .A2(n10452), .ZN(n9456) );
  XNOR2_X1 U11948 ( .A(n12171), .B(n12166), .ZN(n12317) );
  OR2_X1 U11949 ( .A1(n12171), .A2(n13848), .ZN(n9460) );
  NAND2_X1 U11950 ( .A1(n10368), .A2(n12259), .ZN(n9466) );
  NAND2_X1 U11951 ( .A1(n9462), .A2(n9461), .ZN(n9463) );
  NAND2_X1 U11952 ( .A1(n9463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9464) );
  XNOR2_X1 U11953 ( .A(n9464), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U11954 ( .A1(n11312), .A2(n9530), .B1(n12283), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U11955 ( .A1(n9719), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9474) );
  INV_X1 U11956 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9467) );
  OR2_X1 U11957 ( .A1(n12264), .A2(n9467), .ZN(n9473) );
  NAND2_X1 U11958 ( .A1(n9468), .A2(n15429), .ZN(n9469) );
  NAND2_X1 U11959 ( .A1(n9496), .A2(n9469), .ZN(n14510) );
  OR2_X1 U11960 ( .A1(n9598), .A2(n14510), .ZN(n9472) );
  INV_X1 U11961 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9470) );
  OR2_X1 U11962 ( .A1(n12266), .A2(n9470), .ZN(n9471) );
  OR2_X1 U11963 ( .A1(n14513), .A2(n13829), .ZN(n12179) );
  NAND2_X1 U11964 ( .A1(n14513), .A2(n13829), .ZN(n12180) );
  INV_X1 U11965 ( .A(n13829), .ZN(n13847) );
  NAND2_X1 U11966 ( .A1(n14513), .A2(n13847), .ZN(n9477) );
  NOR2_X1 U11967 ( .A1(n9506), .A2(n9287), .ZN(n9478) );
  MUX2_X1 U11968 ( .A(n9287), .B(n9478), .S(P1_IR_REG_15__SCAN_IN), .Z(n9481)
         );
  INV_X1 U11969 ( .A(n9490), .ZN(n9480) );
  OR2_X1 U11970 ( .A1(n9481), .A2(n9480), .ZN(n14578) );
  AOI22_X1 U11971 ( .A1(n12283), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9530), 
        .B2(n11323), .ZN(n9482) );
  NAND2_X1 U11972 ( .A1(n9631), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9489) );
  INV_X1 U11973 ( .A(n9719), .ZN(n12267) );
  INV_X1 U11974 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9483) );
  OR2_X1 U11975 ( .A1(n12267), .A2(n9483), .ZN(n9488) );
  INV_X1 U11976 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9484) );
  XNOR2_X1 U11977 ( .A(n9496), .B(n9484), .ZN(n14243) );
  OR2_X1 U11978 ( .A1(n9598), .A2(n14243), .ZN(n9487) );
  INV_X1 U11979 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9485) );
  OR2_X1 U11980 ( .A1(n12266), .A2(n9485), .ZN(n9486) );
  NAND2_X1 U11981 ( .A1(n14334), .A2(n14217), .ZN(n12186) );
  NAND2_X1 U11982 ( .A1(n12181), .A2(n12186), .ZN(n14235) );
  INV_X1 U11983 ( .A(n14235), .ZN(n14248) );
  INV_X1 U11984 ( .A(n14217), .ZN(n13846) );
  NAND2_X1 U11985 ( .A1(n10332), .A2(n12259), .ZN(n9493) );
  NAND2_X1 U11986 ( .A1(n9490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9491) );
  XNOR2_X1 U11987 ( .A(n9491), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U11988 ( .A1(n12283), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9530), 
        .B2(n11523), .ZN(n9492) );
  NAND2_X1 U11989 ( .A1(n9631), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U11990 ( .A1(n9719), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9500) );
  INV_X1 U11991 ( .A(n9496), .ZN(n9494) );
  AOI21_X1 U11992 ( .B1(n9494), .B2(P1_REG3_REG_15__SCAN_IN), .A(
        P1_REG3_REG_16__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11993 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n9495) );
  NOR2_X1 U11994 ( .A1(n9497), .A2(n9510), .ZN(n14222) );
  NAND2_X1 U11995 ( .A1(n9633), .A2(n14222), .ZN(n9499) );
  NAND2_X1 U11996 ( .A1(n9718), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9498) );
  NAND4_X1 U11997 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(n14208) );
  INV_X1 U11998 ( .A(n14208), .ZN(n13828) );
  XNOR2_X1 U11999 ( .A(n14330), .B(n13828), .ZN(n14228) );
  NAND2_X1 U12000 ( .A1(n14229), .A2(n14228), .ZN(n9503) );
  OR2_X1 U12001 ( .A1(n14330), .A2(n14208), .ZN(n9502) );
  NAND2_X1 U12002 ( .A1(n10388), .A2(n12259), .ZN(n9509) );
  NAND2_X1 U12003 ( .A1(n9646), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9507) );
  XNOR2_X1 U12004 ( .A(n9507), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U12005 ( .A1(n12283), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9530), 
        .B2(n11517), .ZN(n9508) );
  NAND2_X1 U12006 ( .A1(n9631), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U12007 ( .A1(n9719), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9514) );
  OR2_X1 U12008 ( .A1(n9510), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U12009 ( .A1(n9510), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9522) );
  AND2_X1 U12010 ( .A1(n9511), .A2(n9522), .ZN(n14200) );
  NAND2_X1 U12011 ( .A1(n9633), .A2(n14200), .ZN(n9513) );
  NAND2_X1 U12012 ( .A1(n9718), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9512) );
  NAND4_X1 U12013 ( .A1(n9515), .A2(n9514), .A3(n9513), .A4(n9512), .ZN(n13845) );
  OR2_X1 U12014 ( .A1(n14202), .A2(n14220), .ZN(n9516) );
  OR2_X1 U12015 ( .A1(n10574), .A2(n9545), .ZN(n9520) );
  OR2_X1 U12016 ( .A1(n9646), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U12017 ( .A1(n9517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9518) );
  XNOR2_X1 U12018 ( .A(n9518), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14005) );
  AOI22_X1 U12019 ( .A1(n12283), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9530), 
        .B2(n14005), .ZN(n9519) );
  INV_X1 U12020 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9521) );
  NAND2_X1 U12021 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  NAND2_X1 U12022 ( .A1(n9533), .A2(n9523), .ZN(n14190) );
  INV_X1 U12023 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14191) );
  OAI22_X1 U12024 ( .A1(n14190), .A2(n9598), .B1(n12266), .B2(n14191), .ZN(
        n9525) );
  INV_X1 U12025 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14321) );
  INV_X1 U12026 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15270) );
  OAI22_X1 U12027 ( .A1(n12264), .A2(n14321), .B1(n12267), .B2(n15270), .ZN(
        n9524) );
  AND2_X1 U12028 ( .A1(n14193), .A2(n14206), .ZN(n12210) );
  INV_X1 U12029 ( .A(n12210), .ZN(n9526) );
  OR2_X1 U12030 ( .A1(n14193), .A2(n14206), .ZN(n12209) );
  NAND2_X1 U12031 ( .A1(n10852), .A2(n9433), .ZN(n9532) );
  NAND2_X1 U12032 ( .A1(n6670), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9528) );
  MUX2_X1 U12033 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9528), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9529) );
  AOI22_X1 U12034 ( .A1(n12283), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9530), 
        .B2(n14143), .ZN(n9531) );
  AND2_X1 U12035 ( .A1(n9533), .A2(n13732), .ZN(n9534) );
  OR2_X1 U12036 ( .A1(n9534), .A2(n9541), .ZN(n14168) );
  AOI22_X1 U12037 ( .A1(n9631), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n9718), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U12038 ( .A1(n9719), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9535) );
  OAI211_X1 U12039 ( .C1(n14168), .C2(n9598), .A(n9536), .B(n9535), .ZN(n14151) );
  INV_X1 U12040 ( .A(n14151), .ZN(n9537) );
  OR2_X1 U12041 ( .A1(n14313), .A2(n9537), .ZN(n12214) );
  NAND2_X1 U12042 ( .A1(n14313), .A2(n9537), .ZN(n12215) );
  OR2_X1 U12043 ( .A1(n14313), .A2(n14151), .ZN(n9538) );
  OR2_X1 U12044 ( .A1(n11175), .A2(n9545), .ZN(n9540) );
  NAND2_X1 U12045 ( .A1(n12283), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9539) );
  NOR2_X1 U12046 ( .A1(n9541), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9542) );
  OR2_X1 U12047 ( .A1(n9548), .A2(n9542), .ZN(n13788) );
  AOI22_X1 U12048 ( .A1(n9631), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n9718), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U12049 ( .A1(n9719), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9543) );
  OAI211_X1 U12050 ( .C1(n13788), .C2(n9598), .A(n9544), .B(n9543), .ZN(n13844) );
  XNOR2_X1 U12051 ( .A(n14304), .B(n13844), .ZN(n14161) );
  OR2_X1 U12052 ( .A1(n11359), .A2(n9545), .ZN(n9547) );
  NAND2_X1 U12053 ( .A1(n12283), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9546) );
  NOR2_X1 U12054 ( .A1(n9548), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9549) );
  OR2_X1 U12055 ( .A1(n9558), .A2(n9549), .ZN(n14145) );
  INV_X1 U12056 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15438) );
  NAND2_X1 U12057 ( .A1(n9718), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U12058 ( .A1(n9719), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9550) );
  OAI211_X1 U12059 ( .C1(n12264), .C2(n15438), .A(n9551), .B(n9550), .ZN(n9552) );
  INV_X1 U12060 ( .A(n9552), .ZN(n9553) );
  XNOR2_X1 U12061 ( .A(n14299), .B(n14152), .ZN(n14134) );
  INV_X1 U12062 ( .A(n14152), .ZN(n13790) );
  NAND2_X1 U12063 ( .A1(n14149), .A2(n13790), .ZN(n9555) );
  XNOR2_X1 U12064 ( .A(n9557), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14372) );
  OR2_X1 U12065 ( .A1(n9558), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U12066 ( .A1(n9558), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9568) );
  AND2_X1 U12067 ( .A1(n9559), .A2(n9568), .ZN(n14127) );
  NAND2_X1 U12068 ( .A1(n14127), .A2(n9633), .ZN(n9564) );
  INV_X1 U12069 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15271) );
  NAND2_X1 U12070 ( .A1(n9718), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U12071 ( .A1(n9719), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9560) );
  OAI211_X1 U12072 ( .C1(n12264), .C2(n15271), .A(n9561), .B(n9560), .ZN(n9562) );
  INV_X1 U12073 ( .A(n9562), .ZN(n9563) );
  NAND2_X1 U12074 ( .A1(n9564), .A2(n9563), .ZN(n13843) );
  NAND2_X1 U12075 ( .A1(n14298), .A2(n13843), .ZN(n9565) );
  NAND2_X1 U12076 ( .A1(n11669), .A2(n9433), .ZN(n9567) );
  NAND2_X1 U12077 ( .A1(n12283), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9566) );
  OAI21_X1 U12078 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9569), .A(n9577), .ZN(
        n14108) );
  OR2_X1 U12079 ( .A1(n9598), .A2(n14108), .ZN(n9573) );
  NAND2_X1 U12080 ( .A1(n9718), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U12081 ( .A1(n9631), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U12082 ( .A1(n9719), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9570) );
  NAND4_X1 U12083 ( .A1(n9573), .A2(n9572), .A3(n9571), .A4(n9570), .ZN(n14121) );
  NAND2_X1 U12084 ( .A1(n14291), .A2(n14121), .ZN(n9583) );
  OR2_X1 U12085 ( .A1(n14291), .A2(n14121), .ZN(n9574) );
  NAND2_X1 U12086 ( .A1(n9583), .A2(n9574), .ZN(n14105) );
  NAND2_X1 U12087 ( .A1(n11715), .A2(n9433), .ZN(n9576) );
  NAND2_X1 U12088 ( .A1(n12283), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U12089 ( .A1(n9578), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9588) );
  OAI21_X1 U12090 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9578), .A(n9588), .ZN(
        n14095) );
  OR2_X1 U12091 ( .A1(n9598), .A2(n14095), .ZN(n9582) );
  NAND2_X1 U12092 ( .A1(n9631), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U12093 ( .A1(n9719), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U12094 ( .A1(n9718), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9579) );
  NAND4_X1 U12095 ( .A1(n9582), .A2(n9581), .A3(n9580), .A4(n9579), .ZN(n13842) );
  XNOR2_X1 U12096 ( .A(n14097), .B(n13842), .ZN(n14085) );
  INV_X1 U12097 ( .A(n9583), .ZN(n14086) );
  NOR2_X1 U12098 ( .A1(n14085), .A2(n14086), .ZN(n9584) );
  OR2_X1 U12099 ( .A1(n14097), .A2(n13842), .ZN(n9585) );
  NAND2_X1 U12100 ( .A1(n11895), .A2(n12259), .ZN(n9587) );
  NAND2_X1 U12101 ( .A1(n12283), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9586) );
  NAND2_X1 U12102 ( .A1(n9589), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9596) );
  OAI21_X1 U12103 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9589), .A(n9596), .ZN(
        n14075) );
  OR2_X1 U12104 ( .A1(n9598), .A2(n14075), .ZN(n9593) );
  NAND2_X1 U12105 ( .A1(n9718), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9592) );
  NAND2_X1 U12106 ( .A1(n9631), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U12107 ( .A1(n9719), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9590) );
  NAND4_X1 U12108 ( .A1(n9593), .A2(n9592), .A3(n9591), .A4(n9590), .ZN(n13841) );
  XNOR2_X1 U12109 ( .A(n14077), .B(n13841), .ZN(n14072) );
  NAND2_X1 U12110 ( .A1(n11971), .A2(n9433), .ZN(n9595) );
  NAND2_X1 U12111 ( .A1(n12283), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9594) );
  INV_X1 U12112 ( .A(n9596), .ZN(n9597) );
  NAND2_X1 U12113 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9597), .ZN(n9614) );
  OAI21_X1 U12114 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n9597), .A(n9614), .ZN(
        n14052) );
  OR2_X1 U12115 ( .A1(n9598), .A2(n14052), .ZN(n9602) );
  NAND2_X1 U12116 ( .A1(n9718), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U12117 ( .A1(n9631), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U12118 ( .A1(n9719), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9599) );
  NAND4_X1 U12119 ( .A1(n9602), .A2(n9601), .A3(n9600), .A4(n9599), .ZN(n14033) );
  XNOR2_X1 U12120 ( .A(n14275), .B(n13749), .ZN(n14056) );
  NAND2_X1 U12121 ( .A1(n14275), .A2(n14033), .ZN(n9603) );
  NAND2_X1 U12122 ( .A1(n12049), .A2(n9433), .ZN(n9605) );
  NAND2_X1 U12123 ( .A1(n12283), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U12124 ( .A1(n9718), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U12125 ( .A1(n9631), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9608) );
  XNOR2_X1 U12126 ( .A(n9614), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n14039) );
  NAND2_X1 U12127 ( .A1(n9633), .A2(n14039), .ZN(n9607) );
  NAND2_X1 U12128 ( .A1(n9719), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9606) );
  OR2_X1 U12129 ( .A1(n14270), .A2(n13840), .ZN(n9610) );
  NAND2_X1 U12130 ( .A1(n12283), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9611) );
  INV_X1 U12131 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9613) );
  INV_X1 U12132 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9612) );
  OAI21_X1 U12133 ( .B1(n9614), .B2(n9613), .A(n9612), .ZN(n9617) );
  INV_X1 U12134 ( .A(n9614), .ZN(n9616) );
  AND2_X1 U12135 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9615) );
  NAND2_X1 U12136 ( .A1(n9616), .A2(n9615), .ZN(n9632) );
  NAND2_X1 U12137 ( .A1(n9617), .A2(n9632), .ZN(n12470) );
  OR2_X1 U12138 ( .A1(n9598), .A2(n12470), .ZN(n9621) );
  NAND2_X1 U12139 ( .A1(n9718), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U12140 ( .A1(n9631), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U12141 ( .A1(n9719), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12142 ( .A1(n14265), .A2(n14034), .ZN(n9623) );
  INV_X1 U12143 ( .A(n12326), .ZN(n12062) );
  INV_X1 U12144 ( .A(n9624), .ZN(n9625) );
  INV_X1 U12145 ( .A(SI_28_), .ZN(n12363) );
  NAND2_X1 U12146 ( .A1(n9625), .A2(n12363), .ZN(n9626) );
  INV_X1 U12147 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14363) );
  MUX2_X1 U12148 ( .A(n14363), .B(n13695), .S(n10006), .Z(n9886) );
  XNOR2_X1 U12149 ( .A(n9886), .B(SI_29_), .ZN(n9884) );
  NAND2_X1 U12150 ( .A1(n13694), .A2(n9433), .ZN(n9630) );
  NAND2_X1 U12151 ( .A1(n12283), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U12152 ( .A1(n9718), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U12153 ( .A1(n9631), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9636) );
  INV_X1 U12154 ( .A(n9632), .ZN(n9723) );
  NAND2_X1 U12155 ( .A1(n9633), .A2(n9723), .ZN(n9635) );
  NAND2_X1 U12156 ( .A1(n9719), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9634) );
  NAND4_X1 U12157 ( .A1(n9637), .A2(n9636), .A3(n9635), .A4(n9634), .ZN(n13839) );
  XNOR2_X1 U12158 ( .A(n14260), .B(n13839), .ZN(n12328) );
  NAND2_X1 U12159 ( .A1(n9643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12160 ( .A1(n14371), .A2(n12273), .ZN(n12287) );
  INV_X1 U12161 ( .A(n12287), .ZN(n9713) );
  NAND2_X1 U12162 ( .A1(n9641), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9642) );
  MUX2_X1 U12163 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9642), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9644) );
  NAND2_X1 U12164 ( .A1(n12275), .A2(n14014), .ZN(n10355) );
  XNOR2_X2 U12165 ( .A(n9648), .B(P1_IR_REG_25__SCAN_IN), .ZN(n11896) );
  INV_X1 U12166 ( .A(n9649), .ZN(n9650) );
  NAND2_X1 U12167 ( .A1(n9650), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9651) );
  MUX2_X1 U12168 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9651), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9652) );
  OAI21_X2 U12169 ( .B1(n9653), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9654) );
  AOI21_X1 U12170 ( .B1(n9713), .B2(n10355), .A(n10343), .ZN(n10586) );
  NAND2_X1 U12171 ( .A1(n9656), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9658) );
  XNOR2_X1 U12172 ( .A(n9658), .B(n9657), .ZN(n10081) );
  INV_X1 U12173 ( .A(P1_B_REG_SCAN_IN), .ZN(n9716) );
  NOR2_X1 U12174 ( .A1(n11896), .A2(n9716), .ZN(n9659) );
  MUX2_X1 U12175 ( .A(n9659), .B(n9716), .S(n11716), .Z(n9660) );
  NOR4_X1 U12176 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9669) );
  NOR4_X1 U12177 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9668) );
  INV_X1 U12178 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15418) );
  INV_X1 U12179 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15372) );
  INV_X1 U12180 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15229) );
  INV_X1 U12181 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15310) );
  NAND4_X1 U12182 ( .A1(n15418), .A2(n15372), .A3(n15229), .A4(n15310), .ZN(
        n9666) );
  NOR4_X1 U12183 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9664) );
  NOR4_X1 U12184 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9663) );
  NOR4_X1 U12185 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9662) );
  NOR4_X1 U12186 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9661) );
  NAND4_X1 U12187 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9665)
         );
  NOR4_X1 U12188 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9666), .A4(n9665), .ZN(n9667) );
  NAND3_X1 U12189 ( .A1(n9669), .A2(n9668), .A3(n9667), .ZN(n9670) );
  NAND2_X1 U12190 ( .A1(n9676), .A2(n9670), .ZN(n10352) );
  INV_X1 U12191 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9672) );
  NOR2_X1 U12192 ( .A1(n10075), .A2(n11716), .ZN(n9671) );
  INV_X1 U12193 ( .A(n10353), .ZN(n9673) );
  INV_X1 U12194 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9675) );
  NOR2_X1 U12195 ( .A1(n10075), .A2(n11896), .ZN(n9674) );
  NAND2_X1 U12196 ( .A1(n10235), .A2(n10354), .ZN(n9715) );
  NAND2_X1 U12197 ( .A1(n10237), .A2(n12275), .ZN(n12286) );
  INV_X1 U12198 ( .A(n10072), .ZN(n10069) );
  INV_X1 U12199 ( .A(n12288), .ZN(n9677) );
  NAND2_X2 U12200 ( .A1(n9677), .A2(n12088), .ZN(n12450) );
  NAND2_X1 U12201 ( .A1(n12288), .A2(n14371), .ZN(n9678) );
  NAND2_X1 U12202 ( .A1(n10817), .A2(n12302), .ZN(n9680) );
  NAND2_X1 U12203 ( .A1(n9680), .A2(n12110), .ZN(n14608) );
  AND2_X1 U12204 ( .A1(n12114), .A2(n12115), .ZN(n9682) );
  NAND2_X1 U12205 ( .A1(n13857), .A2(n14684), .ZN(n9681) );
  OR2_X1 U12206 ( .A1(n11982), .A2(n12304), .ZN(n11984) );
  NAND2_X1 U12207 ( .A1(n11204), .A2(n14692), .ZN(n9683) );
  NAND2_X1 U12208 ( .A1(n11104), .A2(n12306), .ZN(n11103) );
  INV_X1 U12209 ( .A(n13855), .ZN(n9684) );
  NAND2_X1 U12210 ( .A1(n14696), .A2(n9684), .ZN(n9685) );
  INV_X1 U12211 ( .A(n13854), .ZN(n9687) );
  OR2_X1 U12212 ( .A1(n12129), .A2(n9687), .ZN(n9686) );
  NAND2_X1 U12213 ( .A1(n12129), .A2(n9687), .ZN(n9688) );
  INV_X1 U12214 ( .A(n13853), .ZN(n11266) );
  OR2_X1 U12215 ( .A1(n12132), .A2(n11266), .ZN(n9689) );
  INV_X1 U12216 ( .A(n12311), .ZN(n11263) );
  NAND2_X1 U12217 ( .A1(n12141), .A2(n11555), .ZN(n9690) );
  INV_X1 U12218 ( .A(n13851), .ZN(n11265) );
  OR2_X1 U12219 ( .A1(n12150), .A2(n11265), .ZN(n9691) );
  OR2_X1 U12220 ( .A1(n14530), .A2(n13850), .ZN(n9692) );
  NAND2_X1 U12221 ( .A1(n14530), .A2(n13850), .ZN(n9693) );
  NAND2_X1 U12222 ( .A1(n9694), .A2(n9693), .ZN(n11601) );
  NAND2_X1 U12223 ( .A1(n11601), .A2(n12315), .ZN(n9696) );
  INV_X1 U12224 ( .A(n13849), .ZN(n12167) );
  OR2_X1 U12225 ( .A1(n14401), .A2(n12167), .ZN(n9695) );
  NAND2_X1 U12226 ( .A1(n9696), .A2(n9695), .ZN(n11786) );
  INV_X1 U12227 ( .A(n12317), .ZN(n11790) );
  NAND2_X1 U12228 ( .A1(n11786), .A2(n11790), .ZN(n9698) );
  OR2_X1 U12229 ( .A1(n12171), .A2(n12166), .ZN(n9697) );
  INV_X1 U12230 ( .A(n12179), .ZN(n9699) );
  INV_X1 U12231 ( .A(n14330), .ZN(n14227) );
  XNOR2_X1 U12232 ( .A(n12204), .B(n14220), .ZN(n14203) );
  NAND2_X1 U12233 ( .A1(n14202), .A2(n13845), .ZN(n9701) );
  XNOR2_X1 U12234 ( .A(n14193), .B(n13774), .ZN(n12319) );
  INV_X1 U12235 ( .A(n12319), .ZN(n14185) );
  NAND2_X1 U12236 ( .A1(n14318), .A2(n14206), .ZN(n9702) );
  NAND2_X1 U12237 ( .A1(n14184), .A2(n9702), .ZN(n14172) );
  INV_X1 U12238 ( .A(n13844), .ZN(n13740) );
  OR2_X1 U12239 ( .A1(n14304), .A2(n13740), .ZN(n14140) );
  NAND2_X1 U12240 ( .A1(n9703), .A2(n14134), .ZN(n14142) );
  NAND2_X1 U12241 ( .A1(n14149), .A2(n14152), .ZN(n9704) );
  NAND2_X1 U12242 ( .A1(n14142), .A2(n9704), .ZN(n14117) );
  OR2_X2 U12243 ( .A1(n14117), .A2(n14118), .ZN(n14124) );
  INV_X1 U12244 ( .A(n14121), .ZN(n13802) );
  AND2_X1 U12245 ( .A1(n14291), .A2(n13802), .ZN(n9706) );
  INV_X1 U12246 ( .A(n13842), .ZN(n13721) );
  OR2_X1 U12247 ( .A1(n14097), .A2(n13721), .ZN(n9707) );
  INV_X1 U12248 ( .A(n14077), .ZN(n14282) );
  INV_X1 U12249 ( .A(n14056), .ZN(n14047) );
  INV_X1 U12250 ( .A(n14270), .ZN(n14041) );
  INV_X1 U12251 ( .A(n14034), .ZN(n9709) );
  NAND2_X1 U12252 ( .A1(n14371), .A2(n14143), .ZN(n9712) );
  INV_X1 U12253 ( .A(n12275), .ZN(n12090) );
  NAND2_X1 U12254 ( .A1(n12273), .A2(n12090), .ZN(n9711) );
  NAND2_X2 U12255 ( .A1(n9712), .A2(n9711), .ZN(n14611) );
  AND2_X2 U12256 ( .A1(n14621), .A2(n11995), .ZN(n11991) );
  INV_X1 U12257 ( .A(n14696), .ZN(n11311) );
  NAND2_X1 U12258 ( .A1(n11991), .A2(n11311), .ZN(n11161) );
  NOR2_X1 U12259 ( .A1(n11159), .A2(n12132), .ZN(n11274) );
  INV_X1 U12260 ( .A(n12141), .ZN(n11500) );
  INV_X1 U12261 ( .A(n12150), .ZN(n14603) );
  OR2_X2 U12262 ( .A1(n14513), .A2(n14518), .ZN(n14519) );
  OR2_X2 U12263 ( .A1(n14334), .A2(n14519), .ZN(n14240) );
  AND2_X2 U12264 ( .A1(n14225), .A2(n14202), .ZN(n14198) );
  NAND2_X1 U12265 ( .A1(n14041), .A2(n14051), .ZN(n14036) );
  OR2_X2 U12266 ( .A1(n14036), .A2(n14265), .ZN(n12056) );
  NOR2_X2 U12267 ( .A1(n14260), .A2(n12056), .ZN(n14026) );
  AOI211_X1 U12268 ( .C1(n14260), .C2(n12056), .A(n14242), .B(n14026), .ZN(
        n14258) );
  INV_X1 U12269 ( .A(n14260), .ZN(n9727) );
  INV_X1 U12270 ( .A(n12273), .ZN(n12089) );
  NAND2_X1 U12271 ( .A1(n12089), .A2(n12090), .ZN(n12332) );
  INV_X1 U12272 ( .A(n12332), .ZN(n9714) );
  NAND2_X1 U12273 ( .A1(n10237), .A2(n9714), .ZN(n14630) );
  INV_X1 U12274 ( .A(n9715), .ZN(n9724) );
  NOR2_X1 U12275 ( .A1(n14370), .A2(n9716), .ZN(n9717) );
  NOR2_X1 U12276 ( .A1(n14221), .A2(n9717), .ZN(n14022) );
  INV_X1 U12277 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U12278 ( .A1(n9718), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U12279 ( .A1(n9719), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9720) );
  OAI211_X1 U12280 ( .C1(n12264), .C2(n9722), .A(n9721), .B(n9720), .ZN(n13838) );
  AND2_X1 U12281 ( .A1(n14022), .A2(n13838), .ZN(n14259) );
  AOI22_X1 U12282 ( .A1(n9724), .A2(n14259), .B1(n9723), .B2(n14599), .ZN(
        n9726) );
  NAND2_X1 U12283 ( .A1(n14642), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9725) );
  OAI211_X1 U12284 ( .C1(n9727), .C2(n14616), .A(n9726), .B(n9725), .ZN(n9728)
         );
  NAND2_X1 U12285 ( .A1(n10619), .A2(n10723), .ZN(n9971) );
  NAND2_X1 U12286 ( .A1(n9733), .A2(n9735), .ZN(n9736) );
  NAND2_X1 U12287 ( .A1(n9737), .A2(n9736), .ZN(n9739) );
  NAND3_X1 U12288 ( .A1(n9734), .A2(n10723), .A3(n9906), .ZN(n9738) );
  NAND2_X1 U12289 ( .A1(n13325), .A2(n9749), .ZN(n9742) );
  NAND2_X1 U12290 ( .A1(n9743), .A2(n6560), .ZN(n9741) );
  NAND2_X1 U12291 ( .A1(n9742), .A2(n9741), .ZN(n9746) );
  AOI22_X1 U12292 ( .A1(n13325), .A2(n9743), .B1(n6560), .B2(n9906), .ZN(n9744) );
  INV_X1 U12293 ( .A(n9745), .ZN(n9748) );
  NAND2_X1 U12294 ( .A1(n13323), .A2(n9937), .ZN(n9751) );
  NAND2_X1 U12295 ( .A1(n14831), .A2(n9906), .ZN(n9750) );
  NAND2_X1 U12296 ( .A1(n9751), .A2(n9750), .ZN(n9753) );
  AOI22_X1 U12297 ( .A1(n13323), .A2(n9906), .B1(n9880), .B2(n14831), .ZN(
        n9752) );
  NAND2_X1 U12298 ( .A1(n13322), .A2(n9906), .ZN(n9755) );
  NAND2_X1 U12299 ( .A1(n14837), .A2(n9937), .ZN(n9754) );
  NAND2_X1 U12300 ( .A1(n9755), .A2(n9754), .ZN(n9757) );
  INV_X1 U12301 ( .A(n9906), .ZN(n9800) );
  AOI22_X1 U12302 ( .A1(n13322), .A2(n9937), .B1(n14837), .B2(n9906), .ZN(
        n9756) );
  NAND2_X1 U12303 ( .A1(n14848), .A2(n9906), .ZN(n9759) );
  NAND2_X1 U12304 ( .A1(n13321), .A2(n9937), .ZN(n9758) );
  NAND2_X1 U12305 ( .A1(n9759), .A2(n9758), .ZN(n9764) );
  NAND2_X1 U12306 ( .A1(n9763), .A2(n9764), .ZN(n9762) );
  NAND2_X1 U12307 ( .A1(n14848), .A2(n9937), .ZN(n9760) );
  OAI21_X1 U12308 ( .B1(n10659), .B2(n9800), .A(n9760), .ZN(n9761) );
  NAND2_X1 U12309 ( .A1(n9762), .A2(n9761), .ZN(n9768) );
  INV_X1 U12310 ( .A(n9763), .ZN(n9766) );
  INV_X1 U12311 ( .A(n9764), .ZN(n9765) );
  NAND2_X1 U12312 ( .A1(n9766), .A2(n9765), .ZN(n9767) );
  NAND2_X1 U12313 ( .A1(n9768), .A2(n9767), .ZN(n9773) );
  NAND2_X1 U12314 ( .A1(n10919), .A2(n9937), .ZN(n9770) );
  NAND2_X1 U12315 ( .A1(n13320), .A2(n9906), .ZN(n9769) );
  NAND2_X1 U12316 ( .A1(n9770), .A2(n9769), .ZN(n9772) );
  AOI22_X1 U12317 ( .A1(n10919), .A2(n9906), .B1(n9880), .B2(n13320), .ZN(
        n9771) );
  NAND2_X1 U12318 ( .A1(n10835), .A2(n9906), .ZN(n9775) );
  NAND2_X1 U12319 ( .A1(n13319), .A2(n9937), .ZN(n9774) );
  NAND2_X1 U12320 ( .A1(n9775), .A2(n9774), .ZN(n9778) );
  INV_X1 U12321 ( .A(n13319), .ZN(n10834) );
  NAND2_X1 U12322 ( .A1(n10835), .A2(n9800), .ZN(n9776) );
  OAI21_X1 U12323 ( .B1(n10834), .B2(n9937), .A(n9776), .ZN(n9777) );
  NAND2_X1 U12324 ( .A1(n6661), .A2(n9779), .ZN(n9784) );
  NAND2_X1 U12325 ( .A1(n14796), .A2(n9937), .ZN(n9781) );
  NAND2_X1 U12326 ( .A1(n13318), .A2(n9906), .ZN(n9780) );
  INV_X1 U12327 ( .A(n13318), .ZN(n10972) );
  NAND2_X1 U12328 ( .A1(n14796), .A2(n9906), .ZN(n9782) );
  OAI21_X1 U12329 ( .B1(n10972), .B2(n9906), .A(n9782), .ZN(n9783) );
  NAND2_X1 U12330 ( .A1(n11141), .A2(n9906), .ZN(n9786) );
  NAND2_X1 U12331 ( .A1(n13317), .A2(n9800), .ZN(n9785) );
  NAND2_X1 U12332 ( .A1(n9786), .A2(n9785), .ZN(n9788) );
  INV_X1 U12333 ( .A(n9788), .ZN(n9787) );
  INV_X1 U12334 ( .A(n13317), .ZN(n11140) );
  NAND2_X1 U12335 ( .A1(n11141), .A2(n9937), .ZN(n9789) );
  OAI21_X1 U12336 ( .B1(n11140), .B2(n9937), .A(n9789), .ZN(n9790) );
  NAND2_X1 U12337 ( .A1(n11334), .A2(n9937), .ZN(n9792) );
  NAND2_X1 U12338 ( .A1(n13316), .A2(n9906), .ZN(n9791) );
  NAND2_X1 U12339 ( .A1(n9792), .A2(n9791), .ZN(n9795) );
  AOI22_X1 U12340 ( .A1(n11334), .A2(n9906), .B1(n9880), .B2(n13316), .ZN(
        n9793) );
  NAND2_X1 U12341 ( .A1(n11190), .A2(n9906), .ZN(n9798) );
  NAND2_X1 U12342 ( .A1(n13315), .A2(n9937), .ZN(n9797) );
  NAND2_X1 U12343 ( .A1(n11190), .A2(n9800), .ZN(n9799) );
  OAI21_X1 U12344 ( .B1(n11152), .B2(n9800), .A(n9799), .ZN(n9801) );
  NAND2_X1 U12345 ( .A1(n11389), .A2(n9880), .ZN(n9803) );
  NAND2_X1 U12346 ( .A1(n13314), .A2(n9906), .ZN(n9802) );
  AOI22_X1 U12347 ( .A1(n11389), .A2(n9906), .B1(n9880), .B2(n13314), .ZN(
        n9804) );
  NAND2_X1 U12348 ( .A1(n13667), .A2(n9749), .ZN(n9806) );
  NAND2_X1 U12349 ( .A1(n13313), .A2(n9880), .ZN(n9805) );
  AOI22_X1 U12350 ( .A1(n13667), .A2(n9937), .B1(n13313), .B2(n9906), .ZN(
        n9807) );
  NAND2_X1 U12351 ( .A1(n11692), .A2(n9800), .ZN(n9810) );
  NAND2_X1 U12352 ( .A1(n13312), .A2(n9906), .ZN(n9809) );
  INV_X1 U12353 ( .A(n13312), .ZN(n11691) );
  NAND2_X1 U12354 ( .A1(n11692), .A2(n9906), .ZN(n9811) );
  OAI21_X1 U12355 ( .B1(n11691), .B2(n9906), .A(n9811), .ZN(n9812) );
  NAND2_X1 U12356 ( .A1(n9813), .A2(n9812), .ZN(n9815) );
  NAND2_X1 U12357 ( .A1(n13661), .A2(n9749), .ZN(n9817) );
  NAND2_X1 U12358 ( .A1(n13311), .A2(n9880), .ZN(n9816) );
  AOI22_X1 U12359 ( .A1(n13661), .A2(n9937), .B1(n13311), .B2(n9906), .ZN(
        n9818) );
  NAND2_X1 U12360 ( .A1(n13656), .A2(n9800), .ZN(n9820) );
  NAND2_X1 U12361 ( .A1(n13310), .A2(n9906), .ZN(n9819) );
  NAND2_X1 U12362 ( .A1(n9820), .A2(n9819), .ZN(n9825) );
  AND2_X1 U12363 ( .A1(n13309), .A2(n9800), .ZN(n9821) );
  AOI21_X1 U12364 ( .B1(n11884), .B2(n9906), .A(n9821), .ZN(n9829) );
  NAND2_X1 U12365 ( .A1(n11884), .A2(n9880), .ZN(n9823) );
  NAND2_X1 U12366 ( .A1(n13309), .A2(n9906), .ZN(n9822) );
  NAND2_X1 U12367 ( .A1(n9823), .A2(n9822), .ZN(n9828) );
  AOI22_X1 U12368 ( .A1(n13656), .A2(n9906), .B1(n9880), .B2(n13310), .ZN(
        n9824) );
  AOI22_X1 U12369 ( .A1(n13651), .A2(n9906), .B1(n9880), .B2(n13308), .ZN(
        n9830) );
  NAND2_X1 U12370 ( .A1(n13651), .A2(n9880), .ZN(n9827) );
  NAND2_X1 U12371 ( .A1(n13308), .A2(n9906), .ZN(n9826) );
  NAND2_X1 U12372 ( .A1(n9827), .A2(n9826), .ZN(n9833) );
  AOI22_X1 U12373 ( .A1(n9830), .A2(n9833), .B1(n9829), .B2(n9828), .ZN(n9831)
         );
  NOR2_X1 U12374 ( .A1(n13651), .A2(n13308), .ZN(n9832) );
  NAND2_X1 U12375 ( .A1(n13645), .A2(n9906), .ZN(n9836) );
  NAND2_X1 U12376 ( .A1(n13541), .A2(n9880), .ZN(n9835) );
  NAND2_X1 U12377 ( .A1(n9836), .A2(n9835), .ZN(n9839) );
  INV_X1 U12378 ( .A(n13541), .ZN(n12002) );
  NAND2_X1 U12379 ( .A1(n13645), .A2(n9800), .ZN(n9837) );
  OAI21_X1 U12380 ( .B1(n12002), .B2(n9937), .A(n9837), .ZN(n9838) );
  INV_X1 U12381 ( .A(n9839), .ZN(n9840) );
  NAND2_X1 U12382 ( .A1(n13640), .A2(n9800), .ZN(n9842) );
  NAND2_X1 U12383 ( .A1(n13307), .A2(n9749), .ZN(n9841) );
  AOI22_X1 U12384 ( .A1(n13640), .A2(n9906), .B1(n9880), .B2(n13307), .ZN(
        n9843) );
  NAND2_X1 U12385 ( .A1(n13635), .A2(n9749), .ZN(n9846) );
  NAND2_X1 U12386 ( .A1(n13539), .A2(n9880), .ZN(n9845) );
  NAND2_X1 U12387 ( .A1(n9846), .A2(n9845), .ZN(n9849) );
  AOI22_X1 U12388 ( .A1(n13635), .A2(n9937), .B1(n13539), .B2(n9906), .ZN(
        n9847) );
  INV_X1 U12389 ( .A(n9848), .ZN(n9851) );
  NAND2_X1 U12390 ( .A1(n13629), .A2(n9800), .ZN(n9853) );
  NAND2_X1 U12391 ( .A1(n13485), .A2(n9906), .ZN(n9852) );
  NAND2_X1 U12392 ( .A1(n9853), .A2(n9852), .ZN(n9855) );
  AOI22_X1 U12393 ( .A1(n13629), .A2(n9906), .B1(n9880), .B2(n13485), .ZN(
        n9854) );
  NAND2_X1 U12394 ( .A1(n13621), .A2(n9749), .ZN(n9858) );
  NAND2_X1 U12395 ( .A1(n13502), .A2(n9880), .ZN(n9857) );
  NAND2_X1 U12396 ( .A1(n9858), .A2(n9857), .ZN(n9860) );
  INV_X1 U12397 ( .A(n13502), .ZN(n13237) );
  NAND2_X1 U12398 ( .A1(n13621), .A2(n9880), .ZN(n9859) );
  OAI21_X1 U12399 ( .B1(n13237), .B2(n9937), .A(n9859), .ZN(n9861) );
  NAND2_X1 U12400 ( .A1(n13614), .A2(n9880), .ZN(n9863) );
  NAND2_X1 U12401 ( .A1(n13484), .A2(n9749), .ZN(n9862) );
  AOI22_X1 U12402 ( .A1(n13614), .A2(n9749), .B1(n9880), .B2(n13484), .ZN(
        n9864) );
  INV_X1 U12403 ( .A(n9864), .ZN(n9865) );
  NAND2_X1 U12404 ( .A1(n9866), .A2(n7693), .ZN(n9867) );
  NAND2_X1 U12405 ( .A1(n13607), .A2(n9906), .ZN(n9870) );
  NAND2_X1 U12406 ( .A1(n13471), .A2(n9880), .ZN(n9869) );
  NAND2_X1 U12407 ( .A1(n9870), .A2(n9869), .ZN(n9874) );
  NAND2_X1 U12408 ( .A1(n13607), .A2(n9880), .ZN(n9872) );
  NAND2_X1 U12409 ( .A1(n13471), .A2(n9749), .ZN(n9871) );
  NAND2_X1 U12410 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  NAND2_X1 U12411 ( .A1(n13603), .A2(n9880), .ZN(n9876) );
  NAND2_X1 U12412 ( .A1(n13456), .A2(n9749), .ZN(n9875) );
  NAND2_X1 U12413 ( .A1(n9876), .A2(n9875), .ZN(n9882) );
  AND2_X1 U12414 ( .A1(n13448), .A2(n9800), .ZN(n9877) );
  AOI21_X1 U12415 ( .B1(n13598), .B2(n9906), .A(n9877), .ZN(n9918) );
  NAND2_X1 U12416 ( .A1(n13598), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U12417 ( .A1(n13448), .A2(n9749), .ZN(n9878) );
  NAND2_X1 U12418 ( .A1(n9879), .A2(n9878), .ZN(n9917) );
  OAI22_X1 U12419 ( .A1(n9883), .A2(n9882), .B1(n9918), .B2(n9917), .ZN(n9952)
         );
  AOI22_X1 U12420 ( .A1(n13603), .A2(n9906), .B1(n9880), .B2(n13456), .ZN(
        n9881) );
  AOI21_X1 U12421 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9916) );
  NAND2_X1 U12422 ( .A1(n9885), .A2(n9884), .ZN(n9888) );
  INV_X1 U12423 ( .A(SI_29_), .ZN(n13206) );
  NAND2_X1 U12424 ( .A1(n9886), .A2(n13206), .ZN(n9887) );
  NAND2_X1 U12425 ( .A1(n9888), .A2(n9887), .ZN(n9925) );
  MUX2_X1 U12426 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10025), .Z(n9889) );
  XNOR2_X1 U12427 ( .A(n9889), .B(SI_30_), .ZN(n9923) );
  NAND2_X1 U12428 ( .A1(n9889), .A2(SI_30_), .ZN(n9890) );
  OAI21_X1 U12429 ( .B1(n9925), .B2(n9923), .A(n9890), .ZN(n9893) );
  MUX2_X1 U12430 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10006), .Z(n9891) );
  XNOR2_X1 U12431 ( .A(n9891), .B(SI_31_), .ZN(n9892) );
  XNOR2_X1 U12432 ( .A(n9893), .B(n9892), .ZN(n13690) );
  NAND2_X1 U12433 ( .A1(n13690), .A2(n9894), .ZN(n9896) );
  NAND2_X1 U12434 ( .A1(n9926), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U12435 ( .A1(n9896), .A2(n9895), .ZN(n9921) );
  INV_X1 U12436 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U12437 ( .A1(n8380), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U12438 ( .A1(n6565), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9897) );
  OAI211_X1 U12439 ( .C1(n9900), .C2(n9899), .A(n9898), .B(n9897), .ZN(n13378)
         );
  INV_X1 U12440 ( .A(n13378), .ZN(n9956) );
  XNOR2_X1 U12441 ( .A(n9921), .B(n9956), .ZN(n9944) );
  AND2_X1 U12442 ( .A1(n13414), .A2(n9800), .ZN(n9901) );
  AOI21_X1 U12443 ( .B1(n13586), .B2(n9749), .A(n9901), .ZN(n9947) );
  NAND2_X1 U12444 ( .A1(n13586), .A2(n9937), .ZN(n9903) );
  NAND2_X1 U12445 ( .A1(n13414), .A2(n9906), .ZN(n9902) );
  NAND2_X1 U12446 ( .A1(n9903), .A2(n9902), .ZN(n9945) );
  NAND2_X1 U12447 ( .A1(n13694), .A2(n9894), .ZN(n9905) );
  NAND2_X1 U12448 ( .A1(n9926), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9904) );
  AND2_X1 U12449 ( .A1(n13392), .A2(n9906), .ZN(n9907) );
  AOI21_X1 U12450 ( .B1(n13583), .B2(n9937), .A(n9907), .ZN(n9941) );
  NAND2_X1 U12451 ( .A1(n13583), .A2(n9749), .ZN(n9909) );
  NAND2_X1 U12452 ( .A1(n13392), .A2(n9880), .ZN(n9908) );
  NAND2_X1 U12453 ( .A1(n9909), .A2(n9908), .ZN(n9940) );
  NAND2_X1 U12454 ( .A1(n9941), .A2(n9940), .ZN(n9946) );
  OAI21_X1 U12455 ( .B1(n9947), .B2(n9945), .A(n9946), .ZN(n9910) );
  NAND2_X1 U12456 ( .A1(n13591), .A2(n9880), .ZN(n9912) );
  NAND2_X1 U12457 ( .A1(n13428), .A2(n9749), .ZN(n9911) );
  NAND2_X1 U12458 ( .A1(n9912), .A2(n9911), .ZN(n9919) );
  INV_X1 U12459 ( .A(n9919), .ZN(n9915) );
  AND2_X1 U12460 ( .A1(n13428), .A2(n9880), .ZN(n9913) );
  AOI21_X1 U12461 ( .B1(n13591), .B2(n9906), .A(n9913), .ZN(n9920) );
  INV_X1 U12462 ( .A(n9920), .ZN(n9914) );
  NAND2_X1 U12463 ( .A1(n9920), .A2(n9919), .ZN(n9950) );
  NAND2_X1 U12464 ( .A1(n13378), .A2(n9800), .ZN(n9958) );
  OAI211_X1 U12465 ( .C1(n9921), .C2(n13378), .A(n9958), .B(n9922), .ZN(n9943)
         );
  INV_X1 U12466 ( .A(n9923), .ZN(n9924) );
  NAND2_X1 U12467 ( .A1(n12260), .A2(n9894), .ZN(n9928) );
  NAND2_X1 U12468 ( .A1(n9926), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9927) );
  NAND2_X1 U12469 ( .A1(n13378), .A2(n9906), .ZN(n9930) );
  NOR2_X1 U12470 ( .A1(n12069), .A2(n13373), .ZN(n10629) );
  NAND2_X1 U12471 ( .A1(n10629), .A2(n11176), .ZN(n9964) );
  NAND3_X1 U12472 ( .A1(n9930), .A2(n9929), .A3(n9964), .ZN(n9935) );
  INV_X1 U12473 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U12474 ( .A1(n8380), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U12475 ( .A1(n9931), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9932) );
  OAI211_X1 U12476 ( .C1(n8463), .C2(n9934), .A(n9933), .B(n9932), .ZN(n13306)
         );
  AND2_X1 U12477 ( .A1(n9935), .A2(n13306), .ZN(n9936) );
  AOI21_X1 U12478 ( .B1(n13382), .B2(n9937), .A(n9936), .ZN(n9954) );
  NAND2_X1 U12479 ( .A1(n13382), .A2(n9906), .ZN(n9939) );
  NAND2_X1 U12480 ( .A1(n13306), .A2(n9880), .ZN(n9938) );
  NAND2_X1 U12481 ( .A1(n9939), .A2(n9938), .ZN(n9953) );
  OAI22_X1 U12482 ( .A1(n9954), .A2(n9953), .B1(n9941), .B2(n9940), .ZN(n9942)
         );
  NAND2_X1 U12483 ( .A1(n9943), .A2(n9942), .ZN(n9949) );
  INV_X1 U12484 ( .A(n9944), .ZN(n9984) );
  NAND4_X1 U12485 ( .A1(n9984), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n9948)
         );
  NAND2_X1 U12486 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  NAND2_X1 U12487 ( .A1(n9956), .A2(n9749), .ZN(n9957) );
  MUX2_X1 U12488 ( .A(n9958), .B(n9957), .S(n9921), .Z(n9959) );
  AOI21_X1 U12489 ( .B1(n11360), .B2(n9988), .A(n10646), .ZN(n9961) );
  INV_X1 U12490 ( .A(n9962), .ZN(n9963) );
  AND2_X1 U12491 ( .A1(n8377), .A2(n9988), .ZN(n10628) );
  INV_X1 U12492 ( .A(n9964), .ZN(n9965) );
  AOI21_X1 U12493 ( .B1(n10646), .B2(n10628), .A(n9965), .ZN(n9966) );
  INV_X1 U12494 ( .A(n10142), .ZN(n9996) );
  NAND2_X1 U12495 ( .A1(n9996), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11670) );
  INV_X1 U12496 ( .A(n11670), .ZN(n9967) );
  NAND2_X1 U12497 ( .A1(n13586), .A2(n13414), .ZN(n12038) );
  OR2_X1 U12498 ( .A1(n13586), .A2(n13414), .ZN(n9968) );
  INV_X1 U12499 ( .A(n13428), .ZN(n13298) );
  XNOR2_X1 U12500 ( .A(n13591), .B(n13298), .ZN(n12013) );
  INV_X1 U12501 ( .A(n13456), .ZN(n13294) );
  INV_X1 U12502 ( .A(n13448), .ZN(n9969) );
  OR2_X1 U12503 ( .A1(n13598), .A2(n9969), .ZN(n12010) );
  NAND2_X1 U12504 ( .A1(n13598), .A2(n9969), .ZN(n12011) );
  INV_X1 U12505 ( .A(n13471), .ZN(n12009) );
  XNOR2_X1 U12506 ( .A(n13607), .B(n12009), .ZN(n13459) );
  XNOR2_X1 U12507 ( .A(n13629), .B(n13523), .ZN(n13509) );
  INV_X1 U12508 ( .A(n13539), .ZN(n13236) );
  OR2_X1 U12509 ( .A1(n13635), .A2(n13236), .ZN(n12007) );
  NAND2_X1 U12510 ( .A1(n13635), .A2(n13236), .ZN(n13500) );
  NAND2_X1 U12511 ( .A1(n12007), .A2(n13500), .ZN(n13518) );
  OR2_X1 U12512 ( .A1(n13640), .A2(n13307), .ZN(n12025) );
  NAND2_X1 U12513 ( .A1(n13640), .A2(n13307), .ZN(n12024) );
  NAND2_X1 U12514 ( .A1(n12025), .A2(n12024), .ZN(n13535) );
  INV_X1 U12515 ( .A(n13308), .ZN(n11999) );
  XNOR2_X1 U12516 ( .A(n13651), .B(n11999), .ZN(n12019) );
  INV_X1 U12517 ( .A(n13311), .ZN(n11758) );
  INV_X1 U12518 ( .A(n13309), .ZN(n11883) );
  XNOR2_X1 U12519 ( .A(n11884), .B(n11883), .ZN(n11851) );
  XNOR2_X1 U12520 ( .A(n11692), .B(n13312), .ZN(n11430) );
  XNOR2_X1 U12521 ( .A(n11190), .B(n11152), .ZN(n11179) );
  XNOR2_X1 U12522 ( .A(n11334), .B(n11181), .ZN(n11144) );
  XNOR2_X1 U12523 ( .A(n11141), .B(n11140), .ZN(n10975) );
  XNOR2_X1 U12524 ( .A(n14796), .B(n13318), .ZN(n10838) );
  NAND2_X1 U12525 ( .A1(n10801), .A2(n14831), .ZN(n10782) );
  NAND2_X1 U12526 ( .A1(n13323), .A2(n10776), .ZN(n9970) );
  NAND2_X1 U12527 ( .A1(n9971), .A2(n10607), .ZN(n10722) );
  NAND4_X1 U12528 ( .A1(n10803), .A2(n10768), .A3(n9988), .A4(n10722), .ZN(
        n9973) );
  NAND2_X1 U12529 ( .A1(n10795), .A2(n13322), .ZN(n9972) );
  NOR3_X1 U12530 ( .A1(n9973), .A2(n10752), .A3(n10783), .ZN(n9974) );
  XNOR2_X1 U12531 ( .A(n10835), .B(n13319), .ZN(n10832) );
  XNOR2_X1 U12532 ( .A(n10919), .B(n13320), .ZN(n10921) );
  NAND4_X1 U12533 ( .A1(n10838), .A2(n9974), .A3(n10832), .A4(n10921), .ZN(
        n9975) );
  NOR4_X1 U12534 ( .A1(n11179), .A2(n11144), .A3(n10975), .A4(n9975), .ZN(
        n9976) );
  XNOR2_X1 U12535 ( .A(n13667), .B(n13313), .ZN(n11253) );
  XNOR2_X1 U12536 ( .A(n11389), .B(n13314), .ZN(n11150) );
  NAND4_X1 U12537 ( .A1(n11430), .A2(n9976), .A3(n11253), .A4(n11150), .ZN(
        n9977) );
  NOR4_X1 U12538 ( .A1(n12019), .A2(n11725), .A3(n11851), .A4(n9977), .ZN(
        n9978) );
  XNOR2_X1 U12539 ( .A(n13645), .B(n13541), .ZN(n13565) );
  XNOR2_X1 U12540 ( .A(n13656), .B(n13310), .ZN(n11854) );
  NAND4_X1 U12541 ( .A1(n13535), .A2(n9978), .A3(n13565), .A4(n11854), .ZN(
        n9979) );
  NOR4_X1 U12542 ( .A1(n13459), .A2(n13509), .A3(n13518), .A4(n9979), .ZN(
        n9980) );
  XNOR2_X1 U12543 ( .A(n13614), .B(n13484), .ZN(n13478) );
  XNOR2_X1 U12544 ( .A(n13621), .B(n13502), .ZN(n13495) );
  NAND4_X1 U12545 ( .A1(n13431), .A2(n9980), .A3(n13478), .A4(n13495), .ZN(
        n9981) );
  NOR4_X1 U12546 ( .A1(n13398), .A2(n12013), .A3(n13446), .A4(n9981), .ZN(
        n9983) );
  XNOR2_X1 U12547 ( .A(n13382), .B(n13306), .ZN(n9982) );
  XNOR2_X1 U12548 ( .A(n13583), .B(n13392), .ZN(n12039) );
  NAND4_X1 U12549 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n12039), .ZN(n9985) );
  XOR2_X1 U12550 ( .A(n10646), .B(n9985), .Z(n9986) );
  NOR3_X1 U12551 ( .A1(n9986), .A2(n8377), .A3(n11670), .ZN(n9987) );
  OAI21_X1 U12552 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(n9995) );
  INV_X1 U12553 ( .A(n12050), .ZN(n12015) );
  INV_X1 U12554 ( .A(n9990), .ZN(n9991) );
  NAND4_X1 U12555 ( .A1(n14818), .A2(n12015), .A3(n9991), .A4(n13540), .ZN(
        n9992) );
  OAI211_X1 U12556 ( .C1(n9993), .C2(n11670), .A(n9992), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9994) );
  AOI211_X1 U12557 ( .C1(n10001), .C2(n10000), .A(n14427), .B(n9999), .ZN(
        n10004) );
  MUX2_X1 U12558 ( .A(n14444), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n10003) );
  AOI22_X1 U12559 ( .A1(n15061), .A2(n15063), .B1(n12780), .B2(n15064), .ZN(
        n10869) );
  OAI22_X1 U12560 ( .A1(n12574), .A2(n15089), .B1(n10869), .B2(n14446), .ZN(
        n10002) );
  OR3_X1 U12561 ( .A1(n10004), .A2(n10003), .A3(n10002), .ZN(P3_U3158) );
  NOR2_X1 U12562 ( .A1(n10025), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13698) );
  INV_X2 U12563 ( .A(n13698), .ZN(n12073) );
  INV_X2 U12564 ( .A(n11668), .ZN(n12071) );
  OAI222_X1 U12565 ( .A1(n12073), .A2(n10005), .B1(n12071), .B2(n10051), .C1(
        P2_U3088), .C2(n10331), .ZN(P2_U3326) );
  INV_X2 U12566 ( .A(n14386), .ZN(n15456) );
  AND2_X1 U12567 ( .A1(n6566), .A2(P3_U3151), .ZN(n14387) );
  INV_X2 U12568 ( .A(n14387), .ZN(n15458) );
  OAI222_X1 U12569 ( .A1(P3_U3151), .A2(n6940), .B1(n15456), .B2(n10008), .C1(
        n15458), .C2(n10007), .ZN(P3_U3294) );
  INV_X1 U12570 ( .A(SI_4_), .ZN(n10009) );
  OAI222_X1 U12571 ( .A1(n15458), .A2(n10010), .B1(n15456), .B2(n10009), .C1(
        n11046), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12572 ( .A(SI_5_), .ZN(n10011) );
  OAI222_X1 U12573 ( .A1(n15458), .A2(n10012), .B1(n15456), .B2(n10011), .C1(
        n11053), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12574 ( .A(n14972), .ZN(n11060) );
  INV_X1 U12575 ( .A(SI_6_), .ZN(n10013) );
  OAI222_X1 U12576 ( .A1(n11060), .A2(P3_U3151), .B1(n15458), .B2(n10014), 
        .C1(n10013), .C2(n15456), .ZN(P3_U3289) );
  OAI222_X1 U12577 ( .A1(n11039), .A2(P3_U3151), .B1(n15458), .B2(n10015), 
        .C1(n6966), .C2(n15456), .ZN(P3_U3292) );
  INV_X1 U12578 ( .A(SI_2_), .ZN(n10016) );
  OAI222_X1 U12579 ( .A1(n6564), .A2(P3_U3151), .B1(n15458), .B2(n10017), .C1(
        n10016), .C2(n15456), .ZN(P3_U3293) );
  INV_X1 U12580 ( .A(n6922), .ZN(n10536) );
  INV_X1 U12581 ( .A(n10018), .ZN(n10020) );
  OAI222_X1 U12582 ( .A1(n10536), .A2(P3_U3151), .B1(n15458), .B2(n10020), 
        .C1(n10019), .C2(n15456), .ZN(P3_U3295) );
  OAI222_X1 U12583 ( .A1(n14986), .A2(P3_U3151), .B1(n15458), .B2(n10022), 
        .C1(n10021), .C2(n15456), .ZN(P3_U3288) );
  INV_X1 U12584 ( .A(SI_8_), .ZN(n10023) );
  OAI222_X1 U12585 ( .A1(n15458), .A2(n10024), .B1(n15456), .B2(n10023), .C1(
        n11072), .C2(P3_U3151), .ZN(P3_U3287) );
  NAND2_X1 U12586 ( .A1(n6566), .A2(P1_U3086), .ZN(n14369) );
  INV_X1 U12587 ( .A(n10026), .ZN(n10032) );
  INV_X1 U12588 ( .A(n13902), .ZN(n10027) );
  OAI222_X1 U12589 ( .A1(n14366), .A2(n10028), .B1(n14369), .B2(n10032), .C1(
        n10027), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U12590 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10030) );
  INV_X1 U12591 ( .A(n10029), .ZN(n10043) );
  INV_X1 U12592 ( .A(n10187), .ZN(n10200) );
  OAI222_X1 U12593 ( .A1(n12073), .A2(n10030), .B1(n12071), .B2(n10043), .C1(
        P2_U3088), .C2(n10200), .ZN(P2_U3322) );
  INV_X1 U12594 ( .A(n13335), .ZN(n10031) );
  OAI222_X1 U12595 ( .A1(n12073), .A2(n10033), .B1(n12071), .B2(n10032), .C1(
        P2_U3088), .C2(n10031), .ZN(P2_U3324) );
  INV_X1 U12596 ( .A(n10222), .ZN(n10230) );
  OAI222_X1 U12597 ( .A1(n12073), .A2(n10034), .B1(n12071), .B2(n10054), .C1(
        P2_U3088), .C2(n10230), .ZN(P2_U3325) );
  INV_X1 U12598 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10036) );
  INV_X1 U12599 ( .A(n10035), .ZN(n10041) );
  INV_X1 U12600 ( .A(n10174), .ZN(n10264) );
  OAI222_X1 U12601 ( .A1(n12073), .A2(n10036), .B1(n12071), .B2(n10041), .C1(
        P2_U3088), .C2(n10264), .ZN(P2_U3323) );
  OAI222_X1 U12602 ( .A1(n15458), .A2(n10037), .B1(n15456), .B2(n15294), .C1(
        n11462), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12603 ( .A(n10038), .ZN(n10046) );
  INV_X1 U12604 ( .A(n10176), .ZN(n14723) );
  OAI222_X1 U12605 ( .A1(n12073), .A2(n10039), .B1(n12071), .B2(n10046), .C1(
        P2_U3088), .C2(n14723), .ZN(P2_U3321) );
  INV_X1 U12606 ( .A(n14366), .ZN(n14360) );
  AOI22_X1 U12607 ( .A1(n13917), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n14360), .ZN(n10040) );
  OAI21_X1 U12608 ( .B1(n10041), .B2(n14369), .A(n10040), .ZN(P1_U3351) );
  AOI22_X1 U12609 ( .A1(n13927), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n14360), .ZN(n10042) );
  OAI21_X1 U12610 ( .B1(n10043), .B2(n14369), .A(n10042), .ZN(P1_U3350) );
  INV_X1 U12611 ( .A(n10044), .ZN(n10048) );
  INV_X1 U12612 ( .A(n10274), .ZN(n10186) );
  OAI222_X1 U12613 ( .A1(n12073), .A2(n10045), .B1(n12071), .B2(n10048), .C1(
        P2_U3088), .C2(n10186), .ZN(P2_U3320) );
  INV_X1 U12614 ( .A(n10105), .ZN(n10124) );
  OAI222_X1 U12615 ( .A1(n14366), .A2(n10047), .B1(n14369), .B2(n10046), .C1(
        n10124), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12616 ( .A(n14369), .ZN(n11665) );
  INV_X1 U12617 ( .A(n11665), .ZN(n12362) );
  INV_X1 U12618 ( .A(n13950), .ZN(n10119) );
  OAI222_X1 U12619 ( .A1(n14366), .A2(n10049), .B1(n12362), .B2(n10048), .C1(
        n10119), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U12620 ( .A(n13865), .ZN(n10050) );
  OAI222_X1 U12621 ( .A1(n14366), .A2(n10052), .B1(n12362), .B2(n10051), .C1(
        n10050), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U12622 ( .A(n13890), .ZN(n10055) );
  OAI222_X1 U12623 ( .A1(n10055), .A2(P1_U3086), .B1(n14369), .B2(n10054), 
        .C1(n10053), .C2(n14366), .ZN(P1_U3353) );
  NAND2_X1 U12624 ( .A1(n9734), .A2(P2_U3947), .ZN(n10056) );
  OAI21_X1 U12625 ( .B1(n9302), .B2(P2_U3947), .A(n10056), .ZN(P2_U3531) );
  INV_X1 U12626 ( .A(n10057), .ZN(n10059) );
  INV_X1 U12627 ( .A(n10276), .ZN(n14738) );
  OAI222_X1 U12628 ( .A1(n12073), .A2(n10058), .B1(n12071), .B2(n10059), .C1(
        P2_U3088), .C2(n14738), .ZN(P2_U3319) );
  INV_X1 U12629 ( .A(n10211), .ZN(n10205) );
  OAI222_X1 U12630 ( .A1(n14366), .A2(n10060), .B1(n12362), .B2(n10059), .C1(
        n10205), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U12631 ( .A(n10061), .ZN(n10064) );
  INV_X1 U12632 ( .A(n13968), .ZN(n10062) );
  OAI222_X1 U12633 ( .A1(n14366), .A2(n10063), .B1(n12362), .B2(n10064), .C1(
        n10062), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U12634 ( .A(n10396), .ZN(n10281) );
  OAI222_X1 U12635 ( .A1(n12073), .A2(n10065), .B1(n12071), .B2(n10064), .C1(
        P2_U3088), .C2(n10281), .ZN(P2_U3318) );
  INV_X1 U12636 ( .A(n12085), .ZN(n10067) );
  INV_X1 U12637 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n15307) );
  NOR2_X1 U12638 ( .A1(n10067), .A2(n15307), .ZN(P3_U3236) );
  INV_X1 U12639 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n15435) );
  NOR2_X1 U12640 ( .A1(n10067), .A2(n15435), .ZN(P3_U3235) );
  INV_X1 U12641 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15211) );
  NOR2_X1 U12642 ( .A1(n10067), .A2(n15211), .ZN(P3_U3253) );
  INV_X1 U12643 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n15354) );
  NOR2_X1 U12644 ( .A1(n10067), .A2(n15354), .ZN(P3_U3247) );
  INV_X1 U12645 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n15367) );
  NOR2_X1 U12646 ( .A1(n10067), .A2(n15367), .ZN(P3_U3239) );
  INV_X1 U12647 ( .A(n10363), .ZN(n10357) );
  OR3_X1 U12648 ( .A1(n10069), .A2(n10075), .A3(n11896), .ZN(n10070) );
  OAI21_X1 U12649 ( .B1(n14669), .B2(P1_D_REG_1__SCAN_IN), .A(n10070), .ZN(
        n10071) );
  INV_X1 U12650 ( .A(n10071), .ZN(P1_U3446) );
  INV_X1 U12651 ( .A(n11716), .ZN(n10073) );
  NAND2_X1 U12652 ( .A1(n10073), .A2(n10072), .ZN(n10074) );
  OAI22_X1 U12653 ( .A1(n14669), .A2(P1_D_REG_0__SCAN_IN), .B1(n10075), .B2(
        n10074), .ZN(n10076) );
  INV_X1 U12654 ( .A(n10076), .ZN(P1_U3445) );
  INV_X1 U12655 ( .A(n10077), .ZN(n10079) );
  OAI222_X1 U12656 ( .A1(n14366), .A2(n10078), .B1(n12362), .B2(n10079), .C1(
        n10297), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U12657 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10080) );
  INV_X1 U12658 ( .A(n10428), .ZN(n10403) );
  OAI222_X1 U12659 ( .A1(n12073), .A2(n10080), .B1(n12071), .B2(n10079), .C1(
        P2_U3088), .C2(n10403), .ZN(P2_U3317) );
  INV_X1 U12660 ( .A(n10081), .ZN(n10083) );
  OR2_X1 U12661 ( .A1(n12287), .A2(n10083), .ZN(n10082) );
  AND2_X1 U12662 ( .A1(n10082), .A2(n9305), .ZN(n10112) );
  NAND2_X1 U12663 ( .A1(n10083), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12349) );
  NAND2_X1 U12664 ( .A1(n10363), .A2(n12349), .ZN(n10113) );
  NAND2_X1 U12665 ( .A1(n10112), .A2(n10113), .ZN(n14570) );
  OR2_X1 U12666 ( .A1(n14570), .A2(n13878), .ZN(n14592) );
  MUX2_X1 U12667 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9308), .S(n13890), .Z(
        n10088) );
  MUX2_X1 U12668 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10084), .S(n13865), .Z(
        n10086) );
  AND2_X1 U12669 ( .A1(n14566), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U12670 ( .A1(n10086), .A2(n10085), .ZN(n13869) );
  NAND2_X1 U12671 ( .A1(n13865), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12672 ( .A1(n13869), .A2(n10087), .ZN(n13884) );
  NAND2_X1 U12673 ( .A1(n10088), .A2(n13884), .ZN(n13895) );
  NAND2_X1 U12674 ( .A1(n13890), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13894) );
  NAND2_X1 U12675 ( .A1(n13895), .A2(n13894), .ZN(n10091) );
  MUX2_X1 U12676 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10089), .S(n13902), .Z(
        n10090) );
  NAND2_X1 U12677 ( .A1(n10091), .A2(n10090), .ZN(n13909) );
  NAND2_X1 U12678 ( .A1(n13902), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13908) );
  MUX2_X1 U12679 ( .A(n9330), .B(P1_REG1_REG_4__SCAN_IN), .S(n13917), .Z(
        n13910) );
  AOI21_X1 U12680 ( .B1(n13909), .B2(n13908), .A(n13910), .ZN(n13907) );
  AOI21_X1 U12681 ( .B1(n13917), .B2(P1_REG1_REG_4__SCAN_IN), .A(n13907), .ZN(
        n13929) );
  INV_X1 U12682 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14714) );
  MUX2_X1 U12683 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n14714), .S(n13927), .Z(
        n13930) );
  NAND2_X1 U12684 ( .A1(n13929), .A2(n13930), .ZN(n13928) );
  OAI21_X1 U12685 ( .B1(n13927), .B2(P1_REG1_REG_5__SCAN_IN), .A(n13928), .ZN(
        n10093) );
  INV_X1 U12686 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14716) );
  MUX2_X1 U12687 ( .A(n14716), .B(P1_REG1_REG_6__SCAN_IN), .S(n10105), .Z(
        n10092) );
  NOR2_X1 U12688 ( .A1(n10093), .A2(n10092), .ZN(n13949) );
  INV_X1 U12689 ( .A(n14370), .ZN(n14564) );
  OR2_X1 U12690 ( .A1(n14570), .A2(n14564), .ZN(n14590) );
  AOI211_X1 U12691 ( .C1(n10093), .C2(n10092), .A(n13949), .B(n14590), .ZN(
        n10111) );
  NAND2_X1 U12692 ( .A1(n13878), .A2(n14564), .ZN(n10094) );
  MUX2_X1 U12693 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10095), .S(n13890), .Z(
        n13882) );
  MUX2_X1 U12694 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10096), .S(n13865), .Z(
        n13871) );
  AND2_X1 U12695 ( .A1(n14566), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13877) );
  NAND2_X1 U12696 ( .A1(n13871), .A2(n13877), .ZN(n13870) );
  NAND2_X1 U12697 ( .A1(n13865), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U12698 ( .A1(n13870), .A2(n10097), .ZN(n13881) );
  NAND2_X1 U12699 ( .A1(n13882), .A2(n13881), .ZN(n13899) );
  NAND2_X1 U12700 ( .A1(n13890), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U12701 ( .A1(n13899), .A2(n13898), .ZN(n10099) );
  MUX2_X1 U12702 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10819), .S(n13902), .Z(
        n10098) );
  NAND2_X1 U12703 ( .A1(n10099), .A2(n10098), .ZN(n13914) );
  NAND2_X1 U12704 ( .A1(n13902), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13913) );
  NAND2_X1 U12705 ( .A1(n13914), .A2(n13913), .ZN(n10102) );
  MUX2_X1 U12706 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10100), .S(n13917), .Z(
        n10101) );
  NAND2_X1 U12707 ( .A1(n10102), .A2(n10101), .ZN(n13934) );
  NAND2_X1 U12708 ( .A1(n13917), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13933) );
  INV_X1 U12709 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10103) );
  MUX2_X1 U12710 ( .A(n10103), .B(P1_REG2_REG_5__SCAN_IN), .S(n13927), .Z(
        n13932) );
  AOI21_X1 U12711 ( .B1(n13934), .B2(n13933), .A(n13932), .ZN(n10104) );
  INV_X1 U12712 ( .A(n10104), .ZN(n13936) );
  NAND2_X1 U12713 ( .A1(n13927), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10108) );
  INV_X1 U12714 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U12715 ( .A(n10106), .B(P1_REG2_REG_6__SCAN_IN), .S(n10105), .Z(
        n10107) );
  AOI21_X1 U12716 ( .B1(n13936), .B2(n10108), .A(n10107), .ZN(n13956) );
  AND3_X1 U12717 ( .A1(n13936), .A2(n10108), .A3(n10107), .ZN(n10109) );
  NOR3_X1 U12718 ( .A1(n14588), .A2(n13956), .A3(n10109), .ZN(n10110) );
  NOR2_X1 U12719 ( .A1(n10111), .A2(n10110), .ZN(n10116) );
  INV_X1 U12720 ( .A(n10112), .ZN(n10114) );
  AND2_X1 U12721 ( .A1(n10114), .A2(n10113), .ZN(n14568) );
  NOR2_X1 U12722 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9361), .ZN(n11304) );
  AOI21_X1 U12723 ( .B1(n14568), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11304), .ZN(
        n10115) );
  OAI211_X1 U12724 ( .C1(n10124), .C2(n14592), .A(n10116), .B(n10115), .ZN(
        P1_U3249) );
  INV_X1 U12725 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10117) );
  MUX2_X1 U12726 ( .A(n10117), .B(P1_REG1_REG_8__SCAN_IN), .S(n10211), .Z(
        n10121) );
  INV_X1 U12727 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n13943) );
  NOR2_X1 U12728 ( .A1(n10124), .A2(n14716), .ZN(n13944) );
  MUX2_X1 U12729 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n13943), .S(n13950), .Z(
        n10118) );
  OAI21_X1 U12730 ( .B1(n13949), .B2(n13944), .A(n10118), .ZN(n13947) );
  OAI21_X1 U12731 ( .B1(n13943), .B2(n10119), .A(n13947), .ZN(n10120) );
  NOR2_X1 U12732 ( .A1(n10120), .A2(n10121), .ZN(n13963) );
  AOI21_X1 U12733 ( .B1(n10121), .B2(n10120), .A(n13963), .ZN(n10134) );
  NAND2_X1 U12734 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11582) );
  OAI21_X1 U12735 ( .B1(n14596), .B2(n10122), .A(n11582), .ZN(n10123) );
  AOI21_X1 U12736 ( .B1(n10211), .B2(n13984), .A(n10123), .ZN(n10133) );
  NOR2_X1 U12737 ( .A1(n10124), .A2(n10106), .ZN(n13951) );
  INV_X1 U12738 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10125) );
  MUX2_X1 U12739 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10125), .S(n13950), .Z(
        n10126) );
  OAI21_X1 U12740 ( .B1(n13956), .B2(n13951), .A(n10126), .ZN(n13954) );
  NAND2_X1 U12741 ( .A1(n13950), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10129) );
  INV_X1 U12742 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10127) );
  MUX2_X1 U12743 ( .A(n10127), .B(P1_REG2_REG_8__SCAN_IN), .S(n10211), .Z(
        n10128) );
  AOI21_X1 U12744 ( .B1(n13954), .B2(n10129), .A(n10128), .ZN(n13974) );
  INV_X1 U12745 ( .A(n13974), .ZN(n10131) );
  NAND3_X1 U12746 ( .A1(n13954), .A2(n10129), .A3(n10128), .ZN(n10130) );
  NAND3_X1 U12747 ( .A1(n14012), .A2(n10131), .A3(n10130), .ZN(n10132) );
  OAI211_X1 U12748 ( .C1(n10134), .C2(n14590), .A(n10133), .B(n10132), .ZN(
        P1_U3251) );
  INV_X1 U12749 ( .A(n13985), .ZN(n10303) );
  INV_X1 U12750 ( .A(n10135), .ZN(n10137) );
  OAI222_X1 U12751 ( .A1(n10303), .A2(P1_U3086), .B1(n12362), .B2(n10137), 
        .C1(n10136), .C2(n14366), .ZN(P1_U3344) );
  INV_X1 U12752 ( .A(n11487), .ZN(n10426) );
  OAI222_X1 U12753 ( .A1(n12073), .A2(n10138), .B1(n12071), .B2(n10137), .C1(
        P2_U3088), .C2(n10426), .ZN(P2_U3316) );
  INV_X1 U12754 ( .A(n12801), .ZN(n12790) );
  OAI222_X1 U12755 ( .A1(n15458), .A2(n10140), .B1(n15456), .B2(n10139), .C1(
        n12790), .C2(P3_U3151), .ZN(P3_U3282) );
  AOI21_X1 U12756 ( .B1(n10143), .B2(n10142), .A(n10141), .ZN(n10144) );
  AND2_X1 U12757 ( .A1(n9012), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10146) );
  NOR2_X1 U12758 ( .A1(n9012), .A2(P2_U3088), .ZN(n13697) );
  AND2_X1 U12759 ( .A1(n10169), .A2(n13697), .ZN(n10178) );
  INV_X1 U12760 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10148) );
  MUX2_X1 U12761 ( .A(n10148), .B(P2_REG1_REG_1__SCAN_IN), .S(n10331), .Z(
        n10149) );
  AND2_X1 U12762 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10322) );
  NAND2_X1 U12763 ( .A1(n10149), .A2(n10322), .ZN(n10323) );
  NAND2_X1 U12764 ( .A1(n10170), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10224) );
  NAND2_X1 U12765 ( .A1(n10323), .A2(n10224), .ZN(n10152) );
  INV_X1 U12766 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10150) );
  MUX2_X1 U12767 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10150), .S(n10222), .Z(
        n10151) );
  NAND2_X1 U12768 ( .A1(n10152), .A2(n10151), .ZN(n13338) );
  NAND2_X1 U12769 ( .A1(n10222), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13337) );
  NAND2_X1 U12770 ( .A1(n13338), .A2(n13337), .ZN(n10155) );
  INV_X1 U12771 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10153) );
  MUX2_X1 U12772 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10153), .S(n13335), .Z(
        n10154) );
  NAND2_X1 U12773 ( .A1(n10155), .A2(n10154), .ZN(n13340) );
  NAND2_X1 U12774 ( .A1(n13335), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U12775 ( .A1(n13340), .A2(n10156), .ZN(n10259) );
  INV_X1 U12776 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10157) );
  MUX2_X1 U12777 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10157), .S(n10174), .Z(
        n10258) );
  NAND2_X1 U12778 ( .A1(n10259), .A2(n10258), .ZN(n10257) );
  NAND2_X1 U12779 ( .A1(n10174), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U12780 ( .A1(n10257), .A2(n10189), .ZN(n10160) );
  INV_X1 U12781 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10158) );
  MUX2_X1 U12782 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10158), .S(n10187), .Z(
        n10159) );
  NAND2_X1 U12783 ( .A1(n10160), .A2(n10159), .ZN(n10191) );
  NAND2_X1 U12784 ( .A1(n10187), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U12785 ( .A1(n10191), .A2(n10161), .ZN(n14731) );
  INV_X1 U12786 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10162) );
  MUX2_X1 U12787 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10162), .S(n10176), .Z(
        n14730) );
  NAND2_X1 U12788 ( .A1(n14731), .A2(n14730), .ZN(n14729) );
  NAND2_X1 U12789 ( .A1(n10176), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10167) );
  NAND2_X1 U12790 ( .A1(n14729), .A2(n10167), .ZN(n10165) );
  INV_X1 U12791 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10163) );
  MUX2_X1 U12792 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10163), .S(n10274), .Z(
        n10164) );
  NAND2_X1 U12793 ( .A1(n10165), .A2(n10164), .ZN(n10266) );
  MUX2_X1 U12794 ( .A(n10163), .B(P2_REG1_REG_7__SCAN_IN), .S(n10274), .Z(
        n10166) );
  NAND3_X1 U12795 ( .A1(n14729), .A2(n10167), .A3(n10166), .ZN(n10168) );
  NAND3_X1 U12796 ( .A1(n14782), .A2(n10266), .A3(n10168), .ZN(n10185) );
  NOR2_X2 U12797 ( .A1(n10169), .A2(P2_U3088), .ZN(n14788) );
  NAND2_X1 U12798 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n10906) );
  XNOR2_X1 U12799 ( .A(n10331), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n10321) );
  AND2_X1 U12800 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10320) );
  AOI22_X1 U12801 ( .A1(n10321), .A2(n10320), .B1(n10170), .B2(
        P2_REG2_REG_1__SCAN_IN), .ZN(n10221) );
  INV_X1 U12802 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10171) );
  MUX2_X1 U12803 ( .A(n10171), .B(P2_REG2_REG_2__SCAN_IN), .S(n10222), .Z(
        n10220) );
  NOR2_X1 U12804 ( .A1(n10221), .A2(n10220), .ZN(n13334) );
  NOR2_X1 U12805 ( .A1(n10230), .A2(n10171), .ZN(n13329) );
  INV_X1 U12806 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10790) );
  MUX2_X1 U12807 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10790), .S(n13335), .Z(
        n10172) );
  NAND2_X1 U12808 ( .A1(n13335), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10254) );
  INV_X1 U12809 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10173) );
  MUX2_X1 U12810 ( .A(n10173), .B(P2_REG2_REG_4__SCAN_IN), .S(n10174), .Z(
        n10253) );
  AOI21_X1 U12811 ( .B1(n13332), .B2(n10254), .A(n10253), .ZN(n10252) );
  INV_X1 U12812 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n15349) );
  MUX2_X1 U12813 ( .A(n15349), .B(P2_REG2_REG_5__SCAN_IN), .S(n10187), .Z(
        n10193) );
  NOR2_X1 U12814 ( .A1(n10194), .A2(n10193), .ZN(n10192) );
  AOI21_X1 U12815 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n10187), .A(n10192), .ZN(
        n14727) );
  INV_X1 U12816 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10175) );
  MUX2_X1 U12817 ( .A(n10175), .B(P2_REG2_REG_6__SCAN_IN), .S(n10176), .Z(
        n14726) );
  NOR2_X1 U12818 ( .A1(n14727), .A2(n14726), .ZN(n14725) );
  INV_X1 U12819 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10177) );
  MUX2_X1 U12820 ( .A(n10177), .B(P2_REG2_REG_7__SCAN_IN), .S(n10274), .Z(
        n10179) );
  NOR2_X1 U12821 ( .A1(n10180), .A2(n10179), .ZN(n10273) );
  NAND2_X1 U12822 ( .A1(n10178), .A2(n12015), .ZN(n14744) );
  AOI211_X1 U12823 ( .C1(n10180), .C2(n10179), .A(n10273), .B(n14744), .ZN(
        n10181) );
  INV_X1 U12824 ( .A(n10181), .ZN(n10182) );
  NAND2_X1 U12825 ( .A1(n10906), .A2(n10182), .ZN(n10183) );
  AOI21_X1 U12826 ( .B1(n14788), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n10183), .ZN(
        n10184) );
  OAI211_X1 U12827 ( .C1(n14795), .C2(n10186), .A(n10185), .B(n10184), .ZN(
        P2_U3221) );
  MUX2_X1 U12828 ( .A(n10158), .B(P2_REG1_REG_5__SCAN_IN), .S(n10187), .Z(
        n10188) );
  NAND3_X1 U12829 ( .A1(n10257), .A2(n10189), .A3(n10188), .ZN(n10190) );
  NAND3_X1 U12830 ( .A1(n14782), .A2(n10191), .A3(n10190), .ZN(n10199) );
  NAND2_X1 U12831 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10500) );
  AOI211_X1 U12832 ( .C1(n10194), .C2(n10193), .A(n10192), .B(n14744), .ZN(
        n10195) );
  INV_X1 U12833 ( .A(n10195), .ZN(n10196) );
  NAND2_X1 U12834 ( .A1(n10500), .A2(n10196), .ZN(n10197) );
  AOI21_X1 U12835 ( .B1(n14788), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10197), .ZN(
        n10198) );
  OAI211_X1 U12836 ( .C1(n14795), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        P2_U3219) );
  INV_X1 U12837 ( .A(n10449), .ZN(n10456) );
  INV_X1 U12838 ( .A(n10201), .ZN(n10203) );
  OAI222_X1 U12839 ( .A1(P1_U3086), .A2(n10456), .B1(n12362), .B2(n10203), 
        .C1(n10202), .C2(n14366), .ZN(P1_U3343) );
  INV_X1 U12840 ( .A(n11486), .ZN(n14763) );
  OAI222_X1 U12841 ( .A1(n12073), .A2(n10204), .B1(n12071), .B2(n10203), .C1(
        n14763), .C2(P2_U3088), .ZN(P2_U3315) );
  CLKBUF_X1 U12842 ( .A(P1_U4016), .Z(n13861) );
  NOR2_X1 U12843 ( .A1(n14568), .A2(n13861), .ZN(P1_U3085) );
  NOR2_X1 U12844 ( .A1(n10205), .A2(n10127), .ZN(n13969) );
  INV_X1 U12845 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11273) );
  MUX2_X1 U12846 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11273), .S(n13968), .Z(
        n10206) );
  OAI21_X1 U12847 ( .B1(n13974), .B2(n13969), .A(n10206), .ZN(n13972) );
  NAND2_X1 U12848 ( .A1(n13968), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10209) );
  INV_X1 U12849 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10207) );
  MUX2_X1 U12850 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10207), .S(n10297), .Z(
        n10208) );
  AOI21_X1 U12851 ( .B1(n13972), .B2(n10209), .A(n10208), .ZN(n13988) );
  NAND3_X1 U12852 ( .A1(n13972), .A2(n10209), .A3(n10208), .ZN(n10210) );
  NAND2_X1 U12853 ( .A1(n10210), .A2(n14012), .ZN(n10219) );
  NOR2_X1 U12854 ( .A1(n10211), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n13961) );
  INV_X1 U12855 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11504) );
  MUX2_X1 U12856 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n11504), .S(n13968), .Z(
        n13962) );
  OAI21_X1 U12857 ( .B1(n13963), .B2(n13961), .A(n13962), .ZN(n13960) );
  OAI21_X1 U12858 ( .B1(n13968), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13960), .ZN(
        n10213) );
  INV_X1 U12859 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11410) );
  MUX2_X1 U12860 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11410), .S(n10297), .Z(
        n10212) );
  NOR2_X1 U12861 ( .A1(n10213), .A2(n10212), .ZN(n10301) );
  AOI211_X1 U12862 ( .C1(n10213), .C2(n10212), .A(n14590), .B(n10301), .ZN(
        n10214) );
  INV_X1 U12863 ( .A(n10214), .ZN(n10218) );
  AND2_X1 U12864 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11681) );
  NOR2_X1 U12865 ( .A1(n14596), .A2(n10215), .ZN(n10216) );
  AOI211_X1 U12866 ( .C1(n13984), .C2(n10302), .A(n11681), .B(n10216), .ZN(
        n10217) );
  OAI211_X1 U12867 ( .C1(n13988), .C2(n10219), .A(n10218), .B(n10217), .ZN(
        P1_U3253) );
  AOI211_X1 U12868 ( .C1(n10221), .C2(n10220), .A(n13334), .B(n14744), .ZN(
        n10227) );
  MUX2_X1 U12869 ( .A(n10150), .B(P2_REG1_REG_2__SCAN_IN), .S(n10222), .Z(
        n10223) );
  NAND3_X1 U12870 ( .A1(n10323), .A2(n10224), .A3(n10223), .ZN(n10225) );
  AND3_X1 U12871 ( .A1(n14782), .A2(n13338), .A3(n10225), .ZN(n10226) );
  NOR2_X1 U12872 ( .A1(n10227), .A2(n10226), .ZN(n10229) );
  AOI22_X1 U12873 ( .A1(n14788), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n10228) );
  OAI211_X1 U12874 ( .C1(n10230), .C2(n14795), .A(n10229), .B(n10228), .ZN(
        P2_U3216) );
  INV_X1 U12875 ( .A(n10231), .ZN(n10233) );
  OAI222_X1 U12876 ( .A1(n12787), .A2(P3_U3151), .B1(n15458), .B2(n10233), 
        .C1(n10232), .C2(n15456), .ZN(P3_U3281) );
  INV_X1 U12877 ( .A(n10360), .ZN(n10234) );
  INV_X1 U12878 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U12879 ( .A1(n10342), .A2(n7578), .ZN(n12092) );
  NAND2_X1 U12880 ( .A1(n12093), .A2(n12092), .ZN(n12298) );
  NAND2_X1 U12881 ( .A1(n14404), .A2(n14234), .ZN(n10236) );
  AND2_X1 U12882 ( .A1(n12298), .A2(n10236), .ZN(n14639) );
  INV_X1 U12883 ( .A(n14639), .ZN(n10239) );
  NAND2_X1 U12884 ( .A1(n13860), .A2(n14207), .ZN(n14635) );
  NAND3_X1 U12885 ( .A1(n10237), .A2(n14632), .A3(n12089), .ZN(n10238) );
  NAND3_X1 U12886 ( .A1(n10239), .A2(n14635), .A3(n10238), .ZN(n10248) );
  NAND2_X1 U12887 ( .A1(n14710), .A2(n10248), .ZN(n10240) );
  OAI21_X1 U12888 ( .B1(n14710), .B2(n10241), .A(n10240), .ZN(P1_U3459) );
  INV_X1 U12889 ( .A(n10242), .ZN(n10244) );
  OAI222_X1 U12890 ( .A1(P1_U3086), .A2(n10521), .B1(n12362), .B2(n10244), 
        .C1(n10243), .C2(n14366), .ZN(P1_U3342) );
  INV_X1 U12891 ( .A(n11478), .ZN(n14780) );
  OAI222_X1 U12892 ( .A1(n12073), .A2(n10245), .B1(n12071), .B2(n10244), .C1(
        n14780), .C2(P2_U3088), .ZN(P2_U3314) );
  NAND2_X1 U12893 ( .A1(n14720), .A2(n10248), .ZN(n10249) );
  OAI21_X1 U12894 ( .B1(n14720), .B2(n9296), .A(n10249), .ZN(P1_U3528) );
  OAI222_X1 U12895 ( .A1(n15458), .A2(n10251), .B1(n15456), .B2(n10250), .C1(
        n6753), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12896 ( .A(n10252), .ZN(n10256) );
  NAND3_X1 U12897 ( .A1(n13332), .A2(n10254), .A3(n10253), .ZN(n10255) );
  NAND3_X1 U12898 ( .A1(n14790), .A2(n10256), .A3(n10255), .ZN(n10263) );
  NAND2_X1 U12899 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10510) );
  OAI211_X1 U12900 ( .C1(n10259), .C2(n10258), .A(n14782), .B(n10257), .ZN(
        n10260) );
  NAND2_X1 U12901 ( .A1(n10510), .A2(n10260), .ZN(n10261) );
  AOI21_X1 U12902 ( .B1(n14788), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n10261), .ZN(
        n10262) );
  OAI211_X1 U12903 ( .C1(n14795), .C2(n10264), .A(n10263), .B(n10262), .ZN(
        P2_U3218) );
  NAND2_X1 U12904 ( .A1(n10274), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12905 ( .A1(n10266), .A2(n10265), .ZN(n14742) );
  INV_X1 U12906 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10267) );
  MUX2_X1 U12907 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10267), .S(n10276), .Z(
        n14741) );
  NAND2_X1 U12908 ( .A1(n14742), .A2(n14741), .ZN(n14740) );
  NAND2_X1 U12909 ( .A1(n10276), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U12910 ( .A1(n14740), .A2(n10268), .ZN(n10272) );
  INV_X1 U12911 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10269) );
  MUX2_X1 U12912 ( .A(n10269), .B(P2_REG1_REG_9__SCAN_IN), .S(n10396), .Z(
        n10271) );
  OR2_X1 U12913 ( .A1(n10272), .A2(n10271), .ZN(n10398) );
  INV_X1 U12914 ( .A(n10398), .ZN(n10270) );
  AOI21_X1 U12915 ( .B1(n10272), .B2(n10271), .A(n10270), .ZN(n10285) );
  INV_X1 U12916 ( .A(n14782), .ZN(n13370) );
  AOI21_X1 U12917 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n10274), .A(n10273), .ZN(
        n14746) );
  INV_X1 U12918 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10275) );
  MUX2_X1 U12919 ( .A(n10275), .B(P2_REG2_REG_8__SCAN_IN), .S(n10276), .Z(
        n14745) );
  NOR2_X1 U12920 ( .A1(n14746), .A2(n14745), .ZN(n14743) );
  INV_X1 U12921 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10277) );
  MUX2_X1 U12922 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10277), .S(n10396), .Z(
        n10278) );
  NAND2_X1 U12923 ( .A1(n10279), .A2(n10278), .ZN(n10392) );
  OAI21_X1 U12924 ( .B1(n10279), .B2(n10278), .A(n10392), .ZN(n10280) );
  NAND2_X1 U12925 ( .A1(n10280), .A2(n14790), .ZN(n10284) );
  NAND2_X1 U12926 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10947) );
  OAI21_X1 U12927 ( .B1(n14795), .B2(n10281), .A(n10947), .ZN(n10282) );
  AOI21_X1 U12928 ( .B1(n14788), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n10282), .ZN(
        n10283) );
  OAI211_X1 U12929 ( .C1(n10285), .C2(n13370), .A(n10284), .B(n10283), .ZN(
        P2_U3223) );
  NOR2_X1 U12930 ( .A1(n15060), .A2(n12627), .ZN(n12595) );
  INV_X1 U12931 ( .A(n10286), .ZN(n10287) );
  NAND2_X1 U12932 ( .A1(n10287), .A2(n15124), .ZN(n10288) );
  OAI22_X1 U12933 ( .A1(n12595), .A2(n10288), .B1(n7838), .B2(n15050), .ZN(
        n10493) );
  INV_X1 U12934 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10289) );
  NOR2_X1 U12935 ( .A1(n15144), .A2(n10289), .ZN(n10290) );
  AOI21_X1 U12936 ( .B1(n15144), .B2(n10493), .A(n10290), .ZN(n10291) );
  OAI21_X1 U12937 ( .B1(n10317), .B2(n13136), .A(n10291), .ZN(P3_U3459) );
  NAND2_X1 U12938 ( .A1(n14433), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12357) );
  NAND2_X1 U12939 ( .A1(n12357), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U12940 ( .A1(n14416), .A2(n12782), .B1(n14441), .B2(n10492), .ZN(
        n10292) );
  OAI211_X1 U12941 ( .C1(n12595), .C2(n14427), .A(n10293), .B(n10292), .ZN(
        P3_U3172) );
  OAI222_X1 U12942 ( .A1(n15458), .A2(n10295), .B1(n15456), .B2(n10294), .C1(
        n12845), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12943 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U12944 ( .A1(P3_U3897), .A2(n13049), .ZN(n10296) );
  OAI21_X1 U12945 ( .B1(P3_U3897), .B2(n15385), .A(n10296), .ZN(P3_U3510) );
  NOR2_X1 U12946 ( .A1(n10297), .A2(n10207), .ZN(n13987) );
  MUX2_X1 U12947 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11379), .S(n13985), .Z(
        n13986) );
  OAI21_X1 U12948 ( .B1(n13988), .B2(n13987), .A(n13986), .ZN(n13990) );
  OAI21_X1 U12949 ( .B1(n11379), .B2(n10303), .A(n13990), .ZN(n10300) );
  INV_X1 U12950 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U12951 ( .A1(n10449), .A2(n10298), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10456), .ZN(n10299) );
  NOR2_X1 U12952 ( .A1(n10299), .A2(n10300), .ZN(n10450) );
  AOI21_X1 U12953 ( .B1(n10300), .B2(n10299), .A(n10450), .ZN(n10313) );
  AOI21_X1 U12954 ( .B1(n10302), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10301), 
        .ZN(n13979) );
  MUX2_X1 U12955 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9423), .S(n13985), .Z(
        n13980) );
  NAND2_X1 U12956 ( .A1(n13979), .A2(n13980), .ZN(n13978) );
  NAND2_X1 U12957 ( .A1(n10303), .A2(n9423), .ZN(n10305) );
  INV_X1 U12958 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10304) );
  MUX2_X1 U12959 ( .A(n10304), .B(P1_REG1_REG_12__SCAN_IN), .S(n10449), .Z(
        n10306) );
  AOI21_X1 U12960 ( .B1(n13978), .B2(n10305), .A(n10306), .ZN(n10455) );
  AND3_X1 U12961 ( .A1(n13978), .A2(n10306), .A3(n10305), .ZN(n10307) );
  INV_X1 U12962 ( .A(n14590), .ZN(n14011) );
  OAI21_X1 U12963 ( .B1(n10455), .B2(n10307), .A(n14011), .ZN(n10312) );
  INV_X1 U12964 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10308) );
  NOR2_X1 U12965 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10308), .ZN(n10310) );
  NOR2_X1 U12966 ( .A1(n14592), .A2(n10456), .ZN(n10309) );
  AOI211_X1 U12967 ( .C1(n14568), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10310), 
        .B(n10309), .ZN(n10311) );
  OAI211_X1 U12968 ( .C1(n10313), .C2(n14588), .A(n10312), .B(n10311), .ZN(
        P1_U3255) );
  INV_X1 U12969 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n15356) );
  NAND2_X1 U12970 ( .A1(P3_U3897), .A2(n15063), .ZN(n10314) );
  OAI21_X1 U12971 ( .B1(P3_U3897), .B2(n15356), .A(n10314), .ZN(P3_U3493) );
  NOR2_X1 U12972 ( .A1(n15130), .A2(n7819), .ZN(n10315) );
  AOI21_X1 U12973 ( .B1(n15130), .B2(n10493), .A(n10315), .ZN(n10316) );
  OAI21_X1 U12974 ( .B1(n10317), .B2(n13196), .A(n10316), .ZN(P3_U3390) );
  INV_X1 U12975 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n15324) );
  NAND2_X1 U12976 ( .A1(n12551), .A2(P3_U3897), .ZN(n10318) );
  OAI21_X1 U12977 ( .B1(P3_U3897), .B2(n15324), .A(n10318), .ZN(P3_U3513) );
  INV_X1 U12978 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n15256) );
  NAND2_X1 U12979 ( .A1(n13036), .A2(P3_U3897), .ZN(n10319) );
  OAI21_X1 U12980 ( .B1(P3_U3897), .B2(n15256), .A(n10319), .ZN(P3_U3511) );
  XOR2_X1 U12981 ( .A(n10321), .B(n10320), .Z(n10328) );
  MUX2_X1 U12982 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10148), .S(n10331), .Z(
        n10326) );
  INV_X1 U12983 ( .A(n10322), .ZN(n10325) );
  INV_X1 U12984 ( .A(n10323), .ZN(n10324) );
  AOI211_X1 U12985 ( .C1(n10326), .C2(n10325), .A(n10324), .B(n13370), .ZN(
        n10327) );
  AOI21_X1 U12986 ( .B1(n14790), .B2(n10328), .A(n10327), .ZN(n10330) );
  AOI22_X1 U12987 ( .A1(n14788), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n10329) );
  OAI211_X1 U12988 ( .C1(n10331), .C2(n14795), .A(n10330), .B(n10329), .ZN(
        P2_U3215) );
  INV_X1 U12989 ( .A(n10332), .ZN(n10334) );
  INV_X1 U12990 ( .A(n11611), .ZN(n11868) );
  OAI222_X1 U12991 ( .A1(n12073), .A2(n10333), .B1(n12071), .B2(n10334), .C1(
        n11868), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U12992 ( .A(n11523), .ZN(n11332) );
  OAI222_X1 U12993 ( .A1(P1_U3086), .A2(n11332), .B1(n12362), .B2(n10334), 
        .C1(n15293), .C2(n14366), .ZN(P1_U3339) );
  XOR2_X1 U12994 ( .A(n10336), .B(n10335), .Z(n10341) );
  AOI22_X1 U12995 ( .A1(n14416), .A2(n12781), .B1(n14441), .B2(n10337), .ZN(
        n10338) );
  OAI21_X1 U12996 ( .B1(n7838), .B2(n14418), .A(n10338), .ZN(n10339) );
  AOI21_X1 U12997 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n12357), .A(n10339), .ZN(
        n10340) );
  OAI21_X1 U12998 ( .B1(n10341), .B2(n14427), .A(n10340), .ZN(P3_U3177) );
  INV_X1 U12999 ( .A(n10343), .ZN(n10345) );
  INV_X1 U13000 ( .A(n14242), .ZN(n10344) );
  INV_X1 U13001 ( .A(n14566), .ZN(n13867) );
  NAND3_X1 U13002 ( .A1(n10354), .A2(n10353), .A3(n10352), .ZN(n10361) );
  NAND2_X1 U13003 ( .A1(n12089), .A2(n10355), .ZN(n10356) );
  NAND3_X1 U13004 ( .A1(n10357), .A2(n12287), .A3(n14702), .ZN(n10358) );
  INV_X1 U13005 ( .A(n12346), .ZN(n10359) );
  INV_X1 U13006 ( .A(n13811), .ZN(n13830) );
  NAND2_X1 U13007 ( .A1(n13859), .A2(n14207), .ZN(n10744) );
  INV_X1 U13008 ( .A(n10744), .ZN(n10362) );
  NAND2_X1 U13009 ( .A1(n10361), .A2(n10360), .ZN(n10587) );
  NAND2_X1 U13010 ( .A1(n10587), .A2(n12346), .ZN(n10445) );
  AOI22_X1 U13011 ( .A1(n13830), .A2(n10362), .B1(n10445), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10366) );
  INV_X1 U13012 ( .A(n14209), .ZN(n14218) );
  NOR2_X1 U13013 ( .A1(n13811), .A2(n14218), .ZN(n13799) );
  NOR2_X1 U13014 ( .A1(n14702), .A2(n10363), .ZN(n10364) );
  AOI22_X1 U13015 ( .A1(n13799), .A2(n10342), .B1(n13834), .B2(n12100), .ZN(
        n10365) );
  OAI211_X1 U13016 ( .C1(n10367), .C2(n13836), .A(n10366), .B(n10365), .ZN(
        P1_U3222) );
  INV_X1 U13017 ( .A(n11312), .ZN(n11322) );
  INV_X1 U13018 ( .A(n10368), .ZN(n10369) );
  OAI222_X1 U13019 ( .A1(P1_U3086), .A2(n11322), .B1(n12362), .B2(n10369), 
        .C1(n15357), .C2(n14366), .ZN(P1_U3341) );
  INV_X1 U13020 ( .A(n11482), .ZN(n14794) );
  OAI222_X1 U13021 ( .A1(n12073), .A2(n15428), .B1(n12071), .B2(n10369), .C1(
        n14794), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13022 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13023 ( .A1(n14790), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14782), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10372) );
  INV_X1 U13024 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10656) );
  OAI21_X1 U13025 ( .B1(n13370), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14795), .ZN(
        n10370) );
  AOI21_X1 U13026 ( .B1(n14790), .B2(n10656), .A(n10370), .ZN(n10371) );
  MUX2_X1 U13027 ( .A(n10372), .B(n10371), .S(P2_IR_REG_0__SCAN_IN), .Z(n10374) );
  NAND2_X1 U13028 ( .A1(n14788), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10373) );
  OAI211_X1 U13029 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10652), .A(n10374), .B(
        n10373), .ZN(P2_U3214) );
  INV_X1 U13030 ( .A(n13834), .ZN(n13817) );
  AOI21_X1 U13031 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(n13876) );
  OAI22_X1 U13032 ( .A1(n13876), .A2(n13836), .B1(n13811), .B2(n14635), .ZN(
        n10378) );
  AOI21_X1 U13033 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10445), .A(n10378), .ZN(
        n10379) );
  OAI21_X1 U13034 ( .B1(n7578), .B2(n13817), .A(n10379), .ZN(P1_U3232) );
  INV_X1 U13035 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U13036 ( .A1(n12731), .A2(P3_U3897), .ZN(n10380) );
  OAI21_X1 U13037 ( .B1(P3_U3897), .B2(n15285), .A(n10380), .ZN(P3_U3514) );
  INV_X1 U13038 ( .A(n14466), .ZN(n12857) );
  INV_X1 U13039 ( .A(n10381), .ZN(n10383) );
  OAI222_X1 U13040 ( .A1(n12857), .A2(P3_U3151), .B1(n15458), .B2(n10383), 
        .C1(n10382), .C2(n15456), .ZN(P3_U3278) );
  INV_X1 U13041 ( .A(n10384), .ZN(n10386) );
  OAI222_X1 U13042 ( .A1(n14366), .A2(n10385), .B1(n12362), .B2(n10386), .C1(
        n14578), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13043 ( .A(n11616), .ZN(n11497) );
  OAI222_X1 U13044 ( .A1(n12073), .A2(n10387), .B1(n12071), .B2(n10386), .C1(
        P2_U3088), .C2(n11497), .ZN(P2_U3312) );
  INV_X1 U13045 ( .A(n10388), .ZN(n10391) );
  INV_X1 U13046 ( .A(n13344), .ZN(n13353) );
  OAI222_X1 U13047 ( .A1(n12073), .A2(n10389), .B1(n12071), .B2(n10391), .C1(
        n13353), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13048 ( .A(n11517), .ZN(n14001) );
  OAI222_X1 U13049 ( .A1(P1_U3086), .A2(n14001), .B1(n14369), .B2(n10391), 
        .C1(n10390), .C2(n14366), .ZN(P1_U3338) );
  OAI21_X1 U13050 ( .B1(n10396), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10392), .ZN(
        n10395) );
  INV_X1 U13051 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10393) );
  MUX2_X1 U13052 ( .A(n10393), .B(P2_REG2_REG_10__SCAN_IN), .S(n10428), .Z(
        n10394) );
  NOR2_X1 U13053 ( .A1(n10395), .A2(n10394), .ZN(n10420) );
  AOI211_X1 U13054 ( .C1(n10395), .C2(n10394), .A(n14744), .B(n10420), .ZN(
        n10406) );
  OR2_X1 U13055 ( .A1(n10396), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U13056 ( .A1(n10398), .A2(n10397), .ZN(n10401) );
  INV_X1 U13057 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14889) );
  MUX2_X1 U13058 ( .A(n14889), .B(P2_REG1_REG_10__SCAN_IN), .S(n10428), .Z(
        n10400) );
  INV_X1 U13059 ( .A(n10434), .ZN(n10399) );
  AOI211_X1 U13060 ( .C1(n10401), .C2(n10400), .A(n13370), .B(n10399), .ZN(
        n10405) );
  AOI22_X1 U13061 ( .A1(n14788), .A2(P2_ADDR_REG_10__SCAN_IN), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(P2_U3088), .ZN(n10402) );
  OAI21_X1 U13062 ( .B1(n10403), .B2(n14795), .A(n10402), .ZN(n10404) );
  OR3_X1 U13063 ( .A1(n10406), .A2(n10405), .A3(n10404), .ZN(P2_U3224) );
  OAI222_X1 U13064 ( .A1(n15458), .A2(n10408), .B1(n15456), .B2(n10407), .C1(
        n6926), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13065 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15416) );
  XNOR2_X1 U13066 ( .A(n10409), .B(n10411), .ZN(n10415) );
  XNOR2_X1 U13067 ( .A(n10410), .B(n10411), .ZN(n10413) );
  AOI21_X1 U13068 ( .B1(n10413), .B2(n14707), .A(n10412), .ZN(n10414) );
  OAI21_X1 U13069 ( .B1(n14234), .B2(n10415), .A(n10414), .ZN(n10705) );
  INV_X1 U13070 ( .A(n10705), .ZN(n10416) );
  OAI211_X1 U13071 ( .C1(n10738), .C2(n10441), .A(n14622), .B(n10820), .ZN(
        n10704) );
  OAI211_X1 U13072 ( .C1(n10441), .C2(n14702), .A(n10416), .B(n10704), .ZN(
        n10418) );
  NAND2_X1 U13073 ( .A1(n10418), .A2(n14710), .ZN(n10417) );
  OAI21_X1 U13074 ( .B1(n14710), .B2(n15416), .A(n10417), .ZN(P1_U3465) );
  NAND2_X1 U13075 ( .A1(n10418), .A2(n14720), .ZN(n10419) );
  OAI21_X1 U13076 ( .B1(n14720), .B2(n9308), .A(n10419), .ZN(P1_U3530) );
  AOI21_X1 U13077 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n10428), .A(n10420), 
        .ZN(n10423) );
  INV_X1 U13078 ( .A(n10423), .ZN(n10425) );
  INV_X1 U13079 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10421) );
  MUX2_X1 U13080 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10421), .S(n11487), .Z(
        n10422) );
  INV_X1 U13081 ( .A(n10422), .ZN(n10424) );
  AOI21_X1 U13082 ( .B1(n10425), .B2(n10424), .A(n14753), .ZN(n10438) );
  NOR2_X1 U13083 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15250), .ZN(n11369) );
  NOR2_X1 U13084 ( .A1(n14795), .A2(n10426), .ZN(n10427) );
  AOI211_X1 U13085 ( .C1(n14788), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11369), 
        .B(n10427), .ZN(n10437) );
  NAND2_X1 U13086 ( .A1(n10428), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U13087 ( .A1(n10434), .A2(n10433), .ZN(n10431) );
  INV_X1 U13088 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10429) );
  MUX2_X1 U13089 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10429), .S(n11487), .Z(
        n10430) );
  NAND2_X1 U13090 ( .A1(n10431), .A2(n10430), .ZN(n14758) );
  MUX2_X1 U13091 ( .A(n10429), .B(P2_REG1_REG_11__SCAN_IN), .S(n11487), .Z(
        n10432) );
  NAND3_X1 U13092 ( .A1(n10434), .A2(n10433), .A3(n10432), .ZN(n10435) );
  NAND3_X1 U13093 ( .A1(n14758), .A2(n14782), .A3(n10435), .ZN(n10436) );
  OAI211_X1 U13094 ( .C1(n10438), .C2(n14744), .A(n10437), .B(n10436), .ZN(
        P2_U3225) );
  OAI22_X1 U13095 ( .A1(n12394), .A2(n9318), .B1(n10441), .B2(n10442), .ZN(
        n10591) );
  OAI22_X1 U13096 ( .A1(n9318), .A2(n12391), .B1(n10441), .B2(n12396), .ZN(
        n10443) );
  XNOR2_X1 U13097 ( .A(n10443), .B(n12450), .ZN(n10590) );
  AOI21_X1 U13098 ( .B1(n10444), .B2(n7548), .A(n10594), .ZN(n10448) );
  AOI22_X1 U13099 ( .A1(n13834), .A2(n10708), .B1(n10445), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10447) );
  NOR2_X1 U13100 ( .A1(n13811), .A2(n14221), .ZN(n13758) );
  AOI22_X1 U13101 ( .A1(n13758), .A2(n13858), .B1(n13799), .B2(n13860), .ZN(
        n10446) );
  OAI211_X1 U13102 ( .C1(n10448), .C2(n13836), .A(n10447), .B(n10446), .ZN(
        P1_U3237) );
  NOR2_X1 U13103 ( .A1(n10449), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10451) );
  NOR2_X1 U13104 ( .A1(n10451), .A2(n10450), .ZN(n10454) );
  MUX2_X1 U13105 ( .A(n10452), .B(P1_REG2_REG_13__SCAN_IN), .S(n10521), .Z(
        n10453) );
  NAND2_X1 U13106 ( .A1(n10453), .A2(n10454), .ZN(n10520) );
  OAI211_X1 U13107 ( .C1(n10454), .C2(n10453), .A(n10520), .B(n14012), .ZN(
        n10463) );
  NAND2_X1 U13108 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11958)
         );
  AOI21_X1 U13109 ( .B1(n10304), .B2(n10456), .A(n10455), .ZN(n10459) );
  MUX2_X1 U13110 ( .A(n10457), .B(P1_REG1_REG_13__SCAN_IN), .S(n10521), .Z(
        n10458) );
  NAND2_X1 U13111 ( .A1(n10459), .A2(n10458), .ZN(n10516) );
  OAI211_X1 U13112 ( .C1(n10459), .C2(n10458), .A(n14011), .B(n10516), .ZN(
        n10460) );
  NAND2_X1 U13113 ( .A1(n11958), .A2(n10460), .ZN(n10461) );
  AOI21_X1 U13114 ( .B1(n14568), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10461), 
        .ZN(n10462) );
  OAI211_X1 U13115 ( .C1(n14592), .C2(n10521), .A(n10463), .B(n10462), .ZN(
        P1_U3256) );
  XNOR2_X1 U13116 ( .A(n10465), .B(n10464), .ZN(n10473) );
  INV_X1 U13117 ( .A(n13283), .ZN(n13297) );
  INV_X1 U13118 ( .A(n10466), .ZN(n10714) );
  INV_X1 U13119 ( .A(n13252), .ZN(n10469) );
  NAND2_X1 U13120 ( .A1(n13320), .A2(n13540), .ZN(n10468) );
  NAND2_X1 U13121 ( .A1(n13318), .A2(n13538), .ZN(n10467) );
  NAND2_X1 U13122 ( .A1(n10468), .A2(n10467), .ZN(n10630) );
  NOR2_X1 U13123 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8485), .ZN(n14721) );
  AOI21_X1 U13124 ( .B1(n10469), .B2(n10630), .A(n14721), .ZN(n10470) );
  OAI21_X1 U13125 ( .B1(n13297), .B2(n10714), .A(n10470), .ZN(n10471) );
  AOI21_X1 U13126 ( .B1(n10835), .B2(n13302), .A(n10471), .ZN(n10472) );
  OAI21_X1 U13127 ( .B1(n10473), .B2(n13304), .A(n10472), .ZN(P2_U3211) );
  OAI21_X1 U13128 ( .B1(n10476), .B2(n10475), .A(n10474), .ZN(n10477) );
  NAND2_X1 U13129 ( .A1(n10477), .A2(n14439), .ZN(n10483) );
  NAND2_X1 U13130 ( .A1(n12781), .A2(n15061), .ZN(n10479) );
  NAND2_X1 U13131 ( .A1(n12779), .A2(n15064), .ZN(n10478) );
  AND2_X1 U13132 ( .A1(n10479), .A2(n10478), .ZN(n10861) );
  INV_X1 U13133 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10480) );
  OAI22_X1 U13134 ( .A1(n14446), .A2(n10861), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10480), .ZN(n10481) );
  AOI21_X1 U13135 ( .B1(n15096), .B2(n14441), .A(n10481), .ZN(n10482) );
  OAI211_X1 U13136 ( .C1(n10863), .C2(n14433), .A(n10483), .B(n10482), .ZN(
        P3_U3170) );
  XNOR2_X1 U13137 ( .A(n10485), .B(n10484), .ZN(n10486) );
  NAND3_X1 U13138 ( .A1(n10488), .A2(n10487), .A3(n10486), .ZN(n10491) );
  NAND2_X1 U13139 ( .A1(n15105), .A2(n15071), .ZN(n10490) );
  NOR2_X2 U13140 ( .A1(n10491), .A2(n10490), .ZN(n13026) );
  AOI22_X1 U13141 ( .A1(n13026), .A2(n10492), .B1(n13069), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10495) );
  NAND2_X1 U13142 ( .A1(n15077), .A2(n10493), .ZN(n10494) );
  OAI211_X1 U13143 ( .C1(n10552), .C2(n15077), .A(n10495), .B(n10494), .ZN(
        P3_U3233) );
  INV_X1 U13144 ( .A(n10919), .ZN(n14858) );
  OAI21_X1 U13145 ( .B1(n10498), .B2(n10497), .A(n10496), .ZN(n10499) );
  NAND2_X1 U13146 ( .A1(n10499), .A2(n13278), .ZN(n10503) );
  AOI22_X1 U13147 ( .A1(n13540), .A2(n13321), .B1(n13319), .B2(n13538), .ZN(
        n10923) );
  OAI21_X1 U13148 ( .B1(n13252), .B2(n10923), .A(n10500), .ZN(n10501) );
  AOI21_X1 U13149 ( .B1(n10918), .B2(n13283), .A(n10501), .ZN(n10502) );
  OAI211_X1 U13150 ( .C1(n14858), .C2(n11948), .A(n10503), .B(n10502), .ZN(
        P2_U3199) );
  INV_X1 U13151 ( .A(n14848), .ZN(n10762) );
  OAI21_X1 U13152 ( .B1(n10506), .B2(n10505), .A(n10504), .ZN(n10507) );
  NAND2_X1 U13153 ( .A1(n10507), .A2(n13278), .ZN(n10515) );
  NAND2_X1 U13154 ( .A1(n13322), .A2(n13540), .ZN(n10509) );
  NAND2_X1 U13155 ( .A1(n13320), .A2(n13538), .ZN(n10508) );
  NAND2_X1 U13156 ( .A1(n10509), .A2(n10508), .ZN(n10758) );
  INV_X1 U13157 ( .A(n10758), .ZN(n10511) );
  OAI21_X1 U13158 ( .B1(n13252), .B2(n10511), .A(n10510), .ZN(n10512) );
  AOI21_X1 U13159 ( .B1(n10513), .B2(n13283), .A(n10512), .ZN(n10514) );
  OAI211_X1 U13160 ( .C1(n10762), .C2(n11948), .A(n10515), .B(n10514), .ZN(
        P2_U3202) );
  AOI22_X1 U13161 ( .A1(n11312), .A2(n9467), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11322), .ZN(n10518) );
  OAI21_X1 U13162 ( .B1(n10521), .B2(n10457), .A(n10516), .ZN(n10517) );
  NOR2_X1 U13163 ( .A1(n10518), .A2(n10517), .ZN(n11321) );
  AOI21_X1 U13164 ( .B1(n10518), .B2(n10517), .A(n11321), .ZN(n10528) );
  MUX2_X1 U13165 ( .A(n9470), .B(P1_REG2_REG_14__SCAN_IN), .S(n11312), .Z(
        n10519) );
  INV_X1 U13166 ( .A(n10519), .ZN(n10523) );
  OAI21_X1 U13167 ( .B1(n10521), .B2(n10452), .A(n10520), .ZN(n10522) );
  NAND2_X1 U13168 ( .A1(n10523), .A2(n10522), .ZN(n11313) );
  OAI211_X1 U13169 ( .C1(n10523), .C2(n10522), .A(n14012), .B(n11313), .ZN(
        n10525) );
  AND2_X1 U13170 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13716) );
  AOI21_X1 U13171 ( .B1(n14568), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n13716), 
        .ZN(n10524) );
  OAI211_X1 U13172 ( .C1(n14592), .C2(n11322), .A(n10525), .B(n10524), .ZN(
        n10526) );
  INV_X1 U13173 ( .A(n10526), .ZN(n10527) );
  OAI21_X1 U13174 ( .B1(n10528), .B2(n14590), .A(n10527), .ZN(P1_U3257) );
  OAI222_X1 U13175 ( .A1(P3_U3151), .A2(n12883), .B1(n15456), .B2(n10530), 
        .C1(n15458), .C2(n10529), .ZN(P3_U3276) );
  INV_X1 U13176 ( .A(n10533), .ZN(n10531) );
  NAND2_X1 U13177 ( .A1(n10531), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12764) );
  NAND2_X1 U13178 ( .A1(n10532), .A2(n12764), .ZN(n10542) );
  INV_X1 U13179 ( .A(n10556), .ZN(n10535) );
  MUX2_X1 U13180 ( .A(n10535), .B(n10942), .S(n10534), .Z(n14985) );
  NAND2_X1 U13181 ( .A1(n10556), .A2(n6973), .ZN(n14908) );
  INV_X1 U13182 ( .A(n6940), .ZN(n10545) );
  NAND2_X1 U13183 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10536), .ZN(n10538) );
  INV_X1 U13184 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n15407) );
  NAND3_X1 U13185 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n15407), .A3(n10536), 
        .ZN(n10680) );
  INV_X1 U13186 ( .A(n10680), .ZN(n10537) );
  OAI21_X1 U13187 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10539), .A(n10681), .ZN(
        n10560) );
  INV_X1 U13188 ( .A(n10540), .ZN(n10541) );
  MUX2_X1 U13189 ( .A(n10552), .B(n10289), .S(n6973), .Z(n14892) );
  AND2_X1 U13190 ( .A1(n14892), .A2(n6922), .ZN(n14895) );
  INV_X1 U13191 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10543) );
  MUX2_X1 U13192 ( .A(n10544), .B(n10543), .S(n6973), .Z(n10546) );
  NAND2_X1 U13193 ( .A1(n10546), .A2(n10545), .ZN(n10676) );
  INV_X1 U13194 ( .A(n10546), .ZN(n10547) );
  NAND2_X1 U13195 ( .A1(n10547), .A2(n6940), .ZN(n10548) );
  AND2_X1 U13196 ( .A1(n10676), .A2(n10548), .ZN(n10549) );
  OAI21_X1 U13197 ( .B1(n14895), .B2(n10549), .A(n10678), .ZN(n10550) );
  AOI22_X1 U13198 ( .A1(n15031), .A2(n10550), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10551) );
  OAI21_X1 U13199 ( .B1(n15041), .B2(n15382), .A(n10551), .ZN(n10559) );
  NAND2_X1 U13200 ( .A1(n10553), .A2(n10544), .ZN(n10557) );
  INV_X1 U13201 ( .A(n10554), .ZN(n10555) );
  AOI21_X1 U13202 ( .B1(n10665), .B2(n10557), .A(n15036), .ZN(n10558) );
  AOI211_X1 U13203 ( .C1(n15023), .C2(n10560), .A(n10559), .B(n10558), .ZN(
        n10561) );
  OAI21_X1 U13204 ( .B1(n6940), .B2(n14985), .A(n10561), .ZN(P3_U3183) );
  XNOR2_X1 U13205 ( .A(n10563), .B(n10562), .ZN(n10570) );
  INV_X1 U13206 ( .A(n10697), .ZN(n10568) );
  INV_X1 U13207 ( .A(n14418), .ZN(n12479) );
  AOI22_X1 U13208 ( .A1(n12479), .A2(n12780), .B1(n14416), .B2(n12778), .ZN(
        n10567) );
  OAI22_X1 U13209 ( .A1(n12574), .A2(n15097), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10564), .ZN(n10565) );
  INV_X1 U13210 ( .A(n10565), .ZN(n10566) );
  OAI211_X1 U13211 ( .C1(n10568), .C2(n14433), .A(n10567), .B(n10566), .ZN(
        n10569) );
  AOI21_X1 U13212 ( .B1(n10570), .B2(n14439), .A(n10569), .ZN(n10571) );
  INV_X1 U13213 ( .A(n10571), .ZN(P3_U3167) );
  INV_X1 U13214 ( .A(n14005), .ZN(n14591) );
  OAI222_X1 U13215 ( .A1(n14366), .A2(n10572), .B1(n12362), .B2(n10574), .C1(
        P1_U3086), .C2(n14591), .ZN(P1_U3337) );
  INV_X1 U13216 ( .A(n13364), .ZN(n13350) );
  OAI222_X1 U13217 ( .A1(P2_U3088), .A2(n13350), .B1(n12071), .B2(n10574), 
        .C1(n10573), .C2(n12073), .ZN(P2_U3309) );
  OAI222_X1 U13218 ( .A1(P3_U3151), .A2(n10577), .B1(n15456), .B2(n10576), 
        .C1(n15458), .C2(n10575), .ZN(P3_U3275) );
  OAI21_X1 U13219 ( .B1(n10580), .B2(n10579), .A(n10578), .ZN(n10584) );
  NOR2_X1 U13220 ( .A1(n10581), .A2(n14815), .ZN(n10724) );
  INV_X1 U13221 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10775) );
  OAI22_X1 U13222 ( .A1(n11948), .A2(n10776), .B1(n10724), .B2(n10775), .ZN(
        n10583) );
  INV_X1 U13223 ( .A(n13325), .ZN(n10649) );
  INV_X1 U13224 ( .A(n13282), .ZN(n13295) );
  INV_X1 U13225 ( .A(n13284), .ZN(n13299) );
  OAI22_X1 U13226 ( .A1(n10649), .A2(n13295), .B1(n13299), .B2(n10610), .ZN(
        n10582) );
  AOI211_X1 U13227 ( .C1(n13278), .C2(n10584), .A(n10583), .B(n10582), .ZN(
        n10585) );
  INV_X1 U13228 ( .A(n10585), .ZN(P2_U3209) );
  NAND2_X1 U13229 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  NAND2_X1 U13230 ( .A1(n10588), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10589) );
  INV_X1 U13231 ( .A(n10590), .ZN(n10593) );
  INV_X1 U13232 ( .A(n10591), .ZN(n10592) );
  OAI22_X1 U13233 ( .A1(n10596), .A2(n10442), .B1(n7439), .B2(n12396), .ZN(
        n10595) );
  XOR2_X1 U13234 ( .A(n12450), .B(n10595), .Z(n10930) );
  OAI22_X1 U13235 ( .A1(n12394), .A2(n10596), .B1(n7439), .B2(n12391), .ZN(
        n10928) );
  XNOR2_X1 U13236 ( .A(n10930), .B(n10928), .ZN(n10597) );
  OAI211_X1 U13237 ( .C1(n10598), .C2(n10597), .A(n10932), .B(n13809), .ZN(
        n10601) );
  AND2_X1 U13238 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13901) );
  INV_X1 U13239 ( .A(n13799), .ZN(n13761) );
  INV_X1 U13240 ( .A(n13758), .ZN(n13801) );
  OAI22_X1 U13241 ( .A1(n9318), .A2(n13761), .B1(n13801), .B2(n12114), .ZN(
        n10599) );
  AOI211_X1 U13242 ( .C1(n13834), .C2(n10822), .A(n13901), .B(n10599), .ZN(
        n10600) );
  OAI211_X1 U13243 ( .C1(n13832), .C2(P1_REG3_REG_3__SCAN_IN), .A(n10601), .B(
        n10600), .ZN(P1_U3218) );
  INV_X1 U13244 ( .A(n10640), .ZN(n10602) );
  NOR2_X1 U13245 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  NAND4_X1 U13246 ( .A1(n10605), .A2(n14818), .A3(n10604), .A4(n14817), .ZN(
        n10637) );
  INV_X1 U13247 ( .A(n10642), .ZN(n10606) );
  INV_X1 U13248 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10636) );
  INV_X1 U13249 ( .A(n10607), .ZN(n10802) );
  NAND2_X1 U13250 ( .A1(n10769), .A2(n10771), .ZN(n10609) );
  NAND2_X1 U13251 ( .A1(n10801), .A2(n10776), .ZN(n10608) );
  NAND2_X1 U13252 ( .A1(n10609), .A2(n10608), .ZN(n10781) );
  NAND2_X1 U13253 ( .A1(n10781), .A2(n10783), .ZN(n10612) );
  NAND2_X1 U13254 ( .A1(n10610), .A2(n10795), .ZN(n10611) );
  NAND2_X1 U13255 ( .A1(n10753), .A2(n10752), .ZN(n10614) );
  OR2_X1 U13256 ( .A1(n13321), .A2(n14848), .ZN(n10613) );
  NOR2_X1 U13257 ( .A1(n10919), .A2(n13320), .ZN(n10615) );
  NAND2_X1 U13258 ( .A1(n10919), .A2(n13320), .ZN(n10616) );
  INV_X1 U13259 ( .A(n10829), .ZN(n10617) );
  AOI21_X1 U13260 ( .B1(n10832), .B2(n10618), .A(n10617), .ZN(n10721) );
  INV_X1 U13261 ( .A(n14877), .ZN(n14827) );
  AND2_X1 U13262 ( .A1(n10619), .A2(n10807), .ZN(n10800) );
  NAND2_X1 U13263 ( .A1(n10803), .A2(n10800), .ZN(n10799) );
  NAND2_X1 U13264 ( .A1(n10649), .A2(n6560), .ZN(n10770) );
  NAND2_X1 U13265 ( .A1(n10799), .A2(n10770), .ZN(n10620) );
  NAND2_X1 U13266 ( .A1(n10784), .A2(n10782), .ZN(n10621) );
  INV_X1 U13267 ( .A(n10783), .ZN(n10780) );
  NAND2_X1 U13268 ( .A1(n10621), .A2(n10780), .ZN(n10786) );
  NAND2_X1 U13269 ( .A1(n10786), .A2(n10622), .ZN(n10755) );
  INV_X1 U13270 ( .A(n10752), .ZN(n10754) );
  NAND2_X1 U13271 ( .A1(n10755), .A2(n10754), .ZN(n10757) );
  NAND2_X1 U13272 ( .A1(n14848), .A2(n10659), .ZN(n10623) );
  NAND2_X1 U13273 ( .A1(n10757), .A2(n10623), .ZN(n10922) );
  INV_X1 U13274 ( .A(n13320), .ZN(n10625) );
  OR2_X1 U13275 ( .A1(n10919), .A2(n10625), .ZN(n10624) );
  NAND2_X1 U13276 ( .A1(n10922), .A2(n10624), .ZN(n10627) );
  NAND2_X1 U13277 ( .A1(n10919), .A2(n10625), .ZN(n10626) );
  NAND2_X1 U13278 ( .A1(n10627), .A2(n10626), .ZN(n10833) );
  XNOR2_X1 U13279 ( .A(n10833), .B(n10832), .ZN(n10631) );
  AOI21_X1 U13280 ( .B1(n10631), .B2(n13569), .A(n10630), .ZN(n10718) );
  INV_X1 U13281 ( .A(n10632), .ZN(n10916) );
  INV_X1 U13282 ( .A(n10835), .ZN(n10715) );
  INV_X1 U13283 ( .A(n10843), .ZN(n10633) );
  AOI211_X1 U13284 ( .C1(n10835), .C2(n10916), .A(n6569), .B(n10633), .ZN(
        n10717) );
  AOI21_X1 U13285 ( .B1(n14847), .B2(n10835), .A(n10717), .ZN(n10634) );
  OAI211_X1 U13286 ( .C1(n10721), .C2(n14840), .A(n10718), .B(n10634), .ZN(
        n10638) );
  NAND2_X1 U13287 ( .A1(n10638), .A2(n14880), .ZN(n10635) );
  OAI21_X1 U13288 ( .B1(n14880), .B2(n10636), .A(n10635), .ZN(P2_U3448) );
  NAND2_X1 U13289 ( .A1(n10638), .A2(n14891), .ZN(n10639) );
  OAI21_X1 U13290 ( .B1(n14891), .B2(n10162), .A(n10639), .ZN(P2_U3505) );
  NAND4_X1 U13291 ( .A1(n14818), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10643) );
  INV_X1 U13292 ( .A(n10644), .ZN(n10645) );
  NAND2_X1 U13293 ( .A1(n13562), .A2(n10645), .ZN(n13410) );
  INV_X1 U13294 ( .A(n13410), .ZN(n11341) );
  INV_X1 U13295 ( .A(n10722), .ZN(n14821) );
  NOR2_X4 U13296 ( .A1(n14809), .A2(n10646), .ZN(n14797) );
  INV_X1 U13297 ( .A(n10647), .ZN(n10648) );
  NOR2_X1 U13298 ( .A1(n10648), .A2(n10723), .ZN(n14820) );
  AOI22_X1 U13299 ( .A1(n11341), .A2(n14821), .B1(n14797), .B2(n14820), .ZN(
        n10655) );
  INV_X1 U13300 ( .A(n11185), .ZN(n14862) );
  NOR2_X1 U13301 ( .A1(n14862), .A2(n13569), .ZN(n10650) );
  OAI22_X1 U13302 ( .A1(n10722), .A2(n10650), .B1(n10649), .B2(n13524), .ZN(
        n14819) );
  INV_X1 U13303 ( .A(n14820), .ZN(n10651) );
  OAI22_X1 U13304 ( .A1(n13571), .A2(n10652), .B1(n11176), .B2(n10651), .ZN(
        n10653) );
  OAI21_X1 U13305 ( .B1(n14819), .B2(n10653), .A(n13562), .ZN(n10654) );
  OAI211_X1 U13306 ( .C1(n13562), .C2(n10656), .A(n10655), .B(n10654), .ZN(
        P2_U3265) );
  XNOR2_X1 U13307 ( .A(n10658), .B(n10657), .ZN(n10663) );
  NAND2_X1 U13308 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13326) );
  OAI21_X1 U13309 ( .B1(n13295), .B2(n10801), .A(n13326), .ZN(n10661) );
  OAI22_X1 U13310 ( .A1(n13299), .A2(n10659), .B1(n10795), .B2(n11948), .ZN(
        n10660) );
  AOI211_X1 U13311 ( .C1(n13283), .C2(n8423), .A(n10661), .B(n10660), .ZN(
        n10662) );
  OAI21_X1 U13312 ( .B1(n10663), .B2(n13304), .A(n10662), .ZN(P2_U3190) );
  OAI21_X1 U13313 ( .B1(n10667), .B2(n10666), .A(n11006), .ZN(n10688) );
  NAND2_X1 U13314 ( .A1(n10678), .A2(n10676), .ZN(n10674) );
  INV_X1 U13315 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10668) );
  MUX2_X1 U13316 ( .A(n10669), .B(n10668), .S(n6973), .Z(n10671) );
  NAND2_X1 U13318 ( .A1(n10671), .A2(n6562), .ZN(n14902) );
  INV_X1 U13319 ( .A(n10671), .ZN(n10672) );
  NAND2_X1 U13320 ( .A1(n10672), .A2(n6564), .ZN(n10673) );
  AND2_X1 U13321 ( .A1(n14902), .A2(n10673), .ZN(n10675) );
  NAND2_X1 U13322 ( .A1(n10674), .A2(n10675), .ZN(n14903) );
  INV_X1 U13323 ( .A(n10675), .ZN(n10677) );
  NAND3_X1 U13324 ( .A1(n10678), .A2(n10677), .A3(n10676), .ZN(n10679) );
  AOI21_X1 U13325 ( .B1(n14903), .B2(n10679), .A(n15010), .ZN(n10687) );
  MUX2_X1 U13326 ( .A(n10668), .B(P3_REG1_REG_2__SCAN_IN), .S(n6564), .Z(
        n10683) );
  AOI21_X1 U13327 ( .B1(n10683), .B2(n10682), .A(n11021), .ZN(n10685) );
  AOI22_X1 U13328 ( .A1(n14990), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10684) );
  OAI21_X1 U13329 ( .B1(n10685), .B2(n14908), .A(n10684), .ZN(n10686) );
  AOI211_X1 U13330 ( .C1(n14474), .C2(n10688), .A(n10687), .B(n10686), .ZN(
        n10689) );
  OAI21_X1 U13331 ( .B1(n6564), .B2(n14985), .A(n10689), .ZN(P3_U3184) );
  INV_X1 U13332 ( .A(n10690), .ZN(n10691) );
  AOI21_X1 U13333 ( .B1(n12652), .B2(n10692), .A(n10691), .ZN(n10696) );
  AOI22_X1 U13334 ( .A1(n15061), .A2(n12780), .B1(n12778), .B2(n15064), .ZN(
        n10695) );
  XNOR2_X1 U13335 ( .A(n10693), .B(n12652), .ZN(n15100) );
  NAND2_X1 U13336 ( .A1(n15100), .A2(n15118), .ZN(n10694) );
  OAI211_X1 U13337 ( .C1(n10696), .C2(n13063), .A(n10695), .B(n10694), .ZN(
        n15098) );
  INV_X1 U13338 ( .A(n15098), .ZN(n10702) );
  NOR2_X1 U13339 ( .A1(n15071), .A2(n10827), .ZN(n15057) );
  NAND2_X1 U13340 ( .A1(n15077), .A2(n15057), .ZN(n15074) );
  INV_X1 U13341 ( .A(n15074), .ZN(n11356) );
  AOI22_X1 U13342 ( .A1(n13026), .A2(n10698), .B1(n13069), .B2(n10697), .ZN(
        n10699) );
  OAI21_X1 U13343 ( .B1(n11051), .B2(n15077), .A(n10699), .ZN(n10700) );
  AOI21_X1 U13344 ( .B1(n11356), .B2(n15100), .A(n10700), .ZN(n10701) );
  OAI21_X1 U13345 ( .B1(n10702), .B2(n13011), .A(n10701), .ZN(P3_U3228) );
  OAI22_X1 U13346 ( .A1(n14196), .A2(n10704), .B1(n10703), .B2(n14637), .ZN(
        n10707) );
  MUX2_X1 U13347 ( .A(n10705), .B(P1_REG2_REG_2__SCAN_IN), .S(n14642), .Z(
        n10706) );
  AOI211_X1 U13348 ( .C1(n14512), .C2(n10708), .A(n10707), .B(n10706), .ZN(
        n10709) );
  INV_X1 U13349 ( .A(n10709), .ZN(P1_U3291) );
  NAND2_X1 U13350 ( .A1(n11185), .A2(n13373), .ZN(n10710) );
  NAND2_X1 U13351 ( .A1(n6567), .A2(n10710), .ZN(n10711) );
  INV_X1 U13352 ( .A(n10712), .ZN(n10713) );
  OAI22_X1 U13353 ( .A1(n14803), .A2(n10715), .B1(n13571), .B2(n10714), .ZN(
        n10716) );
  AOI21_X1 U13354 ( .B1(n10717), .B2(n14797), .A(n10716), .ZN(n10720) );
  MUX2_X1 U13355 ( .A(n10175), .B(n10718), .S(n13562), .Z(n10719) );
  OAI211_X1 U13356 ( .C1(n10721), .C2(n13576), .A(n10720), .B(n10719), .ZN(
        P2_U3259) );
  MUX2_X1 U13357 ( .A(n10723), .B(n10722), .S(n6569), .Z(n10727) );
  AOI22_X1 U13358 ( .A1(n13284), .A2(n13325), .B1(n10807), .B2(n13302), .ZN(
        n10726) );
  INV_X1 U13359 ( .A(n10724), .ZN(n10732) );
  NAND2_X1 U13360 ( .A1(n10732), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n10725) );
  OAI211_X1 U13361 ( .C1(n10727), .C2(n13304), .A(n10726), .B(n10725), .ZN(
        P2_U3204) );
  INV_X1 U13362 ( .A(n10728), .ZN(n10729) );
  AOI21_X1 U13363 ( .B1(n10731), .B2(n10730), .A(n10729), .ZN(n10735) );
  AOI22_X1 U13364 ( .A1(n13282), .A2(n9734), .B1(n13284), .B2(n13323), .ZN(
        n10734) );
  AOI22_X1 U13365 ( .A1(n10732), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n6560), .B2(
        n13302), .ZN(n10733) );
  OAI211_X1 U13366 ( .C1(n10735), .C2(n13304), .A(n10734), .B(n10733), .ZN(
        P2_U3194) );
  XNOR2_X1 U13367 ( .A(n10736), .B(n10737), .ZN(n14675) );
  NOR2_X1 U13368 ( .A1(n10736), .A2(n14209), .ZN(n10743) );
  INV_X1 U13369 ( .A(n10738), .ZN(n10740) );
  NAND2_X1 U13370 ( .A1(n14632), .A2(n12100), .ZN(n10739) );
  NAND2_X1 U13371 ( .A1(n10740), .A2(n10739), .ZN(n10747) );
  MUX2_X1 U13372 ( .A(n10743), .B(n10742), .S(n10741), .Z(n10746) );
  AOI21_X1 U13373 ( .B1(n10342), .B2(n14209), .A(n14611), .ZN(n10745) );
  OAI21_X1 U13374 ( .B1(n10746), .B2(n10745), .A(n10744), .ZN(n14673) );
  MUX2_X1 U13375 ( .A(n14673), .B(P1_REG2_REG_1__SCAN_IN), .S(n14642), .Z(
        n10750) );
  NOR2_X1 U13376 ( .A1(n10747), .A2(n14242), .ZN(n14670) );
  AOI22_X1 U13377 ( .A1(n14626), .A2(n14670), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14599), .ZN(n10748) );
  OAI21_X1 U13378 ( .B1(n14672), .B2(n14616), .A(n10748), .ZN(n10749) );
  AOI211_X1 U13379 ( .C1(n14627), .C2(n14675), .A(n10750), .B(n10749), .ZN(
        n10751) );
  INV_X1 U13380 ( .A(n10751), .ZN(P1_U3292) );
  XNOR2_X1 U13381 ( .A(n10753), .B(n10752), .ZN(n14846) );
  INV_X1 U13382 ( .A(n14846), .ZN(n10767) );
  OR2_X1 U13383 ( .A1(n10755), .A2(n10754), .ZN(n10756) );
  NAND2_X1 U13384 ( .A1(n10757), .A2(n10756), .ZN(n10759) );
  AOI21_X1 U13385 ( .B1(n10759), .B2(n13569), .A(n10758), .ZN(n14854) );
  MUX2_X1 U13386 ( .A(n14854), .B(n10173), .S(n14809), .Z(n10766) );
  OAI21_X1 U13387 ( .B1(n10794), .B2(n10762), .A(n11860), .ZN(n10760) );
  OR2_X1 U13388 ( .A1(n10917), .A2(n10760), .ZN(n14850) );
  INV_X1 U13389 ( .A(n14850), .ZN(n10764) );
  OAI22_X1 U13390 ( .A1(n14803), .A2(n10762), .B1(n13571), .B2(n10761), .ZN(
        n10763) );
  AOI21_X1 U13391 ( .B1(n14797), .B2(n10764), .A(n10763), .ZN(n10765) );
  OAI211_X1 U13392 ( .C1(n13576), .C2(n10767), .A(n10766), .B(n10765), .ZN(
        P2_U3261) );
  XNOR2_X1 U13393 ( .A(n10769), .B(n10768), .ZN(n14834) );
  NAND3_X1 U13394 ( .A1(n10771), .A2(n10770), .A3(n10799), .ZN(n10772) );
  NAND2_X1 U13395 ( .A1(n10772), .A2(n10784), .ZN(n10773) );
  AOI222_X1 U13396 ( .A1(n13569), .A2(n10773), .B1(n13322), .B2(n13538), .C1(
        n13325), .C2(n13540), .ZN(n14833) );
  MUX2_X1 U13397 ( .A(n10171), .B(n14833), .S(n13562), .Z(n10779) );
  XNOR2_X1 U13398 ( .A(n10808), .B(n14831), .ZN(n10774) );
  NOR2_X1 U13399 ( .A1(n10774), .A2(n6569), .ZN(n14830) );
  OAI22_X1 U13400 ( .A1(n14803), .A2(n10776), .B1(n13571), .B2(n10775), .ZN(
        n10777) );
  AOI21_X1 U13401 ( .B1(n14797), .B2(n14830), .A(n10777), .ZN(n10778) );
  OAI211_X1 U13402 ( .C1(n14834), .C2(n13576), .A(n10779), .B(n10778), .ZN(
        P2_U3263) );
  XNOR2_X1 U13403 ( .A(n10781), .B(n10780), .ZN(n14841) );
  NAND3_X1 U13404 ( .A1(n10784), .A2(n10783), .A3(n10782), .ZN(n10785) );
  NAND2_X1 U13405 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  NAND2_X1 U13406 ( .A1(n10787), .A2(n13569), .ZN(n10789) );
  AOI22_X1 U13407 ( .A1(n13540), .A2(n13323), .B1(n13321), .B2(n13538), .ZN(
        n10788) );
  AND2_X1 U13408 ( .A1(n10789), .A2(n10788), .ZN(n14844) );
  MUX2_X1 U13409 ( .A(n14844), .B(n10790), .S(n14809), .Z(n10798) );
  NAND2_X1 U13410 ( .A1(n10791), .A2(n14837), .ZN(n10792) );
  NAND2_X1 U13411 ( .A1(n10792), .A2(n11860), .ZN(n10793) );
  NOR2_X1 U13412 ( .A1(n10794), .A2(n10793), .ZN(n14839) );
  OAI22_X1 U13413 ( .A1(n14803), .A2(n10795), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13571), .ZN(n10796) );
  AOI21_X1 U13414 ( .B1(n14797), .B2(n14839), .A(n10796), .ZN(n10797) );
  OAI211_X1 U13415 ( .C1(n14841), .C2(n13576), .A(n10798), .B(n10797), .ZN(
        P2_U3262) );
  OAI21_X1 U13416 ( .B1(n10800), .B2(n10803), .A(n10799), .ZN(n10806) );
  OAI22_X1 U13417 ( .A1(n10801), .A2(n13524), .B1(n10619), .B2(n13522), .ZN(
        n10805) );
  XNOR2_X1 U13418 ( .A(n10802), .B(n10803), .ZN(n10814) );
  INV_X1 U13419 ( .A(n10814), .ZN(n14826) );
  NOR2_X1 U13420 ( .A1(n14826), .A2(n11185), .ZN(n10804) );
  AOI211_X1 U13421 ( .C1(n13569), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        n14825) );
  AOI21_X1 U13422 ( .B1(n10807), .B2(n6560), .A(n8811), .ZN(n10809) );
  AND2_X1 U13423 ( .A1(n10809), .A2(n10808), .ZN(n14823) );
  NAND2_X1 U13424 ( .A1(n14797), .A2(n14823), .ZN(n10811) );
  AOI22_X1 U13425 ( .A1(n13469), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n14800), 
        .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10810) );
  OAI211_X1 U13426 ( .C1(n14803), .C2(n10812), .A(n10811), .B(n10810), .ZN(
        n10813) );
  AOI21_X1 U13427 ( .B1(n11341), .B2(n10814), .A(n10813), .ZN(n10815) );
  OAI21_X1 U13428 ( .B1(n14825), .B2(n13469), .A(n10815), .ZN(P2_U3264) );
  XNOR2_X1 U13429 ( .A(n10816), .B(n12302), .ZN(n14676) );
  XNOR2_X1 U13430 ( .A(n10817), .B(n12302), .ZN(n10818) );
  AOI222_X1 U13431 ( .A1(n13859), .A2(n14209), .B1(n13857), .B2(n14207), .C1(
        n14611), .C2(n10818), .ZN(n14678) );
  MUX2_X1 U13432 ( .A(n10819), .B(n14678), .S(n14226), .Z(n10824) );
  OAI211_X1 U13433 ( .C1(n7440), .C2(n7439), .A(n14622), .B(n14620), .ZN(
        n14677) );
  OAI22_X1 U13434 ( .A1(n14196), .A2(n14677), .B1(n14637), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n10821) );
  AOI21_X1 U13435 ( .B1(n14512), .B2(n10822), .A(n10821), .ZN(n10823) );
  OAI211_X1 U13436 ( .C1(n14676), .C2(n14249), .A(n10824), .B(n10823), .ZN(
        P1_U3290) );
  INV_X1 U13437 ( .A(SI_21_), .ZN(n10826) );
  OAI222_X1 U13438 ( .A1(P3_U3151), .A2(n10827), .B1(n15456), .B2(n10826), 
        .C1(n15458), .C2(n10825), .ZN(P3_U3274) );
  OR2_X1 U13439 ( .A1(n10835), .A2(n13319), .ZN(n10828) );
  INV_X1 U13440 ( .A(n10838), .ZN(n10830) );
  OAI21_X1 U13441 ( .B1(n10831), .B2(n10830), .A(n10968), .ZN(n14805) );
  INV_X1 U13442 ( .A(n14805), .ZN(n10845) );
  NAND2_X1 U13443 ( .A1(n10833), .A2(n10832), .ZN(n10837) );
  NAND2_X1 U13444 ( .A1(n10835), .A2(n10834), .ZN(n10836) );
  NAND2_X1 U13445 ( .A1(n10837), .A2(n10836), .ZN(n10974) );
  XNOR2_X1 U13446 ( .A(n10974), .B(n10838), .ZN(n10841) );
  NAND2_X1 U13447 ( .A1(n13319), .A2(n13540), .ZN(n10840) );
  NAND2_X1 U13448 ( .A1(n13317), .A2(n13538), .ZN(n10839) );
  NAND2_X1 U13449 ( .A1(n10840), .A2(n10839), .ZN(n10905) );
  AOI21_X1 U13450 ( .B1(n10841), .B2(n13569), .A(n10905), .ZN(n14808) );
  INV_X1 U13451 ( .A(n10982), .ZN(n10842) );
  AOI211_X1 U13452 ( .C1(n14796), .C2(n10843), .A(n6569), .B(n10842), .ZN(
        n14798) );
  AOI21_X1 U13453 ( .B1(n14847), .B2(n14796), .A(n14798), .ZN(n10844) );
  OAI211_X1 U13454 ( .C1(n10845), .C2(n14840), .A(n14808), .B(n10844), .ZN(
        n10847) );
  NAND2_X1 U13455 ( .A1(n10847), .A2(n14891), .ZN(n10846) );
  OAI21_X1 U13456 ( .B1(n14891), .B2(n10163), .A(n10846), .ZN(P2_U3506) );
  INV_X1 U13457 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10849) );
  NAND2_X1 U13458 ( .A1(n10847), .A2(n14880), .ZN(n10848) );
  OAI21_X1 U13459 ( .B1(n14880), .B2(n10849), .A(n10848), .ZN(P2_U3451) );
  OAI22_X1 U13460 ( .A1(n12761), .A2(P3_U3151), .B1(SI_22_), .B2(n15456), .ZN(
        n10850) );
  AOI21_X1 U13461 ( .B1(n10851), .B2(n14387), .A(n10850), .ZN(P3_U3273) );
  INV_X1 U13462 ( .A(n10852), .ZN(n10854) );
  OAI222_X1 U13463 ( .A1(n14014), .A2(P1_U3086), .B1(n14369), .B2(n10854), 
        .C1(n10853), .C2(n14366), .ZN(P1_U3336) );
  OAI222_X1 U13464 ( .A1(n12073), .A2(n10855), .B1(n12071), .B2(n10854), .C1(
        n13373), .C2(P2_U3088), .ZN(P2_U3308) );
  OR2_X1 U13465 ( .A1(n15118), .A2(n15057), .ZN(n10856) );
  XNOR2_X1 U13466 ( .A(n10857), .B(n10859), .ZN(n15092) );
  OAI211_X1 U13467 ( .C1(n10860), .C2(n10859), .A(n10858), .B(n15067), .ZN(
        n10862) );
  AND2_X1 U13468 ( .A1(n10862), .A2(n10861), .ZN(n15093) );
  MUX2_X1 U13469 ( .A(n15093), .B(n11044), .S(n15079), .Z(n10866) );
  INV_X1 U13470 ( .A(n10863), .ZN(n10864) );
  AOI22_X1 U13471 ( .A1(n13026), .A2(n15096), .B1(n13069), .B2(n10864), .ZN(
        n10865) );
  OAI211_X1 U13472 ( .C1(n13029), .C2(n15092), .A(n10866), .B(n10865), .ZN(
        P3_U3229) );
  XNOR2_X1 U13473 ( .A(n10867), .B(n12593), .ZN(n15091) );
  INV_X1 U13474 ( .A(n15091), .ZN(n10877) );
  AOI21_X1 U13475 ( .B1(n10868), .B2(n12593), .A(n13063), .ZN(n10872) );
  INV_X1 U13476 ( .A(n10869), .ZN(n10870) );
  AOI21_X1 U13477 ( .B1(n10872), .B2(n10871), .A(n10870), .ZN(n15088) );
  MUX2_X1 U13478 ( .A(n15088), .B(n11037), .S(n15079), .Z(n10876) );
  INV_X1 U13479 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13480 ( .A1(n13026), .A2(n10874), .B1(n13069), .B2(n10873), .ZN(
        n10875) );
  OAI211_X1 U13481 ( .C1(n13029), .C2(n10877), .A(n10876), .B(n10875), .ZN(
        P3_U3230) );
  INV_X1 U13482 ( .A(n11141), .ZN(n14865) );
  OAI21_X1 U13483 ( .B1(n10880), .B2(n10879), .A(n10878), .ZN(n10881) );
  NAND2_X1 U13484 ( .A1(n10881), .A2(n13278), .ZN(n10885) );
  AND2_X1 U13485 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14735) );
  INV_X1 U13486 ( .A(n10984), .ZN(n10882) );
  OAI22_X1 U13487 ( .A1(n13299), .A2(n11181), .B1(n13297), .B2(n10882), .ZN(
        n10883) );
  AOI211_X1 U13488 ( .C1(n13282), .C2(n13318), .A(n14735), .B(n10883), .ZN(
        n10884) );
  OAI211_X1 U13489 ( .C1(n14865), .C2(n11948), .A(n10885), .B(n10884), .ZN(
        P2_U3193) );
  OAI211_X1 U13490 ( .C1(n10888), .C2(n10887), .A(n10886), .B(n14439), .ZN(
        n10893) );
  NAND2_X1 U13491 ( .A1(n12778), .A2(n15061), .ZN(n10890) );
  NAND2_X1 U13492 ( .A1(n12776), .A2(n15064), .ZN(n10889) );
  AND2_X1 U13493 ( .A1(n10890), .A2(n10889), .ZN(n11115) );
  INV_X1 U13494 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n14978) );
  OAI22_X1 U13495 ( .A1(n14446), .A2(n11115), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14978), .ZN(n10891) );
  AOI21_X1 U13496 ( .B1(n12661), .B2(n14441), .A(n10891), .ZN(n10892) );
  OAI211_X1 U13497 ( .C1(n11118), .C2(n14433), .A(n10893), .B(n10892), .ZN(
        P3_U3153) );
  XNOR2_X1 U13498 ( .A(n10894), .B(n10896), .ZN(n15101) );
  OAI211_X1 U13499 ( .C1(n10897), .C2(n10896), .A(n10895), .B(n15067), .ZN(
        n10901) );
  NAND2_X1 U13500 ( .A1(n12779), .A2(n15061), .ZN(n10899) );
  NAND2_X1 U13501 ( .A1(n12777), .A2(n15064), .ZN(n10898) );
  NAND2_X1 U13502 ( .A1(n10899), .A2(n10898), .ZN(n10989) );
  INV_X1 U13503 ( .A(n10989), .ZN(n10900) );
  NAND2_X1 U13504 ( .A1(n10901), .A2(n10900), .ZN(n15102) );
  MUX2_X1 U13505 ( .A(n15102), .B(P3_REG2_REG_6__SCAN_IN), .S(n15079), .Z(
        n10902) );
  INV_X1 U13506 ( .A(n10902), .ZN(n10904) );
  AOI22_X1 U13507 ( .A1(n13026), .A2(n15104), .B1(n13069), .B2(n10996), .ZN(
        n10903) );
  OAI211_X1 U13508 ( .C1(n13029), .C2(n15101), .A(n10904), .B(n10903), .ZN(
        P3_U3227) );
  INV_X1 U13509 ( .A(n10905), .ZN(n10908) );
  NAND2_X1 U13510 ( .A1(n13283), .A2(n14799), .ZN(n10907) );
  OAI211_X1 U13511 ( .C1(n10908), .C2(n13252), .A(n10907), .B(n10906), .ZN(
        n10913) );
  XNOR2_X1 U13512 ( .A(n10910), .B(n10909), .ZN(n10911) );
  NOR2_X1 U13513 ( .A1(n10911), .A2(n13304), .ZN(n10912) );
  AOI211_X1 U13514 ( .C1(n14796), .C2(n13302), .A(n10913), .B(n10912), .ZN(
        n10914) );
  INV_X1 U13515 ( .A(n10914), .ZN(P2_U3185) );
  XOR2_X1 U13516 ( .A(n10915), .B(n10921), .Z(n14861) );
  OAI211_X1 U13517 ( .C1(n14858), .C2(n10917), .A(n10916), .B(n11860), .ZN(
        n14856) );
  AOI22_X1 U13518 ( .A1(n13547), .A2(n10919), .B1(n14800), .B2(n10918), .ZN(
        n10920) );
  OAI21_X1 U13519 ( .B1(n13494), .B2(n14856), .A(n10920), .ZN(n10926) );
  XOR2_X1 U13520 ( .A(n10922), .B(n10921), .Z(n10924) );
  OAI21_X1 U13521 ( .B1(n10924), .B2(n13520), .A(n10923), .ZN(n14860) );
  MUX2_X1 U13522 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n14860), .S(n13562), .Z(
        n10925) );
  AOI211_X1 U13523 ( .C1(n14861), .C2(n14806), .A(n10926), .B(n10925), .ZN(
        n10927) );
  INV_X1 U13524 ( .A(n10927), .ZN(P2_U3260) );
  INV_X1 U13525 ( .A(n10928), .ZN(n10929) );
  OAI22_X1 U13526 ( .A1(n12394), .A2(n12114), .B1(n14684), .B2(n12395), .ZN(
        n11207) );
  INV_X1 U13527 ( .A(n11207), .ZN(n10933) );
  XNOR2_X1 U13528 ( .A(n11208), .B(n10933), .ZN(n11211) );
  OAI22_X1 U13529 ( .A1(n12114), .A2(n12395), .B1(n14684), .B2(n12396), .ZN(
        n10934) );
  XNOR2_X1 U13530 ( .A(n10934), .B(n12450), .ZN(n11210) );
  XNOR2_X1 U13531 ( .A(n11211), .B(n11210), .ZN(n10940) );
  NAND2_X1 U13532 ( .A1(n13858), .A2(n14209), .ZN(n10936) );
  NAND2_X1 U13533 ( .A1(n14207), .A2(n13856), .ZN(n10935) );
  AND2_X1 U13534 ( .A1(n10936), .A2(n10935), .ZN(n14609) );
  NAND2_X1 U13535 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13919) );
  OAI21_X1 U13536 ( .B1(n13811), .B2(n14609), .A(n13919), .ZN(n10938) );
  NOR2_X1 U13537 ( .A1(n13832), .A2(n14613), .ZN(n10937) );
  AOI211_X1 U13538 ( .C1(n13834), .C2(n12115), .A(n10938), .B(n10937), .ZN(
        n10939) );
  OAI21_X1 U13539 ( .B1(n10940), .B2(n13836), .A(n10939), .ZN(P1_U3230) );
  NAND2_X1 U13540 ( .A1(n10942), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10941) );
  OAI21_X1 U13541 ( .B1(n10942), .B2(n12588), .A(n10941), .ZN(P3_U3521) );
  INV_X1 U13542 ( .A(n11334), .ZN(n11239) );
  OAI21_X1 U13543 ( .B1(n10945), .B2(n10944), .A(n10943), .ZN(n10946) );
  NAND2_X1 U13544 ( .A1(n10946), .A2(n13278), .ZN(n10952) );
  INV_X1 U13545 ( .A(n10947), .ZN(n10950) );
  INV_X1 U13546 ( .A(n11333), .ZN(n10948) );
  OAI22_X1 U13547 ( .A1(n13299), .A2(n11152), .B1(n13297), .B2(n10948), .ZN(
        n10949) );
  AOI211_X1 U13548 ( .C1(n13282), .C2(n13317), .A(n10950), .B(n10949), .ZN(
        n10951) );
  OAI211_X1 U13549 ( .C1(n11239), .C2(n11948), .A(n10952), .B(n10951), .ZN(
        P2_U3203) );
  INV_X1 U13550 ( .A(n10953), .ZN(n11231) );
  OAI211_X1 U13551 ( .C1(n10956), .C2(n10955), .A(n10954), .B(n14439), .ZN(
        n10963) );
  NAND2_X1 U13552 ( .A1(n12777), .A2(n15061), .ZN(n10958) );
  NAND2_X1 U13553 ( .A1(n12775), .A2(n15064), .ZN(n10957) );
  AND2_X1 U13554 ( .A1(n10958), .A2(n10957), .ZN(n11229) );
  OAI22_X1 U13555 ( .A1(n14446), .A2(n11229), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10959), .ZN(n10960) );
  AOI21_X1 U13556 ( .B1(n14441), .B2(n10961), .A(n10960), .ZN(n10962) );
  OAI211_X1 U13557 ( .C1(n11231), .C2(n14433), .A(n10963), .B(n10962), .ZN(
        P3_U3161) );
  INV_X1 U13558 ( .A(n10964), .ZN(n10966) );
  NAND2_X1 U13559 ( .A1(n14386), .A2(SI_23_), .ZN(n10965) );
  OAI211_X1 U13560 ( .C1(n10966), .C2(n15458), .A(n12764), .B(n10965), .ZN(
        P3_U3272) );
  OR2_X1 U13561 ( .A1(n14796), .A2(n13318), .ZN(n10967) );
  INV_X1 U13562 ( .A(n10970), .ZN(n10969) );
  INV_X1 U13563 ( .A(n10975), .ZN(n11138) );
  NAND2_X1 U13564 ( .A1(n10970), .A2(n11138), .ZN(n10971) );
  NAND2_X1 U13565 ( .A1(n11136), .A2(n10971), .ZN(n10980) );
  AOI22_X1 U13566 ( .A1(n13540), .A2(n13318), .B1(n13316), .B2(n13538), .ZN(
        n10978) );
  AND2_X1 U13567 ( .A1(n14796), .A2(n10972), .ZN(n10973) );
  XNOR2_X1 U13568 ( .A(n11139), .B(n10975), .ZN(n10976) );
  NAND2_X1 U13569 ( .A1(n10976), .A2(n13569), .ZN(n10977) );
  OAI211_X1 U13570 ( .C1(n10980), .C2(n11185), .A(n10978), .B(n10977), .ZN(
        n14866) );
  MUX2_X1 U13571 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n14866), .S(n13562), .Z(
        n10979) );
  INV_X1 U13572 ( .A(n10979), .ZN(n10988) );
  INV_X1 U13573 ( .A(n10980), .ZN(n14868) );
  NAND2_X1 U13574 ( .A1(n10982), .A2(n11141), .ZN(n10981) );
  NAND2_X1 U13575 ( .A1(n10981), .A2(n11860), .ZN(n10983) );
  OR2_X1 U13576 ( .A1(n10983), .A2(n11238), .ZN(n14864) );
  AOI22_X1 U13577 ( .A1(n13547), .A2(n11141), .B1(n14800), .B2(n10984), .ZN(
        n10985) );
  OAI21_X1 U13578 ( .B1(n14864), .B2(n13494), .A(n10985), .ZN(n10986) );
  AOI21_X1 U13579 ( .B1(n14868), .B2(n11341), .A(n10986), .ZN(n10987) );
  NAND2_X1 U13580 ( .A1(n10988), .A2(n10987), .ZN(P2_U3257) );
  AOI22_X1 U13581 ( .A1(n12510), .A2(n10989), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10990) );
  OAI21_X1 U13582 ( .B1(n10991), .B2(n12574), .A(n10990), .ZN(n10995) );
  AOI211_X1 U13583 ( .C1(n10993), .C2(n10992), .A(n14427), .B(n6735), .ZN(
        n10994) );
  AOI211_X1 U13584 ( .C1(n10996), .C2(n14444), .A(n10995), .B(n10994), .ZN(
        n10997) );
  INV_X1 U13585 ( .A(n10997), .ZN(P3_U3179) );
  XNOR2_X1 U13586 ( .A(n10999), .B(n10998), .ZN(n11004) );
  OAI22_X1 U13587 ( .A1(n13295), .A2(n11181), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8573), .ZN(n11002) );
  INV_X1 U13588 ( .A(n13314), .ZN(n11250) );
  INV_X1 U13589 ( .A(n11000), .ZN(n11186) );
  OAI22_X1 U13590 ( .A1(n13299), .A2(n11250), .B1(n13297), .B2(n11186), .ZN(
        n11001) );
  AOI211_X1 U13591 ( .C1(n11190), .C2(n13302), .A(n11002), .B(n11001), .ZN(
        n11003) );
  OAI21_X1 U13592 ( .B1(n11004), .B2(n13304), .A(n11003), .ZN(P2_U3189) );
  INV_X1 U13593 ( .A(n14384), .ZN(n15022) );
  INV_X1 U13594 ( .A(n14986), .ZN(n11065) );
  NAND2_X1 U13595 ( .A1(n6564), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11005) );
  XNOR2_X1 U13596 ( .A(n11046), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n14923) );
  NOR2_X1 U13597 ( .A1(n14951), .A2(n11009), .ZN(n11010) );
  NAND2_X1 U13598 ( .A1(n14972), .A2(n11058), .ZN(n11011) );
  NAND2_X1 U13599 ( .A1(n11012), .A2(n11011), .ZN(n14957) );
  NOR2_X1 U13600 ( .A1(n11065), .A2(n11013), .ZN(n11014) );
  NAND2_X1 U13601 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11072), .ZN(n11015) );
  OAI21_X1 U13602 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11072), .A(n11015), .ZN(
        n14997) );
  NOR2_X1 U13603 ( .A1(n15022), .A2(n11016), .ZN(n11017) );
  NAND2_X1 U13604 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11462), .ZN(n11018) );
  OAI21_X1 U13605 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11462), .A(n11018), 
        .ZN(n11019) );
  AOI21_X1 U13606 ( .B1(n11020), .B2(n11019), .A(n11456), .ZN(n11095) );
  INV_X1 U13607 ( .A(n11462), .ZN(n11083) );
  INV_X1 U13608 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U13609 ( .A1(n11083), .A2(n15142), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11462), .ZN(n11034) );
  NAND2_X1 U13610 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11072), .ZN(n11030) );
  INV_X1 U13611 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U13612 ( .A1(n15002), .A2(n15138), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n11072), .ZN(n15001) );
  NAND2_X1 U13613 ( .A1(n11060), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11027) );
  INV_X1 U13614 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11057) );
  MUX2_X1 U13615 ( .A(n11057), .B(P3_REG1_REG_6__SCAN_IN), .S(n14972), .Z(
        n14960) );
  NAND2_X1 U13616 ( .A1(n11046), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n11024) );
  INV_X1 U13617 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11043) );
  MUX2_X1 U13618 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n11043), .S(n11046), .Z(
        n14926) );
  AOI21_X1 U13619 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n6564), .A(n11021), .ZN(
        n11023) );
  INV_X1 U13620 ( .A(n11039), .ZN(n14913) );
  XNOR2_X1 U13621 ( .A(n11023), .B(n14913), .ZN(n14907) );
  INV_X1 U13622 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11036) );
  OAI22_X1 U13623 ( .A1(n14907), .A2(n11036), .B1(n14913), .B2(n11023), .ZN(
        n14927) );
  NAND2_X1 U13624 ( .A1(n11053), .A2(n11025), .ZN(n11026) );
  NAND2_X1 U13625 ( .A1(n14960), .A2(n14961), .ZN(n14959) );
  NAND2_X1 U13626 ( .A1(n14986), .A2(n11028), .ZN(n11029) );
  NAND2_X1 U13627 ( .A1(n15001), .A2(n15000), .ZN(n14999) );
  NAND2_X1 U13628 ( .A1(n14384), .A2(n11031), .ZN(n11032) );
  OAI21_X1 U13629 ( .B1(n11034), .B2(n11033), .A(n11463), .ZN(n11093) );
  NAND2_X1 U13630 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11532)
         );
  NAND2_X1 U13631 ( .A1(n14990), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11035) );
  OAI211_X1 U13632 ( .C1(n14985), .C2(n11462), .A(n11532), .B(n11035), .ZN(
        n11092) );
  NAND2_X1 U13633 ( .A1(n14903), .A2(n14902), .ZN(n11042) );
  MUX2_X1 U13634 ( .A(n11037), .B(n11036), .S(n6973), .Z(n11038) );
  NAND2_X1 U13635 ( .A1(n11038), .A2(n14913), .ZN(n14919) );
  INV_X1 U13636 ( .A(n11038), .ZN(n11040) );
  NAND2_X1 U13637 ( .A1(n11040), .A2(n11039), .ZN(n11041) );
  AND2_X1 U13638 ( .A1(n14919), .A2(n11041), .ZN(n14900) );
  NAND2_X1 U13639 ( .A1(n14920), .A2(n14919), .ZN(n11049) );
  MUX2_X1 U13640 ( .A(n11044), .B(n11043), .S(n6973), .Z(n11045) );
  INV_X1 U13641 ( .A(n11046), .ZN(n14933) );
  NAND2_X1 U13642 ( .A1(n11045), .A2(n14933), .ZN(n14939) );
  INV_X1 U13643 ( .A(n11045), .ZN(n11047) );
  NAND2_X1 U13644 ( .A1(n11047), .A2(n11046), .ZN(n11048) );
  AND2_X1 U13645 ( .A1(n14939), .A2(n11048), .ZN(n14917) );
  NAND2_X1 U13646 ( .A1(n11049), .A2(n14917), .ZN(n14940) );
  NAND2_X1 U13647 ( .A1(n14940), .A2(n14939), .ZN(n11056) );
  INV_X1 U13648 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11050) );
  MUX2_X1 U13649 ( .A(n11051), .B(n11050), .S(n6973), .Z(n11052) );
  NAND2_X1 U13650 ( .A1(n11052), .A2(n14951), .ZN(n14967) );
  INV_X1 U13651 ( .A(n11052), .ZN(n11054) );
  NAND2_X1 U13652 ( .A1(n11054), .A2(n11053), .ZN(n11055) );
  AND2_X1 U13653 ( .A1(n14967), .A2(n11055), .ZN(n14937) );
  NAND2_X1 U13654 ( .A1(n14968), .A2(n14967), .ZN(n11063) );
  MUX2_X1 U13655 ( .A(n11058), .B(n11057), .S(n6973), .Z(n11059) );
  NAND2_X1 U13656 ( .A1(n11059), .A2(n14972), .ZN(n14979) );
  INV_X1 U13657 ( .A(n11059), .ZN(n11061) );
  NAND2_X1 U13658 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  AND2_X1 U13659 ( .A1(n14979), .A2(n11062), .ZN(n14965) );
  NAND2_X1 U13660 ( .A1(n14983), .A2(n14979), .ZN(n11069) );
  INV_X1 U13661 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11064) );
  MUX2_X1 U13662 ( .A(n11117), .B(n11064), .S(n6973), .Z(n11066) );
  NAND2_X1 U13663 ( .A1(n11066), .A2(n11065), .ZN(n15008) );
  INV_X1 U13664 ( .A(n11066), .ZN(n11067) );
  NAND2_X1 U13665 ( .A1(n11067), .A2(n14986), .ZN(n11068) );
  AND2_X1 U13666 ( .A1(n15008), .A2(n11068), .ZN(n14981) );
  NAND2_X1 U13667 ( .A1(n11069), .A2(n14981), .ZN(n15009) );
  NAND2_X1 U13668 ( .A1(n15009), .A2(n15008), .ZN(n11075) );
  MUX2_X1 U13669 ( .A(n11070), .B(n15138), .S(n6973), .Z(n11071) );
  NAND2_X1 U13670 ( .A1(n11071), .A2(n15002), .ZN(n15026) );
  INV_X1 U13671 ( .A(n11071), .ZN(n11073) );
  NAND2_X1 U13672 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  AND2_X1 U13673 ( .A1(n15026), .A2(n11074), .ZN(n15006) );
  NAND2_X1 U13674 ( .A1(n15025), .A2(n15026), .ZN(n11081) );
  INV_X1 U13675 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11076) );
  MUX2_X1 U13676 ( .A(n11077), .B(n11076), .S(n6973), .Z(n11078) );
  NAND2_X1 U13677 ( .A1(n11078), .A2(n15022), .ZN(n11089) );
  INV_X1 U13678 ( .A(n11078), .ZN(n11079) );
  NAND2_X1 U13679 ( .A1(n11079), .A2(n14384), .ZN(n11080) );
  AND2_X1 U13680 ( .A1(n11089), .A2(n11080), .ZN(n15027) );
  NAND2_X1 U13681 ( .A1(n11081), .A2(n15027), .ZN(n15030) );
  MUX2_X1 U13682 ( .A(n11082), .B(n15142), .S(n6973), .Z(n11084) );
  NAND2_X1 U13683 ( .A1(n11084), .A2(n11083), .ZN(n11458) );
  INV_X1 U13684 ( .A(n11084), .ZN(n11085) );
  NAND2_X1 U13685 ( .A1(n11085), .A2(n11462), .ZN(n11086) );
  AND2_X1 U13686 ( .A1(n11458), .A2(n11086), .ZN(n11087) );
  INV_X1 U13687 ( .A(n11087), .ZN(n11088) );
  NAND3_X1 U13688 ( .A1(n15030), .A2(n11089), .A3(n11088), .ZN(n11090) );
  AOI21_X1 U13689 ( .B1(n11459), .B2(n11090), .A(n15010), .ZN(n11091) );
  AOI211_X1 U13690 ( .C1(n15023), .C2(n11093), .A(n11092), .B(n11091), .ZN(
        n11094) );
  OAI21_X1 U13691 ( .B1(n11095), .B2(n15036), .A(n11094), .ZN(P3_U3192) );
  INV_X1 U13692 ( .A(n11991), .ZN(n11097) );
  INV_X1 U13693 ( .A(n11161), .ZN(n11096) );
  AOI211_X1 U13694 ( .C1(n14696), .C2(n11097), .A(n14242), .B(n11096), .ZN(
        n14695) );
  INV_X1 U13695 ( .A(n11098), .ZN(n11307) );
  OAI22_X1 U13696 ( .A1(n14616), .A2(n11311), .B1(n11307), .B2(n14637), .ZN(
        n11110) );
  OAI21_X1 U13697 ( .B1(n11101), .B2(n11100), .A(n11099), .ZN(n11102) );
  NAND2_X1 U13698 ( .A1(n11102), .A2(n14707), .ZN(n11108) );
  OAI21_X1 U13699 ( .B1(n11104), .B2(n12306), .A(n11103), .ZN(n11105) );
  NAND2_X1 U13700 ( .A1(n11105), .A2(n14611), .ZN(n11107) );
  AOI22_X1 U13701 ( .A1(n14207), .A2(n13854), .B1(n14209), .B2(n13856), .ZN(
        n11106) );
  NAND3_X1 U13702 ( .A1(n11108), .A2(n11107), .A3(n11106), .ZN(n14694) );
  MUX2_X1 U13703 ( .A(n14694), .B(P1_REG2_REG_6__SCAN_IN), .S(n14642), .Z(
        n11109) );
  AOI211_X1 U13704 ( .C1(n14626), .C2(n14695), .A(n11110), .B(n11109), .ZN(
        n11111) );
  INV_X1 U13705 ( .A(n11111), .ZN(P1_U3287) );
  XNOR2_X1 U13706 ( .A(n11112), .B(n12596), .ZN(n15109) );
  OAI211_X1 U13707 ( .C1(n11114), .C2(n12596), .A(n11113), .B(n15067), .ZN(
        n11116) );
  AND2_X1 U13708 ( .A1(n11116), .A2(n11115), .ZN(n15112) );
  MUX2_X1 U13709 ( .A(n15112), .B(n11117), .S(n15079), .Z(n11121) );
  INV_X1 U13710 ( .A(n11118), .ZN(n11119) );
  AOI22_X1 U13711 ( .A1(n13026), .A2(n12661), .B1(n13069), .B2(n11119), .ZN(
        n11120) );
  OAI211_X1 U13712 ( .C1(n13029), .C2(n15109), .A(n11121), .B(n11120), .ZN(
        P3_U3226) );
  NAND2_X1 U13713 ( .A1(n14207), .A2(n13852), .ZN(n11123) );
  NAND2_X1 U13714 ( .A1(n14209), .A2(n13854), .ZN(n11122) );
  AND2_X1 U13715 ( .A1(n11123), .A2(n11122), .ZN(n14700) );
  INV_X1 U13716 ( .A(n14700), .ZN(n11125) );
  AOI211_X1 U13717 ( .C1(n11130), .C2(n11124), .A(n14234), .B(n6736), .ZN(
        n14704) );
  AOI211_X1 U13718 ( .C1(n14599), .C2(n11584), .A(n11125), .B(n14704), .ZN(
        n11134) );
  NAND2_X1 U13719 ( .A1(n11159), .A2(n12132), .ZN(n11126) );
  NAND2_X1 U13720 ( .A1(n11126), .A2(n14622), .ZN(n11127) );
  NOR2_X1 U13721 ( .A1(n11274), .A2(n11127), .ZN(n14699) );
  INV_X1 U13722 ( .A(n12132), .ZN(n14703) );
  OAI22_X1 U13723 ( .A1(n14703), .A2(n14616), .B1(n14226), .B2(n10127), .ZN(
        n11128) );
  AOI21_X1 U13724 ( .B1(n14626), .B2(n14699), .A(n11128), .ZN(n11133) );
  OAI21_X1 U13725 ( .B1(n11131), .B2(n11130), .A(n11129), .ZN(n14706) );
  NAND2_X1 U13726 ( .A1(n14706), .A2(n14627), .ZN(n11132) );
  OAI211_X1 U13727 ( .C1(n11134), .C2(n14642), .A(n11133), .B(n11132), .ZN(
        P1_U3285) );
  NAND2_X1 U13728 ( .A1(n11141), .A2(n13317), .ZN(n11135) );
  NAND2_X1 U13729 ( .A1(n11190), .A2(n13315), .ZN(n11137) );
  XNOR2_X1 U13730 ( .A(n11248), .B(n7311), .ZN(n11391) );
  INV_X1 U13731 ( .A(n13313), .ZN(n11424) );
  NAND2_X1 U13732 ( .A1(n11139), .A2(n11138), .ZN(n11143) );
  OR2_X1 U13733 ( .A1(n11141), .A2(n11140), .ZN(n11142) );
  NAND2_X1 U13734 ( .A1(n11143), .A2(n11142), .ZN(n11241) );
  INV_X1 U13735 ( .A(n11144), .ZN(n11240) );
  NAND2_X1 U13736 ( .A1(n11241), .A2(n11240), .ZN(n11146) );
  OR2_X1 U13737 ( .A1(n11334), .A2(n11181), .ZN(n11145) );
  NAND2_X1 U13738 ( .A1(n11146), .A2(n11145), .ZN(n11180) );
  INV_X1 U13739 ( .A(n11179), .ZN(n11147) );
  NAND2_X1 U13740 ( .A1(n11180), .A2(n11147), .ZN(n11149) );
  OR2_X1 U13741 ( .A1(n11190), .A2(n11152), .ZN(n11148) );
  NAND2_X1 U13742 ( .A1(n11149), .A2(n11148), .ZN(n11252) );
  XNOR2_X1 U13743 ( .A(n11252), .B(n11150), .ZN(n11151) );
  OAI222_X1 U13744 ( .A1(n13524), .A2(n11424), .B1(n13522), .B2(n11152), .C1(
        n11151), .C2(n13520), .ZN(n11387) );
  NAND2_X1 U13745 ( .A1(n11387), .A2(n13562), .ZN(n11158) );
  INV_X1 U13746 ( .A(n11190), .ZN(n14873) );
  NAND2_X1 U13747 ( .A1(n11236), .A2(n14873), .ZN(n11187) );
  OR2_X1 U13748 ( .A1(n11187), .A2(n11389), .ZN(n11255) );
  INV_X1 U13749 ( .A(n11255), .ZN(n11153) );
  AOI211_X1 U13750 ( .C1(n11389), .C2(n11187), .A(n8811), .B(n11153), .ZN(
        n11388) );
  INV_X1 U13751 ( .A(n11389), .ZN(n11155) );
  AOI22_X1 U13752 ( .A1(n13469), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n14800), 
        .B2(n11366), .ZN(n11154) );
  OAI21_X1 U13753 ( .B1(n11155), .B2(n14803), .A(n11154), .ZN(n11156) );
  AOI21_X1 U13754 ( .B1(n11388), .B2(n14797), .A(n11156), .ZN(n11157) );
  OAI211_X1 U13755 ( .C1(n11391), .C2(n13576), .A(n11158), .B(n11157), .ZN(
        P2_U3254) );
  INV_X1 U13756 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11171) );
  INV_X1 U13757 ( .A(n11159), .ZN(n11160) );
  AOI211_X1 U13758 ( .C1(n12129), .C2(n11161), .A(n14242), .B(n11160), .ZN(
        n11224) );
  XNOR2_X1 U13759 ( .A(n11162), .B(n11165), .ZN(n11169) );
  AOI22_X1 U13760 ( .A1(n14207), .A2(n13853), .B1(n14209), .B2(n13855), .ZN(
        n11168) );
  OAI21_X1 U13761 ( .B1(n11165), .B2(n11164), .A(n11163), .ZN(n11166) );
  NAND2_X1 U13762 ( .A1(n11166), .A2(n14707), .ZN(n11167) );
  OAI211_X1 U13763 ( .C1(n11169), .C2(n14234), .A(n11168), .B(n11167), .ZN(
        n11221) );
  AOI211_X1 U13764 ( .C1(n14697), .C2(n12129), .A(n11224), .B(n11221), .ZN(
        n11172) );
  OR2_X1 U13765 ( .A1(n11172), .A2(n14708), .ZN(n11170) );
  OAI21_X1 U13766 ( .B1(n14710), .B2(n11171), .A(n11170), .ZN(P1_U3480) );
  OR2_X1 U13767 ( .A1(n11172), .A2(n14718), .ZN(n11173) );
  OAI21_X1 U13768 ( .B1(n14720), .B2(n13943), .A(n11173), .ZN(P1_U3535) );
  OAI222_X1 U13769 ( .A1(P1_U3086), .A2(n12275), .B1(n12362), .B2(n11175), 
        .C1(n11174), .C2(n14366), .ZN(P1_U3335) );
  OAI222_X1 U13770 ( .A1(n12073), .A2(n11177), .B1(P2_U3088), .B2(n11176), 
        .C1(n12071), .C2(n11175), .ZN(P2_U3307) );
  XNOR2_X1 U13771 ( .A(n11178), .B(n11179), .ZN(n14870) );
  XNOR2_X1 U13772 ( .A(n11180), .B(n11179), .ZN(n11183) );
  OAI22_X1 U13773 ( .A1(n11181), .A2(n13522), .B1(n11250), .B2(n13524), .ZN(
        n11182) );
  AOI21_X1 U13774 ( .B1(n11183), .B2(n13569), .A(n11182), .ZN(n11184) );
  OAI21_X1 U13775 ( .B1(n14870), .B2(n11185), .A(n11184), .ZN(n14874) );
  NAND2_X1 U13776 ( .A1(n14874), .A2(n13562), .ZN(n11192) );
  OAI22_X1 U13777 ( .A1(n13562), .A2(n10393), .B1(n11186), .B2(n13571), .ZN(
        n11189) );
  OAI211_X1 U13778 ( .C1(n11236), .C2(n14873), .A(n11860), .B(n11187), .ZN(
        n14871) );
  NOR2_X1 U13779 ( .A1(n14871), .A2(n13494), .ZN(n11188) );
  AOI211_X1 U13780 ( .C1(n13547), .C2(n11190), .A(n11189), .B(n11188), .ZN(
        n11191) );
  OAI211_X1 U13781 ( .C1(n14870), .C2(n13410), .A(n11192), .B(n11191), .ZN(
        P2_U3255) );
  INV_X1 U13782 ( .A(n11193), .ZN(n11194) );
  AOI21_X1 U13783 ( .B1(n11196), .B2(n11195), .A(n11194), .ZN(n11201) );
  OAI22_X1 U13784 ( .A1(n12574), .A2(n15120), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15369), .ZN(n11199) );
  INV_X1 U13785 ( .A(n14416), .ZN(n12526) );
  OAI22_X1 U13786 ( .A1(n12526), .A2(n11448), .B1(n11197), .B2(n14418), .ZN(
        n11198) );
  AOI211_X1 U13787 ( .C1(n11287), .C2(n14444), .A(n11199), .B(n11198), .ZN(
        n11200) );
  OAI21_X1 U13788 ( .B1(n11201), .B2(n14427), .A(n11200), .ZN(P3_U3171) );
  NAND2_X1 U13789 ( .A1(n6962), .A2(n14692), .ZN(n11202) );
  OAI21_X1 U13790 ( .B1(n11204), .B2(n12391), .A(n11202), .ZN(n11203) );
  XNOR2_X1 U13791 ( .A(n11203), .B(n12450), .ZN(n11294) );
  OR2_X1 U13792 ( .A1(n12394), .A2(n11204), .ZN(n11206) );
  NAND2_X1 U13793 ( .A1(n12455), .A2(n14692), .ZN(n11205) );
  NAND2_X1 U13794 ( .A1(n11206), .A2(n11205), .ZN(n11293) );
  XOR2_X1 U13795 ( .A(n11294), .B(n11293), .Z(n11213) );
  NAND2_X1 U13796 ( .A1(n11212), .A2(n11213), .ZN(n11301) );
  OAI21_X1 U13797 ( .B1(n11213), .B2(n11212), .A(n11301), .ZN(n11214) );
  NAND2_X1 U13798 ( .A1(n11214), .A2(n13809), .ZN(n11219) );
  NAND2_X1 U13799 ( .A1(n13857), .A2(n14209), .ZN(n11216) );
  NAND2_X1 U13800 ( .A1(n14207), .A2(n13855), .ZN(n11215) );
  AND2_X1 U13801 ( .A1(n11216), .A2(n11215), .ZN(n11986) );
  NAND2_X1 U13802 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13925) );
  OAI21_X1 U13803 ( .B1(n13811), .B2(n11986), .A(n13925), .ZN(n11217) );
  AOI21_X1 U13804 ( .B1(n13834), .B2(n14692), .A(n11217), .ZN(n11218) );
  OAI211_X1 U13805 ( .C1(n13832), .C2(n11989), .A(n11219), .B(n11218), .ZN(
        P1_U3227) );
  INV_X1 U13806 ( .A(n12129), .ZN(n11220) );
  OAI22_X1 U13807 ( .A1(n14616), .A2(n11220), .B1(n14637), .B2(n11572), .ZN(
        n11223) );
  MUX2_X1 U13808 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11221), .S(n14226), .Z(
        n11222) );
  AOI211_X1 U13809 ( .C1(n14626), .C2(n11224), .A(n11223), .B(n11222), .ZN(
        n11225) );
  INV_X1 U13810 ( .A(n11225), .ZN(P1_U3286) );
  XOR2_X1 U13811 ( .A(n12665), .B(n11226), .Z(n15115) );
  INV_X1 U13812 ( .A(n11281), .ZN(n11227) );
  AOI21_X1 U13813 ( .B1(n12665), .B2(n11228), .A(n11227), .ZN(n11230) );
  OAI21_X1 U13814 ( .B1(n11230), .B2(n13063), .A(n11229), .ZN(n15116) );
  NAND2_X1 U13815 ( .A1(n15116), .A2(n15077), .ZN(n11234) );
  OAI22_X1 U13816 ( .A1(n13071), .A2(n15113), .B1(n11231), .B2(n15072), .ZN(
        n11232) );
  AOI21_X1 U13817 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15079), .A(n11232), .ZN(
        n11233) );
  OAI211_X1 U13818 ( .C1(n13029), .C2(n15115), .A(n11234), .B(n11233), .ZN(
        P3_U3225) );
  XNOR2_X1 U13819 ( .A(n11235), .B(n11240), .ZN(n11340) );
  INV_X1 U13820 ( .A(n11236), .ZN(n11237) );
  OAI211_X1 U13821 ( .C1(n11239), .C2(n11238), .A(n11237), .B(n11860), .ZN(
        n11336) );
  OAI21_X1 U13822 ( .B1(n11239), .B2(n14872), .A(n11336), .ZN(n11245) );
  XNOR2_X1 U13823 ( .A(n11241), .B(n11240), .ZN(n11244) );
  NAND2_X1 U13824 ( .A1(n11340), .A2(n14862), .ZN(n11243) );
  AOI22_X1 U13825 ( .A1(n13540), .A2(n13317), .B1(n13315), .B2(n13538), .ZN(
        n11242) );
  OAI211_X1 U13826 ( .C1(n13520), .C2(n11244), .A(n11243), .B(n11242), .ZN(
        n11337) );
  AOI211_X1 U13827 ( .C1(n14877), .C2(n11340), .A(n11245), .B(n11337), .ZN(
        n11343) );
  NAND2_X1 U13828 ( .A1(n14888), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11246) );
  OAI21_X1 U13829 ( .B1(n11343), .B2(n14888), .A(n11246), .ZN(P2_U3508) );
  AND2_X1 U13830 ( .A1(n11389), .A2(n13314), .ZN(n11247) );
  OR2_X1 U13831 ( .A1(n11389), .A2(n13314), .ZN(n11249) );
  XNOR2_X1 U13832 ( .A(n11429), .B(n11253), .ZN(n13669) );
  NAND2_X1 U13833 ( .A1(n11389), .A2(n11250), .ZN(n11251) );
  INV_X1 U13834 ( .A(n11253), .ZN(n11428) );
  OAI211_X1 U13835 ( .C1(n6721), .C2(n11253), .A(n13569), .B(n11425), .ZN(
        n11254) );
  AOI22_X1 U13836 ( .A1(n13540), .A2(n13314), .B1(n13312), .B2(n13538), .ZN(
        n11415) );
  NAND2_X1 U13837 ( .A1(n11254), .A2(n11415), .ZN(n13665) );
  INV_X1 U13838 ( .A(n13667), .ZN(n11420) );
  NAND2_X1 U13839 ( .A1(n13667), .A2(n11255), .ZN(n11256) );
  NAND2_X1 U13840 ( .A1(n11256), .A2(n11860), .ZN(n11257) );
  NOR2_X1 U13841 ( .A1(n11431), .A2(n11257), .ZN(n13666) );
  NAND2_X1 U13842 ( .A1(n13666), .A2(n14797), .ZN(n11259) );
  AOI22_X1 U13843 ( .A1(n13469), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n14800), 
        .B2(n11417), .ZN(n11258) );
  OAI211_X1 U13844 ( .C1(n11420), .C2(n14803), .A(n11259), .B(n11258), .ZN(
        n11260) );
  AOI21_X1 U13845 ( .B1(n13665), .B2(n13562), .A(n11260), .ZN(n11261) );
  OAI21_X1 U13846 ( .B1(n13576), .B2(n13669), .A(n11261), .ZN(P2_U3253) );
  OAI21_X1 U13847 ( .B1(n11264), .B2(n11263), .A(n11262), .ZN(n11272) );
  OAI22_X1 U13848 ( .A1(n14218), .A2(n11266), .B1(n11265), .B2(n14221), .ZN(
        n11271) );
  OAI21_X1 U13849 ( .B1(n12311), .B2(n11268), .A(n11267), .ZN(n11269) );
  AND2_X1 U13850 ( .A1(n11269), .A2(n14707), .ZN(n11270) );
  AOI211_X1 U13851 ( .C1(n14611), .C2(n11272), .A(n11271), .B(n11270), .ZN(
        n11499) );
  OAI22_X1 U13852 ( .A1(n14226), .A2(n11273), .B1(n11565), .B2(n14637), .ZN(
        n11277) );
  OAI21_X1 U13853 ( .B1(n11274), .B2(n11500), .A(n14622), .ZN(n11275) );
  OR2_X1 U13854 ( .A1(n11275), .A2(n11403), .ZN(n11498) );
  NOR2_X1 U13855 ( .A1(n11498), .A2(n14196), .ZN(n11276) );
  AOI211_X1 U13856 ( .C1(n14512), .C2(n12141), .A(n11277), .B(n11276), .ZN(
        n11278) );
  OAI21_X1 U13857 ( .B1(n11499), .B2(n14642), .A(n11278), .ZN(P1_U3284) );
  INV_X1 U13858 ( .A(n15118), .ZN(n15108) );
  XNOR2_X1 U13859 ( .A(n11279), .B(n12598), .ZN(n11286) );
  AND2_X1 U13860 ( .A1(n11281), .A2(n11280), .ZN(n11283) );
  OAI211_X1 U13861 ( .C1(n11283), .C2(n12598), .A(n11282), .B(n15067), .ZN(
        n11285) );
  AOI22_X1 U13862 ( .A1(n15061), .A2(n12776), .B1(n12774), .B2(n15064), .ZN(
        n11284) );
  OAI211_X1 U13863 ( .C1(n15108), .C2(n11286), .A(n11285), .B(n11284), .ZN(
        n15121) );
  INV_X1 U13864 ( .A(n15121), .ZN(n11292) );
  INV_X1 U13865 ( .A(n11286), .ZN(n15123) );
  AOI22_X1 U13866 ( .A1(n13026), .A2(n11288), .B1(n13069), .B2(n11287), .ZN(
        n11289) );
  OAI21_X1 U13867 ( .B1(n11077), .B2(n15077), .A(n11289), .ZN(n11290) );
  AOI21_X1 U13868 ( .B1(n15123), .B2(n11356), .A(n11290), .ZN(n11291) );
  OAI21_X1 U13869 ( .B1(n11292), .B2(n13011), .A(n11291), .ZN(P3_U3224) );
  INV_X1 U13870 ( .A(n11293), .ZN(n11296) );
  INV_X1 U13871 ( .A(n11294), .ZN(n11295) );
  NAND2_X1 U13872 ( .A1(n11296), .A2(n11295), .ZN(n11300) );
  AND2_X1 U13873 ( .A1(n11301), .A2(n11300), .ZN(n11303) );
  AOI22_X1 U13874 ( .A1(n12462), .A2(n13855), .B1(n12455), .B2(n14696), .ZN(
        n11540) );
  NAND2_X1 U13875 ( .A1(n14696), .A2(n6962), .ZN(n11298) );
  NAND2_X1 U13876 ( .A1(n12455), .A2(n13855), .ZN(n11297) );
  NAND2_X1 U13877 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  XNOR2_X1 U13878 ( .A(n11299), .B(n12450), .ZN(n11539) );
  XNOR2_X1 U13879 ( .A(n11540), .B(n11539), .ZN(n11302) );
  OAI211_X1 U13880 ( .C1(n11303), .C2(n11302), .A(n13809), .B(n11543), .ZN(
        n11310) );
  AOI21_X1 U13881 ( .B1(n13799), .B2(n13856), .A(n11304), .ZN(n11306) );
  NAND2_X1 U13882 ( .A1(n13758), .A2(n13854), .ZN(n11305) );
  OAI211_X1 U13883 ( .C1(n13832), .C2(n11307), .A(n11306), .B(n11305), .ZN(
        n11308) );
  INV_X1 U13884 ( .A(n11308), .ZN(n11309) );
  OAI211_X1 U13885 ( .C1(n11311), .C2(n13817), .A(n11310), .B(n11309), .ZN(
        P1_U3239) );
  NAND2_X1 U13886 ( .A1(n11312), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U13887 ( .A1(n11314), .A2(n11313), .ZN(n11315) );
  INV_X1 U13888 ( .A(n11315), .ZN(n11316) );
  XNOR2_X1 U13889 ( .A(n11315), .B(n11323), .ZN(n14575) );
  NOR2_X1 U13890 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14575), .ZN(n14574) );
  AOI21_X1 U13891 ( .B1(n11316), .B2(n14578), .A(n14574), .ZN(n11320) );
  INV_X1 U13892 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11317) );
  MUX2_X1 U13893 ( .A(n11317), .B(P1_REG2_REG_16__SCAN_IN), .S(n11523), .Z(
        n11318) );
  INV_X1 U13894 ( .A(n11318), .ZN(n11319) );
  NAND2_X1 U13895 ( .A1(n11319), .A2(n11320), .ZN(n11513) );
  OAI211_X1 U13896 ( .C1(n11320), .C2(n11319), .A(n14012), .B(n11513), .ZN(
        n11331) );
  NAND2_X1 U13897 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13760)
         );
  AOI21_X1 U13898 ( .B1(n9467), .B2(n11322), .A(n11321), .ZN(n11324) );
  INV_X1 U13899 ( .A(n11324), .ZN(n11325) );
  XNOR2_X1 U13900 ( .A(n11324), .B(n11323), .ZN(n14573) );
  NOR2_X1 U13901 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14573), .ZN(n14572) );
  AOI21_X1 U13902 ( .B1(n14578), .B2(n11325), .A(n14572), .ZN(n11327) );
  XOR2_X1 U13903 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11523), .Z(n11326) );
  NAND2_X1 U13904 ( .A1(n11326), .A2(n11327), .ZN(n11521) );
  OAI211_X1 U13905 ( .C1(n11327), .C2(n11326), .A(n14011), .B(n11521), .ZN(
        n11328) );
  NAND2_X1 U13906 ( .A1(n13760), .A2(n11328), .ZN(n11329) );
  AOI21_X1 U13907 ( .B1(n14568), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11329), 
        .ZN(n11330) );
  OAI211_X1 U13908 ( .C1(n14592), .C2(n11332), .A(n11331), .B(n11330), .ZN(
        P1_U3259) );
  AOI22_X1 U13909 ( .A1(n11334), .A2(n13547), .B1(n14800), .B2(n11333), .ZN(
        n11335) );
  OAI21_X1 U13910 ( .B1(n11336), .B2(n13494), .A(n11335), .ZN(n11339) );
  MUX2_X1 U13911 ( .A(n11337), .B(P2_REG2_REG_9__SCAN_IN), .S(n14809), .Z(
        n11338) );
  AOI211_X1 U13912 ( .C1(n11341), .C2(n11340), .A(n11339), .B(n11338), .ZN(
        n11342) );
  INV_X1 U13913 ( .A(n11342), .ZN(P2_U3256) );
  OAI222_X1 U13914 ( .A1(P1_U3086), .A2(n12089), .B1(n14369), .B2(n11359), 
        .C1(n15421), .C2(n14366), .ZN(P1_U3334) );
  INV_X1 U13915 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11345) );
  OR2_X1 U13916 ( .A1(n11343), .A2(n14878), .ZN(n11344) );
  OAI21_X1 U13917 ( .B1(n14880), .B2(n11345), .A(n11344), .ZN(P2_U3457) );
  XNOR2_X1 U13918 ( .A(n11346), .B(n7373), .ZN(n11352) );
  OAI211_X1 U13919 ( .C1(n11349), .C2(n11348), .A(n11347), .B(n15067), .ZN(
        n11351) );
  AOI22_X1 U13920 ( .A1(n15061), .A2(n12775), .B1(n12773), .B2(n15064), .ZN(
        n11350) );
  OAI211_X1 U13921 ( .C1(n15108), .C2(n11352), .A(n11351), .B(n11350), .ZN(
        n15126) );
  INV_X1 U13922 ( .A(n15126), .ZN(n11358) );
  INV_X1 U13923 ( .A(n11352), .ZN(n15128) );
  AOI22_X1 U13924 ( .A1(n13026), .A2(n11353), .B1(n13069), .B2(n11531), .ZN(
        n11354) );
  OAI21_X1 U13925 ( .B1(n11082), .B2(n15077), .A(n11354), .ZN(n11355) );
  AOI21_X1 U13926 ( .B1(n15128), .B2(n11356), .A(n11355), .ZN(n11357) );
  OAI21_X1 U13927 ( .B1(n11358), .B2(n13011), .A(n11357), .ZN(P3_U3223) );
  OAI222_X1 U13928 ( .A1(n12073), .A2(n11361), .B1(P2_U3088), .B2(n11360), 
        .C1(n12071), .C2(n11359), .ZN(P2_U3306) );
  INV_X1 U13929 ( .A(n11362), .ZN(n11363) );
  AOI21_X1 U13930 ( .B1(n11365), .B2(n11364), .A(n11363), .ZN(n11372) );
  INV_X1 U13931 ( .A(n11366), .ZN(n11367) );
  OAI22_X1 U13932 ( .A1(n13299), .A2(n11424), .B1(n13297), .B2(n11367), .ZN(
        n11368) );
  AOI211_X1 U13933 ( .C1(n13282), .C2(n13315), .A(n11369), .B(n11368), .ZN(
        n11371) );
  NAND2_X1 U13934 ( .A1(n11389), .A2(n13302), .ZN(n11370) );
  OAI211_X1 U13935 ( .C1(n11372), .C2(n13304), .A(n11371), .B(n11370), .ZN(
        P2_U3208) );
  XNOR2_X1 U13936 ( .A(n12159), .B(n13850), .ZN(n12313) );
  INV_X1 U13937 ( .A(n12313), .ZN(n11376) );
  XNOR2_X1 U13938 ( .A(n11373), .B(n11376), .ZN(n11375) );
  NAND2_X1 U13939 ( .A1(n14209), .A2(n13851), .ZN(n11374) );
  OAI21_X1 U13940 ( .B1(n12167), .B2(n14221), .A(n11374), .ZN(n11846) );
  AOI21_X1 U13941 ( .B1(n11375), .B2(n14611), .A(n11846), .ZN(n14536) );
  XNOR2_X1 U13942 ( .A(n11377), .B(n11376), .ZN(n14533) );
  AOI21_X1 U13943 ( .B1(n11402), .B2(n12159), .A(n14242), .ZN(n11378) );
  NAND2_X1 U13944 ( .A1(n11378), .A2(n11597), .ZN(n14532) );
  OAI22_X1 U13945 ( .A1(n14226), .A2(n11379), .B1(n11843), .B2(n14637), .ZN(
        n11380) );
  AOI21_X1 U13946 ( .B1(n14512), .B2(n12159), .A(n11380), .ZN(n11381) );
  OAI21_X1 U13947 ( .B1(n14532), .B2(n14196), .A(n11381), .ZN(n11382) );
  AOI21_X1 U13948 ( .B1(n14533), .B2(n14627), .A(n11382), .ZN(n11383) );
  OAI21_X1 U13949 ( .B1(n14536), .B2(n14642), .A(n11383), .ZN(P1_U3282) );
  INV_X1 U13950 ( .A(SI_24_), .ZN(n11386) );
  INV_X1 U13951 ( .A(n11384), .ZN(n11385) );
  OAI222_X1 U13952 ( .A1(n8294), .A2(P3_U3151), .B1(n15456), .B2(n11386), .C1(
        n15458), .C2(n11385), .ZN(P3_U3271) );
  INV_X1 U13953 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11393) );
  AOI211_X1 U13954 ( .C1(n14847), .C2(n11389), .A(n11388), .B(n11387), .ZN(
        n11390) );
  OAI21_X1 U13955 ( .B1(n14840), .B2(n11391), .A(n11390), .ZN(n11394) );
  NAND2_X1 U13956 ( .A1(n11394), .A2(n14880), .ZN(n11392) );
  OAI21_X1 U13957 ( .B1(n14880), .B2(n11393), .A(n11392), .ZN(P2_U3463) );
  NAND2_X1 U13958 ( .A1(n11394), .A2(n14891), .ZN(n11395) );
  OAI21_X1 U13959 ( .B1(n14891), .B2(n10429), .A(n11395), .ZN(P2_U3510) );
  INV_X1 U13960 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15248) );
  OAI21_X1 U13961 ( .B1(n11398), .B2(n11397), .A(n11396), .ZN(n14605) );
  INV_X1 U13962 ( .A(n14605), .ZN(n11406) );
  OAI211_X1 U13963 ( .C1(n11400), .C2(n12312), .A(n11399), .B(n14611), .ZN(
        n11401) );
  NAND2_X1 U13964 ( .A1(n14209), .A2(n13852), .ZN(n11679) );
  AND2_X1 U13965 ( .A1(n11401), .A2(n11679), .ZN(n14607) );
  OAI211_X1 U13966 ( .C1(n14603), .C2(n11403), .A(n11402), .B(n14622), .ZN(
        n11404) );
  NAND2_X1 U13967 ( .A1(n13850), .A2(n14207), .ZN(n11678) );
  NAND2_X1 U13968 ( .A1(n11404), .A2(n11678), .ZN(n14598) );
  AOI21_X1 U13969 ( .B1(n14697), .B2(n12150), .A(n14598), .ZN(n11405) );
  OAI211_X1 U13970 ( .C1(n11406), .C2(n14404), .A(n14607), .B(n11405), .ZN(
        n11408) );
  NAND2_X1 U13971 ( .A1(n11408), .A2(n14710), .ZN(n11407) );
  OAI21_X1 U13972 ( .B1(n14710), .B2(n15248), .A(n11407), .ZN(P1_U3489) );
  NAND2_X1 U13973 ( .A1(n11408), .A2(n14720), .ZN(n11409) );
  OAI21_X1 U13974 ( .B1(n14720), .B2(n11410), .A(n11409), .ZN(P1_U3538) );
  OAI21_X1 U13975 ( .B1(n11413), .B2(n11412), .A(n11411), .ZN(n11414) );
  NAND2_X1 U13976 ( .A1(n11414), .A2(n13278), .ZN(n11419) );
  NAND2_X1 U13977 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14765)
         );
  OAI21_X1 U13978 ( .B1(n13252), .B2(n11415), .A(n14765), .ZN(n11416) );
  AOI21_X1 U13979 ( .B1(n11417), .B2(n13283), .A(n11416), .ZN(n11418) );
  OAI211_X1 U13980 ( .C1(n11420), .C2(n11948), .A(n11419), .B(n11418), .ZN(
        P2_U3196) );
  OAI222_X1 U13981 ( .A1(n15458), .A2(n11423), .B1(P3_U3151), .B2(n11422), 
        .C1(n11421), .C2(n15456), .ZN(P3_U3270) );
  XNOR2_X1 U13982 ( .A(n11690), .B(n11430), .ZN(n11426) );
  AOI22_X1 U13983 ( .A1(n13311), .A2(n13538), .B1(n13313), .B2(n13540), .ZN(
        n11441) );
  OAI21_X1 U13984 ( .B1(n11426), .B2(n13520), .A(n11441), .ZN(n11507) );
  INV_X1 U13985 ( .A(n11507), .ZN(n11436) );
  NOR2_X1 U13986 ( .A1(n13667), .A2(n13313), .ZN(n11427) );
  XNOR2_X1 U13987 ( .A(n11686), .B(n11430), .ZN(n11509) );
  INV_X1 U13988 ( .A(n11692), .ZN(n11506) );
  OAI211_X1 U13989 ( .C1(n11506), .C2(n11431), .A(n11860), .B(n11721), .ZN(
        n11505) );
  AOI22_X1 U13990 ( .A1(n13469), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n14800), 
        .B2(n11439), .ZN(n11433) );
  NAND2_X1 U13991 ( .A1(n11692), .A2(n13547), .ZN(n11432) );
  OAI211_X1 U13992 ( .C1(n11505), .C2(n13494), .A(n11433), .B(n11432), .ZN(
        n11434) );
  AOI21_X1 U13993 ( .B1(n11509), .B2(n14806), .A(n11434), .ZN(n11435) );
  OAI21_X1 U13994 ( .B1(n11436), .B2(n13469), .A(n11435), .ZN(P2_U3252) );
  XNOR2_X1 U13995 ( .A(n11438), .B(n11437), .ZN(n11444) );
  NAND2_X1 U13996 ( .A1(n13283), .A2(n11439), .ZN(n11440) );
  NAND2_X1 U13997 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14773)
         );
  OAI211_X1 U13998 ( .C1(n11441), .C2(n13252), .A(n11440), .B(n14773), .ZN(
        n11442) );
  AOI21_X1 U13999 ( .B1(n11692), .B2(n13302), .A(n11442), .ZN(n11443) );
  OAI21_X1 U14000 ( .B1(n11444), .B2(n13304), .A(n11443), .ZN(P2_U3206) );
  XNOR2_X1 U14001 ( .A(n11445), .B(n12676), .ZN(n14499) );
  OAI211_X1 U14002 ( .C1(n11447), .C2(n12676), .A(n11446), .B(n15067), .ZN(
        n11450) );
  OAI22_X1 U14003 ( .A1(n11448), .A2(n15049), .B1(n11803), .B2(n15050), .ZN(
        n11633) );
  INV_X1 U14004 ( .A(n11633), .ZN(n11449) );
  NAND2_X1 U14005 ( .A1(n11450), .A2(n11449), .ZN(n14501) );
  NAND2_X1 U14006 ( .A1(n14501), .A2(n15077), .ZN(n11455) );
  INV_X1 U14007 ( .A(n11451), .ZN(n14497) );
  INV_X1 U14008 ( .A(n11636), .ZN(n11452) );
  OAI22_X1 U14009 ( .A1(n13071), .A2(n14497), .B1(n11452), .B2(n15072), .ZN(
        n11453) );
  AOI21_X1 U14010 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n15079), .A(n11453), 
        .ZN(n11454) );
  OAI211_X1 U14011 ( .C1(n14499), .C2(n13029), .A(n11455), .B(n11454), .ZN(
        P3_U3222) );
  INV_X1 U14012 ( .A(n11652), .ZN(n15454) );
  AOI21_X1 U14013 ( .B1(n7982), .B2(n11457), .A(n11640), .ZN(n11473) );
  NAND2_X1 U14014 ( .A1(n11459), .A2(n11458), .ZN(n11461) );
  MUX2_X1 U14015 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6973), .Z(n11651) );
  XNOR2_X1 U14016 ( .A(n11651), .B(n11652), .ZN(n11460) );
  OAI21_X1 U14017 ( .B1(n11461), .B2(n11460), .A(n11657), .ZN(n11471) );
  NAND2_X1 U14018 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11462), .ZN(n11464) );
  XNOR2_X1 U14019 ( .A(n11644), .B(n11652), .ZN(n11465) );
  NAND2_X1 U14020 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11465), .ZN(n11645) );
  OAI21_X1 U14021 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11465), .A(n11645), 
        .ZN(n11466) );
  NAND2_X1 U14022 ( .A1(n11466), .A2(n15023), .ZN(n11469) );
  NOR2_X1 U14023 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15291), .ZN(n11467) );
  AOI21_X1 U14024 ( .B1(n14990), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11467), 
        .ZN(n11468) );
  OAI211_X1 U14025 ( .C1(n14985), .C2(n15454), .A(n11469), .B(n11468), .ZN(
        n11470) );
  AOI21_X1 U14026 ( .B1(n15031), .B2(n11471), .A(n11470), .ZN(n11472) );
  OAI21_X1 U14027 ( .B1(n11473), .B2(n15036), .A(n11472), .ZN(P3_U3193) );
  NAND2_X1 U14028 ( .A1(n11478), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11481) );
  INV_X1 U14029 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11477) );
  NOR2_X1 U14030 ( .A1(n11487), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n14751) );
  INV_X1 U14031 ( .A(n14751), .ZN(n11475) );
  MUX2_X1 U14032 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11477), .S(n11486), .Z(
        n14752) );
  INV_X1 U14033 ( .A(n14752), .ZN(n11474) );
  AOI21_X1 U14034 ( .B1(n11476), .B2(n11475), .A(n11474), .ZN(n14754) );
  AOI21_X1 U14035 ( .B1(n14763), .B2(n11477), .A(n14754), .ZN(n14777) );
  INV_X1 U14036 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11479) );
  MUX2_X1 U14037 ( .A(n11479), .B(P2_REG2_REG_13__SCAN_IN), .S(n11478), .Z(
        n11480) );
  INV_X1 U14038 ( .A(n11480), .ZN(n14776) );
  NAND2_X1 U14039 ( .A1(n14777), .A2(n14776), .ZN(n14775) );
  NAND2_X1 U14040 ( .A1(n11481), .A2(n14775), .ZN(n11483) );
  NAND2_X1 U14041 ( .A1(n11482), .A2(n11483), .ZN(n11484) );
  XNOR2_X1 U14042 ( .A(n11483), .B(n14794), .ZN(n14791) );
  NAND2_X1 U14043 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14791), .ZN(n14789) );
  NAND2_X1 U14044 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11485), .ZN(n11609) );
  OAI211_X1 U14045 ( .C1(n11485), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14790), 
        .B(n11609), .ZN(n11496) );
  NAND2_X1 U14046 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n11757)
         );
  INV_X1 U14047 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11491) );
  XNOR2_X1 U14048 ( .A(n14794), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14783) );
  INV_X1 U14049 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11490) );
  INV_X1 U14050 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11489) );
  XNOR2_X1 U14051 ( .A(n11486), .B(n11489), .ZN(n14756) );
  NAND2_X1 U14052 ( .A1(n11487), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n14757) );
  AND2_X1 U14053 ( .A1(n14756), .A2(n14757), .ZN(n11488) );
  AOI21_X1 U14054 ( .B1(n14763), .B2(n11489), .A(n14759), .ZN(n14771) );
  XNOR2_X1 U14055 ( .A(n14780), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14770) );
  NAND2_X1 U14056 ( .A1(n14771), .A2(n14770), .ZN(n14769) );
  OAI21_X1 U14057 ( .B1(n11490), .B2(n14780), .A(n14769), .ZN(n14784) );
  NAND2_X1 U14058 ( .A1(n14783), .A2(n14784), .ZN(n14781) );
  OAI21_X1 U14059 ( .B1(n11491), .B2(n14794), .A(n14781), .ZN(n11615) );
  XNOR2_X1 U14060 ( .A(n11615), .B(n11497), .ZN(n11492) );
  NAND2_X1 U14061 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n11492), .ZN(n11617) );
  OAI211_X1 U14062 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n11492), .A(n14782), 
        .B(n11617), .ZN(n11493) );
  NAND2_X1 U14063 ( .A1(n11757), .A2(n11493), .ZN(n11494) );
  AOI21_X1 U14064 ( .B1(n14788), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n11494), 
        .ZN(n11495) );
  OAI211_X1 U14065 ( .C1(n14795), .C2(n11497), .A(n11496), .B(n11495), .ZN(
        P2_U3229) );
  INV_X1 U14066 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15268) );
  OAI211_X1 U14067 ( .C1(n11500), .C2(n14702), .A(n11499), .B(n11498), .ZN(
        n11502) );
  NAND2_X1 U14068 ( .A1(n11502), .A2(n14710), .ZN(n11501) );
  OAI21_X1 U14069 ( .B1(n14710), .B2(n15268), .A(n11501), .ZN(P1_U3486) );
  NAND2_X1 U14070 ( .A1(n11502), .A2(n14720), .ZN(n11503) );
  OAI21_X1 U14071 ( .B1(n14720), .B2(n11504), .A(n11503), .ZN(P1_U3537) );
  INV_X1 U14072 ( .A(n14840), .ZN(n13618) );
  OAI21_X1 U14073 ( .B1(n11506), .B2(n14872), .A(n11505), .ZN(n11508) );
  AOI211_X1 U14074 ( .C1(n11509), .C2(n13618), .A(n11508), .B(n11507), .ZN(
        n11512) );
  NAND2_X1 U14075 ( .A1(n14888), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11510) );
  OAI21_X1 U14076 ( .B1(n11512), .B2(n14888), .A(n11510), .ZN(P2_U3512) );
  NAND2_X1 U14077 ( .A1(n14878), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11511) );
  OAI21_X1 U14078 ( .B1(n11512), .B2(n14878), .A(n11511), .ZN(P2_U3469) );
  NAND2_X1 U14079 ( .A1(n11523), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11514) );
  NAND2_X1 U14080 ( .A1(n11514), .A2(n11513), .ZN(n11520) );
  INV_X1 U14081 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U14082 ( .A1(n14001), .A2(n11515), .ZN(n11518) );
  INV_X1 U14083 ( .A(n11518), .ZN(n11516) );
  AOI21_X1 U14084 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n11517), .A(n11516), 
        .ZN(n11519) );
  NAND2_X1 U14085 ( .A1(n11517), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13995) );
  NAND3_X1 U14086 ( .A1(n11520), .A2(n13995), .A3(n11518), .ZN(n13994) );
  OAI211_X1 U14087 ( .C1(n11520), .C2(n11519), .A(n13994), .B(n14012), .ZN(
        n11528) );
  NAND2_X1 U14088 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13772)
         );
  INV_X1 U14089 ( .A(n11521), .ZN(n11522) );
  AOI21_X1 U14090 ( .B1(n11523), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11522), 
        .ZN(n14002) );
  XNOR2_X1 U14091 ( .A(n14001), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13999) );
  XNOR2_X1 U14092 ( .A(n14002), .B(n13999), .ZN(n11524) );
  NAND2_X1 U14093 ( .A1(n14011), .A2(n11524), .ZN(n11525) );
  NAND2_X1 U14094 ( .A1(n13772), .A2(n11525), .ZN(n11526) );
  AOI21_X1 U14095 ( .B1(n14568), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11526), 
        .ZN(n11527) );
  OAI211_X1 U14096 ( .C1(n14592), .C2(n14001), .A(n11528), .B(n11527), .ZN(
        P1_U3260) );
  AOI211_X1 U14097 ( .C1(n11530), .C2(n11529), .A(n14427), .B(n6734), .ZN(
        n11538) );
  INV_X1 U14098 ( .A(n11531), .ZN(n11536) );
  AOI22_X1 U14099 ( .A1(n12479), .A2(n12775), .B1(n14416), .B2(n12773), .ZN(
        n11535) );
  OAI21_X1 U14100 ( .B1(n12574), .B2(n15125), .A(n11532), .ZN(n11533) );
  INV_X1 U14101 ( .A(n11533), .ZN(n11534) );
  OAI211_X1 U14102 ( .C1(n11536), .C2(n14433), .A(n11535), .B(n11534), .ZN(
        n11537) );
  OR2_X1 U14103 ( .A1(n11538), .A2(n11537), .ZN(P3_U3157) );
  INV_X1 U14104 ( .A(n11540), .ZN(n11541) );
  NAND2_X1 U14105 ( .A1(n11539), .A2(n11541), .ZN(n11542) );
  NAND2_X1 U14106 ( .A1(n12129), .A2(n6962), .ZN(n11545) );
  NAND2_X1 U14107 ( .A1(n12455), .A2(n13854), .ZN(n11544) );
  NAND2_X1 U14108 ( .A1(n11545), .A2(n11544), .ZN(n11546) );
  XNOR2_X1 U14109 ( .A(n11546), .B(n12450), .ZN(n11547) );
  AOI22_X1 U14110 ( .A1(n12462), .A2(n13854), .B1(n12129), .B2(n12455), .ZN(
        n11548) );
  XNOR2_X1 U14111 ( .A(n11547), .B(n11548), .ZN(n11573) );
  NOR2_X1 U14112 ( .A1(n11549), .A2(n11548), .ZN(n11550) );
  AOI22_X1 U14113 ( .A1(n12132), .A2(n12455), .B1(n12462), .B2(n13853), .ZN(
        n11557) );
  AOI22_X1 U14114 ( .A1(n12132), .A2(n6962), .B1(n12455), .B2(n13853), .ZN(
        n11551) );
  XNOR2_X1 U14115 ( .A(n11551), .B(n12450), .ZN(n11558) );
  XOR2_X1 U14116 ( .A(n11557), .B(n11558), .Z(n11580) );
  NAND2_X1 U14117 ( .A1(n12141), .A2(n6962), .ZN(n11553) );
  NAND2_X1 U14118 ( .A1(n12455), .A2(n13852), .ZN(n11552) );
  NAND2_X1 U14119 ( .A1(n11553), .A2(n11552), .ZN(n11554) );
  XNOR2_X1 U14120 ( .A(n11554), .B(n12450), .ZN(n11672) );
  NOR2_X1 U14121 ( .A1(n12394), .A2(n11555), .ZN(n11556) );
  AOI21_X1 U14122 ( .B1(n12141), .B2(n12455), .A(n11556), .ZN(n11674) );
  XNOR2_X1 U14123 ( .A(n11672), .B(n11674), .ZN(n11560) );
  NAND2_X1 U14124 ( .A1(n11558), .A2(n11557), .ZN(n11561) );
  NAND2_X1 U14125 ( .A1(n11673), .A2(n13809), .ZN(n11569) );
  AOI21_X1 U14126 ( .B1(n11559), .B2(n11561), .A(n11560), .ZN(n11568) );
  NAND2_X1 U14127 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n13966) );
  INV_X1 U14128 ( .A(n13966), .ZN(n11562) );
  AOI21_X1 U14129 ( .B1(n13799), .B2(n13853), .A(n11562), .ZN(n11564) );
  NAND2_X1 U14130 ( .A1(n13758), .A2(n13851), .ZN(n11563) );
  OAI211_X1 U14131 ( .C1(n13832), .C2(n11565), .A(n11564), .B(n11563), .ZN(
        n11566) );
  AOI21_X1 U14132 ( .B1(n13834), .B2(n12141), .A(n11566), .ZN(n11567) );
  OAI21_X1 U14133 ( .B1(n11569), .B2(n11568), .A(n11567), .ZN(P1_U3231) );
  AND2_X1 U14134 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13942) );
  AOI21_X1 U14135 ( .B1(n13799), .B2(n13855), .A(n13942), .ZN(n11571) );
  NAND2_X1 U14136 ( .A1(n13758), .A2(n13853), .ZN(n11570) );
  OAI211_X1 U14137 ( .C1(n13832), .C2(n11572), .A(n11571), .B(n11570), .ZN(
        n11577) );
  XNOR2_X1 U14138 ( .A(n11574), .B(n11573), .ZN(n11575) );
  NOR2_X1 U14139 ( .A1(n11575), .A2(n13836), .ZN(n11576) );
  AOI211_X1 U14140 ( .C1(n13834), .C2(n12129), .A(n11577), .B(n11576), .ZN(
        n11578) );
  INV_X1 U14141 ( .A(n11578), .ZN(P1_U3213) );
  OAI21_X1 U14142 ( .B1(n11580), .B2(n11579), .A(n11559), .ZN(n11581) );
  NAND2_X1 U14143 ( .A1(n11581), .A2(n13809), .ZN(n11586) );
  OAI21_X1 U14144 ( .B1(n13811), .B2(n14700), .A(n11582), .ZN(n11583) );
  AOI21_X1 U14145 ( .B1(n13814), .B2(n11584), .A(n11583), .ZN(n11585) );
  OAI211_X1 U14146 ( .C1(n14703), .C2(n13817), .A(n11586), .B(n11585), .ZN(
        P1_U3221) );
  XNOR2_X1 U14147 ( .A(n11588), .B(n12604), .ZN(n14493) );
  XNOR2_X1 U14148 ( .A(n11589), .B(n12604), .ZN(n11590) );
  AOI22_X1 U14149 ( .A1(n15061), .A2(n12773), .B1(n12771), .B2(n15064), .ZN(
        n11734) );
  OAI21_X1 U14150 ( .B1(n11590), .B2(n13063), .A(n11734), .ZN(n14495) );
  NAND2_X1 U14151 ( .A1(n14495), .A2(n15077), .ZN(n11595) );
  INV_X1 U14152 ( .A(n14492), .ZN(n11736) );
  INV_X1 U14153 ( .A(n11591), .ZN(n11739) );
  OAI22_X1 U14154 ( .A1(n15077), .A2(n11592), .B1(n11739), .B2(n15072), .ZN(
        n11593) );
  AOI21_X1 U14155 ( .B1(n11736), .B2(n13026), .A(n11593), .ZN(n11594) );
  OAI211_X1 U14156 ( .C1(n13029), .C2(n14493), .A(n11595), .B(n11594), .ZN(
        P3_U3221) );
  XNOR2_X1 U14157 ( .A(n11596), .B(n12315), .ZN(n14405) );
  NAND2_X1 U14158 ( .A1(n11597), .A2(n14401), .ZN(n11598) );
  NAND2_X1 U14159 ( .A1(n11598), .A2(n14622), .ZN(n11599) );
  OR2_X1 U14160 ( .A1(n6729), .A2(n11599), .ZN(n14403) );
  XNOR2_X1 U14161 ( .A(n11601), .B(n11600), .ZN(n11603) );
  NAND2_X1 U14162 ( .A1(n13850), .A2(n14209), .ZN(n11602) );
  OAI21_X1 U14163 ( .B1(n12166), .B2(n14221), .A(n11602), .ZN(n11827) );
  AOI21_X1 U14164 ( .B1(n11603), .B2(n14611), .A(n11827), .ZN(n14408) );
  OAI21_X1 U14165 ( .B1(n14143), .B2(n14403), .A(n14408), .ZN(n11604) );
  NAND2_X1 U14166 ( .A1(n11604), .A2(n14226), .ZN(n11607) );
  OAI22_X1 U14167 ( .A1(n14226), .A2(n10298), .B1(n11829), .B2(n14637), .ZN(
        n11605) );
  AOI21_X1 U14168 ( .B1(n14512), .B2(n14401), .A(n11605), .ZN(n11606) );
  OAI211_X1 U14169 ( .C1(n14249), .C2(n14405), .A(n11607), .B(n11606), .ZN(
        P1_U3281) );
  NAND2_X1 U14170 ( .A1(n11616), .A2(n11608), .ZN(n11610) );
  NAND2_X1 U14171 ( .A1(n11610), .A2(n11609), .ZN(n11614) );
  NAND2_X1 U14172 ( .A1(n11611), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11872) );
  INV_X1 U14173 ( .A(n11872), .ZN(n11612) );
  AOI21_X1 U14174 ( .B1(n8740), .B2(n11868), .A(n11612), .ZN(n11613) );
  NAND2_X1 U14175 ( .A1(n11613), .A2(n11614), .ZN(n11871) );
  OAI211_X1 U14176 ( .C1(n11614), .C2(n11613), .A(n14790), .B(n11871), .ZN(
        n11624) );
  NAND2_X1 U14177 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11942)
         );
  NAND2_X1 U14178 ( .A1(n11616), .A2(n11615), .ZN(n11618) );
  NAND2_X1 U14179 ( .A1(n11618), .A2(n11617), .ZN(n11620) );
  XNOR2_X1 U14180 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n11868), .ZN(n11619) );
  NAND2_X1 U14181 ( .A1(n11619), .A2(n11620), .ZN(n11866) );
  OAI211_X1 U14182 ( .C1(n11620), .C2(n11619), .A(n14782), .B(n11866), .ZN(
        n11621) );
  NAND2_X1 U14183 ( .A1(n11942), .A2(n11621), .ZN(n11622) );
  AOI21_X1 U14184 ( .B1(n14788), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11622), 
        .ZN(n11623) );
  OAI211_X1 U14185 ( .C1(n14795), .C2(n11868), .A(n11624), .B(n11623), .ZN(
        P2_U3230) );
  INV_X1 U14186 ( .A(n11625), .ZN(n11627) );
  OAI222_X1 U14187 ( .A1(P3_U3151), .A2(n11628), .B1(n15458), .B2(n11627), 
        .C1(n11626), .C2(n15456), .ZN(P3_U3269) );
  NAND2_X1 U14188 ( .A1(n11630), .A2(n11629), .ZN(n11632) );
  XNOR2_X1 U14189 ( .A(n11632), .B(n11631), .ZN(n11638) );
  AOI22_X1 U14190 ( .A1(n12510), .A2(n11633), .B1(P3_REG3_REG_11__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11634) );
  OAI21_X1 U14191 ( .B1(n14497), .B2(n12574), .A(n11634), .ZN(n11635) );
  AOI21_X1 U14192 ( .B1(n14444), .B2(n11636), .A(n11635), .ZN(n11637) );
  OAI21_X1 U14193 ( .B1(n11638), .B2(n14427), .A(n11637), .ZN(P3_U3176) );
  NOR2_X1 U14194 ( .A1(n11652), .A2(n11639), .ZN(n11641) );
  INV_X1 U14195 ( .A(n14390), .ZN(n11908) );
  AOI22_X1 U14196 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11908), .B1(n14390), 
        .B2(n11592), .ZN(n11642) );
  AOI21_X1 U14197 ( .B1(n11643), .B2(n11642), .A(n11905), .ZN(n11664) );
  INV_X1 U14198 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U14199 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n14390), .B1(n11908), 
        .B2(n14496), .ZN(n11648) );
  NAND2_X1 U14200 ( .A1(n15454), .A2(n11644), .ZN(n11646) );
  NAND2_X1 U14201 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  NAND2_X1 U14202 ( .A1(n11648), .A2(n11647), .ZN(n11907) );
  OAI21_X1 U14203 ( .B1(n11648), .B2(n11647), .A(n11907), .ZN(n11662) );
  NOR2_X1 U14204 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11733), .ZN(n11649) );
  AOI21_X1 U14205 ( .B1(n14990), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11649), 
        .ZN(n11650) );
  OAI21_X1 U14206 ( .B1(n14985), .B2(n14390), .A(n11650), .ZN(n11661) );
  MUX2_X1 U14207 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6973), .Z(n11910) );
  XNOR2_X1 U14208 ( .A(n11910), .B(n11908), .ZN(n11655) );
  INV_X1 U14209 ( .A(n11651), .ZN(n11653) );
  NAND2_X1 U14210 ( .A1(n11653), .A2(n11652), .ZN(n11656) );
  AND2_X1 U14211 ( .A1(n11655), .A2(n11656), .ZN(n11654) );
  NAND2_X1 U14212 ( .A1(n11657), .A2(n11654), .ZN(n11914) );
  INV_X1 U14213 ( .A(n11914), .ZN(n11659) );
  AOI21_X1 U14214 ( .B1(n11657), .B2(n11656), .A(n11655), .ZN(n11658) );
  NOR3_X1 U14215 ( .A1(n11659), .A2(n11658), .A3(n15010), .ZN(n11660) );
  AOI211_X1 U14216 ( .C1(n15023), .C2(n11662), .A(n11661), .B(n11660), .ZN(
        n11663) );
  OAI21_X1 U14217 ( .B1(n11664), .B2(n15036), .A(n11663), .ZN(P3_U3194) );
  NAND2_X1 U14218 ( .A1(n11669), .A2(n11665), .ZN(n11666) );
  OAI211_X1 U14219 ( .C1(n11667), .C2(n14366), .A(n11666), .B(n12349), .ZN(
        P1_U3332) );
  NAND2_X1 U14220 ( .A1(n11669), .A2(n11668), .ZN(n11671) );
  OAI211_X1 U14221 ( .C1(n15238), .C2(n12073), .A(n11671), .B(n11670), .ZN(
        P2_U3304) );
  NAND2_X1 U14222 ( .A1(n12150), .A2(n6962), .ZN(n11676) );
  NAND2_X1 U14223 ( .A1(n12455), .A2(n13851), .ZN(n11675) );
  NAND2_X1 U14224 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  XNOR2_X1 U14225 ( .A(n11677), .B(n12450), .ZN(n11811) );
  AOI22_X1 U14226 ( .A1(n12150), .A2(n12455), .B1(n12462), .B2(n13851), .ZN(
        n11809) );
  XNOR2_X1 U14227 ( .A(n11811), .B(n11809), .ZN(n11812) );
  XNOR2_X1 U14228 ( .A(n11813), .B(n11812), .ZN(n11684) );
  AOI21_X1 U14229 ( .B1(n11679), .B2(n11678), .A(n13811), .ZN(n11680) );
  AOI211_X1 U14230 ( .C1(n13814), .C2(n14600), .A(n11681), .B(n11680), .ZN(
        n11683) );
  NAND2_X1 U14231 ( .A1(n12150), .A2(n13834), .ZN(n11682) );
  OAI211_X1 U14232 ( .C1(n11684), .C2(n13836), .A(n11683), .B(n11682), .ZN(
        P1_U3217) );
  OR2_X1 U14233 ( .A1(n11692), .A2(n13312), .ZN(n11685) );
  NAND2_X1 U14234 ( .A1(n11692), .A2(n13312), .ZN(n11687) );
  NAND2_X1 U14235 ( .A1(n13661), .A2(n13311), .ZN(n11688) );
  XOR2_X1 U14236 ( .A(n11855), .B(n11854), .Z(n13659) );
  NOR2_X1 U14237 ( .A1(n11692), .A2(n11691), .ZN(n11689) );
  NAND2_X1 U14238 ( .A1(n11692), .A2(n11691), .ZN(n11693) );
  NAND2_X1 U14239 ( .A1(n11694), .A2(n11693), .ZN(n11718) );
  AND2_X1 U14240 ( .A1(n13661), .A2(n11758), .ZN(n11695) );
  OR2_X1 U14241 ( .A1(n13661), .A2(n11758), .ZN(n11696) );
  XOR2_X1 U14242 ( .A(n11854), .B(n11849), .Z(n11697) );
  NAND2_X1 U14243 ( .A1(n11697), .A2(n13569), .ZN(n13657) );
  INV_X1 U14244 ( .A(n13657), .ZN(n11700) );
  NAND2_X1 U14245 ( .A1(n13309), .A2(n13538), .ZN(n11699) );
  NAND2_X1 U14246 ( .A1(n13311), .A2(n13540), .ZN(n11698) );
  NAND2_X1 U14247 ( .A1(n11699), .A2(n11698), .ZN(n13655) );
  OAI21_X1 U14248 ( .B1(n11700), .B2(n13655), .A(n13562), .ZN(n11704) );
  INV_X1 U14249 ( .A(n11859), .ZN(n11861) );
  AOI211_X1 U14250 ( .C1(n13656), .C2(n11720), .A(n8811), .B(n11861), .ZN(
        n13654) );
  NOR2_X1 U14251 ( .A1(n7125), .A2(n14803), .ZN(n11702) );
  INV_X1 U14252 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15235) );
  OAI22_X1 U14253 ( .A1(n13562), .A2(n15235), .B1(n11759), .B2(n13571), .ZN(
        n11701) );
  AOI211_X1 U14254 ( .C1(n13654), .C2(n14797), .A(n11702), .B(n11701), .ZN(
        n11703) );
  OAI211_X1 U14255 ( .C1(n13659), .C2(n13576), .A(n11704), .B(n11703), .ZN(
        P2_U3250) );
  OAI21_X1 U14256 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(n11708) );
  NAND2_X1 U14257 ( .A1(n11708), .A2(n13278), .ZN(n11712) );
  NAND2_X1 U14258 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14786)
         );
  INV_X1 U14259 ( .A(n14786), .ZN(n11710) );
  INV_X1 U14260 ( .A(n13310), .ZN(n11850) );
  OAI22_X1 U14261 ( .A1(n13299), .A2(n11850), .B1(n11722), .B2(n13297), .ZN(
        n11709) );
  AOI211_X1 U14262 ( .C1(n13282), .C2(n13312), .A(n11710), .B(n11709), .ZN(
        n11711) );
  OAI211_X1 U14263 ( .C1(n7127), .C2(n11948), .A(n11712), .B(n11711), .ZN(
        P2_U3187) );
  INV_X1 U14264 ( .A(n11713), .ZN(n11714) );
  INV_X1 U14265 ( .A(SI_27_), .ZN(n15348) );
  OAI222_X1 U14266 ( .A1(n6973), .A2(P3_U3151), .B1(n15458), .B2(n11714), .C1(
        n15348), .C2(n15456), .ZN(P3_U3268) );
  INV_X1 U14267 ( .A(n11715), .ZN(n11741) );
  AOI22_X1 U14268 ( .A1(n11716), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n14360), .ZN(n11717) );
  OAI21_X1 U14269 ( .B1(n11741), .B2(n14369), .A(n11717), .ZN(P1_U3331) );
  XOR2_X1 U14270 ( .A(n11725), .B(n11718), .Z(n11719) );
  AOI222_X1 U14271 ( .A1(n13569), .A2(n11719), .B1(n13312), .B2(n13540), .C1(
        n13310), .C2(n13538), .ZN(n13663) );
  AOI211_X1 U14272 ( .C1(n13661), .C2(n11721), .A(n6569), .B(n7126), .ZN(
        n13660) );
  INV_X1 U14273 ( .A(n11722), .ZN(n11723) );
  AOI22_X1 U14274 ( .A1(n13469), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14800), 
        .B2(n11723), .ZN(n11724) );
  OAI21_X1 U14275 ( .B1(n7127), .B2(n14803), .A(n11724), .ZN(n11728) );
  XNOR2_X1 U14276 ( .A(n11726), .B(n11725), .ZN(n13664) );
  NOR2_X1 U14277 ( .A1(n13664), .A2(n13576), .ZN(n11727) );
  AOI211_X1 U14278 ( .C1(n13660), .C2(n14797), .A(n11728), .B(n11727), .ZN(
        n11729) );
  OAI21_X1 U14279 ( .B1(n13663), .B2(n13469), .A(n11729), .ZN(P2_U3251) );
  NAND2_X1 U14280 ( .A1(n11730), .A2(n11731), .ZN(n11765) );
  OAI21_X1 U14281 ( .B1(n11731), .B2(n11730), .A(n11765), .ZN(n11732) );
  NAND2_X1 U14282 ( .A1(n11732), .A2(n14439), .ZN(n11738) );
  OAI22_X1 U14283 ( .A1(n14446), .A2(n11734), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11733), .ZN(n11735) );
  AOI21_X1 U14284 ( .B1(n11736), .B2(n14441), .A(n11735), .ZN(n11737) );
  OAI211_X1 U14285 ( .C1(n11739), .C2(n14433), .A(n11738), .B(n11737), .ZN(
        P3_U3164) );
  OAI222_X1 U14286 ( .A1(n11742), .A2(P2_U3088), .B1(n12071), .B2(n11741), 
        .C1(n11740), .C2(n12073), .ZN(P2_U3303) );
  INV_X1 U14287 ( .A(n11778), .ZN(n11743) );
  AOI21_X1 U14288 ( .B1(n11744), .B2(n12592), .A(n11743), .ZN(n14483) );
  NAND2_X1 U14289 ( .A1(n11745), .A2(n15067), .ZN(n11749) );
  AOI21_X1 U14290 ( .B1(n11800), .B2(n11746), .A(n12592), .ZN(n11748) );
  AOI22_X1 U14291 ( .A1(n15061), .A2(n12771), .B1(n14415), .B2(n15064), .ZN(
        n11747) );
  OAI21_X1 U14292 ( .B1(n11749), .B2(n11748), .A(n11747), .ZN(n14485) );
  NAND2_X1 U14293 ( .A1(n14485), .A2(n15077), .ZN(n11753) );
  OAI22_X1 U14294 ( .A1(n15077), .A2(n11750), .B1(n14434), .B2(n15072), .ZN(
        n11751) );
  AOI21_X1 U14295 ( .B1(n13026), .B2(n14481), .A(n11751), .ZN(n11752) );
  OAI211_X1 U14296 ( .C1(n14483), .C2(n13029), .A(n11753), .B(n11752), .ZN(
        P3_U3219) );
  XNOR2_X1 U14297 ( .A(n11755), .B(n11754), .ZN(n11756) );
  XNOR2_X1 U14298 ( .A(n6709), .B(n11756), .ZN(n11763) );
  OAI21_X1 U14299 ( .B1(n13295), .B2(n11758), .A(n11757), .ZN(n11761) );
  OAI22_X1 U14300 ( .A1(n13299), .A2(n11883), .B1(n13297), .B2(n11759), .ZN(
        n11760) );
  AOI211_X1 U14301 ( .C1(n13656), .C2(n13302), .A(n11761), .B(n11760), .ZN(
        n11762) );
  OAI21_X1 U14302 ( .B1(n11763), .B2(n13304), .A(n11762), .ZN(P2_U3213) );
  NAND2_X1 U14303 ( .A1(n11765), .A2(n11764), .ZN(n14421) );
  XNOR2_X1 U14304 ( .A(n11766), .B(n12771), .ZN(n11767) );
  XNOR2_X1 U14305 ( .A(n14421), .B(n11767), .ZN(n11772) );
  AND2_X1 U14306 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11917) );
  AOI21_X1 U14307 ( .B1(n14416), .B2(n12770), .A(n11917), .ZN(n11769) );
  NAND2_X1 U14308 ( .A1(n12479), .A2(n12772), .ZN(n11768) );
  OAI211_X1 U14309 ( .C1(n14433), .C2(n11804), .A(n11769), .B(n11768), .ZN(
        n11770) );
  AOI21_X1 U14310 ( .B1(n14490), .B2(n14441), .A(n11770), .ZN(n11771) );
  OAI21_X1 U14311 ( .B1(n11772), .B2(n14427), .A(n11771), .ZN(P3_U3174) );
  XNOR2_X1 U14312 ( .A(n11773), .B(n12698), .ZN(n11774) );
  NAND2_X1 U14313 ( .A1(n11774), .A2(n15067), .ZN(n11776) );
  AOI22_X1 U14314 ( .A1(n15061), .A2(n12770), .B1(n12769), .B2(n15064), .ZN(
        n11775) );
  NAND2_X1 U14315 ( .A1(n11776), .A2(n11775), .ZN(n13142) );
  INV_X1 U14316 ( .A(n13142), .ZN(n11784) );
  NAND3_X1 U14317 ( .A1(n11778), .A2(n12694), .A3(n11777), .ZN(n11779) );
  NAND2_X1 U14318 ( .A1(n11780), .A2(n11779), .ZN(n13139) );
  INV_X1 U14319 ( .A(n13137), .ZN(n12084) );
  AOI22_X1 U14320 ( .A1(n15079), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13069), 
        .B2(n12081), .ZN(n11781) );
  OAI21_X1 U14321 ( .B1(n12084), .B2(n13071), .A(n11781), .ZN(n11782) );
  AOI21_X1 U14322 ( .B1(n13139), .B2(n13073), .A(n11782), .ZN(n11783) );
  OAI21_X1 U14323 ( .B1(n11784), .B2(n15079), .A(n11783), .ZN(P3_U3218) );
  NAND2_X1 U14324 ( .A1(n11785), .A2(n14707), .ZN(n11788) );
  NAND2_X1 U14325 ( .A1(n11789), .A2(n14611), .ZN(n11787) );
  NAND2_X1 U14326 ( .A1(n11788), .A2(n11787), .ZN(n11792) );
  OAI22_X1 U14327 ( .A1(n14404), .A2(n11785), .B1(n11789), .B2(n14234), .ZN(
        n11791) );
  MUX2_X1 U14328 ( .A(n11792), .B(n11791), .S(n11790), .Z(n11795) );
  NAND2_X1 U14329 ( .A1(n14209), .A2(n13849), .ZN(n11793) );
  OAI21_X1 U14330 ( .B1(n13829), .B2(n14221), .A(n11793), .ZN(n11794) );
  OR2_X1 U14331 ( .A1(n11795), .A2(n11794), .ZN(n11836) );
  OAI211_X1 U14332 ( .C1(n6729), .C2(n12170), .A(n14518), .B(n14622), .ZN(
        n11834) );
  OAI22_X1 U14333 ( .A1(n11834), .A2(n14143), .B1(n14637), .B2(n11961), .ZN(
        n11796) );
  OAI21_X1 U14334 ( .B1(n11836), .B2(n11796), .A(n14226), .ZN(n11798) );
  NAND2_X1 U14335 ( .A1(n12171), .A2(n14512), .ZN(n11797) );
  OAI211_X1 U14336 ( .C1(n10452), .C2(n14226), .A(n11798), .B(n11797), .ZN(
        P1_U3280) );
  XNOR2_X1 U14337 ( .A(n11799), .B(n8019), .ZN(n14487) );
  AOI21_X1 U14338 ( .B1(n12685), .B2(n11801), .A(n7036), .ZN(n11802) );
  OAI222_X1 U14339 ( .A1(n15050), .A2(n12079), .B1(n15049), .B2(n11803), .C1(
        n13063), .C2(n11802), .ZN(n14488) );
  NAND2_X1 U14340 ( .A1(n14488), .A2(n15077), .ZN(n11808) );
  OAI22_X1 U14341 ( .A1(n15077), .A2(n11805), .B1(n11804), .B2(n15072), .ZN(
        n11806) );
  AOI21_X1 U14342 ( .B1(n14490), .B2(n13026), .A(n11806), .ZN(n11807) );
  OAI211_X1 U14343 ( .C1(n13029), .C2(n14487), .A(n11808), .B(n11807), .ZN(
        P3_U3220) );
  INV_X1 U14344 ( .A(n11809), .ZN(n11810) );
  OAI22_X1 U14345 ( .A1(n14530), .A2(n12395), .B1(n12158), .B2(n12394), .ZN(
        n11820) );
  OAI22_X1 U14346 ( .A1(n14530), .A2(n12396), .B1(n12158), .B2(n12395), .ZN(
        n11814) );
  XNOR2_X1 U14347 ( .A(n11814), .B(n12450), .ZN(n11819) );
  XOR2_X1 U14348 ( .A(n11820), .B(n11819), .Z(n11841) );
  NAND2_X1 U14349 ( .A1(n14401), .A2(n6962), .ZN(n11816) );
  NAND2_X1 U14350 ( .A1(n12455), .A2(n13849), .ZN(n11815) );
  NAND2_X1 U14351 ( .A1(n11816), .A2(n11815), .ZN(n11817) );
  XNOR2_X1 U14352 ( .A(n11817), .B(n12450), .ZN(n11950) );
  NOR2_X1 U14353 ( .A1(n12394), .A2(n12167), .ZN(n11818) );
  AOI21_X1 U14354 ( .B1(n14401), .B2(n12455), .A(n11818), .ZN(n11951) );
  XNOR2_X1 U14355 ( .A(n11950), .B(n11951), .ZN(n11825) );
  INV_X1 U14356 ( .A(n11819), .ZN(n11822) );
  INV_X1 U14357 ( .A(n11820), .ZN(n11821) );
  NAND2_X1 U14358 ( .A1(n11822), .A2(n11821), .ZN(n11826) );
  NAND2_X1 U14359 ( .A1(n11954), .A2(n13809), .ZN(n11833) );
  AOI21_X1 U14360 ( .B1(n11824), .B2(n11826), .A(n11825), .ZN(n11832) );
  AOI22_X1 U14361 ( .A1(n13830), .A2(n11827), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11828) );
  OAI21_X1 U14362 ( .B1(n13832), .B2(n11829), .A(n11828), .ZN(n11830) );
  AOI21_X1 U14363 ( .B1(n14401), .B2(n13834), .A(n11830), .ZN(n11831) );
  OAI21_X1 U14364 ( .B1(n11833), .B2(n11832), .A(n11831), .ZN(P1_U3224) );
  OAI21_X1 U14365 ( .B1(n12170), .B2(n14702), .A(n11834), .ZN(n11835) );
  NOR2_X1 U14366 ( .A1(n11836), .A2(n11835), .ZN(n11838) );
  MUX2_X1 U14367 ( .A(n10457), .B(n11838), .S(n14720), .Z(n11837) );
  INV_X1 U14368 ( .A(n11837), .ZN(P1_U3541) );
  INV_X1 U14369 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15228) );
  MUX2_X1 U14370 ( .A(n15228), .B(n11838), .S(n14710), .Z(n11839) );
  INV_X1 U14371 ( .A(n11839), .ZN(P1_U3498) );
  OAI21_X1 U14372 ( .B1(n11841), .B2(n11840), .A(n11824), .ZN(n11842) );
  NAND2_X1 U14373 ( .A1(n11842), .A2(n13809), .ZN(n11848) );
  NAND2_X1 U14374 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n13982)
         );
  INV_X1 U14375 ( .A(n13982), .ZN(n11845) );
  NOR2_X1 U14376 ( .A1(n13832), .A2(n11843), .ZN(n11844) );
  AOI211_X1 U14377 ( .C1(n13830), .C2(n11846), .A(n11845), .B(n11844), .ZN(
        n11847) );
  OAI211_X1 U14378 ( .C1(n14530), .C2(n13817), .A(n11848), .B(n11847), .ZN(
        P1_U3236) );
  AOI22_X1 U14379 ( .A1(n13308), .A2(n13538), .B1(n13540), .B2(n13310), .ZN(
        n11943) );
  INV_X1 U14380 ( .A(n11943), .ZN(n11853) );
  XNOR2_X1 U14381 ( .A(n11887), .B(n7361), .ZN(n11852) );
  NOR2_X1 U14382 ( .A1(n11852), .A2(n13520), .ZN(n11899) );
  AOI211_X1 U14383 ( .C1(n14800), .C2(n11945), .A(n11853), .B(n11899), .ZN(
        n11865) );
  OR2_X1 U14384 ( .A1(n13656), .A2(n13310), .ZN(n11856) );
  INV_X1 U14385 ( .A(n11882), .ZN(n11857) );
  AOI21_X1 U14386 ( .B1(n7361), .B2(n11858), .A(n11857), .ZN(n11901) );
  INV_X1 U14387 ( .A(n11884), .ZN(n11949) );
  OAI211_X1 U14388 ( .C1(n11949), .C2(n11861), .A(n11889), .B(n11860), .ZN(
        n11898) );
  AOI22_X1 U14389 ( .A1(n11884), .A2(n13547), .B1(n14809), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n11862) );
  OAI21_X1 U14390 ( .B1(n11898), .B2(n13494), .A(n11862), .ZN(n11863) );
  AOI21_X1 U14391 ( .B1(n11901), .B2(n14806), .A(n11863), .ZN(n11864) );
  OAI21_X1 U14392 ( .B1(n11865), .B2(n13469), .A(n11864), .ZN(P2_U3249) );
  XNOR2_X1 U14393 ( .A(n13353), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11870) );
  INV_X1 U14394 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11867) );
  OAI21_X1 U14395 ( .B1(n11868), .B2(n11867), .A(n11866), .ZN(n11869) );
  NAND2_X1 U14396 ( .A1(n11870), .A2(n11869), .ZN(n13352) );
  OAI211_X1 U14397 ( .C1(n11870), .C2(n11869), .A(n14782), .B(n13352), .ZN(
        n11880) );
  NAND2_X1 U14398 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13250)
         );
  NAND2_X1 U14399 ( .A1(n11872), .A2(n11871), .ZN(n11876) );
  INV_X1 U14400 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11873) );
  MUX2_X1 U14401 ( .A(n11873), .B(P2_REG2_REG_17__SCAN_IN), .S(n13344), .Z(
        n11874) );
  INV_X1 U14402 ( .A(n11874), .ZN(n11875) );
  NAND2_X1 U14403 ( .A1(n11875), .A2(n11876), .ZN(n13345) );
  OAI211_X1 U14404 ( .C1(n11876), .C2(n11875), .A(n14790), .B(n13345), .ZN(
        n11877) );
  NAND2_X1 U14405 ( .A1(n13250), .A2(n11877), .ZN(n11878) );
  AOI21_X1 U14406 ( .B1(n14788), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n11878), 
        .ZN(n11879) );
  OAI211_X1 U14407 ( .C1(n14795), .C2(n13353), .A(n11880), .B(n11879), .ZN(
        P2_U3231) );
  NAND2_X1 U14408 ( .A1(n11884), .A2(n13309), .ZN(n11881) );
  XNOR2_X1 U14409 ( .A(n12020), .B(n12019), .ZN(n13653) );
  NOR2_X1 U14410 ( .A1(n11884), .A2(n11883), .ZN(n11886) );
  NAND2_X1 U14411 ( .A1(n11884), .A2(n11883), .ZN(n11885) );
  OAI21_X2 U14412 ( .B1(n11887), .B2(n11886), .A(n11885), .ZN(n11998) );
  XNOR2_X1 U14413 ( .A(n11998), .B(n12019), .ZN(n11888) );
  AOI22_X1 U14414 ( .A1(n13541), .A2(n13538), .B1(n13540), .B2(n13309), .ZN(
        n13253) );
  OAI21_X1 U14415 ( .B1(n11888), .B2(n13520), .A(n13253), .ZN(n13649) );
  NAND2_X1 U14416 ( .A1(n13649), .A2(n13562), .ZN(n11894) );
  AOI211_X1 U14417 ( .C1(n13651), .C2(n11889), .A(n6569), .B(n13557), .ZN(
        n13650) );
  INV_X1 U14418 ( .A(n13651), .ZN(n11891) );
  AOI22_X1 U14419 ( .A1(n13469), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14800), 
        .B2(n13249), .ZN(n11890) );
  OAI21_X1 U14420 ( .B1(n11891), .B2(n14803), .A(n11890), .ZN(n11892) );
  AOI21_X1 U14421 ( .B1(n13650), .B2(n14797), .A(n11892), .ZN(n11893) );
  OAI211_X1 U14422 ( .C1(n13653), .C2(n13576), .A(n11894), .B(n11893), .ZN(
        P2_U3248) );
  INV_X1 U14423 ( .A(n11895), .ZN(n11925) );
  AOI22_X1 U14424 ( .A1(n11896), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n14360), .ZN(n11897) );
  OAI21_X1 U14425 ( .B1(n11925), .B2(n14369), .A(n11897), .ZN(P1_U3330) );
  OAI211_X1 U14426 ( .C1(n11949), .C2(n14872), .A(n11898), .B(n11943), .ZN(
        n11900) );
  AOI211_X1 U14427 ( .C1(n11901), .C2(n13618), .A(n11900), .B(n11899), .ZN(
        n11904) );
  NAND2_X1 U14428 ( .A1(n14888), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11902) );
  OAI21_X1 U14429 ( .B1(n11904), .B2(n14888), .A(n11902), .ZN(P2_U3515) );
  NAND2_X1 U14430 ( .A1(n14878), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n11903) );
  OAI21_X1 U14431 ( .B1(n11904), .B2(n14878), .A(n11903), .ZN(P2_U3478) );
  AOI21_X1 U14432 ( .B1(n11906), .B2(n11805), .A(n12785), .ZN(n11923) );
  XNOR2_X1 U14433 ( .A(n12789), .B(n12801), .ZN(n11909) );
  NAND2_X1 U14434 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11909), .ZN(n12791) );
  OAI21_X1 U14435 ( .B1(n11909), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12791), 
        .ZN(n11921) );
  MUX2_X1 U14436 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6973), .Z(n12800) );
  XNOR2_X1 U14437 ( .A(n12800), .B(n12801), .ZN(n11912) );
  NAND2_X1 U14438 ( .A1(n11910), .A2(n14390), .ZN(n11913) );
  AND2_X1 U14439 ( .A1(n11912), .A2(n11913), .ZN(n11911) );
  NAND2_X1 U14440 ( .A1(n11914), .A2(n11911), .ZN(n12812) );
  INV_X1 U14441 ( .A(n12812), .ZN(n11916) );
  AOI21_X1 U14442 ( .B1(n11914), .B2(n11913), .A(n11912), .ZN(n11915) );
  OAI21_X1 U14443 ( .B1(n11916), .B2(n11915), .A(n15031), .ZN(n11919) );
  AOI21_X1 U14444 ( .B1(n14990), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11917), 
        .ZN(n11918) );
  OAI211_X1 U14445 ( .C1(n14985), .C2(n12790), .A(n11919), .B(n11918), .ZN(
        n11920) );
  AOI21_X1 U14446 ( .B1(n11921), .B2(n15023), .A(n11920), .ZN(n11922) );
  OAI21_X1 U14447 ( .B1(n11923), .B2(n15036), .A(n11922), .ZN(P3_U3195) );
  OAI222_X1 U14448 ( .A1(n12073), .A2(n15247), .B1(n12071), .B2(n11925), .C1(
        n11924), .C2(P2_U3088), .ZN(P2_U3302) );
  XNOR2_X1 U14449 ( .A(n11926), .B(n12606), .ZN(n11929) );
  NAND2_X1 U14450 ( .A1(n13050), .A2(n15064), .ZN(n11928) );
  NAND2_X1 U14451 ( .A1(n14415), .A2(n15061), .ZN(n11927) );
  AND2_X1 U14452 ( .A1(n11928), .A2(n11927), .ZN(n14447) );
  OAI21_X1 U14453 ( .B1(n11929), .B2(n13063), .A(n14447), .ZN(n13132) );
  INV_X1 U14454 ( .A(n13132), .ZN(n11934) );
  XNOR2_X1 U14455 ( .A(n11930), .B(n12606), .ZN(n13133) );
  INV_X1 U14456 ( .A(n14442), .ZN(n13197) );
  AOI22_X1 U14457 ( .A1(n15079), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13069), 
        .B2(n14443), .ZN(n11931) );
  OAI21_X1 U14458 ( .B1(n13197), .B2(n13071), .A(n11931), .ZN(n11932) );
  AOI21_X1 U14459 ( .B1(n13133), .B2(n13073), .A(n11932), .ZN(n11933) );
  OAI21_X1 U14460 ( .B1(n11934), .B2(n15079), .A(n11933), .ZN(P3_U3217) );
  INV_X1 U14461 ( .A(n13254), .ZN(n11936) );
  NOR2_X1 U14462 ( .A1(n11936), .A2(n11935), .ZN(n11940) );
  AND2_X1 U14463 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  NAND2_X1 U14464 ( .A1(n11939), .A2(n11940), .ZN(n13256) );
  OAI21_X1 U14465 ( .B1(n11940), .B2(n11939), .A(n13256), .ZN(n11941) );
  NAND2_X1 U14466 ( .A1(n11941), .A2(n13278), .ZN(n11947) );
  OAI21_X1 U14467 ( .B1(n13252), .B2(n11943), .A(n11942), .ZN(n11944) );
  AOI21_X1 U14468 ( .B1(n11945), .B2(n13283), .A(n11944), .ZN(n11946) );
  OAI211_X1 U14469 ( .C1(n11949), .C2(n11948), .A(n11947), .B(n11946), .ZN(
        P2_U3198) );
  INV_X1 U14470 ( .A(n11951), .ZN(n11952) );
  NAND2_X1 U14471 ( .A1(n11950), .A2(n11952), .ZN(n11953) );
  OAI22_X1 U14472 ( .A1(n12170), .A2(n12395), .B1(n12166), .B2(n12394), .ZN(
        n12369) );
  NAND2_X1 U14473 ( .A1(n12171), .A2(n6962), .ZN(n11956) );
  NAND2_X1 U14474 ( .A1(n13848), .A2(n12455), .ZN(n11955) );
  NAND2_X1 U14475 ( .A1(n11956), .A2(n11955), .ZN(n11957) );
  XNOR2_X1 U14476 ( .A(n11957), .B(n12450), .ZN(n12370) );
  XOR2_X1 U14477 ( .A(n12369), .B(n12370), .Z(n12372) );
  XNOR2_X1 U14478 ( .A(n12373), .B(n12372), .ZN(n11964) );
  OAI21_X1 U14479 ( .B1(n13761), .B2(n12167), .A(n11958), .ZN(n11959) );
  AOI21_X1 U14480 ( .B1(n13758), .B2(n13847), .A(n11959), .ZN(n11960) );
  OAI21_X1 U14481 ( .B1(n13832), .B2(n11961), .A(n11960), .ZN(n11962) );
  AOI21_X1 U14482 ( .B1(n13834), .B2(n12171), .A(n11962), .ZN(n11963) );
  OAI21_X1 U14483 ( .B1(n11964), .B2(n13836), .A(n11963), .ZN(P1_U3234) );
  XNOR2_X1 U14484 ( .A(n11966), .B(n11965), .ZN(n11970) );
  NOR2_X1 U14485 ( .A1(n13297), .A2(n13572), .ZN(n11968) );
  AOI22_X1 U14486 ( .A1(n13307), .A2(n13538), .B1(n13540), .B2(n13308), .ZN(
        n13567) );
  NAND2_X1 U14487 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13348)
         );
  OAI21_X1 U14488 ( .B1(n13567), .B2(n13252), .A(n13348), .ZN(n11967) );
  AOI211_X1 U14489 ( .C1(n13645), .C2(n13302), .A(n11968), .B(n11967), .ZN(
        n11969) );
  OAI21_X1 U14490 ( .B1(n11970), .B2(n13304), .A(n11969), .ZN(P2_U3210) );
  INV_X1 U14491 ( .A(n11971), .ZN(n11975) );
  OAI222_X1 U14492 ( .A1(n11973), .A2(P2_U3088), .B1(n12071), .B2(n11975), 
        .C1(n11972), .C2(n12073), .ZN(P2_U3301) );
  OAI222_X1 U14493 ( .A1(P1_U3086), .A2(n11976), .B1(n14369), .B2(n11975), 
        .C1(n11974), .C2(n14366), .ZN(P1_U3329) );
  NAND2_X1 U14494 ( .A1(n11978), .A2(n11977), .ZN(n11979) );
  NAND2_X1 U14495 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  NAND2_X1 U14496 ( .A1(n11981), .A2(n14707), .ZN(n11988) );
  NAND2_X1 U14497 ( .A1(n11982), .A2(n12304), .ZN(n11983) );
  NAND2_X1 U14498 ( .A1(n11984), .A2(n11983), .ZN(n11985) );
  NAND2_X1 U14499 ( .A1(n11985), .A2(n14611), .ZN(n11987) );
  NAND3_X1 U14500 ( .A1(n11988), .A2(n11987), .A3(n11986), .ZN(n14690) );
  MUX2_X1 U14501 ( .A(n14690), .B(P1_REG2_REG_5__SCAN_IN), .S(n14642), .Z(
        n11997) );
  INV_X1 U14502 ( .A(n11989), .ZN(n11990) );
  NAND2_X1 U14503 ( .A1(n14599), .A2(n11990), .ZN(n11994) );
  OAI21_X1 U14504 ( .B1(n14621), .B2(n11995), .A(n14622), .ZN(n11992) );
  NOR2_X1 U14505 ( .A1(n11992), .A2(n11991), .ZN(n14691) );
  NAND2_X1 U14506 ( .A1(n14626), .A2(n14691), .ZN(n11993) );
  OAI211_X1 U14507 ( .C1(n14616), .C2(n11995), .A(n11994), .B(n11993), .ZN(
        n11996) );
  OR2_X1 U14508 ( .A1(n11997), .A2(n11996), .ZN(P1_U3288) );
  NAND2_X1 U14509 ( .A1(n13651), .A2(n11999), .ZN(n12000) );
  AND2_X1 U14510 ( .A1(n13645), .A2(n12002), .ZN(n12001) );
  OR2_X1 U14511 ( .A1(n13645), .A2(n12002), .ZN(n12003) );
  INV_X1 U14512 ( .A(n13307), .ZN(n13521) );
  NAND2_X1 U14513 ( .A1(n13640), .A2(n13521), .ZN(n12004) );
  NAND2_X1 U14514 ( .A1(n13536), .A2(n12004), .ZN(n12006) );
  OR2_X1 U14515 ( .A1(n13640), .A2(n13521), .ZN(n12005) );
  NAND2_X1 U14516 ( .A1(n13629), .A2(n13523), .ZN(n12008) );
  INV_X1 U14517 ( .A(n13614), .ZN(n13475) );
  INV_X1 U14518 ( .A(n13459), .ZN(n13454) );
  NAND2_X1 U14519 ( .A1(n13607), .A2(n12009), .ZN(n13445) );
  INV_X1 U14520 ( .A(n12010), .ZN(n12012) );
  NAND2_X1 U14521 ( .A1(n13414), .A2(n13540), .ZN(n12017) );
  AOI21_X1 U14522 ( .B1(n12015), .B2(P2_B_REG_SCAN_IN), .A(n13524), .ZN(n13379) );
  NAND2_X1 U14523 ( .A1(n13306), .A2(n13379), .ZN(n12016) );
  NAND2_X1 U14524 ( .A1(n13651), .A2(n13308), .ZN(n12021) );
  OR2_X1 U14525 ( .A1(n13645), .A2(n13541), .ZN(n12023) );
  NAND2_X1 U14526 ( .A1(n13635), .A2(n13539), .ZN(n12026) );
  OR2_X1 U14527 ( .A1(n13635), .A2(n13539), .ZN(n12027) );
  NAND2_X1 U14528 ( .A1(n13510), .A2(n13509), .ZN(n12030) );
  INV_X1 U14529 ( .A(n13629), .ZN(n13508) );
  NAND2_X1 U14530 ( .A1(n13508), .A2(n13523), .ZN(n12029) );
  NAND2_X1 U14531 ( .A1(n13621), .A2(n13502), .ZN(n12032) );
  NAND2_X1 U14532 ( .A1(n13607), .A2(n13471), .ZN(n12033) );
  OR2_X1 U14533 ( .A1(n13603), .A2(n13456), .ZN(n12034) );
  NAND2_X1 U14534 ( .A1(n13440), .A2(n12034), .ZN(n12036) );
  NAND2_X1 U14535 ( .A1(n13603), .A2(n13456), .ZN(n12035) );
  AND2_X1 U14536 ( .A1(n13598), .A2(n13448), .ZN(n12037) );
  INV_X1 U14537 ( .A(n13585), .ZN(n12046) );
  INV_X1 U14538 ( .A(n13583), .ZN(n12044) );
  INV_X1 U14539 ( .A(n13645), .ZN(n13563) );
  INV_X1 U14540 ( .A(n13607), .ZN(n13462) );
  AOI21_X1 U14541 ( .B1(n13396), .B2(n13583), .A(n8811), .ZN(n12040) );
  NAND2_X1 U14542 ( .A1(n13582), .A2(n14797), .ZN(n12043) );
  AOI22_X1 U14543 ( .A1(n13469), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n14800), 
        .B2(n12041), .ZN(n12042) );
  OAI211_X1 U14544 ( .C1(n12044), .C2(n14803), .A(n12043), .B(n12042), .ZN(
        n12045) );
  AOI21_X1 U14545 ( .B1(n12046), .B2(n14806), .A(n12045), .ZN(n12047) );
  OAI21_X1 U14546 ( .B1(n6623), .B2(n13469), .A(n12047), .ZN(P2_U3236) );
  INV_X1 U14547 ( .A(n12048), .ZN(n13700) );
  OAI222_X1 U14548 ( .A1(n13875), .A2(P1_U3086), .B1(n12362), .B2(n13700), 
        .C1(n15279), .C2(n14366), .ZN(P1_U3327) );
  INV_X1 U14549 ( .A(n12049), .ZN(n14368) );
  OAI222_X1 U14550 ( .A1(n12073), .A2(n12051), .B1(n12071), .B2(n14368), .C1(
        n12050), .C2(P2_U3088), .ZN(P2_U3300) );
  AND2_X1 U14551 ( .A1(n13839), .A2(n14207), .ZN(n12054) );
  AOI211_X2 U14552 ( .C1(n12055), .C2(n14611), .A(n12054), .B(n12053), .ZN(
        n14267) );
  INV_X1 U14553 ( .A(n12056), .ZN(n12057) );
  AOI211_X1 U14554 ( .C1(n14265), .C2(n14036), .A(n14242), .B(n12057), .ZN(
        n14264) );
  INV_X1 U14555 ( .A(n14265), .ZN(n12060) );
  INV_X1 U14556 ( .A(n12470), .ZN(n12058) );
  AOI22_X1 U14557 ( .A1(n14642), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n12058), 
        .B2(n14599), .ZN(n12059) );
  OAI21_X1 U14558 ( .B1(n12060), .B2(n14616), .A(n12059), .ZN(n12065) );
  OAI21_X1 U14559 ( .B1(n12063), .B2(n12062), .A(n12061), .ZN(n14268) );
  NOR2_X1 U14560 ( .A1(n14268), .A2(n14249), .ZN(n12064) );
  OAI21_X1 U14561 ( .B1(n14267), .B2(n14642), .A(n12066), .ZN(P1_U3265) );
  INV_X1 U14562 ( .A(n12260), .ZN(n12361) );
  INV_X1 U14563 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n15415) );
  OAI222_X1 U14564 ( .A1(n12071), .A2(n12361), .B1(P2_U3088), .B2(n12067), 
        .C1(n15415), .C2(n12073), .ZN(P2_U3297) );
  INV_X1 U14565 ( .A(n12068), .ZN(n12070) );
  OAI222_X1 U14566 ( .A1(n12073), .A2(n12072), .B1(n12071), .B2(n12070), .C1(
        n12069), .C2(P2_U3088), .ZN(P2_U3305) );
  AOI21_X1 U14567 ( .B1(n12074), .B2(n12075), .A(n14427), .ZN(n12077) );
  NAND2_X1 U14568 ( .A1(n12077), .A2(n12076), .ZN(n12083) );
  AND2_X1 U14569 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12831) );
  AOI21_X1 U14570 ( .B1(n14416), .B2(n12769), .A(n12831), .ZN(n12078) );
  OAI21_X1 U14571 ( .B1(n12079), .B2(n14418), .A(n12078), .ZN(n12080) );
  AOI21_X1 U14572 ( .B1(n12081), .B2(n14444), .A(n12080), .ZN(n12082) );
  OAI211_X1 U14573 ( .C1(n12084), .C2(n12574), .A(n12083), .B(n12082), .ZN(
        P3_U3181) );
  AND2_X1 U14574 ( .A1(n12085), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14575 ( .A1(n12085), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U14576 ( .A1(n12085), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14577 ( .A1(n12085), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14578 ( .A1(n12085), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14579 ( .A1(n12085), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14580 ( .A1(n12085), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14581 ( .A1(n12085), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14582 ( .A1(n12085), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14583 ( .A1(n12085), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U14584 ( .A1(n12085), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U14585 ( .A1(n12085), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14586 ( .A1(n12085), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14587 ( .A1(n12085), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14588 ( .A1(n12085), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14589 ( .A1(n12085), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14590 ( .A1(n12085), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14591 ( .A1(n12085), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14592 ( .A1(n12085), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14593 ( .A1(n12085), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14594 ( .A1(n12085), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U14595 ( .A1(n12085), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U14596 ( .A1(n12085), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14597 ( .A1(n12085), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U14598 ( .A1(n12085), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  NAND2_X1 U14599 ( .A1(n12088), .A2(n12087), .ZN(n12271) );
  INV_X4 U14600 ( .A(n12165), .ZN(n12189) );
  AND2_X1 U14601 ( .A1(n12092), .A2(n12288), .ZN(n12096) );
  INV_X1 U14602 ( .A(n12093), .ZN(n12094) );
  NAND2_X1 U14603 ( .A1(n12099), .A2(n12098), .ZN(n12103) );
  MUX2_X1 U14604 ( .A(n13860), .B(n12100), .S(n12189), .Z(n12102) );
  NAND2_X1 U14605 ( .A1(n12103), .A2(n7704), .ZN(n12105) );
  MUX2_X1 U14606 ( .A(n12106), .B(n12107), .S(n12189), .Z(n12104) );
  NAND2_X1 U14607 ( .A1(n12105), .A2(n12104), .ZN(n12109) );
  MUX2_X1 U14608 ( .A(n12107), .B(n12106), .S(n12189), .Z(n12108) );
  NAND3_X1 U14609 ( .A1(n12109), .A2(n12302), .A3(n12108), .ZN(n12113) );
  MUX2_X1 U14610 ( .A(n12111), .B(n12110), .S(n12189), .Z(n12112) );
  NAND2_X1 U14611 ( .A1(n12113), .A2(n12112), .ZN(n12118) );
  MUX2_X1 U14612 ( .A(n12114), .B(n14684), .S(n12165), .Z(n12117) );
  MUX2_X1 U14613 ( .A(n12115), .B(n13857), .S(n12165), .Z(n12116) );
  NAND2_X1 U14614 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  MUX2_X1 U14615 ( .A(n13856), .B(n14692), .S(n12189), .Z(n12122) );
  MUX2_X1 U14616 ( .A(n14692), .B(n13856), .S(n12189), .Z(n12121) );
  BUF_X1 U14617 ( .A(n12165), .Z(n12256) );
  MUX2_X1 U14618 ( .A(n14696), .B(n13855), .S(n12293), .Z(n12125) );
  NAND2_X1 U14619 ( .A1(n12126), .A2(n12125), .ZN(n12124) );
  MUX2_X1 U14620 ( .A(n13855), .B(n14696), .S(n12293), .Z(n12123) );
  NAND2_X1 U14621 ( .A1(n12124), .A2(n12123), .ZN(n12128) );
  MUX2_X1 U14622 ( .A(n13854), .B(n12129), .S(n12189), .Z(n12131) );
  MUX2_X1 U14623 ( .A(n12129), .B(n13854), .S(n12293), .Z(n12130) );
  MUX2_X1 U14624 ( .A(n13853), .B(n12132), .S(n12165), .Z(n12136) );
  NAND2_X1 U14625 ( .A1(n12135), .A2(n12136), .ZN(n12134) );
  MUX2_X1 U14626 ( .A(n13853), .B(n12132), .S(n12293), .Z(n12133) );
  NAND2_X1 U14627 ( .A1(n12134), .A2(n12133), .ZN(n12140) );
  INV_X1 U14628 ( .A(n12135), .ZN(n12138) );
  INV_X1 U14629 ( .A(n12136), .ZN(n12137) );
  NAND2_X1 U14630 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  NAND2_X1 U14631 ( .A1(n12140), .A2(n12139), .ZN(n12144) );
  MUX2_X1 U14632 ( .A(n13852), .B(n12141), .S(n12293), .Z(n12145) );
  NAND2_X1 U14633 ( .A1(n12144), .A2(n12145), .ZN(n12143) );
  MUX2_X1 U14634 ( .A(n13852), .B(n12141), .S(n12165), .Z(n12142) );
  NAND2_X1 U14635 ( .A1(n12143), .A2(n12142), .ZN(n12149) );
  INV_X1 U14636 ( .A(n12144), .ZN(n12147) );
  INV_X1 U14637 ( .A(n12145), .ZN(n12146) );
  NAND2_X1 U14638 ( .A1(n12149), .A2(n12148), .ZN(n12152) );
  MUX2_X1 U14639 ( .A(n13851), .B(n12150), .S(n12165), .Z(n12153) );
  MUX2_X1 U14640 ( .A(n13851), .B(n12150), .S(n12293), .Z(n12151) );
  NAND2_X1 U14641 ( .A1(n12181), .A2(n12166), .ZN(n12157) );
  MUX2_X1 U14642 ( .A(n13849), .B(n14401), .S(n12256), .Z(n12173) );
  NAND2_X1 U14643 ( .A1(n12171), .A2(n12166), .ZN(n12154) );
  OAI21_X1 U14644 ( .B1(n12173), .B2(n12155), .A(n12154), .ZN(n12156) );
  AOI21_X1 U14645 ( .B1(n12177), .B2(n12157), .A(n12156), .ZN(n12162) );
  MUX2_X1 U14646 ( .A(n12158), .B(n14530), .S(n12256), .Z(n12164) );
  MUX2_X1 U14647 ( .A(n13850), .B(n12159), .S(n12293), .Z(n12163) );
  NAND2_X1 U14648 ( .A1(n12164), .A2(n12163), .ZN(n12160) );
  AOI22_X1 U14649 ( .A1(n12173), .A2(n12167), .B1(n12165), .B2(n12166), .ZN(
        n12176) );
  NAND2_X1 U14650 ( .A1(n12189), .A2(n13848), .ZN(n12168) );
  AOI21_X1 U14651 ( .B1(n12171), .B2(n14401), .A(n12168), .ZN(n12169) );
  OAI21_X1 U14652 ( .B1(n12173), .B2(n12170), .A(n12169), .ZN(n12175) );
  OAI22_X1 U14653 ( .A1(n12171), .A2(n14401), .B1(n13848), .B2(n13849), .ZN(
        n12172) );
  NAND3_X1 U14654 ( .A1(n12181), .A2(n12173), .A3(n12172), .ZN(n12174) );
  OAI211_X1 U14655 ( .C1(n12177), .C2(n12176), .A(n12175), .B(n12174), .ZN(
        n12178) );
  NAND2_X1 U14656 ( .A1(n12181), .A2(n12179), .ZN(n12184) );
  NAND2_X1 U14657 ( .A1(n12186), .A2(n12180), .ZN(n12182) );
  AND2_X1 U14658 ( .A1(n12182), .A2(n12181), .ZN(n12183) );
  MUX2_X1 U14659 ( .A(n12184), .B(n12183), .S(n12256), .Z(n12185) );
  MUX2_X1 U14660 ( .A(n14208), .B(n14330), .S(n12189), .Z(n12202) );
  NAND2_X1 U14661 ( .A1(n12202), .A2(n13845), .ZN(n12187) );
  NAND2_X1 U14662 ( .A1(n12189), .A2(n13828), .ZN(n12200) );
  AOI21_X1 U14663 ( .B1(n12187), .B2(n12200), .A(n14202), .ZN(n12193) );
  NAND2_X1 U14664 ( .A1(n12202), .A2(n14220), .ZN(n12188) );
  OR2_X1 U14665 ( .A1(n14330), .A2(n12189), .ZN(n12194) );
  AOI21_X1 U14666 ( .B1(n12188), .B2(n12194), .A(n12204), .ZN(n12192) );
  NAND2_X1 U14667 ( .A1(n12165), .A2(n13845), .ZN(n12196) );
  OR2_X1 U14668 ( .A1(n14330), .A2(n12196), .ZN(n12191) );
  NAND3_X1 U14669 ( .A1(n12189), .A2(n13828), .A3(n14220), .ZN(n12190) );
  NAND2_X1 U14670 ( .A1(n12191), .A2(n12190), .ZN(n12198) );
  INV_X1 U14671 ( .A(n12194), .ZN(n12195) );
  NAND2_X1 U14672 ( .A1(n12202), .A2(n12195), .ZN(n12197) );
  NAND2_X1 U14673 ( .A1(n12197), .A2(n12196), .ZN(n12199) );
  AOI22_X1 U14674 ( .A1(n12199), .A2(n14202), .B1(n12202), .B2(n12198), .ZN(
        n12207) );
  INV_X1 U14675 ( .A(n12200), .ZN(n12201) );
  AOI22_X1 U14676 ( .A1(n12202), .A2(n12201), .B1(n14220), .B2(n12189), .ZN(
        n12203) );
  INV_X1 U14677 ( .A(n12203), .ZN(n12205) );
  NAND2_X1 U14678 ( .A1(n12205), .A2(n12204), .ZN(n12206) );
  MUX2_X1 U14679 ( .A(n13774), .B(n14318), .S(n12165), .Z(n12208) );
  OAI21_X1 U14680 ( .B1(n12211), .B2(n12209), .A(n12208), .ZN(n12213) );
  NAND2_X1 U14681 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  MUX2_X1 U14682 ( .A(n12215), .B(n12214), .S(n12293), .Z(n12216) );
  MUX2_X1 U14683 ( .A(n13844), .B(n14304), .S(n12293), .Z(n12217) );
  INV_X1 U14684 ( .A(n12217), .ZN(n12219) );
  MUX2_X1 U14685 ( .A(n14304), .B(n13844), .S(n12293), .Z(n12218) );
  MUX2_X1 U14686 ( .A(n14152), .B(n14299), .S(n12256), .Z(n12222) );
  MUX2_X1 U14687 ( .A(n14299), .B(n14152), .S(n12256), .Z(n12220) );
  NAND2_X1 U14688 ( .A1(n12221), .A2(n12220), .ZN(n12224) );
  MUX2_X1 U14689 ( .A(n13843), .B(n14128), .S(n12293), .Z(n12226) );
  MUX2_X1 U14690 ( .A(n13843), .B(n14128), .S(n12165), .Z(n12225) );
  INV_X1 U14691 ( .A(n12226), .ZN(n12227) );
  MUX2_X1 U14692 ( .A(n14121), .B(n14291), .S(n12165), .Z(n12230) );
  NAND2_X1 U14693 ( .A1(n12231), .A2(n12230), .ZN(n12229) );
  MUX2_X1 U14694 ( .A(n14121), .B(n14291), .S(n12293), .Z(n12228) );
  NAND2_X1 U14695 ( .A1(n12229), .A2(n12228), .ZN(n12233) );
  MUX2_X1 U14696 ( .A(n14097), .B(n13842), .S(n12256), .Z(n12235) );
  MUX2_X1 U14697 ( .A(n14097), .B(n13842), .S(n12293), .Z(n12234) );
  MUX2_X1 U14698 ( .A(n13841), .B(n14077), .S(n12256), .Z(n12238) );
  MUX2_X1 U14699 ( .A(n13841), .B(n14077), .S(n12293), .Z(n12236) );
  INV_X1 U14700 ( .A(n12238), .ZN(n12239) );
  MUX2_X1 U14701 ( .A(n14033), .B(n14275), .S(n12189), .Z(n12243) );
  MUX2_X1 U14702 ( .A(n14033), .B(n14275), .S(n12165), .Z(n12240) );
  NAND2_X1 U14703 ( .A1(n12241), .A2(n12240), .ZN(n12247) );
  INV_X1 U14704 ( .A(n12242), .ZN(n12245) );
  INV_X1 U14705 ( .A(n12243), .ZN(n12244) );
  NAND2_X1 U14706 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  MUX2_X1 U14707 ( .A(n14270), .B(n13840), .S(n12189), .Z(n12249) );
  MUX2_X1 U14708 ( .A(n14270), .B(n13840), .S(n12256), .Z(n12248) );
  MUX2_X1 U14709 ( .A(n14034), .B(n14265), .S(n12189), .Z(n12253) );
  NAND2_X1 U14710 ( .A1(n12252), .A2(n12253), .ZN(n12251) );
  MUX2_X1 U14711 ( .A(n14034), .B(n14265), .S(n12256), .Z(n12250) );
  INV_X1 U14712 ( .A(n12252), .ZN(n12255) );
  INV_X1 U14713 ( .A(n12253), .ZN(n12254) );
  MUX2_X1 U14714 ( .A(n13839), .B(n14260), .S(n12256), .Z(n12257) );
  MUX2_X1 U14715 ( .A(n13839), .B(n14260), .S(n12189), .Z(n12258) );
  NAND2_X1 U14716 ( .A1(n12260), .A2(n12259), .ZN(n12262) );
  NAND2_X1 U14717 ( .A1(n12283), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12261) );
  INV_X1 U14718 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n12263) );
  OR2_X1 U14719 ( .A1(n12264), .A2(n12263), .ZN(n12270) );
  INV_X1 U14720 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n12265) );
  OR2_X1 U14721 ( .A1(n12266), .A2(n12265), .ZN(n12269) );
  INV_X1 U14722 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15419) );
  OR2_X1 U14723 ( .A1(n12267), .A2(n15419), .ZN(n12268) );
  INV_X1 U14724 ( .A(n12271), .ZN(n12272) );
  OAI22_X1 U14725 ( .A1(n12293), .A2(n12291), .B1(n12273), .B2(n12272), .ZN(
        n12274) );
  AOI22_X1 U14726 ( .A1(n14029), .A2(n12189), .B1(n13838), .B2(n12274), .ZN(
        n12278) );
  NAND2_X1 U14727 ( .A1(n12277), .A2(n12278), .ZN(n12282) );
  OAI21_X1 U14728 ( .B1(n14021), .B2(n12275), .A(n13838), .ZN(n12276) );
  MUX2_X1 U14729 ( .A(n14257), .B(n12276), .S(n12189), .Z(n12281) );
  INV_X1 U14730 ( .A(n12277), .ZN(n12280) );
  INV_X1 U14731 ( .A(n12278), .ZN(n12279) );
  AOI22_X1 U14732 ( .A1(n12282), .A2(n12281), .B1(n12280), .B2(n12279), .ZN(
        n12297) );
  NAND2_X1 U14733 ( .A1(n13690), .A2(n9433), .ZN(n12285) );
  NAND2_X1 U14734 ( .A1(n12283), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12284) );
  XNOR2_X1 U14735 ( .A(n12292), .B(n12291), .ZN(n12335) );
  NAND2_X1 U14736 ( .A1(n12287), .A2(n12286), .ZN(n12290) );
  NAND2_X1 U14737 ( .A1(n12288), .A2(n14143), .ZN(n12289) );
  NAND2_X1 U14738 ( .A1(n12290), .A2(n12289), .ZN(n12334) );
  NOR3_X1 U14739 ( .A1(n12297), .A2(n12335), .A3(n12334), .ZN(n12345) );
  NOR2_X1 U14740 ( .A1(n14254), .A2(n14021), .ZN(n12295) );
  NOR2_X1 U14741 ( .A1(n12292), .A2(n12291), .ZN(n12294) );
  MUX2_X1 U14742 ( .A(n12295), .B(n12294), .S(n12293), .Z(n12338) );
  NAND2_X1 U14743 ( .A1(n12334), .A2(n12332), .ZN(n12336) );
  INV_X1 U14744 ( .A(n12336), .ZN(n12296) );
  XOR2_X1 U14745 ( .A(n13838), .B(n14029), .Z(n12330) );
  NOR2_X1 U14746 ( .A1(n10736), .A2(n12298), .ZN(n12303) );
  NAND2_X1 U14747 ( .A1(n12300), .A2(n12299), .ZN(n14618) );
  NAND4_X1 U14748 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n14618), .ZN(
        n12305) );
  NOR2_X1 U14749 ( .A1(n12305), .A2(n12304), .ZN(n12308) );
  NAND4_X1 U14750 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12310) );
  NOR2_X1 U14751 ( .A1(n12311), .A2(n12310), .ZN(n12314) );
  NAND4_X1 U14752 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n12312), .ZN(
        n12316) );
  OR4_X1 U14753 ( .A1(n9475), .A2(n12317), .A3(n14228), .A4(n12316), .ZN(
        n12318) );
  OR4_X1 U14754 ( .A1(n12319), .A2(n14203), .A3(n14235), .A4(n12318), .ZN(
        n12320) );
  NOR2_X1 U14755 ( .A1(n12321), .A2(n12320), .ZN(n12322) );
  AND4_X1 U14756 ( .A1(n14105), .A2(n12322), .A3(n14134), .A4(n14161), .ZN(
        n12323) );
  NAND4_X1 U14757 ( .A1(n14072), .A2(n12324), .A3(n12323), .A4(n14085), .ZN(
        n12325) );
  NOR2_X1 U14758 ( .A1(n14056), .A2(n12325), .ZN(n12327) );
  NAND4_X1 U14759 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n7328), .ZN(
        n12329) );
  NOR3_X1 U14760 ( .A1(n12335), .A2(n12330), .A3(n12329), .ZN(n12331) );
  XOR2_X1 U14761 ( .A(n14014), .B(n12331), .Z(n12333) );
  NOR2_X1 U14762 ( .A1(n12333), .A2(n12332), .ZN(n12343) );
  INV_X1 U14763 ( .A(n12334), .ZN(n12341) );
  INV_X1 U14764 ( .A(n12335), .ZN(n12337) );
  NOR2_X1 U14765 ( .A1(n12337), .A2(n12336), .ZN(n12340) );
  INV_X1 U14766 ( .A(n12338), .ZN(n12339) );
  MUX2_X1 U14767 ( .A(n12341), .B(n12340), .S(n12339), .Z(n12342) );
  NAND3_X1 U14768 ( .A1(n12346), .A2(n14564), .A3(n14209), .ZN(n12347) );
  OAI211_X1 U14769 ( .C1(n14371), .C2(n12349), .A(n12347), .B(P1_B_REG_SCAN_IN), .ZN(n12348) );
  OAI21_X1 U14770 ( .B1(n12350), .B2(n12349), .A(n12348), .ZN(P1_U3242) );
  INV_X1 U14771 ( .A(n15065), .ZN(n12354) );
  INV_X1 U14772 ( .A(n15066), .ZN(n12599) );
  NOR3_X1 U14773 ( .A1(n12599), .A2(n12352), .A3(n15060), .ZN(n12353) );
  OAI22_X1 U14774 ( .A1(n12526), .A2(n12355), .B1(n15059), .B2(n12574), .ZN(
        n12356) );
  AOI21_X1 U14775 ( .B1(n12479), .B2(n15062), .A(n12356), .ZN(n12359) );
  NAND2_X1 U14776 ( .A1(n12357), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n12358) );
  OAI211_X1 U14777 ( .C1(n12360), .C2(n14427), .A(n12359), .B(n12358), .ZN(
        P3_U3162) );
  INV_X1 U14778 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12577) );
  OAI222_X1 U14779 ( .A1(n12362), .A2(n12361), .B1(n9282), .B2(P1_U3086), .C1(
        n12577), .C2(n14366), .ZN(P1_U3325) );
  OAI222_X1 U14780 ( .A1(n15458), .A2(n12364), .B1(n12759), .B2(P3_U3151), 
        .C1(n12363), .C2(n15456), .ZN(P3_U3267) );
  INV_X1 U14781 ( .A(SI_30_), .ZN(n12586) );
  NAND2_X1 U14782 ( .A1(n13695), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12366) );
  XOR2_X1 U14783 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .Z(n12368) );
  XNOR2_X1 U14784 ( .A(n12575), .B(n12368), .ZN(n12587) );
  OAI222_X1 U14785 ( .A1(P3_U3151), .A2(n12365), .B1(n15456), .B2(n12586), 
        .C1(n15458), .C2(n12587), .ZN(P3_U3265) );
  OAI22_X1 U14786 ( .A1(n14525), .A2(n12396), .B1(n13829), .B2(n12395), .ZN(
        n12374) );
  XNOR2_X1 U14787 ( .A(n12374), .B(n12450), .ZN(n12376) );
  OAI22_X1 U14788 ( .A1(n14525), .A2(n12395), .B1(n13829), .B2(n12394), .ZN(
        n12375) );
  NOR2_X1 U14789 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  AOI21_X1 U14790 ( .B1(n12376), .B2(n12375), .A(n12377), .ZN(n13712) );
  INV_X1 U14791 ( .A(n12377), .ZN(n12378) );
  NAND2_X1 U14792 ( .A1(n14334), .A2(n6962), .ZN(n12380) );
  NAND2_X1 U14793 ( .A1(n13846), .A2(n12455), .ZN(n12379) );
  NAND2_X1 U14794 ( .A1(n12380), .A2(n12379), .ZN(n12381) );
  XNOR2_X1 U14795 ( .A(n12381), .B(n12450), .ZN(n12383) );
  INV_X1 U14796 ( .A(n14334), .ZN(n14246) );
  OAI22_X1 U14797 ( .A1(n14246), .A2(n12395), .B1(n14217), .B2(n12394), .ZN(
        n13827) );
  INV_X1 U14798 ( .A(n12382), .ZN(n12384) );
  AOI22_X1 U14799 ( .A1(n14330), .A2(n6962), .B1(n12455), .B2(n14208), .ZN(
        n12385) );
  XOR2_X1 U14800 ( .A(n12450), .B(n12385), .Z(n12387) );
  OAI22_X1 U14801 ( .A1(n14227), .A2(n12395), .B1(n13828), .B2(n12394), .ZN(
        n12386) );
  NOR2_X1 U14802 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  AOI21_X1 U14803 ( .B1(n12387), .B2(n12386), .A(n12388), .ZN(n13756) );
  INV_X1 U14804 ( .A(n12388), .ZN(n12389) );
  OAI22_X1 U14805 ( .A1(n14202), .A2(n12396), .B1(n14220), .B2(n12395), .ZN(
        n12390) );
  XNOR2_X1 U14806 ( .A(n12390), .B(n12450), .ZN(n12393) );
  OAI22_X1 U14807 ( .A1(n14202), .A2(n12395), .B1(n14220), .B2(n12394), .ZN(
        n12392) );
  NAND2_X1 U14808 ( .A1(n12393), .A2(n12392), .ZN(n13769) );
  OR2_X1 U14809 ( .A1(n12393), .A2(n12392), .ZN(n13768) );
  OAI22_X1 U14810 ( .A1(n14318), .A2(n12395), .B1(n13774), .B2(n12394), .ZN(
        n12398) );
  OAI22_X1 U14811 ( .A1(n14318), .A2(n12396), .B1(n13774), .B2(n12395), .ZN(
        n12397) );
  XNOR2_X1 U14812 ( .A(n12397), .B(n12450), .ZN(n12399) );
  XOR2_X1 U14813 ( .A(n12398), .B(n12399), .Z(n13808) );
  AOI22_X1 U14814 ( .A1(n14313), .A2(n6962), .B1(n12455), .B2(n14151), .ZN(
        n12401) );
  XNOR2_X1 U14815 ( .A(n12401), .B(n12450), .ZN(n12402) );
  AOI22_X1 U14816 ( .A1(n14313), .A2(n12455), .B1(n12462), .B2(n14151), .ZN(
        n12403) );
  XNOR2_X1 U14817 ( .A(n12402), .B(n12403), .ZN(n13726) );
  INV_X1 U14818 ( .A(n12402), .ZN(n12405) );
  INV_X1 U14819 ( .A(n12403), .ZN(n12404) );
  AND2_X1 U14820 ( .A1(n12462), .A2(n13844), .ZN(n12406) );
  AOI21_X1 U14821 ( .B1(n14304), .B2(n12455), .A(n12406), .ZN(n12409) );
  AOI22_X1 U14822 ( .A1(n14304), .A2(n6962), .B1(n12455), .B2(n13844), .ZN(
        n12407) );
  XNOR2_X1 U14823 ( .A(n12407), .B(n12450), .ZN(n12408) );
  XOR2_X1 U14824 ( .A(n12409), .B(n12408), .Z(n13786) );
  INV_X1 U14825 ( .A(n12408), .ZN(n12411) );
  INV_X1 U14826 ( .A(n12409), .ZN(n12410) );
  NAND2_X1 U14827 ( .A1(n12411), .A2(n12410), .ZN(n12412) );
  AOI22_X1 U14828 ( .A1(n14299), .A2(n6962), .B1(n12455), .B2(n14152), .ZN(
        n12413) );
  XNOR2_X1 U14829 ( .A(n12413), .B(n12450), .ZN(n12416) );
  AOI22_X1 U14830 ( .A1(n14299), .A2(n12455), .B1(n12462), .B2(n14152), .ZN(
        n12415) );
  XNOR2_X1 U14831 ( .A(n12416), .B(n12415), .ZN(n13739) );
  INV_X1 U14832 ( .A(n13739), .ZN(n12414) );
  NAND2_X1 U14833 ( .A1(n12416), .A2(n12415), .ZN(n12417) );
  NAND2_X1 U14834 ( .A1(n14128), .A2(n6962), .ZN(n12419) );
  NAND2_X1 U14835 ( .A1(n13843), .A2(n12463), .ZN(n12418) );
  NAND2_X1 U14836 ( .A1(n12419), .A2(n12418), .ZN(n12420) );
  XNOR2_X1 U14837 ( .A(n12420), .B(n12450), .ZN(n12421) );
  AOI22_X1 U14838 ( .A1(n14128), .A2(n12463), .B1(n12462), .B2(n13843), .ZN(
        n12422) );
  XNOR2_X1 U14839 ( .A(n12421), .B(n12422), .ZN(n13797) );
  INV_X1 U14840 ( .A(n12421), .ZN(n12423) );
  NAND2_X1 U14841 ( .A1(n12423), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U14842 ( .A1(n14291), .A2(n6962), .ZN(n12426) );
  NAND2_X1 U14843 ( .A1(n12463), .A2(n14121), .ZN(n12425) );
  NAND2_X1 U14844 ( .A1(n12426), .A2(n12425), .ZN(n12427) );
  XNOR2_X1 U14845 ( .A(n12427), .B(n12450), .ZN(n12428) );
  AOI22_X1 U14846 ( .A1(n14291), .A2(n12463), .B1(n12462), .B2(n14121), .ZN(
        n12429) );
  XNOR2_X1 U14847 ( .A(n12428), .B(n12429), .ZN(n13720) );
  INV_X1 U14848 ( .A(n12428), .ZN(n12430) );
  NAND2_X1 U14849 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  NAND2_X1 U14850 ( .A1(n14097), .A2(n6962), .ZN(n12434) );
  NAND2_X1 U14851 ( .A1(n12463), .A2(n13842), .ZN(n12433) );
  NAND2_X1 U14852 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  XNOR2_X1 U14853 ( .A(n12435), .B(n12450), .ZN(n12436) );
  AOI22_X1 U14854 ( .A1(n14097), .A2(n12463), .B1(n12462), .B2(n13842), .ZN(
        n12437) );
  XNOR2_X1 U14855 ( .A(n12436), .B(n12437), .ZN(n13779) );
  INV_X1 U14856 ( .A(n12436), .ZN(n12438) );
  NAND2_X1 U14857 ( .A1(n12438), .A2(n12437), .ZN(n12439) );
  NAND2_X1 U14858 ( .A1(n14077), .A2(n6962), .ZN(n12442) );
  NAND2_X1 U14859 ( .A1(n12455), .A2(n13841), .ZN(n12441) );
  NAND2_X1 U14860 ( .A1(n12442), .A2(n12441), .ZN(n12443) );
  XNOR2_X1 U14861 ( .A(n12443), .B(n12450), .ZN(n12444) );
  AOI22_X1 U14862 ( .A1(n14077), .A2(n12463), .B1(n12462), .B2(n13841), .ZN(
        n12445) );
  XNOR2_X1 U14863 ( .A(n12444), .B(n12445), .ZN(n13747) );
  INV_X1 U14864 ( .A(n12444), .ZN(n12446) );
  NAND2_X1 U14865 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  NAND2_X1 U14866 ( .A1(n14275), .A2(n6962), .ZN(n12449) );
  NAND2_X1 U14867 ( .A1(n12463), .A2(n14033), .ZN(n12448) );
  NAND2_X1 U14868 ( .A1(n12449), .A2(n12448), .ZN(n12451) );
  XNOR2_X1 U14869 ( .A(n12451), .B(n12450), .ZN(n12452) );
  AOI22_X1 U14870 ( .A1(n14275), .A2(n12463), .B1(n12462), .B2(n14033), .ZN(
        n12453) );
  XNOR2_X1 U14871 ( .A(n12452), .B(n12453), .ZN(n13819) );
  INV_X1 U14872 ( .A(n12452), .ZN(n12454) );
  NAND2_X1 U14873 ( .A1(n14270), .A2(n6962), .ZN(n12457) );
  NAND2_X1 U14874 ( .A1(n12463), .A2(n13840), .ZN(n12456) );
  NAND2_X1 U14875 ( .A1(n12457), .A2(n12456), .ZN(n12458) );
  XNOR2_X1 U14876 ( .A(n12458), .B(n12450), .ZN(n12459) );
  AOI22_X1 U14877 ( .A1(n14270), .A2(n12463), .B1(n12462), .B2(n13840), .ZN(
        n12460) );
  XNOR2_X1 U14878 ( .A(n12459), .B(n12460), .ZN(n13704) );
  INV_X1 U14879 ( .A(n12459), .ZN(n12461) );
  AOI22_X1 U14880 ( .A1(n14265), .A2(n12463), .B1(n12462), .B2(n14034), .ZN(
        n12467) );
  AOI22_X1 U14881 ( .A1(n14265), .A2(n6962), .B1(n12463), .B2(n14034), .ZN(
        n12465) );
  XNOR2_X1 U14882 ( .A(n12465), .B(n12450), .ZN(n12466) );
  AOI22_X1 U14883 ( .A1(n13758), .A2(n13839), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12469) );
  NAND2_X1 U14884 ( .A1(n13799), .A2(n13840), .ZN(n12468) );
  OAI211_X1 U14885 ( .C1(n13832), .C2(n12470), .A(n12469), .B(n12468), .ZN(
        n12471) );
  AOI21_X1 U14886 ( .B1(n14265), .B2(n13834), .A(n12471), .ZN(n12472) );
  OAI21_X1 U14887 ( .B1(n12473), .B2(n13836), .A(n12472), .ZN(P1_U3220) );
  XNOR2_X1 U14888 ( .A(n12475), .B(n12474), .ZN(n12483) );
  INV_X1 U14889 ( .A(n12483), .ZN(n12476) );
  NAND2_X1 U14890 ( .A1(n12476), .A2(n14439), .ZN(n12487) );
  INV_X1 U14891 ( .A(n12477), .ZN(n12478) );
  NAND2_X1 U14892 ( .A1(n14444), .A2(n12921), .ZN(n12481) );
  AOI22_X1 U14893 ( .A1(n12479), .A2(n12913), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12480) );
  OAI211_X1 U14894 ( .C1(n12765), .C2(n12526), .A(n12481), .B(n12480), .ZN(
        n12485) );
  NOR4_X1 U14895 ( .A1(n12483), .A2(n12482), .A3(n12913), .A4(n14427), .ZN(
        n12484) );
  AOI211_X1 U14896 ( .C1(n14441), .C2(n12920), .A(n12485), .B(n12484), .ZN(
        n12486) );
  AOI21_X1 U14897 ( .B1(n12731), .B2(n12488), .A(n6604), .ZN(n12493) );
  AOI22_X1 U14898 ( .A1(n12767), .A2(n14416), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12490) );
  NAND2_X1 U14899 ( .A1(n14444), .A2(n12982), .ZN(n12489) );
  OAI211_X1 U14900 ( .C1(n13002), .C2(n14418), .A(n12490), .B(n12489), .ZN(
        n12491) );
  AOI21_X1 U14901 ( .B1(n12986), .B2(n14441), .A(n12491), .ZN(n12492) );
  OAI21_X1 U14902 ( .B1(n12493), .B2(n14427), .A(n12492), .ZN(P3_U3156) );
  XNOR2_X1 U14903 ( .A(n12495), .B(n12494), .ZN(n12500) );
  NAND2_X1 U14904 ( .A1(n14416), .A2(n13036), .ZN(n12496) );
  NAND2_X1 U14905 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12882)
         );
  OAI211_X1 U14906 ( .C1(n14418), .C2(n13065), .A(n12496), .B(n12882), .ZN(
        n12498) );
  NOR2_X1 U14907 ( .A1(n13184), .A2(n12574), .ZN(n12497) );
  AOI211_X1 U14908 ( .C1(n13043), .C2(n14444), .A(n12498), .B(n12497), .ZN(
        n12499) );
  OAI21_X1 U14909 ( .B1(n12500), .B2(n14427), .A(n12499), .ZN(P3_U3159) );
  AOI21_X1 U14910 ( .B1(n12502), .B2(n12501), .A(n6719), .ZN(n12507) );
  NAND2_X1 U14911 ( .A1(n14444), .A2(n13007), .ZN(n12504) );
  AOI22_X1 U14912 ( .A1(n14416), .A2(n12551), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12503) );
  OAI211_X1 U14913 ( .C1(n13003), .C2(n14418), .A(n12504), .B(n12503), .ZN(
        n12505) );
  AOI21_X1 U14914 ( .B1(n13006), .B2(n14441), .A(n12505), .ZN(n12506) );
  OAI21_X1 U14915 ( .B1(n12507), .B2(n14427), .A(n12506), .ZN(P3_U3163) );
  INV_X1 U14916 ( .A(n12961), .ZN(n12512) );
  OR2_X1 U14917 ( .A1(n12978), .A2(n15049), .ZN(n12509) );
  NAND2_X1 U14918 ( .A1(n12928), .A2(n15064), .ZN(n12508) );
  NAND2_X1 U14919 ( .A1(n12509), .A2(n12508), .ZN(n12954) );
  AOI22_X1 U14920 ( .A1(n12954), .A2(n12510), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12511) );
  OAI21_X1 U14921 ( .B1(n12512), .B2(n14433), .A(n12511), .ZN(n12520) );
  INV_X1 U14922 ( .A(n12514), .ZN(n12515) );
  NAND3_X1 U14923 ( .A1(n12513), .A2(n12516), .A3(n12515), .ZN(n12517) );
  AOI21_X1 U14924 ( .B1(n12518), .B2(n12517), .A(n14427), .ZN(n12519) );
  INV_X1 U14925 ( .A(n12521), .ZN(n13192) );
  AOI21_X1 U14926 ( .B1(n12523), .B2(n12522), .A(n14427), .ZN(n12525) );
  NAND2_X1 U14927 ( .A1(n12525), .A2(n12524), .ZN(n12530) );
  NOR2_X1 U14928 ( .A1(n14418), .A2(n13066), .ZN(n12528) );
  OAI22_X1 U14929 ( .A1(n12526), .A2(n13065), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8080), .ZN(n12527) );
  AOI211_X1 U14930 ( .C1(n13068), .C2(n14444), .A(n12528), .B(n12527), .ZN(
        n12529) );
  OAI211_X1 U14931 ( .C1(n13192), .C2(n12574), .A(n12530), .B(n12529), .ZN(
        P3_U3168) );
  INV_X1 U14932 ( .A(n12532), .ZN(n12534) );
  NOR3_X1 U14933 ( .A1(n6604), .A2(n12534), .A3(n12533), .ZN(n12536) );
  INV_X1 U14934 ( .A(n12513), .ZN(n12535) );
  OAI21_X1 U14935 ( .B1(n12536), .B2(n12535), .A(n14439), .ZN(n12540) );
  AOI22_X1 U14936 ( .A1(n12766), .A2(n15064), .B1(n15061), .B2(n12731), .ZN(
        n12966) );
  INV_X1 U14937 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12537) );
  OAI22_X1 U14938 ( .A1(n12966), .A2(n14446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12537), .ZN(n12538) );
  AOI21_X1 U14939 ( .B1(n12970), .B2(n14444), .A(n12538), .ZN(n12539) );
  OAI211_X1 U14940 ( .C1(n13165), .C2(n12574), .A(n12540), .B(n12539), .ZN(
        P3_U3169) );
  XNOR2_X1 U14941 ( .A(n12542), .B(n12541), .ZN(n12547) );
  NAND2_X1 U14942 ( .A1(n14444), .A2(n13022), .ZN(n12544) );
  AOI22_X1 U14943 ( .A1(n14416), .A2(n12768), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12543) );
  OAI211_X1 U14944 ( .C1(n13020), .C2(n14418), .A(n12544), .B(n12543), .ZN(
        n12545) );
  AOI21_X1 U14945 ( .B1(n13113), .B2(n14441), .A(n12545), .ZN(n12546) );
  OAI21_X1 U14946 ( .B1(n12547), .B2(n14427), .A(n12546), .ZN(P3_U3173) );
  INV_X1 U14947 ( .A(n12548), .ZN(n12549) );
  AOI21_X1 U14948 ( .B1(n12551), .B2(n12550), .A(n12549), .ZN(n12556) );
  AOI22_X1 U14949 ( .A1(n15064), .A2(n12731), .B1(n12768), .B2(n15061), .ZN(
        n12991) );
  OAI22_X1 U14950 ( .A1(n12991), .A2(n14446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12552), .ZN(n12554) );
  NOR2_X1 U14951 ( .A1(n13172), .A2(n12574), .ZN(n12553) );
  AOI211_X1 U14952 ( .C1(n12995), .C2(n14444), .A(n12554), .B(n12553), .ZN(
        n12555) );
  OAI21_X1 U14953 ( .B1(n12556), .B2(n14427), .A(n12555), .ZN(P3_U3175) );
  XNOR2_X1 U14954 ( .A(n12558), .B(n12557), .ZN(n12565) );
  NAND2_X1 U14955 ( .A1(n14444), .A2(n13057), .ZN(n12561) );
  NOR2_X1 U14956 ( .A1(n12559), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12862) );
  AOI21_X1 U14957 ( .B1(n14416), .B2(n13049), .A(n12862), .ZN(n12560) );
  OAI211_X1 U14958 ( .C1(n12562), .C2(n14418), .A(n12561), .B(n12560), .ZN(
        n12563) );
  AOI21_X1 U14959 ( .B1(n13056), .B2(n14441), .A(n12563), .ZN(n12564) );
  OAI21_X1 U14960 ( .B1(n12565), .B2(n14427), .A(n12564), .ZN(P3_U3178) );
  OAI21_X1 U14961 ( .B1(n12568), .B2(n12567), .A(n12566), .ZN(n12569) );
  INV_X1 U14962 ( .A(n12946), .ZN(n12572) );
  AOI22_X1 U14963 ( .A1(n12766), .A2(n15061), .B1(n15064), .B2(n12913), .ZN(
        n12944) );
  INV_X1 U14964 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12570) );
  OAI22_X1 U14965 ( .A1(n12944), .A2(n14446), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12570), .ZN(n12571) );
  AOI21_X1 U14966 ( .B1(n12572), .B2(n14444), .A(n12571), .ZN(n12573) );
  OAI21_X1 U14967 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(n15415), .A(n12575), 
        .ZN(n12576) );
  OAI21_X1 U14968 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(n12577), .A(n12576), 
        .ZN(n12579) );
  XNOR2_X1 U14969 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12578) );
  XNOR2_X1 U14970 ( .A(n12579), .B(n12578), .ZN(n13201) );
  INV_X1 U14971 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U14972 ( .A1(n12580), .A2(P3_REG2_REG_31__SCAN_IN), .B1(n7887), 
        .B2(P3_REG0_REG_31__SCAN_IN), .ZN(n12581) );
  OAI211_X1 U14973 ( .C1(n12584), .C2(n12583), .A(n12582), .B(n12581), .ZN(
        n12892) );
  INV_X1 U14974 ( .A(n12942), .ZN(n12741) );
  INV_X1 U14975 ( .A(n12624), .ZN(n12591) );
  INV_X1 U14976 ( .A(n13017), .ZN(n12721) );
  INV_X1 U14977 ( .A(n12592), .ZN(n12692) );
  NAND4_X1 U14978 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12652), .ZN(
        n12597) );
  NOR2_X1 U14979 ( .A1(n12597), .A2(n12596), .ZN(n12602) );
  INV_X1 U14980 ( .A(n12598), .ZN(n12669) );
  AND4_X1 U14981 ( .A1(n12600), .A2(n12645), .A3(n12599), .A4(n12665), .ZN(
        n12601) );
  NAND4_X1 U14982 ( .A1(n12602), .A2(n7373), .A3(n12669), .A4(n12601), .ZN(
        n12603) );
  NOR4_X1 U14983 ( .A1(n12676), .A2(n12604), .A3(n8019), .A4(n12603), .ZN(
        n12605) );
  NAND4_X1 U14984 ( .A1(n12606), .A2(n12692), .A3(n12698), .A4(n12605), .ZN(
        n12607) );
  NOR4_X1 U14985 ( .A1(n8122), .A2(n13055), .A3(n13061), .A4(n12607), .ZN(
        n12608) );
  NAND4_X1 U14986 ( .A1(n13005), .A2(n12993), .A3(n12721), .A4(n12608), .ZN(
        n12609) );
  NOR4_X1 U14987 ( .A1(n8200), .A2(n12976), .A3(n12968), .A4(n12609), .ZN(
        n12610) );
  INV_X1 U14988 ( .A(n12612), .ZN(n12752) );
  AND2_X1 U14989 ( .A1(n12615), .A2(n12614), .ZN(n12751) );
  INV_X1 U14990 ( .A(n12751), .ZN(n12616) );
  INV_X1 U14991 ( .A(n12896), .ZN(n13143) );
  NAND2_X1 U14992 ( .A1(n12620), .A2(n13143), .ZN(n12754) );
  OAI21_X1 U14993 ( .B1(n12617), .B2(n12616), .A(n12754), .ZN(n12618) );
  INV_X1 U14994 ( .A(n12620), .ZN(n12755) );
  OAI21_X1 U14995 ( .B1(n12622), .B2(n12750), .A(n12621), .ZN(n12749) );
  INV_X1 U14996 ( .A(n12986), .ZN(n13168) );
  MUX2_X1 U14997 ( .A(n12624), .B(n7009), .S(n12746), .Z(n12730) );
  INV_X1 U14998 ( .A(n12680), .ZN(n12625) );
  AOI21_X1 U14999 ( .B1(n14497), .B2(n12773), .A(n12625), .ZN(n12684) );
  AND2_X1 U15000 ( .A1(n12626), .A2(n12640), .ZN(n12644) );
  INV_X1 U15001 ( .A(n12638), .ZN(n12628) );
  NOR2_X1 U15002 ( .A1(n12628), .A2(n12627), .ZN(n12632) );
  OAI21_X1 U15003 ( .B1(n15060), .B2(n12630), .A(n12629), .ZN(n12631) );
  MUX2_X1 U15004 ( .A(n12632), .B(n12631), .S(n12750), .Z(n12633) );
  AOI21_X1 U15005 ( .B1(n12633), .B2(n12634), .A(n15047), .ZN(n12642) );
  AOI21_X1 U15006 ( .B1(n12647), .B2(n12635), .A(n12750), .ZN(n12641) );
  INV_X1 U15007 ( .A(n12634), .ZN(n12636) );
  NAND3_X1 U15008 ( .A1(n12636), .A2(n12635), .A3(n12647), .ZN(n12637) );
  MUX2_X1 U15009 ( .A(n12638), .B(n12637), .S(n12746), .Z(n12639) );
  OAI211_X1 U15010 ( .C1(n12642), .C2(n12641), .A(n12640), .B(n12639), .ZN(
        n12643) );
  OAI21_X1 U15011 ( .B1(n12746), .B2(n12644), .A(n12643), .ZN(n12646) );
  OAI211_X1 U15012 ( .C1(n12746), .C2(n12647), .A(n12646), .B(n12645), .ZN(
        n12653) );
  NAND3_X1 U15013 ( .A1(n12653), .A2(n12652), .A3(n12648), .ZN(n12650) );
  NAND3_X1 U15014 ( .A1(n12650), .A2(n12649), .A3(n12656), .ZN(n12658) );
  NAND3_X1 U15015 ( .A1(n12653), .A2(n12652), .A3(n12651), .ZN(n12655) );
  NAND3_X1 U15016 ( .A1(n12655), .A2(n12660), .A3(n12654), .ZN(n12657) );
  INV_X1 U15017 ( .A(n12661), .ZN(n15106) );
  NAND2_X1 U15018 ( .A1(n12777), .A2(n15106), .ZN(n12663) );
  MUX2_X1 U15019 ( .A(n12663), .B(n12662), .S(n12746), .Z(n12664) );
  MUX2_X1 U15020 ( .A(n12667), .B(n12666), .S(n12750), .Z(n12668) );
  NAND3_X1 U15021 ( .A1(n12670), .A2(n12669), .A3(n12668), .ZN(n12673) );
  MUX2_X1 U15022 ( .A(n12746), .B(n12775), .S(n15120), .Z(n12671) );
  OAI21_X1 U15023 ( .B1(n9159), .B2(n12750), .A(n12671), .ZN(n12672) );
  NAND3_X1 U15024 ( .A1(n12673), .A2(n7373), .A3(n12672), .ZN(n12678) );
  MUX2_X1 U15025 ( .A(n12675), .B(n12674), .S(n12750), .Z(n12677) );
  AOI21_X1 U15026 ( .B1(n12678), .B2(n12677), .A(n12676), .ZN(n12682) );
  AOI21_X1 U15027 ( .B1(n12687), .B2(n12679), .A(n12746), .ZN(n12681) );
  OAI21_X1 U15028 ( .B1(n12682), .B2(n12681), .A(n12680), .ZN(n12683) );
  OAI21_X1 U15029 ( .B1(n12684), .B2(n12750), .A(n12683), .ZN(n12686) );
  OAI211_X1 U15030 ( .C1(n12687), .C2(n12750), .A(n12686), .B(n12685), .ZN(
        n12693) );
  NAND3_X1 U15031 ( .A1(n12693), .A2(n12692), .A3(n12688), .ZN(n12690) );
  NAND3_X1 U15032 ( .A1(n12693), .A2(n12692), .A3(n12691), .ZN(n12695) );
  AOI21_X1 U15033 ( .B1(n12702), .B2(n12696), .A(n12746), .ZN(n12697) );
  INV_X1 U15034 ( .A(n12701), .ZN(n12699) );
  AOI21_X1 U15035 ( .B1(n12701), .B2(n12700), .A(n12750), .ZN(n12703) );
  OAI22_X1 U15036 ( .A1(n12704), .A2(n12703), .B1(n12750), .B2(n12702), .ZN(
        n12711) );
  INV_X1 U15037 ( .A(n12705), .ZN(n12710) );
  INV_X1 U15038 ( .A(n12706), .ZN(n12707) );
  OAI21_X1 U15039 ( .B1(n12708), .B2(n12707), .A(n12712), .ZN(n12709) );
  NAND3_X1 U15040 ( .A1(n12709), .A2(n12746), .A3(n12719), .ZN(n12715) );
  AOI22_X1 U15041 ( .A1(n12711), .A2(n7051), .B1(n12710), .B2(n12715), .ZN(
        n12718) );
  INV_X1 U15042 ( .A(n12712), .ZN(n12713) );
  NOR3_X1 U15043 ( .A1(n12714), .A2(n12746), .A3(n12713), .ZN(n12717) );
  INV_X1 U15044 ( .A(n12715), .ZN(n12716) );
  MUX2_X1 U15045 ( .A(n12719), .B(n13013), .S(n12746), .Z(n12720) );
  MUX2_X1 U15046 ( .A(n12723), .B(n12722), .S(n12746), .Z(n12724) );
  INV_X1 U15047 ( .A(n12725), .ZN(n12726) );
  MUX2_X1 U15048 ( .A(n12727), .B(n12726), .S(n12750), .Z(n12728) );
  OAI33_X1 U15049 ( .A1(n12750), .A2(n13168), .A3(n12731), .B1(n12976), .B2(
        n12730), .B3(n12729), .ZN(n12732) );
  INV_X1 U15050 ( .A(n12732), .ZN(n12733) );
  INV_X1 U15051 ( .A(n12734), .ZN(n12738) );
  AOI21_X1 U15052 ( .B1(n12736), .B2(n12735), .A(n12738), .ZN(n12737) );
  MUX2_X1 U15053 ( .A(n12738), .B(n12737), .S(n12750), .Z(n12742) );
  MUX2_X1 U15054 ( .A(n12739), .B(n12938), .S(n12750), .Z(n12740) );
  MUX2_X1 U15055 ( .A(n12744), .B(n12743), .S(n12750), .Z(n12745) );
  MUX2_X1 U15056 ( .A(n12750), .B(n12749), .S(n12748), .Z(n12753) );
  NOR3_X1 U15057 ( .A1(n12760), .A2(n12759), .A3(n15049), .ZN(n12763) );
  OAI21_X1 U15058 ( .B1(n12764), .B2(n12761), .A(P3_B_REG_SCAN_IN), .ZN(n12762) );
  MUX2_X1 U15059 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12892), .S(P3_U3897), .Z(
        P3_U3522) );
  INV_X1 U15060 ( .A(n12765), .ZN(n12914) );
  MUX2_X1 U15061 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12914), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15062 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12927), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15063 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12913), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15064 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12928), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15065 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12766), .S(n12783), .Z(
        P3_U3516) );
  MUX2_X1 U15066 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12767), .S(n12783), .Z(
        P3_U3515) );
  MUX2_X1 U15067 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12768), .S(n12783), .Z(
        P3_U3512) );
  MUX2_X1 U15068 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13035), .S(n12783), .Z(
        P3_U3509) );
  MUX2_X1 U15069 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13050), .S(n12783), .Z(
        P3_U3508) );
  MUX2_X1 U15070 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12769), .S(n12783), .Z(
        P3_U3507) );
  MUX2_X1 U15071 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n14415), .S(n12783), .Z(
        P3_U3506) );
  MUX2_X1 U15072 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12770), .S(n12783), .Z(
        P3_U3505) );
  MUX2_X1 U15073 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12771), .S(n12783), .Z(
        P3_U3504) );
  MUX2_X1 U15074 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12772), .S(n12783), .Z(
        P3_U3503) );
  MUX2_X1 U15075 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12773), .S(n12783), .Z(
        P3_U3502) );
  MUX2_X1 U15076 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12774), .S(n12783), .Z(
        P3_U3501) );
  MUX2_X1 U15077 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12775), .S(n12783), .Z(
        P3_U3500) );
  MUX2_X1 U15078 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12776), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15079 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12777), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15080 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12778), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15081 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12779), .S(n12783), .Z(
        P3_U3496) );
  MUX2_X1 U15082 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12780), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15083 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12781), .S(n12783), .Z(
        P3_U3494) );
  MUX2_X1 U15084 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12782), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15085 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15062), .S(n12783), .Z(
        P3_U3491) );
  NAND2_X1 U15086 ( .A1(n12787), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12822) );
  OAI21_X1 U15087 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12787), .A(n12822), 
        .ZN(n12806) );
  AOI21_X1 U15088 ( .B1(n12786), .B2(n12806), .A(n12821), .ZN(n12816) );
  INV_X1 U15089 ( .A(n14985), .ZN(n15021) );
  OR2_X1 U15090 ( .A1(n12787), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U15091 ( .A1(n12787), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12828) );
  AND2_X1 U15092 ( .A1(n12788), .A2(n12828), .ZN(n12804) );
  NAND2_X1 U15093 ( .A1(n12790), .A2(n12789), .ZN(n12792) );
  OAI21_X1 U15094 ( .B1(n12804), .B2(n12793), .A(n12827), .ZN(n12794) );
  INV_X1 U15095 ( .A(n12794), .ZN(n12797) );
  NOR2_X1 U15096 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12795), .ZN(n14414) );
  AOI21_X1 U15097 ( .B1(n14990), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n14414), 
        .ZN(n12796) );
  OAI21_X1 U15098 ( .B1(n14908), .B2(n12797), .A(n12796), .ZN(n12798) );
  AOI21_X1 U15099 ( .B1(n15021), .B2(n12799), .A(n12798), .ZN(n12815) );
  INV_X1 U15100 ( .A(n12800), .ZN(n12802) );
  AND2_X1 U15101 ( .A1(n12802), .A2(n12801), .ZN(n12809) );
  INV_X1 U15102 ( .A(n12809), .ZN(n12803) );
  NAND2_X1 U15103 ( .A1(n12812), .A2(n12803), .ZN(n12808) );
  INV_X1 U15104 ( .A(n12804), .ZN(n12807) );
  MUX2_X1 U15105 ( .A(n12807), .B(n12806), .S(n12805), .Z(n12810) );
  NAND2_X1 U15106 ( .A1(n12808), .A2(n12810), .ZN(n12813) );
  NOR2_X1 U15107 ( .A1(n12810), .A2(n12809), .ZN(n12811) );
  NAND2_X1 U15108 ( .A1(n12812), .A2(n12811), .ZN(n12818) );
  NAND3_X1 U15109 ( .A1(n12813), .A2(n15031), .A3(n12818), .ZN(n12814) );
  OAI211_X1 U15110 ( .C1(n12816), .C2(n15036), .A(n12815), .B(n12814), .ZN(
        P3_U3196) );
  MUX2_X1 U15111 ( .A(n12822), .B(n12828), .S(n6973), .Z(n12817) );
  NAND2_X1 U15112 ( .A1(n12818), .A2(n12817), .ZN(n12851) );
  XOR2_X1 U15113 ( .A(n12853), .B(n12851), .Z(n12820) );
  MUX2_X1 U15114 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6973), .Z(n12819) );
  NOR2_X1 U15115 ( .A1(n12820), .A2(n12819), .ZN(n12852) );
  AOI21_X1 U15116 ( .B1(n12820), .B2(n12819), .A(n12852), .ZN(n12837) );
  NOR2_X1 U15117 ( .A1(n6625), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n12826) );
  OAI21_X1 U15118 ( .B1(n12826), .B2(n12838), .A(n14474), .ZN(n12836) );
  NAND2_X1 U15119 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12829), .ZN(n12847) );
  OAI21_X1 U15120 ( .B1(n12829), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12847), 
        .ZN(n12830) );
  NAND2_X1 U15121 ( .A1(n15023), .A2(n12830), .ZN(n12833) );
  INV_X1 U15122 ( .A(n12831), .ZN(n12832) );
  OAI211_X1 U15123 ( .C1(n15281), .C2(n15041), .A(n12833), .B(n12832), .ZN(
        n12834) );
  AOI21_X1 U15124 ( .B1(n15021), .B2(n12853), .A(n12834), .ZN(n12835) );
  OAI211_X1 U15125 ( .C1(n12837), .C2(n15010), .A(n12836), .B(n12835), .ZN(
        P3_U3197) );
  NAND2_X1 U15126 ( .A1(n12845), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12840) );
  OAI21_X1 U15127 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12845), .A(n12840), 
        .ZN(n14459) );
  INV_X1 U15128 ( .A(n12840), .ZN(n12841) );
  INV_X1 U15129 ( .A(n12842), .ZN(n12843) );
  NAND2_X1 U15130 ( .A1(n6926), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12869) );
  OAI21_X1 U15131 ( .B1(n6926), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12869), .ZN(
        n12844) );
  AOI21_X1 U15132 ( .B1(n6638), .B2(n12844), .A(n12871), .ZN(n12868) );
  NAND2_X1 U15133 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12845), .ZN(n12849) );
  INV_X1 U15134 ( .A(n12845), .ZN(n14448) );
  INV_X1 U15135 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U15136 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12845), .B1(n14448), 
        .B2(n13134), .ZN(n14451) );
  NAND2_X1 U15137 ( .A1(n6753), .A2(n12846), .ZN(n12848) );
  AOI22_X1 U15138 ( .A1(n14467), .A2(P3_REG1_REG_17__SCAN_IN), .B1(n12850), 
        .B2(n12857), .ZN(n12886) );
  XOR2_X1 U15139 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12884), .Z(n12885) );
  XNOR2_X1 U15140 ( .A(n12886), .B(n12885), .ZN(n12866) );
  MUX2_X1 U15141 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6973), .Z(n12860) );
  MUX2_X1 U15142 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6973), .Z(n12858) );
  INV_X1 U15143 ( .A(n12851), .ZN(n12854) );
  MUX2_X1 U15144 ( .A(n12855), .B(n13134), .S(n6973), .Z(n12856) );
  NOR2_X1 U15145 ( .A1(n14448), .A2(n12856), .ZN(n14452) );
  NAND2_X1 U15146 ( .A1(n14448), .A2(n12856), .ZN(n14453) );
  OAI21_X1 U15147 ( .B1(n14456), .B2(n14452), .A(n14453), .ZN(n14469) );
  XOR2_X1 U15148 ( .A(n12858), .B(n14466), .Z(n14470) );
  NOR2_X1 U15149 ( .A1(n14469), .A2(n14470), .ZN(n14468) );
  NOR2_X1 U15150 ( .A1(n12859), .A2(n12860), .ZN(n12874) );
  AOI21_X1 U15151 ( .B1(n12860), .B2(n12859), .A(n12874), .ZN(n12864) );
  NOR2_X1 U15152 ( .A1(n14985), .A2(n6926), .ZN(n12861) );
  AOI211_X1 U15153 ( .C1(n14990), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n12862), 
        .B(n12861), .ZN(n12863) );
  OAI21_X1 U15154 ( .B1(n12864), .B2(n15010), .A(n12863), .ZN(n12865) );
  AOI21_X1 U15155 ( .B1(n15023), .B2(n12866), .A(n12865), .ZN(n12867) );
  OAI21_X1 U15156 ( .B1(n12868), .B2(n15036), .A(n12867), .ZN(P3_U3200) );
  INV_X1 U15157 ( .A(n12869), .ZN(n12870) );
  NOR2_X1 U15158 ( .A1(n12871), .A2(n12870), .ZN(n12873) );
  XNOR2_X1 U15159 ( .A(n12872), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12876) );
  XNOR2_X1 U15160 ( .A(n12873), .B(n12876), .ZN(n12891) );
  AOI21_X1 U15161 ( .B1(n12875), .B2(n12884), .A(n12874), .ZN(n12880) );
  INV_X1 U15162 ( .A(n12876), .ZN(n12878) );
  XNOR2_X1 U15163 ( .A(n12883), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12887) );
  MUX2_X1 U15164 ( .A(n12878), .B(n12887), .S(n6973), .Z(n12879) );
  XNOR2_X1 U15165 ( .A(n12880), .B(n12879), .ZN(n12890) );
  NAND2_X1 U15166 ( .A1(n14990), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12881) );
  OAI211_X1 U15167 ( .C1(n14985), .C2(n12883), .A(n12882), .B(n12881), .ZN(
        n12889) );
  INV_X1 U15168 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13126) );
  OAI22_X1 U15169 ( .A1(n12886), .A2(n12885), .B1(n12884), .B2(n13126), .ZN(
        n12888) );
  NOR2_X1 U15170 ( .A1(n15072), .A2(n12894), .ZN(n12903) );
  AOI21_X1 U15171 ( .B1(n15077), .B2(n13144), .A(n12903), .ZN(n12897) );
  NAND2_X1 U15172 ( .A1(n13011), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12895) );
  OAI211_X1 U15173 ( .C1(n12896), .C2(n13071), .A(n12897), .B(n12895), .ZN(
        P3_U3202) );
  NAND2_X1 U15174 ( .A1(n13147), .A2(n13026), .ZN(n12898) );
  OAI211_X1 U15175 ( .C1(n15077), .C2(n12899), .A(n12898), .B(n12897), .ZN(
        P3_U3203) );
  INV_X1 U15176 ( .A(n12900), .ZN(n12908) );
  NAND2_X1 U15177 ( .A1(n12901), .A2(n15077), .ZN(n12907) );
  NOR2_X1 U15178 ( .A1(n15077), .A2(n12902), .ZN(n12904) );
  AOI211_X1 U15179 ( .C1(n12905), .C2(n13026), .A(n12904), .B(n12903), .ZN(
        n12906) );
  OAI211_X1 U15180 ( .C1(n12908), .C2(n13029), .A(n12907), .B(n12906), .ZN(
        P3_U3204) );
  NAND2_X1 U15181 ( .A1(n12909), .A2(n12918), .ZN(n12910) );
  NAND2_X1 U15182 ( .A1(n12910), .A2(n15067), .ZN(n12911) );
  OR2_X1 U15183 ( .A1(n12912), .A2(n12911), .ZN(n12916) );
  AOI22_X1 U15184 ( .A1(n12914), .A2(n15064), .B1(n15061), .B2(n12913), .ZN(
        n12915) );
  XNOR2_X1 U15185 ( .A(n12919), .B(n12918), .ZN(n13081) );
  AOI22_X1 U15186 ( .A1(n13011), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n13069), 
        .B2(n12921), .ZN(n12922) );
  OAI21_X1 U15187 ( .B1(n13153), .B2(n13071), .A(n12922), .ZN(n12923) );
  AOI21_X1 U15188 ( .B1(n13081), .B2(n13073), .A(n12923), .ZN(n12924) );
  OAI21_X1 U15189 ( .B1(n6627), .B2(n13011), .A(n12924), .ZN(P3_U3205) );
  OAI21_X1 U15190 ( .B1(n12926), .B2(n12934), .A(n12925), .ZN(n12929) );
  AOI222_X1 U15191 ( .A1(n12929), .A2(n15067), .B1(n12928), .B2(n15061), .C1(
        n12927), .C2(n15064), .ZN(n13086) );
  INV_X1 U15192 ( .A(n12930), .ZN(n12931) );
  OAI22_X1 U15193 ( .A1(n15077), .A2(n12932), .B1(n12931), .B2(n15072), .ZN(
        n12936) );
  AOI21_X1 U15194 ( .B1(n12934), .B2(n12933), .A(n6695), .ZN(n13087) );
  NOR2_X1 U15195 ( .A1(n13087), .A2(n13029), .ZN(n12935) );
  AOI211_X1 U15196 ( .C1(n13026), .C2(n13084), .A(n12936), .B(n12935), .ZN(
        n12937) );
  OAI21_X1 U15197 ( .B1(n13086), .B2(n13011), .A(n12937), .ZN(P3_U3206) );
  NAND2_X1 U15198 ( .A1(n12957), .A2(n12938), .ZN(n12939) );
  NAND2_X1 U15199 ( .A1(n12939), .A2(n12942), .ZN(n12940) );
  INV_X1 U15200 ( .A(n13089), .ZN(n12952) );
  XNOR2_X1 U15201 ( .A(n12942), .B(n12943), .ZN(n12945) );
  OAI21_X1 U15202 ( .B1(n12945), .B2(n13063), .A(n12944), .ZN(n13088) );
  NAND2_X1 U15203 ( .A1(n13088), .A2(n15077), .ZN(n12951) );
  OAI22_X1 U15204 ( .A1(n15077), .A2(n12947), .B1(n12946), .B2(n15072), .ZN(
        n12948) );
  AOI21_X1 U15205 ( .B1(n12949), .B2(n13026), .A(n12948), .ZN(n12950) );
  OAI211_X1 U15206 ( .C1(n12952), .C2(n13029), .A(n12951), .B(n12950), .ZN(
        P3_U3207) );
  AOI21_X1 U15207 ( .B1(n12953), .B2(n12958), .A(n13063), .ZN(n12956) );
  AOI21_X1 U15208 ( .B1(n12956), .B2(n12955), .A(n12954), .ZN(n13094) );
  OAI21_X1 U15209 ( .B1(n12959), .B2(n12958), .A(n12957), .ZN(n13092) );
  INV_X1 U15210 ( .A(n12960), .ZN(n13161) );
  AOI22_X1 U15211 ( .A1(n13011), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13069), 
        .B2(n12961), .ZN(n12962) );
  OAI21_X1 U15212 ( .B1(n13161), .B2(n13071), .A(n12962), .ZN(n12963) );
  AOI21_X1 U15213 ( .B1(n13092), .B2(n13073), .A(n12963), .ZN(n12964) );
  OAI21_X1 U15214 ( .B1(n13094), .B2(n13011), .A(n12964), .ZN(P3_U3208) );
  XNOR2_X1 U15215 ( .A(n12965), .B(n12968), .ZN(n12967) );
  OAI21_X1 U15216 ( .B1(n12967), .B2(n13063), .A(n12966), .ZN(n13097) );
  INV_X1 U15217 ( .A(n13097), .ZN(n12974) );
  OAI21_X1 U15218 ( .B1(n6639), .B2(n7005), .A(n12969), .ZN(n13098) );
  AOI22_X1 U15219 ( .A1(n15079), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n13069), 
        .B2(n12970), .ZN(n12971) );
  OAI21_X1 U15220 ( .B1(n13165), .B2(n13071), .A(n12971), .ZN(n12972) );
  AOI21_X1 U15221 ( .B1(n13098), .B2(n13073), .A(n12972), .ZN(n12973) );
  OAI21_X1 U15222 ( .B1(n12974), .B2(n13011), .A(n12973), .ZN(P3_U3209) );
  XNOR2_X1 U15223 ( .A(n12975), .B(n12976), .ZN(n13102) );
  INV_X1 U15224 ( .A(n13102), .ZN(n12989) );
  XNOR2_X1 U15225 ( .A(n12977), .B(n12976), .ZN(n12981) );
  OAI22_X1 U15226 ( .A1(n12978), .A2(n15050), .B1(n13002), .B2(n15049), .ZN(
        n12979) );
  AOI21_X1 U15227 ( .B1(n13102), .B2(n15118), .A(n12979), .ZN(n12980) );
  OAI21_X1 U15228 ( .B1(n12981), .B2(n13063), .A(n12980), .ZN(n13101) );
  NAND2_X1 U15229 ( .A1(n13101), .A2(n15077), .ZN(n12988) );
  INV_X1 U15230 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12984) );
  INV_X1 U15231 ( .A(n12982), .ZN(n12983) );
  OAI22_X1 U15232 ( .A1(n15077), .A2(n12984), .B1(n12983), .B2(n15072), .ZN(
        n12985) );
  AOI21_X1 U15233 ( .B1(n12986), .B2(n13026), .A(n12985), .ZN(n12987) );
  OAI211_X1 U15234 ( .C1(n12989), .C2(n15074), .A(n12988), .B(n12987), .ZN(
        P3_U3210) );
  XNOR2_X1 U15235 ( .A(n12990), .B(n12993), .ZN(n12992) );
  OAI21_X1 U15236 ( .B1(n12992), .B2(n13063), .A(n12991), .ZN(n13105) );
  INV_X1 U15237 ( .A(n13105), .ZN(n12999) );
  XNOR2_X1 U15238 ( .A(n12994), .B(n12993), .ZN(n13106) );
  AOI22_X1 U15239 ( .A1(n15079), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13069), 
        .B2(n12995), .ZN(n12996) );
  OAI21_X1 U15240 ( .B1(n13172), .B2(n13071), .A(n12996), .ZN(n12997) );
  AOI21_X1 U15241 ( .B1(n13106), .B2(n13073), .A(n12997), .ZN(n12998) );
  OAI21_X1 U15242 ( .B1(n12999), .B2(n13011), .A(n12998), .ZN(P3_U3211) );
  XOR2_X1 U15243 ( .A(n13005), .B(n13000), .Z(n13001) );
  OAI222_X1 U15244 ( .A1(n15049), .A2(n13003), .B1(n15050), .B2(n13002), .C1(
        n13063), .C2(n13001), .ZN(n13109) );
  INV_X1 U15245 ( .A(n13109), .ZN(n13012) );
  XOR2_X1 U15246 ( .A(n13005), .B(n13004), .Z(n13110) );
  INV_X1 U15247 ( .A(n13006), .ZN(n13176) );
  AOI22_X1 U15248 ( .A1(n13011), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13069), 
        .B2(n13007), .ZN(n13008) );
  OAI21_X1 U15249 ( .B1(n13176), .B2(n13071), .A(n13008), .ZN(n13009) );
  AOI21_X1 U15250 ( .B1(n13110), .B2(n13073), .A(n13009), .ZN(n13010) );
  OAI21_X1 U15251 ( .B1(n13012), .B2(n13011), .A(n13010), .ZN(P3_U3212) );
  NAND2_X1 U15252 ( .A1(n13041), .A2(n13013), .ZN(n13014) );
  NAND2_X1 U15253 ( .A1(n13014), .A2(n13017), .ZN(n13016) );
  INV_X1 U15254 ( .A(n13115), .ZN(n13030) );
  XNOR2_X1 U15255 ( .A(n13018), .B(n13017), .ZN(n13019) );
  OAI222_X1 U15256 ( .A1(n15050), .A2(n13021), .B1(n15049), .B2(n13020), .C1(
        n13019), .C2(n13063), .ZN(n13114) );
  NAND2_X1 U15257 ( .A1(n13114), .A2(n15077), .ZN(n13028) );
  INV_X1 U15258 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13024) );
  INV_X1 U15259 ( .A(n13022), .ZN(n13023) );
  OAI22_X1 U15260 ( .A1(n15077), .A2(n13024), .B1(n13023), .B2(n15072), .ZN(
        n13025) );
  AOI21_X1 U15261 ( .B1(n13113), .B2(n13026), .A(n13025), .ZN(n13027) );
  OAI211_X1 U15262 ( .C1(n13030), .C2(n13029), .A(n13028), .B(n13027), .ZN(
        P3_U3213) );
  NAND2_X1 U15263 ( .A1(n13033), .A2(n13032), .ZN(n13034) );
  NAND3_X1 U15264 ( .A1(n13031), .A2(n15067), .A3(n13034), .ZN(n13038) );
  AOI22_X1 U15265 ( .A1(n13036), .A2(n15064), .B1(n15061), .B2(n13035), .ZN(
        n13037) );
  NAND2_X1 U15266 ( .A1(n13052), .A2(n13039), .ZN(n13040) );
  NAND2_X1 U15267 ( .A1(n13040), .A2(n8122), .ZN(n13042) );
  NAND2_X1 U15268 ( .A1(n13042), .A2(n13041), .ZN(n13118) );
  AOI22_X1 U15269 ( .A1(n15079), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13043), 
        .B2(n13069), .ZN(n13044) );
  OAI21_X1 U15270 ( .B1(n13184), .B2(n13071), .A(n13044), .ZN(n13045) );
  AOI21_X1 U15271 ( .B1(n13118), .B2(n13073), .A(n13045), .ZN(n13046) );
  OAI21_X1 U15272 ( .B1(n13120), .B2(n15079), .A(n13046), .ZN(P3_U3214) );
  OAI21_X1 U15273 ( .B1(n13048), .B2(n13055), .A(n13047), .ZN(n13051) );
  AOI222_X1 U15274 ( .A1(n15067), .A2(n13051), .B1(n13050), .B2(n15061), .C1(
        n13049), .C2(n15064), .ZN(n13123) );
  INV_X1 U15275 ( .A(n13052), .ZN(n13053) );
  AOI21_X1 U15276 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(n13125) );
  INV_X1 U15277 ( .A(n13056), .ZN(n13188) );
  AOI22_X1 U15278 ( .A1(n15079), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n13069), 
        .B2(n13057), .ZN(n13058) );
  OAI21_X1 U15279 ( .B1(n13188), .B2(n13071), .A(n13058), .ZN(n13059) );
  AOI21_X1 U15280 ( .B1(n13125), .B2(n13073), .A(n13059), .ZN(n13060) );
  OAI21_X1 U15281 ( .B1(n13123), .B2(n15079), .A(n13060), .ZN(P3_U3215) );
  XNOR2_X1 U15282 ( .A(n13062), .B(n13061), .ZN(n13064) );
  OAI222_X1 U15283 ( .A1(n15049), .A2(n13066), .B1(n15050), .B2(n13065), .C1(
        n13064), .C2(n13063), .ZN(n13128) );
  INV_X1 U15284 ( .A(n13128), .ZN(n13075) );
  XNOR2_X1 U15285 ( .A(n13067), .B(n7051), .ZN(n13129) );
  AOI22_X1 U15286 ( .A1(n13011), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13069), 
        .B2(n13068), .ZN(n13070) );
  OAI21_X1 U15287 ( .B1(n13192), .B2(n13071), .A(n13070), .ZN(n13072) );
  AOI21_X1 U15288 ( .B1(n13129), .B2(n13073), .A(n13072), .ZN(n13074) );
  OAI21_X1 U15289 ( .B1(n13075), .B2(n15079), .A(n13074), .ZN(P3_U3216) );
  INV_X1 U15290 ( .A(n13136), .ZN(n13077) );
  NAND2_X1 U15291 ( .A1(n13143), .A2(n13077), .ZN(n13076) );
  NAND2_X1 U15292 ( .A1(n15144), .A2(n13144), .ZN(n13078) );
  OAI211_X1 U15293 ( .C1(n15144), .C2(n12583), .A(n13076), .B(n13078), .ZN(
        P3_U3490) );
  INV_X1 U15294 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n13080) );
  NAND2_X1 U15295 ( .A1(n13147), .A2(n13077), .ZN(n13079) );
  OAI211_X1 U15296 ( .C1(n15144), .C2(n13080), .A(n13079), .B(n13078), .ZN(
        P3_U3489) );
  INV_X1 U15297 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13082) );
  MUX2_X1 U15298 ( .A(n13082), .B(n13151), .S(n15144), .Z(n13083) );
  OAI21_X1 U15299 ( .B1(n13153), .B2(n13136), .A(n13083), .ZN(P3_U3487) );
  NAND2_X1 U15300 ( .A1(n13084), .A2(n15105), .ZN(n13085) );
  OAI211_X1 U15301 ( .C1(n14498), .C2(n13087), .A(n13086), .B(n13085), .ZN(
        n13154) );
  MUX2_X1 U15302 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13154), .S(n15144), .Z(
        P3_U3486) );
  INV_X1 U15303 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13090) );
  AOI21_X1 U15304 ( .B1(n13089), .B2(n13138), .A(n13088), .ZN(n13155) );
  MUX2_X1 U15305 ( .A(n13090), .B(n13155), .S(n15144), .Z(n13091) );
  OAI21_X1 U15306 ( .B1(n13157), .B2(n13136), .A(n13091), .ZN(P3_U3485) );
  NAND2_X1 U15307 ( .A1(n13092), .A2(n13138), .ZN(n13093) );
  AND2_X1 U15308 ( .A1(n13094), .A2(n13093), .ZN(n13159) );
  INV_X1 U15309 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13095) );
  MUX2_X1 U15310 ( .A(n13159), .B(n13095), .S(n15141), .Z(n13096) );
  OAI21_X1 U15311 ( .B1(n13161), .B2(n13136), .A(n13096), .ZN(P3_U3484) );
  INV_X1 U15312 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13099) );
  AOI21_X1 U15313 ( .B1(n13138), .B2(n13098), .A(n13097), .ZN(n13162) );
  MUX2_X1 U15314 ( .A(n13099), .B(n13162), .S(n15144), .Z(n13100) );
  OAI21_X1 U15315 ( .B1(n13165), .B2(n13136), .A(n13100), .ZN(P3_U3483) );
  INV_X1 U15316 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13103) );
  AOI21_X1 U15317 ( .B1(n15129), .B2(n13102), .A(n13101), .ZN(n13166) );
  MUX2_X1 U15318 ( .A(n13103), .B(n13166), .S(n15144), .Z(n13104) );
  OAI21_X1 U15319 ( .B1(n13168), .B2(n13136), .A(n13104), .ZN(P3_U3482) );
  INV_X1 U15320 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13107) );
  AOI21_X1 U15321 ( .B1(n13106), .B2(n13138), .A(n13105), .ZN(n13169) );
  MUX2_X1 U15322 ( .A(n13107), .B(n13169), .S(n15144), .Z(n13108) );
  OAI21_X1 U15323 ( .B1(n13172), .B2(n13136), .A(n13108), .ZN(P3_U3481) );
  INV_X1 U15324 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13111) );
  AOI21_X1 U15325 ( .B1(n13110), .B2(n13138), .A(n13109), .ZN(n13173) );
  MUX2_X1 U15326 ( .A(n13111), .B(n13173), .S(n15144), .Z(n13112) );
  OAI21_X1 U15327 ( .B1(n13176), .B2(n13136), .A(n13112), .ZN(P3_U3480) );
  INV_X1 U15328 ( .A(n13113), .ZN(n13180) );
  INV_X1 U15329 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13116) );
  AOI21_X1 U15330 ( .B1(n13115), .B2(n13138), .A(n13114), .ZN(n13177) );
  MUX2_X1 U15331 ( .A(n13116), .B(n13177), .S(n15144), .Z(n13117) );
  OAI21_X1 U15332 ( .B1(n13180), .B2(n13136), .A(n13117), .ZN(P3_U3479) );
  NAND2_X1 U15333 ( .A1(n13118), .A2(n13138), .ZN(n13119) );
  NAND2_X1 U15334 ( .A1(n13120), .A2(n13119), .ZN(n13181) );
  MUX2_X1 U15335 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13181), .S(n15144), .Z(
        n13121) );
  INV_X1 U15336 ( .A(n13121), .ZN(n13122) );
  OAI21_X1 U15337 ( .B1(n13136), .B2(n13184), .A(n13122), .ZN(P3_U3478) );
  INV_X1 U15338 ( .A(n13123), .ZN(n13124) );
  AOI21_X1 U15339 ( .B1(n13125), .B2(n13138), .A(n13124), .ZN(n13185) );
  MUX2_X1 U15340 ( .A(n13126), .B(n13185), .S(n15144), .Z(n13127) );
  OAI21_X1 U15341 ( .B1(n13188), .B2(n13136), .A(n13127), .ZN(P3_U3477) );
  INV_X1 U15342 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13130) );
  AOI21_X1 U15343 ( .B1(n13129), .B2(n13138), .A(n13128), .ZN(n13189) );
  MUX2_X1 U15344 ( .A(n13130), .B(n13189), .S(n15144), .Z(n13131) );
  OAI21_X1 U15345 ( .B1(n13192), .B2(n13136), .A(n13131), .ZN(P3_U3476) );
  AOI21_X1 U15346 ( .B1(n13133), .B2(n13138), .A(n13132), .ZN(n13193) );
  MUX2_X1 U15347 ( .A(n13134), .B(n13193), .S(n15144), .Z(n13135) );
  OAI21_X1 U15348 ( .B1(n13197), .B2(n13136), .A(n13135), .ZN(P3_U3475) );
  AND2_X1 U15349 ( .A1(n13137), .A2(n15105), .ZN(n13141) );
  AND2_X1 U15350 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  OR3_X1 U15351 ( .A1(n13142), .A2(n13141), .A3(n13140), .ZN(n13198) );
  MUX2_X1 U15352 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13198), .S(n15144), .Z(
        P3_U3474) );
  INV_X1 U15353 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13146) );
  NAND2_X1 U15354 ( .A1(n13143), .A2(n7028), .ZN(n13145) );
  NAND2_X1 U15355 ( .A1(n15130), .A2(n13144), .ZN(n13148) );
  OAI211_X1 U15356 ( .C1(n15130), .C2(n13146), .A(n13145), .B(n13148), .ZN(
        P3_U3458) );
  INV_X1 U15357 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U15358 ( .A1(n13147), .A2(n7028), .ZN(n13149) );
  OAI211_X1 U15359 ( .C1(n15130), .C2(n13150), .A(n13149), .B(n13148), .ZN(
        P3_U3457) );
  MUX2_X1 U15360 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13154), .S(n15130), .Z(
        P3_U3454) );
  MUX2_X1 U15361 ( .A(n15254), .B(n13155), .S(n15130), .Z(n13156) );
  OAI21_X1 U15362 ( .B1(n13157), .B2(n13196), .A(n13156), .ZN(P3_U3453) );
  INV_X1 U15363 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13158) );
  MUX2_X1 U15364 ( .A(n13159), .B(n13158), .S(n8319), .Z(n13160) );
  OAI21_X1 U15365 ( .B1(n13161), .B2(n13196), .A(n13160), .ZN(P3_U3452) );
  INV_X1 U15366 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13163) );
  MUX2_X1 U15367 ( .A(n13163), .B(n13162), .S(n15130), .Z(n13164) );
  OAI21_X1 U15368 ( .B1(n13165), .B2(n13196), .A(n13164), .ZN(P3_U3451) );
  MUX2_X1 U15369 ( .A(n15364), .B(n13166), .S(n15130), .Z(n13167) );
  OAI21_X1 U15370 ( .B1(n13168), .B2(n13196), .A(n13167), .ZN(P3_U3450) );
  INV_X1 U15371 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13170) );
  MUX2_X1 U15372 ( .A(n13170), .B(n13169), .S(n15130), .Z(n13171) );
  OAI21_X1 U15373 ( .B1(n13172), .B2(n13196), .A(n13171), .ZN(P3_U3449) );
  INV_X1 U15374 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13174) );
  MUX2_X1 U15375 ( .A(n13174), .B(n13173), .S(n15130), .Z(n13175) );
  OAI21_X1 U15376 ( .B1(n13176), .B2(n13196), .A(n13175), .ZN(P3_U3448) );
  MUX2_X1 U15377 ( .A(n13178), .B(n13177), .S(n15130), .Z(n13179) );
  OAI21_X1 U15378 ( .B1(n13180), .B2(n13196), .A(n13179), .ZN(P3_U3447) );
  MUX2_X1 U15379 ( .A(n13181), .B(P3_REG0_REG_19__SCAN_IN), .S(n8319), .Z(
        n13182) );
  INV_X1 U15380 ( .A(n13182), .ZN(n13183) );
  OAI21_X1 U15381 ( .B1(n13196), .B2(n13184), .A(n13183), .ZN(P3_U3446) );
  MUX2_X1 U15382 ( .A(n13186), .B(n13185), .S(n15130), .Z(n13187) );
  OAI21_X1 U15383 ( .B1(n13188), .B2(n13196), .A(n13187), .ZN(P3_U3444) );
  MUX2_X1 U15384 ( .A(n13190), .B(n13189), .S(n15130), .Z(n13191) );
  OAI21_X1 U15385 ( .B1(n13192), .B2(n13196), .A(n13191), .ZN(P3_U3441) );
  MUX2_X1 U15386 ( .A(n13194), .B(n13193), .S(n15130), .Z(n13195) );
  OAI21_X1 U15387 ( .B1(n13197), .B2(n13196), .A(n13195), .ZN(P3_U3438) );
  MUX2_X1 U15388 ( .A(n13198), .B(P3_REG0_REG_15__SCAN_IN), .S(n8319), .Z(
        P3_U3435) );
  MUX2_X1 U15389 ( .A(n13199), .B(P3_D_REG_1__SCAN_IN), .S(n13200), .Z(
        P3_U3377) );
  MUX2_X1 U15390 ( .A(n9129), .B(P3_D_REG_0__SCAN_IN), .S(n13200), .Z(P3_U3376) );
  INV_X1 U15391 ( .A(n13201), .ZN(n13204) );
  NOR4_X1 U15392 ( .A1(n7395), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n8285), .ZN(n13202) );
  AOI21_X1 U15393 ( .B1(n14386), .B2(SI_31_), .A(n13202), .ZN(n13203) );
  OAI21_X1 U15394 ( .B1(n13204), .B2(n15458), .A(n13203), .ZN(P3_U3264) );
  INV_X1 U15395 ( .A(n13205), .ZN(n13208) );
  OAI222_X1 U15396 ( .A1(n15458), .A2(n13208), .B1(n13207), .B2(P3_U3151), 
        .C1(n13206), .C2(n15456), .ZN(P3_U3266) );
  NAND2_X1 U15397 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  NAND3_X1 U15398 ( .A1(n13212), .A2(n13278), .A3(n13211), .ZN(n13216) );
  AOI22_X1 U15399 ( .A1(n13282), .A2(n13448), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13215) );
  AOI22_X1 U15400 ( .A1(n13284), .A2(n13414), .B1(n13419), .B2(n13283), .ZN(
        n13214) );
  NAND2_X1 U15401 ( .A1(n13591), .A2(n13302), .ZN(n13213) );
  NAND4_X1 U15402 ( .A1(n13216), .A2(n13215), .A3(n13214), .A4(n13213), .ZN(
        P2_U3186) );
  OAI211_X1 U15403 ( .C1(n13219), .C2(n13218), .A(n13217), .B(n13278), .ZN(
        n13223) );
  AOI22_X1 U15404 ( .A1(n13282), .A2(n13502), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13222) );
  AOI22_X1 U15405 ( .A1(n13284), .A2(n13471), .B1(n13283), .B2(n13473), .ZN(
        n13221) );
  NAND2_X1 U15406 ( .A1(n13614), .A2(n13302), .ZN(n13220) );
  NAND4_X1 U15407 ( .A1(n13223), .A2(n13222), .A3(n13221), .A4(n13220), .ZN(
        P2_U3188) );
  NAND2_X1 U15408 ( .A1(n13225), .A2(n13224), .ZN(n13227) );
  XOR2_X1 U15409 ( .A(n13227), .B(n13226), .Z(n13231) );
  AOI22_X1 U15410 ( .A1(n13282), .A2(n13541), .B1(n13283), .B2(n13548), .ZN(
        n13228) );
  NAND2_X1 U15411 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13376)
         );
  OAI211_X1 U15412 ( .C1(n13299), .C2(n13236), .A(n13228), .B(n13376), .ZN(
        n13229) );
  AOI21_X1 U15413 ( .B1(n13640), .B2(n13302), .A(n13229), .ZN(n13230) );
  OAI21_X1 U15414 ( .B1(n13231), .B2(n13304), .A(n13230), .ZN(P2_U3191) );
  OAI211_X1 U15415 ( .C1(n13234), .C2(n13233), .A(n13232), .B(n13278), .ZN(
        n13241) );
  OAI22_X1 U15416 ( .A1(n13295), .A2(n13236), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13235), .ZN(n13239) );
  OAI22_X1 U15417 ( .A1(n13299), .A2(n13237), .B1(n13505), .B2(n13297), .ZN(
        n13238) );
  AOI211_X1 U15418 ( .C1(n13629), .C2(n13302), .A(n13239), .B(n13238), .ZN(
        n13240) );
  NAND2_X1 U15419 ( .A1(n13241), .A2(n13240), .ZN(P2_U3195) );
  OAI211_X1 U15420 ( .C1(n13244), .C2(n13243), .A(n13242), .B(n13278), .ZN(
        n13248) );
  AOI22_X1 U15421 ( .A1(n13282), .A2(n13471), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13247) );
  AOI22_X1 U15422 ( .A1(n13284), .A2(n13448), .B1(n13283), .B2(n13442), .ZN(
        n13246) );
  NAND2_X1 U15423 ( .A1(n13603), .A2(n13302), .ZN(n13245) );
  NAND4_X1 U15424 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        P2_U3197) );
  NAND2_X1 U15425 ( .A1(n13283), .A2(n13249), .ZN(n13251) );
  OAI211_X1 U15426 ( .C1(n13253), .C2(n13252), .A(n13251), .B(n13250), .ZN(
        n13260) );
  NAND3_X1 U15427 ( .A1(n13256), .A2(n13255), .A3(n13254), .ZN(n13258) );
  AOI21_X1 U15428 ( .B1(n13258), .B2(n13257), .A(n13304), .ZN(n13259) );
  AOI211_X1 U15429 ( .C1(n13651), .C2(n13302), .A(n13260), .B(n13259), .ZN(
        n13261) );
  INV_X1 U15430 ( .A(n13261), .ZN(P2_U3200) );
  OAI211_X1 U15431 ( .C1(n13264), .C2(n13263), .A(n13262), .B(n13278), .ZN(
        n13268) );
  AOI22_X1 U15432 ( .A1(n13282), .A2(n13484), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13267) );
  AOI22_X1 U15433 ( .A1(n13284), .A2(n13456), .B1(n13283), .B2(n13463), .ZN(
        n13266) );
  NAND2_X1 U15434 ( .A1(n13607), .A2(n13302), .ZN(n13265) );
  NAND4_X1 U15435 ( .A1(n13268), .A2(n13267), .A3(n13266), .A4(n13265), .ZN(
        P2_U3201) );
  AOI21_X1 U15436 ( .B1(n13271), .B2(n13270), .A(n13269), .ZN(n13277) );
  INV_X1 U15437 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13272) );
  OAI22_X1 U15438 ( .A1(n13295), .A2(n13521), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13272), .ZN(n13275) );
  INV_X1 U15439 ( .A(n13528), .ZN(n13273) );
  OAI22_X1 U15440 ( .A1(n13299), .A2(n13523), .B1(n13297), .B2(n13273), .ZN(
        n13274) );
  AOI211_X1 U15441 ( .C1(n13635), .C2(n13302), .A(n13275), .B(n13274), .ZN(
        n13276) );
  OAI21_X1 U15442 ( .B1(n13277), .B2(n13304), .A(n13276), .ZN(P2_U3205) );
  OAI211_X1 U15443 ( .C1(n13281), .C2(n13280), .A(n13279), .B(n13278), .ZN(
        n13288) );
  AOI22_X1 U15444 ( .A1(n13282), .A2(n13485), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13287) );
  AOI22_X1 U15445 ( .A1(n13284), .A2(n13484), .B1(n13491), .B2(n13283), .ZN(
        n13286) );
  NAND2_X1 U15446 ( .A1(n13621), .A2(n13302), .ZN(n13285) );
  NAND4_X1 U15447 ( .A1(n13288), .A2(n13287), .A3(n13286), .A4(n13285), .ZN(
        P2_U3207) );
  INV_X1 U15448 ( .A(n6977), .ZN(n13290) );
  AOI21_X1 U15449 ( .B1(n13292), .B2(n13291), .A(n13290), .ZN(n13305) );
  OAI22_X1 U15450 ( .A1(n13295), .A2(n13294), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13293), .ZN(n13301) );
  INV_X1 U15451 ( .A(n13434), .ZN(n13296) );
  OAI22_X1 U15452 ( .A1(n13299), .A2(n13298), .B1(n13297), .B2(n13296), .ZN(
        n13300) );
  AOI211_X1 U15453 ( .C1(n13598), .C2(n13302), .A(n13301), .B(n13300), .ZN(
        n13303) );
  OAI21_X1 U15454 ( .B1(n13305), .B2(n13304), .A(n13303), .ZN(P2_U3212) );
  INV_X2 U15455 ( .A(P2_U3947), .ZN(n13324) );
  MUX2_X1 U15456 ( .A(n13378), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13324), .Z(
        P2_U3562) );
  MUX2_X1 U15457 ( .A(n13306), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13324), .Z(
        P2_U3561) );
  MUX2_X1 U15458 ( .A(n13392), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13324), .Z(
        P2_U3560) );
  MUX2_X1 U15459 ( .A(n13414), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13324), .Z(
        P2_U3559) );
  MUX2_X1 U15460 ( .A(n13428), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13324), .Z(
        P2_U3558) );
  MUX2_X1 U15461 ( .A(n13448), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13324), .Z(
        P2_U3557) );
  MUX2_X1 U15462 ( .A(n13456), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13324), .Z(
        P2_U3556) );
  MUX2_X1 U15463 ( .A(n13471), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13324), .Z(
        P2_U3555) );
  MUX2_X1 U15464 ( .A(n13484), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13324), .Z(
        P2_U3554) );
  MUX2_X1 U15465 ( .A(n13502), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13324), .Z(
        P2_U3553) );
  MUX2_X1 U15466 ( .A(n13485), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13324), .Z(
        P2_U3552) );
  MUX2_X1 U15467 ( .A(n13539), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13324), .Z(
        P2_U3551) );
  MUX2_X1 U15468 ( .A(n13307), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13324), .Z(
        P2_U3550) );
  MUX2_X1 U15469 ( .A(n13541), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13324), .Z(
        P2_U3549) );
  MUX2_X1 U15470 ( .A(n13308), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13324), .Z(
        P2_U3548) );
  MUX2_X1 U15471 ( .A(n13309), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13324), .Z(
        P2_U3547) );
  MUX2_X1 U15472 ( .A(n13310), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13324), .Z(
        P2_U3546) );
  MUX2_X1 U15473 ( .A(n13311), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13324), .Z(
        P2_U3545) );
  MUX2_X1 U15474 ( .A(n13312), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13324), .Z(
        P2_U3544) );
  MUX2_X1 U15475 ( .A(n13313), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13324), .Z(
        P2_U3543) );
  MUX2_X1 U15476 ( .A(n13314), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13324), .Z(
        P2_U3542) );
  MUX2_X1 U15477 ( .A(n13315), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13324), .Z(
        P2_U3541) );
  MUX2_X1 U15478 ( .A(n13316), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13324), .Z(
        P2_U3540) );
  MUX2_X1 U15479 ( .A(n13317), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13324), .Z(
        P2_U3539) );
  MUX2_X1 U15480 ( .A(n13318), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13324), .Z(
        P2_U3538) );
  MUX2_X1 U15481 ( .A(n13319), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13324), .Z(
        P2_U3537) );
  MUX2_X1 U15482 ( .A(n13320), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13324), .Z(
        P2_U3536) );
  MUX2_X1 U15483 ( .A(n13321), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13324), .Z(
        P2_U3535) );
  MUX2_X1 U15484 ( .A(n13322), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13324), .Z(
        P2_U3534) );
  MUX2_X1 U15485 ( .A(n13323), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13324), .Z(
        P2_U3533) );
  MUX2_X1 U15486 ( .A(n13325), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13324), .Z(
        P2_U3532) );
  INV_X1 U15487 ( .A(n14795), .ZN(n13328) );
  INV_X1 U15488 ( .A(n14788), .ZN(n14767) );
  OAI21_X1 U15489 ( .B1(n14767), .B2(n9051), .A(n13326), .ZN(n13327) );
  AOI21_X1 U15490 ( .B1(n13335), .B2(n13328), .A(n13327), .ZN(n13343) );
  INV_X1 U15491 ( .A(n13329), .ZN(n13331) );
  MUX2_X1 U15492 ( .A(n10790), .B(P2_REG2_REG_3__SCAN_IN), .S(n13335), .Z(
        n13330) );
  NAND2_X1 U15493 ( .A1(n13331), .A2(n13330), .ZN(n13333) );
  OAI211_X1 U15494 ( .C1(n13334), .C2(n13333), .A(n14790), .B(n13332), .ZN(
        n13342) );
  MUX2_X1 U15495 ( .A(n10153), .B(P2_REG1_REG_3__SCAN_IN), .S(n13335), .Z(
        n13336) );
  NAND3_X1 U15496 ( .A1(n13338), .A2(n13337), .A3(n13336), .ZN(n13339) );
  NAND3_X1 U15497 ( .A1(n14782), .A2(n13340), .A3(n13339), .ZN(n13341) );
  NAND3_X1 U15498 ( .A1(n13343), .A2(n13342), .A3(n13341), .ZN(P2_U3217) );
  NAND2_X1 U15499 ( .A1(n13344), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13346) );
  NAND2_X1 U15500 ( .A1(n13346), .A2(n13345), .ZN(n13359) );
  AOI21_X1 U15501 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13347), .A(n13360), 
        .ZN(n13358) );
  NAND2_X1 U15502 ( .A1(n14788), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n13349) );
  OAI211_X1 U15503 ( .C1(n13350), .C2(n14795), .A(n13349), .B(n13348), .ZN(
        n13351) );
  INV_X1 U15504 ( .A(n13351), .ZN(n13357) );
  OAI21_X1 U15505 ( .B1(n13354), .B2(n13353), .A(n13352), .ZN(n13363) );
  XOR2_X1 U15506 ( .A(n13363), .B(n13364), .Z(n13355) );
  NAND2_X1 U15507 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n13355), .ZN(n13366) );
  OAI211_X1 U15508 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13355), .A(n14782), 
        .B(n13366), .ZN(n13356) );
  OAI211_X1 U15509 ( .C1(n13358), .C2(n14744), .A(n13357), .B(n13356), .ZN(
        P2_U3232) );
  NOR2_X1 U15510 ( .A1(n13364), .A2(n13359), .ZN(n13361) );
  NOR2_X1 U15511 ( .A1(n13361), .A2(n13360), .ZN(n13362) );
  NAND2_X1 U15512 ( .A1(n13364), .A2(n13363), .ZN(n13365) );
  NAND2_X1 U15513 ( .A1(n13366), .A2(n13365), .ZN(n13367) );
  XNOR2_X1 U15514 ( .A(n13367), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U15515 ( .A1(n13371), .A2(n14782), .ZN(n13368) );
  OAI211_X1 U15516 ( .C1(n13369), .C2(n14744), .A(n14795), .B(n13368), .ZN(
        n13375) );
  OAI22_X1 U15517 ( .A1(n13372), .A2(n14744), .B1(n13371), .B2(n13370), .ZN(
        n13374) );
  XNOR2_X1 U15518 ( .A(n13384), .B(n9921), .ZN(n13377) );
  NAND2_X1 U15519 ( .A1(n13377), .A2(n11860), .ZN(n13577) );
  NAND2_X1 U15520 ( .A1(n13379), .A2(n13378), .ZN(n13579) );
  NOR2_X1 U15521 ( .A1(n14809), .A2(n13579), .ZN(n13388) );
  INV_X1 U15522 ( .A(n9921), .ZN(n13578) );
  NOR2_X1 U15523 ( .A1(n13578), .A2(n14803), .ZN(n13380) );
  AOI211_X1 U15524 ( .C1(n14809), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13388), 
        .B(n13380), .ZN(n13381) );
  OAI21_X1 U15525 ( .B1(n13494), .B2(n13577), .A(n13381), .ZN(P2_U3234) );
  INV_X1 U15526 ( .A(n13383), .ZN(n13386) );
  OAI211_X1 U15527 ( .C1(n13581), .C2(n13386), .A(n13385), .B(n11860), .ZN(
        n13580) );
  NOR2_X1 U15528 ( .A1(n13581), .A2(n14803), .ZN(n13387) );
  AOI211_X1 U15529 ( .C1(n14809), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13388), 
        .B(n13387), .ZN(n13389) );
  OAI21_X1 U15530 ( .B1(n13494), .B2(n13580), .A(n13389), .ZN(P2_U3235) );
  INV_X1 U15531 ( .A(n13418), .ZN(n13390) );
  AOI21_X1 U15532 ( .B1(n13586), .B2(n13390), .A(n6569), .ZN(n13397) );
  OAI21_X1 U15533 ( .B1(n13391), .B2(n7288), .A(n13569), .ZN(n13395) );
  AOI22_X1 U15534 ( .A1(n13538), .A2(n13392), .B1(n13428), .B2(n13540), .ZN(
        n13393) );
  INV_X1 U15535 ( .A(n13589), .ZN(n13403) );
  NAND2_X1 U15536 ( .A1(n13403), .A2(n13402), .ZN(n13406) );
  AOI21_X1 U15537 ( .B1(n13404), .B2(n13562), .A(n14797), .ZN(n13405) );
  AOI21_X1 U15538 ( .B1(n13588), .B2(n13406), .A(n13405), .ZN(n13412) );
  AOI22_X1 U15539 ( .A1(n14809), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n14800), 
        .B2(n13407), .ZN(n13409) );
  NAND2_X1 U15540 ( .A1(n13586), .A2(n13547), .ZN(n13408) );
  OAI211_X1 U15541 ( .C1(n13589), .C2(n13410), .A(n13409), .B(n13408), .ZN(
        n13411) );
  OR2_X1 U15542 ( .A1(n13412), .A2(n13411), .ZN(P2_U3237) );
  XNOR2_X1 U15543 ( .A(n13413), .B(n13423), .ZN(n13415) );
  AOI222_X1 U15544 ( .A1(n13569), .A2(n13415), .B1(n13448), .B2(n13540), .C1(
        n13414), .C2(n13538), .ZN(n13596) );
  NAND2_X1 U15545 ( .A1(n13591), .A2(n13432), .ZN(n13416) );
  NAND2_X1 U15546 ( .A1(n13416), .A2(n11860), .ZN(n13417) );
  NOR2_X1 U15547 ( .A1(n13418), .A2(n13417), .ZN(n13590) );
  NAND2_X1 U15548 ( .A1(n13591), .A2(n13547), .ZN(n13421) );
  AOI22_X1 U15549 ( .A1(n14809), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n14800), 
        .B2(n13419), .ZN(n13420) );
  NAND2_X1 U15550 ( .A1(n13421), .A2(n13420), .ZN(n13422) );
  AOI21_X1 U15551 ( .B1(n13590), .B2(n14797), .A(n13422), .ZN(n13426) );
  NAND2_X1 U15552 ( .A1(n13424), .A2(n13423), .ZN(n13592) );
  NAND3_X1 U15553 ( .A1(n13593), .A2(n13592), .A3(n14806), .ZN(n13425) );
  OAI211_X1 U15554 ( .C1(n13596), .C2(n14809), .A(n13426), .B(n13425), .ZN(
        P2_U3238) );
  XOR2_X1 U15555 ( .A(n13431), .B(n13427), .Z(n13429) );
  AOI222_X1 U15556 ( .A1(n13569), .A2(n13429), .B1(n13428), .B2(n13538), .C1(
        n13456), .C2(n13540), .ZN(n13600) );
  XOR2_X1 U15557 ( .A(n13430), .B(n13431), .Z(n13601) );
  INV_X1 U15558 ( .A(n13601), .ZN(n13438) );
  AOI21_X1 U15559 ( .B1(n13598), .B2(n13441), .A(n8811), .ZN(n13433) );
  AND2_X1 U15560 ( .A1(n13433), .A2(n13432), .ZN(n13597) );
  NAND2_X1 U15561 ( .A1(n13597), .A2(n14797), .ZN(n13436) );
  AOI22_X1 U15562 ( .A1(n13469), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14800), 
        .B2(n13434), .ZN(n13435) );
  OAI211_X1 U15563 ( .C1(n7122), .C2(n14803), .A(n13436), .B(n13435), .ZN(
        n13437) );
  AOI21_X1 U15564 ( .B1(n13438), .B2(n14806), .A(n13437), .ZN(n13439) );
  OAI21_X1 U15565 ( .B1(n13600), .B2(n13469), .A(n13439), .ZN(P2_U3239) );
  XNOR2_X1 U15566 ( .A(n13440), .B(n13446), .ZN(n13606) );
  AOI211_X1 U15567 ( .C1(n13603), .C2(n13461), .A(n8811), .B(n7123), .ZN(
        n13602) );
  INV_X1 U15568 ( .A(n13603), .ZN(n13444) );
  AOI22_X1 U15569 ( .A1(n13469), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n14800), 
        .B2(n13442), .ZN(n13443) );
  OAI21_X1 U15570 ( .B1(n13444), .B2(n14803), .A(n13443), .ZN(n13451) );
  NAND3_X1 U15571 ( .A1(n13453), .A2(n13446), .A3(n13445), .ZN(n13447) );
  NAND2_X1 U15572 ( .A1(n6665), .A2(n13447), .ZN(n13449) );
  AOI222_X1 U15573 ( .A1(n13569), .A2(n13449), .B1(n13448), .B2(n13538), .C1(
        n13471), .C2(n13540), .ZN(n13605) );
  NOR2_X1 U15574 ( .A1(n13605), .A2(n13469), .ZN(n13450) );
  AOI211_X1 U15575 ( .C1(n13602), .C2(n14797), .A(n13451), .B(n13450), .ZN(
        n13452) );
  OAI21_X1 U15576 ( .B1(n13606), .B2(n13576), .A(n13452), .ZN(P2_U3240) );
  OAI21_X1 U15577 ( .B1(n13455), .B2(n13454), .A(n13453), .ZN(n13457) );
  AOI222_X1 U15578 ( .A1(n13569), .A2(n13457), .B1(n13456), .B2(n13538), .C1(
        n13484), .C2(n13540), .ZN(n13612) );
  OAI21_X1 U15579 ( .B1(n13460), .B2(n13459), .A(n13458), .ZN(n13608) );
  INV_X1 U15580 ( .A(n13608), .ZN(n13467) );
  OAI211_X1 U15581 ( .C1(n6573), .C2(n13462), .A(n11860), .B(n13461), .ZN(
        n13609) );
  AOI22_X1 U15582 ( .A1(n14809), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n14800), 
        .B2(n13463), .ZN(n13465) );
  NAND2_X1 U15583 ( .A1(n13607), .A2(n13547), .ZN(n13464) );
  OAI211_X1 U15584 ( .C1(n13609), .C2(n13494), .A(n13465), .B(n13464), .ZN(
        n13466) );
  AOI21_X1 U15585 ( .B1(n13467), .B2(n14806), .A(n13466), .ZN(n13468) );
  OAI21_X1 U15586 ( .B1(n13612), .B2(n13469), .A(n13468), .ZN(P2_U3241) );
  XOR2_X1 U15587 ( .A(n13470), .B(n13478), .Z(n13472) );
  AOI222_X1 U15588 ( .A1(n13569), .A2(n13472), .B1(n13471), .B2(n13538), .C1(
        n13502), .C2(n13540), .ZN(n13616) );
  AOI211_X1 U15589 ( .C1(n13614), .C2(n13489), .A(n8811), .B(n6573), .ZN(
        n13613) );
  AOI22_X1 U15590 ( .A1(n13469), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14800), 
        .B2(n13473), .ZN(n13474) );
  OAI21_X1 U15591 ( .B1(n13475), .B2(n14803), .A(n13474), .ZN(n13480) );
  AOI21_X1 U15592 ( .B1(n13478), .B2(n13477), .A(n13476), .ZN(n13617) );
  NOR2_X1 U15593 ( .A1(n13617), .A2(n13576), .ZN(n13479) );
  AOI211_X1 U15594 ( .C1(n13613), .C2(n14797), .A(n13480), .B(n13479), .ZN(
        n13481) );
  OAI21_X1 U15595 ( .B1(n14809), .B2(n13616), .A(n13481), .ZN(P2_U3242) );
  XNOR2_X1 U15596 ( .A(n13482), .B(n13495), .ZN(n13483) );
  NAND2_X1 U15597 ( .A1(n13483), .A2(n13569), .ZN(n13487) );
  AOI22_X1 U15598 ( .A1(n13485), .A2(n13540), .B1(n13538), .B2(n13484), .ZN(
        n13486) );
  NAND2_X1 U15599 ( .A1(n13487), .A2(n13486), .ZN(n13626) );
  AOI21_X1 U15600 ( .B1(n13621), .B2(n13488), .A(n6569), .ZN(n13490) );
  NAND2_X1 U15601 ( .A1(n13490), .A2(n13489), .ZN(n13622) );
  AOI22_X1 U15602 ( .A1(n13469), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14800), 
        .B2(n13491), .ZN(n13493) );
  NAND2_X1 U15603 ( .A1(n13621), .A2(n13547), .ZN(n13492) );
  OAI211_X1 U15604 ( .C1(n13622), .C2(n13494), .A(n13493), .B(n13492), .ZN(
        n13498) );
  NAND2_X1 U15605 ( .A1(n13496), .A2(n13495), .ZN(n13619) );
  AND3_X1 U15606 ( .A1(n13620), .A2(n14806), .A3(n13619), .ZN(n13497) );
  AOI211_X1 U15607 ( .C1(n13562), .C2(n13626), .A(n13498), .B(n13497), .ZN(
        n13499) );
  INV_X1 U15608 ( .A(n13499), .ZN(P2_U3243) );
  OR2_X1 U15609 ( .A1(n13517), .A2(n13518), .ZN(n13515) );
  NAND2_X1 U15610 ( .A1(n13515), .A2(n13500), .ZN(n13501) );
  XOR2_X1 U15611 ( .A(n13509), .B(n13501), .Z(n13503) );
  AOI222_X1 U15612 ( .A1(n13569), .A2(n13503), .B1(n13539), .B2(n13540), .C1(
        n13502), .C2(n13538), .ZN(n13631) );
  XNOR2_X1 U15613 ( .A(n13508), .B(n6710), .ZN(n13504) );
  NOR2_X1 U15614 ( .A1(n13504), .A2(n6569), .ZN(n13628) );
  INV_X1 U15615 ( .A(n13505), .ZN(n13506) );
  AOI22_X1 U15616 ( .A1(n13506), .A2(n14800), .B1(n14809), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13507) );
  OAI21_X1 U15617 ( .B1(n13508), .B2(n14803), .A(n13507), .ZN(n13512) );
  XOR2_X1 U15618 ( .A(n13510), .B(n13509), .Z(n13632) );
  NOR2_X1 U15619 ( .A1(n13632), .A2(n13576), .ZN(n13511) );
  AOI211_X1 U15620 ( .C1(n13628), .C2(n14797), .A(n13512), .B(n13511), .ZN(
        n13513) );
  OAI21_X1 U15621 ( .B1(n14809), .B2(n13631), .A(n13513), .ZN(P2_U3244) );
  XOR2_X1 U15622 ( .A(n13514), .B(n13518), .Z(n13637) );
  INV_X1 U15623 ( .A(n13515), .ZN(n13516) );
  AOI21_X1 U15624 ( .B1(n13518), .B2(n13517), .A(n13516), .ZN(n13519) );
  OAI222_X1 U15625 ( .A1(n13524), .A2(n13523), .B1(n13522), .B2(n13521), .C1(
        n13520), .C2(n13519), .ZN(n13633) );
  INV_X1 U15626 ( .A(n13635), .ZN(n13531) );
  NAND2_X1 U15627 ( .A1(n13635), .A2(n13545), .ZN(n13526) );
  NAND2_X1 U15628 ( .A1(n13526), .A2(n11860), .ZN(n13527) );
  NOR2_X1 U15629 ( .A1(n6710), .A2(n13527), .ZN(n13634) );
  NAND2_X1 U15630 ( .A1(n13634), .A2(n14797), .ZN(n13530) );
  AOI22_X1 U15631 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(n13469), .B1(n13528), 
        .B2(n14800), .ZN(n13529) );
  OAI211_X1 U15632 ( .C1(n13531), .C2(n14803), .A(n13530), .B(n13529), .ZN(
        n13532) );
  AOI21_X1 U15633 ( .B1(n13633), .B2(n13562), .A(n13532), .ZN(n13533) );
  OAI21_X1 U15634 ( .B1(n13637), .B2(n13576), .A(n13533), .ZN(P2_U3245) );
  XNOR2_X1 U15635 ( .A(n13534), .B(n13535), .ZN(n13643) );
  XOR2_X1 U15636 ( .A(n13536), .B(n13535), .Z(n13537) );
  NAND2_X1 U15637 ( .A1(n13537), .A2(n13569), .ZN(n13641) );
  INV_X1 U15638 ( .A(n13641), .ZN(n13544) );
  NAND2_X1 U15639 ( .A1(n13539), .A2(n13538), .ZN(n13543) );
  NAND2_X1 U15640 ( .A1(n13541), .A2(n13540), .ZN(n13542) );
  NAND2_X1 U15641 ( .A1(n13543), .A2(n13542), .ZN(n13639) );
  OAI21_X1 U15642 ( .B1(n13544), .B2(n13639), .A(n13562), .ZN(n13553) );
  AOI21_X1 U15643 ( .B1(n13640), .B2(n13558), .A(n6569), .ZN(n13546) );
  AND2_X1 U15644 ( .A1(n13546), .A2(n13545), .ZN(n13638) );
  NAND2_X1 U15645 ( .A1(n13640), .A2(n13547), .ZN(n13550) );
  AOI22_X1 U15646 ( .A1(n14809), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14800), 
        .B2(n13548), .ZN(n13549) );
  NAND2_X1 U15647 ( .A1(n13550), .A2(n13549), .ZN(n13551) );
  AOI21_X1 U15648 ( .B1(n13638), .B2(n14797), .A(n13551), .ZN(n13552) );
  OAI211_X1 U15649 ( .C1(n13643), .C2(n13576), .A(n13553), .B(n13552), .ZN(
        P2_U3246) );
  INV_X1 U15650 ( .A(n13554), .ZN(n13555) );
  AOI21_X1 U15651 ( .B1(n13565), .B2(n13556), .A(n13555), .ZN(n13648) );
  INV_X1 U15652 ( .A(n13557), .ZN(n13560) );
  INV_X1 U15653 ( .A(n13558), .ZN(n13559) );
  AOI211_X1 U15654 ( .C1(n13645), .C2(n13560), .A(n6569), .B(n13559), .ZN(
        n13644) );
  INV_X1 U15655 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13561) );
  OAI22_X1 U15656 ( .A1(n13563), .A2(n14803), .B1(n13562), .B2(n13561), .ZN(
        n13564) );
  AOI21_X1 U15657 ( .B1(n13644), .B2(n14797), .A(n13564), .ZN(n13575) );
  XNOR2_X1 U15658 ( .A(n13566), .B(n13565), .ZN(n13570) );
  INV_X1 U15659 ( .A(n13567), .ZN(n13568) );
  AOI21_X1 U15660 ( .B1(n13570), .B2(n13569), .A(n13568), .ZN(n13647) );
  OAI21_X1 U15661 ( .B1(n13572), .B2(n13571), .A(n13647), .ZN(n13573) );
  NAND2_X1 U15662 ( .A1(n13573), .A2(n13562), .ZN(n13574) );
  OAI211_X1 U15663 ( .C1(n13648), .C2(n13576), .A(n13575), .B(n13574), .ZN(
        P2_U3247) );
  OAI211_X1 U15664 ( .C1(n13578), .C2(n14872), .A(n13577), .B(n13579), .ZN(
        n13670) );
  MUX2_X1 U15665 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13670), .S(n14891), .Z(
        P2_U3530) );
  OAI211_X1 U15666 ( .C1(n13581), .C2(n14872), .A(n13580), .B(n13579), .ZN(
        n13671) );
  MUX2_X1 U15667 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13671), .S(n14891), .Z(
        P2_U3529) );
  AOI21_X1 U15668 ( .B1(n14847), .B2(n13583), .A(n13582), .ZN(n13584) );
  MUX2_X1 U15669 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13672), .S(n14891), .Z(
        P2_U3528) );
  NAND2_X1 U15670 ( .A1(n13586), .A2(n14847), .ZN(n13587) );
  MUX2_X1 U15671 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13673), .S(n14891), .Z(
        P2_U3527) );
  AOI21_X1 U15672 ( .B1(n14847), .B2(n13591), .A(n13590), .ZN(n13595) );
  NAND3_X1 U15673 ( .A1(n13593), .A2(n13618), .A3(n13592), .ZN(n13594) );
  NAND3_X1 U15674 ( .A1(n13596), .A2(n13595), .A3(n13594), .ZN(n13674) );
  MUX2_X1 U15675 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13674), .S(n14891), .Z(
        P2_U3526) );
  AOI21_X1 U15676 ( .B1(n14847), .B2(n13598), .A(n13597), .ZN(n13599) );
  OAI211_X1 U15677 ( .C1(n14840), .C2(n13601), .A(n13600), .B(n13599), .ZN(
        n13675) );
  MUX2_X1 U15678 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13675), .S(n14891), .Z(
        P2_U3525) );
  AOI21_X1 U15679 ( .B1(n14847), .B2(n13603), .A(n13602), .ZN(n13604) );
  OAI211_X1 U15680 ( .C1(n14840), .C2(n13606), .A(n13605), .B(n13604), .ZN(
        n13676) );
  MUX2_X1 U15681 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13676), .S(n14891), .Z(
        P2_U3524) );
  NAND2_X1 U15682 ( .A1(n13607), .A2(n14847), .ZN(n13611) );
  OR2_X1 U15683 ( .A1(n13608), .A2(n14840), .ZN(n13610) );
  NAND4_X1 U15684 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13609), .ZN(
        n13677) );
  MUX2_X1 U15685 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13677), .S(n14891), .Z(
        P2_U3523) );
  AOI21_X1 U15686 ( .B1(n14847), .B2(n13614), .A(n13613), .ZN(n13615) );
  OAI211_X1 U15687 ( .C1(n14840), .C2(n13617), .A(n13616), .B(n13615), .ZN(
        n13678) );
  MUX2_X1 U15688 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13678), .S(n14891), .Z(
        P2_U3522) );
  INV_X1 U15689 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15437) );
  NAND3_X1 U15690 ( .A1(n13620), .A2(n13619), .A3(n13618), .ZN(n13624) );
  NAND2_X1 U15691 ( .A1(n13621), .A2(n14847), .ZN(n13623) );
  NAND3_X1 U15692 ( .A1(n13624), .A2(n13623), .A3(n13622), .ZN(n13625) );
  NOR2_X1 U15693 ( .A1(n13626), .A2(n13625), .ZN(n13679) );
  MUX2_X1 U15694 ( .A(n15437), .B(n13679), .S(n14891), .Z(n13627) );
  INV_X1 U15695 ( .A(n13627), .ZN(P2_U3521) );
  AOI21_X1 U15696 ( .B1(n14847), .B2(n13629), .A(n13628), .ZN(n13630) );
  OAI211_X1 U15697 ( .C1(n14840), .C2(n13632), .A(n13631), .B(n13630), .ZN(
        n13682) );
  MUX2_X1 U15698 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13682), .S(n14891), .Z(
        P2_U3520) );
  AOI211_X1 U15699 ( .C1(n14847), .C2(n13635), .A(n13634), .B(n13633), .ZN(
        n13636) );
  OAI21_X1 U15700 ( .B1(n14840), .B2(n13637), .A(n13636), .ZN(n13683) );
  MUX2_X1 U15701 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13683), .S(n14891), .Z(
        P2_U3519) );
  AOI211_X1 U15702 ( .C1(n14847), .C2(n13640), .A(n13639), .B(n13638), .ZN(
        n13642) );
  OAI211_X1 U15703 ( .C1(n13643), .C2(n14840), .A(n13642), .B(n13641), .ZN(
        n13684) );
  MUX2_X1 U15704 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13684), .S(n14891), .Z(
        P2_U3518) );
  AOI21_X1 U15705 ( .B1(n14847), .B2(n13645), .A(n13644), .ZN(n13646) );
  OAI211_X1 U15706 ( .C1(n13648), .C2(n14840), .A(n13647), .B(n13646), .ZN(
        n13685) );
  MUX2_X1 U15707 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13685), .S(n14891), .Z(
        P2_U3517) );
  AOI211_X1 U15708 ( .C1(n14847), .C2(n13651), .A(n13650), .B(n13649), .ZN(
        n13652) );
  OAI21_X1 U15709 ( .B1(n14840), .B2(n13653), .A(n13652), .ZN(n13686) );
  MUX2_X1 U15710 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13686), .S(n14891), .Z(
        P2_U3516) );
  AOI211_X1 U15711 ( .C1(n14847), .C2(n13656), .A(n13655), .B(n13654), .ZN(
        n13658) );
  OAI211_X1 U15712 ( .C1(n13659), .C2(n14840), .A(n13658), .B(n13657), .ZN(
        n13687) );
  MUX2_X1 U15713 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13687), .S(n14891), .Z(
        P2_U3514) );
  AOI21_X1 U15714 ( .B1(n14847), .B2(n13661), .A(n13660), .ZN(n13662) );
  OAI211_X1 U15715 ( .C1(n14840), .C2(n13664), .A(n13663), .B(n13662), .ZN(
        n13688) );
  MUX2_X1 U15716 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13688), .S(n14891), .Z(
        P2_U3513) );
  AOI211_X1 U15717 ( .C1(n14847), .C2(n13667), .A(n13666), .B(n13665), .ZN(
        n13668) );
  OAI21_X1 U15718 ( .B1(n14840), .B2(n13669), .A(n13668), .ZN(n13689) );
  MUX2_X1 U15719 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13689), .S(n14891), .Z(
        P2_U3511) );
  MUX2_X1 U15720 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13670), .S(n14880), .Z(
        P2_U3498) );
  MUX2_X1 U15721 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13671), .S(n14880), .Z(
        P2_U3497) );
  MUX2_X1 U15722 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13674), .S(n14880), .Z(
        P2_U3494) );
  MUX2_X1 U15723 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13675), .S(n14880), .Z(
        P2_U3493) );
  MUX2_X1 U15724 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13676), .S(n14880), .Z(
        P2_U3492) );
  MUX2_X1 U15725 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13677), .S(n14880), .Z(
        P2_U3491) );
  MUX2_X1 U15726 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13678), .S(n14880), .Z(
        P2_U3490) );
  INV_X1 U15727 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13680) );
  MUX2_X1 U15728 ( .A(n13680), .B(n13679), .S(n14880), .Z(n13681) );
  INV_X1 U15729 ( .A(n13681), .ZN(P2_U3489) );
  MUX2_X1 U15730 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13682), .S(n14880), .Z(
        P2_U3488) );
  MUX2_X1 U15731 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13683), .S(n14880), .Z(
        P2_U3487) );
  MUX2_X1 U15732 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13684), .S(n14880), .Z(
        P2_U3486) );
  MUX2_X1 U15733 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13685), .S(n14880), .Z(
        P2_U3484) );
  MUX2_X1 U15734 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13686), .S(n14880), .Z(
        P2_U3481) );
  MUX2_X1 U15735 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13687), .S(n14880), .Z(
        P2_U3475) );
  MUX2_X1 U15736 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13688), .S(n14880), .Z(
        P2_U3472) );
  MUX2_X1 U15737 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n13689), .S(n14880), .Z(
        P2_U3466) );
  INV_X1 U15738 ( .A(n13690), .ZN(n14362) );
  NOR4_X1 U15739 ( .A1(n13691), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8568), .A4(
        P2_U3088), .ZN(n13692) );
  AOI21_X1 U15740 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13698), .A(n13692), 
        .ZN(n13693) );
  OAI21_X1 U15741 ( .B1(n14362), .B2(n12071), .A(n13693), .ZN(P2_U3296) );
  INV_X1 U15742 ( .A(n13694), .ZN(n14365) );
  OAI222_X1 U15743 ( .A1(n12071), .A2(n14365), .B1(P2_U3088), .B2(n13696), 
        .C1(n13695), .C2(n12073), .ZN(P2_U3298) );
  AOI21_X1 U15744 ( .B1(n13698), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13697), 
        .ZN(n13699) );
  OAI21_X1 U15745 ( .B1(n13700), .B2(n12071), .A(n13699), .ZN(P2_U3299) );
  INV_X1 U15746 ( .A(n13701), .ZN(n13702) );
  MUX2_X1 U15747 ( .A(n13702), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15748 ( .A(n13704), .B(n13703), .Z(n13709) );
  NAND2_X1 U15749 ( .A1(n13814), .A2(n14039), .ZN(n13706) );
  AOI22_X1 U15750 ( .A1(n13758), .A2(n14034), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13705) );
  OAI211_X1 U15751 ( .C1(n13749), .C2(n13761), .A(n13706), .B(n13705), .ZN(
        n13707) );
  AOI21_X1 U15752 ( .B1(n14270), .B2(n13834), .A(n13707), .ZN(n13708) );
  OAI21_X1 U15753 ( .B1(n13709), .B2(n13836), .A(n13708), .ZN(P1_U3214) );
  OAI21_X1 U15754 ( .B1(n13712), .B2(n13711), .A(n13710), .ZN(n13713) );
  NAND2_X1 U15755 ( .A1(n13713), .A2(n13809), .ZN(n13718) );
  NAND2_X1 U15756 ( .A1(n13848), .A2(n14209), .ZN(n13714) );
  OAI21_X1 U15757 ( .B1(n14217), .B2(n14221), .A(n13714), .ZN(n14508) );
  NOR2_X1 U15758 ( .A1(n13832), .A2(n14510), .ZN(n13715) );
  AOI211_X1 U15759 ( .C1(n13830), .C2(n14508), .A(n13716), .B(n13715), .ZN(
        n13717) );
  OAI211_X1 U15760 ( .C1(n14525), .C2(n13817), .A(n13718), .B(n13717), .ZN(
        P1_U3215) );
  XOR2_X1 U15761 ( .A(n13720), .B(n13719), .Z(n13725) );
  INV_X1 U15762 ( .A(n13843), .ZN(n13741) );
  OAI22_X1 U15763 ( .A1(n13741), .A2(n14218), .B1(n13721), .B2(n14221), .ZN(
        n14290) );
  AOI22_X1 U15764 ( .A1(n14290), .A2(n13830), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13722) );
  OAI21_X1 U15765 ( .B1(n13832), .B2(n14108), .A(n13722), .ZN(n13723) );
  AOI21_X1 U15766 ( .B1(n14291), .B2(n13834), .A(n13723), .ZN(n13724) );
  OAI21_X1 U15767 ( .B1(n13725), .B2(n13836), .A(n13724), .ZN(P1_U3216) );
  AOI21_X1 U15768 ( .B1(n13727), .B2(n13726), .A(n13836), .ZN(n13729) );
  NAND2_X1 U15769 ( .A1(n13729), .A2(n13728), .ZN(n13735) );
  NAND2_X1 U15770 ( .A1(n13844), .A2(n14207), .ZN(n13731) );
  NAND2_X1 U15771 ( .A1(n14209), .A2(n14206), .ZN(n13730) );
  NAND2_X1 U15772 ( .A1(n13731), .A2(n13730), .ZN(n14312) );
  NOR2_X1 U15773 ( .A1(n13732), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14017) );
  NOR2_X1 U15774 ( .A1(n13832), .A2(n14168), .ZN(n13733) );
  AOI211_X1 U15775 ( .C1(n13830), .C2(n14312), .A(n14017), .B(n13733), .ZN(
        n13734) );
  OAI211_X1 U15776 ( .C1(n7450), .C2(n13817), .A(n13735), .B(n13734), .ZN(
        P1_U3219) );
  INV_X1 U15777 ( .A(n13736), .ZN(n13737) );
  AOI21_X1 U15778 ( .B1(n13739), .B2(n13738), .A(n13737), .ZN(n13745) );
  OAI22_X1 U15779 ( .A1(n13741), .A2(n14221), .B1(n13740), .B2(n14218), .ZN(
        n14137) );
  AOI22_X1 U15780 ( .A1(n14137), .A2(n13830), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13742) );
  OAI21_X1 U15781 ( .B1(n13832), .B2(n14145), .A(n13742), .ZN(n13743) );
  AOI21_X1 U15782 ( .B1(n14299), .B2(n13834), .A(n13743), .ZN(n13744) );
  OAI21_X1 U15783 ( .B1(n13745), .B2(n13836), .A(n13744), .ZN(P1_U3223) );
  XOR2_X1 U15784 ( .A(n13747), .B(n13746), .Z(n13753) );
  NAND2_X1 U15785 ( .A1(n14209), .A2(n13842), .ZN(n13748) );
  OAI21_X1 U15786 ( .B1(n13749), .B2(n14221), .A(n13748), .ZN(n14068) );
  AOI22_X1 U15787 ( .A1(n13830), .A2(n14068), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13750) );
  OAI21_X1 U15788 ( .B1(n13832), .B2(n14075), .A(n13750), .ZN(n13751) );
  AOI21_X1 U15789 ( .B1(n14077), .B2(n13834), .A(n13751), .ZN(n13752) );
  OAI21_X1 U15790 ( .B1(n13753), .B2(n13836), .A(n13752), .ZN(P1_U3225) );
  OAI21_X1 U15791 ( .B1(n13756), .B2(n13755), .A(n13754), .ZN(n13757) );
  NAND2_X1 U15792 ( .A1(n13757), .A2(n13809), .ZN(n13764) );
  NAND2_X1 U15793 ( .A1(n13758), .A2(n13845), .ZN(n13759) );
  OAI211_X1 U15794 ( .C1(n13761), .C2(n14217), .A(n13760), .B(n13759), .ZN(
        n13762) );
  AOI21_X1 U15795 ( .B1(n14222), .B2(n13814), .A(n13762), .ZN(n13763) );
  OAI211_X1 U15796 ( .C1(n14227), .C2(n13817), .A(n13764), .B(n13763), .ZN(
        P1_U3226) );
  INV_X1 U15797 ( .A(n13768), .ZN(n13765) );
  NOR2_X1 U15798 ( .A1(n13766), .A2(n13765), .ZN(n13771) );
  AOI21_X1 U15799 ( .B1(n13769), .B2(n13768), .A(n13767), .ZN(n13770) );
  OAI21_X1 U15800 ( .B1(n13771), .B2(n13770), .A(n13809), .ZN(n13777) );
  NAND2_X1 U15801 ( .A1(n13799), .A2(n14208), .ZN(n13773) );
  OAI211_X1 U15802 ( .C1(n13801), .C2(n13774), .A(n13773), .B(n13772), .ZN(
        n13775) );
  AOI21_X1 U15803 ( .B1(n14200), .B2(n13814), .A(n13775), .ZN(n13776) );
  OAI211_X1 U15804 ( .C1(n14202), .C2(n13817), .A(n13777), .B(n13776), .ZN(
        P1_U3228) );
  XOR2_X1 U15805 ( .A(n13779), .B(n13778), .Z(n13784) );
  INV_X1 U15806 ( .A(n13841), .ZN(n13780) );
  OAI22_X1 U15807 ( .A1(n14218), .A2(n13802), .B1(n13780), .B2(n14221), .ZN(
        n14091) );
  AOI22_X1 U15808 ( .A1(n13830), .A2(n14091), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13781) );
  OAI21_X1 U15809 ( .B1(n13832), .B2(n14095), .A(n13781), .ZN(n13782) );
  AOI21_X1 U15810 ( .B1(n14097), .B2(n13834), .A(n13782), .ZN(n13783) );
  OAI21_X1 U15811 ( .B1(n13784), .B2(n13836), .A(n13783), .ZN(P1_U3229) );
  INV_X1 U15812 ( .A(n14304), .ZN(n13794) );
  OAI211_X1 U15813 ( .C1(n13787), .C2(n13786), .A(n13785), .B(n13809), .ZN(
        n13793) );
  INV_X1 U15814 ( .A(n13788), .ZN(n14157) );
  AOI22_X1 U15815 ( .A1(n13799), .A2(n14151), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13789) );
  OAI21_X1 U15816 ( .B1(n13790), .B2(n13801), .A(n13789), .ZN(n13791) );
  AOI21_X1 U15817 ( .B1(n14157), .B2(n13814), .A(n13791), .ZN(n13792) );
  OAI211_X1 U15818 ( .C1(n13794), .C2(n13817), .A(n13793), .B(n13792), .ZN(
        P1_U3233) );
  OAI21_X1 U15819 ( .B1(n13797), .B2(n13796), .A(n13795), .ZN(n13798) );
  NAND2_X1 U15820 ( .A1(n13798), .A2(n13809), .ZN(n13805) );
  AOI22_X1 U15821 ( .A1(n13799), .A2(n14152), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13800) );
  OAI21_X1 U15822 ( .B1(n13802), .B2(n13801), .A(n13800), .ZN(n13803) );
  AOI21_X1 U15823 ( .B1(n14127), .B2(n13814), .A(n13803), .ZN(n13804) );
  OAI211_X1 U15824 ( .C1(n13817), .C2(n14298), .A(n13805), .B(n13804), .ZN(
        P1_U3235) );
  OAI21_X1 U15825 ( .B1(n13808), .B2(n13807), .A(n13806), .ZN(n13810) );
  NAND2_X1 U15826 ( .A1(n13810), .A2(n13809), .ZN(n13816) );
  INV_X1 U15827 ( .A(n14190), .ZN(n13813) );
  AOI22_X1 U15828 ( .A1(n14151), .A2(n14207), .B1(n14209), .B2(n13845), .ZN(
        n14187) );
  NAND2_X1 U15829 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14594)
         );
  OAI21_X1 U15830 ( .B1(n13811), .B2(n14187), .A(n14594), .ZN(n13812) );
  AOI21_X1 U15831 ( .B1(n13814), .B2(n13813), .A(n13812), .ZN(n13815) );
  OAI211_X1 U15832 ( .C1(n14318), .C2(n13817), .A(n13816), .B(n13815), .ZN(
        P1_U3238) );
  XOR2_X1 U15833 ( .A(n13819), .B(n13818), .Z(n13825) );
  INV_X1 U15834 ( .A(n13840), .ZN(n13821) );
  NAND2_X1 U15835 ( .A1(n14209), .A2(n13841), .ZN(n13820) );
  OAI21_X1 U15836 ( .B1(n13821), .B2(n14221), .A(n13820), .ZN(n14049) );
  AOI22_X1 U15837 ( .A1(n13830), .A2(n14049), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13822) );
  OAI21_X1 U15838 ( .B1(n13832), .B2(n14052), .A(n13822), .ZN(n13823) );
  AOI21_X1 U15839 ( .B1(n14275), .B2(n13834), .A(n13823), .ZN(n13824) );
  OAI21_X1 U15840 ( .B1(n13825), .B2(n13836), .A(n13824), .ZN(P1_U3240) );
  XNOR2_X1 U15841 ( .A(n13826), .B(n13827), .ZN(n13837) );
  NAND2_X1 U15842 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14580)
         );
  OAI22_X1 U15843 ( .A1(n14218), .A2(n13829), .B1(n13828), .B2(n14221), .ZN(
        n14237) );
  NAND2_X1 U15844 ( .A1(n13830), .A2(n14237), .ZN(n13831) );
  OAI211_X1 U15845 ( .C1(n13832), .C2(n14243), .A(n14580), .B(n13831), .ZN(
        n13833) );
  AOI21_X1 U15846 ( .B1(n14334), .B2(n13834), .A(n13833), .ZN(n13835) );
  OAI21_X1 U15847 ( .B1(n13837), .B2(n13836), .A(n13835), .ZN(P1_U3241) );
  MUX2_X1 U15848 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14021), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15849 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13838), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15850 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13839), .S(n13861), .Z(
        P1_U3589) );
  MUX2_X1 U15851 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14034), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15852 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13840), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15853 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14033), .S(n13861), .Z(
        P1_U3586) );
  MUX2_X1 U15854 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13841), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15855 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13842), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15856 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14121), .S(n13861), .Z(
        P1_U3583) );
  MUX2_X1 U15857 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13843), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15858 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14152), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15859 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13844), .S(n13861), .Z(
        P1_U3580) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14151), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15861 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14206), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15862 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13845), .S(n13861), .Z(
        P1_U3577) );
  MUX2_X1 U15863 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14208), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15864 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13846), .S(n13861), .Z(
        P1_U3575) );
  MUX2_X1 U15865 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13847), .S(n13861), .Z(
        P1_U3574) );
  MUX2_X1 U15866 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13848), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15867 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13849), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15868 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13850), .S(n13861), .Z(
        P1_U3571) );
  MUX2_X1 U15869 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13851), .S(n13861), .Z(
        P1_U3570) );
  MUX2_X1 U15870 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13852), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15871 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13853), .S(n13861), .Z(
        P1_U3568) );
  MUX2_X1 U15872 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13854), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15873 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13855), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15874 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13856), .S(n13861), .Z(
        P1_U3565) );
  MUX2_X1 U15875 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13857), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15876 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13858), .S(n13861), .Z(
        P1_U3563) );
  MUX2_X1 U15877 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13859), .S(n13861), .Z(
        P1_U3562) );
  MUX2_X1 U15878 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13860), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15879 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10342), .S(n13861), .Z(
        P1_U3560) );
  OAI22_X1 U15880 ( .A1(n14596), .A2(n13863), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13862), .ZN(n13864) );
  AOI21_X1 U15881 ( .B1(n13865), .B2(n13984), .A(n13864), .ZN(n13874) );
  MUX2_X1 U15882 ( .A(n10084), .B(P1_REG1_REG_1__SCAN_IN), .S(n13865), .Z(
        n13866) );
  OAI21_X1 U15883 ( .B1(n9296), .B2(n13867), .A(n13866), .ZN(n13868) );
  NAND3_X1 U15884 ( .A1(n14011), .A2(n13869), .A3(n13868), .ZN(n13873) );
  OAI211_X1 U15885 ( .C1(n13877), .C2(n13871), .A(n14012), .B(n13870), .ZN(
        n13872) );
  NAND3_X1 U15886 ( .A1(n13874), .A2(n13873), .A3(n13872), .ZN(P1_U3244) );
  AOI21_X1 U15887 ( .B1(n14564), .B2(n9297), .A(n13875), .ZN(n14563) );
  MUX2_X1 U15888 ( .A(n13877), .B(n13876), .S(n14370), .Z(n13879) );
  NAND2_X1 U15889 ( .A1(n13879), .A2(n13878), .ZN(n13880) );
  OAI211_X1 U15890 ( .C1(n14566), .C2(n14563), .A(n13880), .B(P1_U4016), .ZN(
        n13924) );
  AOI22_X1 U15891 ( .A1(n14568), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13892) );
  OAI21_X1 U15892 ( .B1(n13882), .B2(n13881), .A(n13899), .ZN(n13883) );
  NOR2_X1 U15893 ( .A1(n14588), .A2(n13883), .ZN(n13889) );
  INV_X1 U15894 ( .A(n13884), .ZN(n13887) );
  MUX2_X1 U15895 ( .A(n9308), .B(P1_REG1_REG_2__SCAN_IN), .S(n13890), .Z(
        n13886) );
  INV_X1 U15896 ( .A(n13895), .ZN(n13885) );
  AOI211_X1 U15897 ( .C1(n13887), .C2(n13886), .A(n13885), .B(n14590), .ZN(
        n13888) );
  AOI211_X1 U15898 ( .C1(n13984), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        n13891) );
  NAND3_X1 U15899 ( .A1(n13924), .A2(n13892), .A3(n13891), .ZN(P1_U3245) );
  MUX2_X1 U15900 ( .A(n10089), .B(P1_REG1_REG_3__SCAN_IN), .S(n13902), .Z(
        n13893) );
  NAND3_X1 U15901 ( .A1(n13895), .A2(n13894), .A3(n13893), .ZN(n13896) );
  NAND3_X1 U15902 ( .A1(n14011), .A2(n13909), .A3(n13896), .ZN(n13906) );
  MUX2_X1 U15903 ( .A(n10819), .B(P1_REG2_REG_3__SCAN_IN), .S(n13902), .Z(
        n13897) );
  NAND3_X1 U15904 ( .A1(n13899), .A2(n13898), .A3(n13897), .ZN(n13900) );
  NAND3_X1 U15905 ( .A1(n14012), .A2(n13914), .A3(n13900), .ZN(n13905) );
  AOI21_X1 U15906 ( .B1(n14568), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n13901), .ZN(
        n13904) );
  NAND2_X1 U15907 ( .A1(n13984), .A2(n13902), .ZN(n13903) );
  NAND4_X1 U15908 ( .A1(n13906), .A2(n13905), .A3(n13904), .A4(n13903), .ZN(
        P1_U3246) );
  NAND2_X1 U15909 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14568), .ZN(n13923) );
  INV_X1 U15910 ( .A(n13907), .ZN(n13912) );
  NAND3_X1 U15911 ( .A1(n13910), .A2(n13909), .A3(n13908), .ZN(n13911) );
  NAND3_X1 U15912 ( .A1(n14011), .A2(n13912), .A3(n13911), .ZN(n13921) );
  MUX2_X1 U15913 ( .A(n10100), .B(P1_REG2_REG_4__SCAN_IN), .S(n13917), .Z(
        n13915) );
  NAND3_X1 U15914 ( .A1(n13915), .A2(n13914), .A3(n13913), .ZN(n13916) );
  NAND3_X1 U15915 ( .A1(n14012), .A2(n13934), .A3(n13916), .ZN(n13920) );
  NAND2_X1 U15916 ( .A1(n13984), .A2(n13917), .ZN(n13918) );
  AND4_X1 U15917 ( .A1(n13921), .A2(n13920), .A3(n13919), .A4(n13918), .ZN(
        n13922) );
  NAND3_X1 U15918 ( .A1(n13924), .A2(n13923), .A3(n13922), .ZN(P1_U3247) );
  OAI21_X1 U15919 ( .B1(n14596), .B2(n6948), .A(n13925), .ZN(n13926) );
  AOI21_X1 U15920 ( .B1(n13927), .B2(n13984), .A(n13926), .ZN(n13939) );
  OAI21_X1 U15921 ( .B1(n13930), .B2(n13929), .A(n13928), .ZN(n13931) );
  NAND2_X1 U15922 ( .A1(n14011), .A2(n13931), .ZN(n13938) );
  NAND3_X1 U15923 ( .A1(n13934), .A2(n13933), .A3(n13932), .ZN(n13935) );
  NAND3_X1 U15924 ( .A1(n14012), .A2(n13936), .A3(n13935), .ZN(n13937) );
  NAND3_X1 U15925 ( .A1(n13939), .A2(n13938), .A3(n13937), .ZN(P1_U3248) );
  NOR2_X1 U15926 ( .A1(n14596), .A2(n13940), .ZN(n13941) );
  AOI211_X1 U15927 ( .C1(n13984), .C2(n13950), .A(n13942), .B(n13941), .ZN(
        n13959) );
  MUX2_X1 U15928 ( .A(n13943), .B(P1_REG1_REG_7__SCAN_IN), .S(n13950), .Z(
        n13946) );
  INV_X1 U15929 ( .A(n13944), .ZN(n13945) );
  NAND2_X1 U15930 ( .A1(n13946), .A2(n13945), .ZN(n13948) );
  OAI211_X1 U15931 ( .C1(n13949), .C2(n13948), .A(n14011), .B(n13947), .ZN(
        n13958) );
  MUX2_X1 U15932 ( .A(n10125), .B(P1_REG2_REG_7__SCAN_IN), .S(n13950), .Z(
        n13953) );
  INV_X1 U15933 ( .A(n13951), .ZN(n13952) );
  NAND2_X1 U15934 ( .A1(n13953), .A2(n13952), .ZN(n13955) );
  OAI211_X1 U15935 ( .C1(n13956), .C2(n13955), .A(n14012), .B(n13954), .ZN(
        n13957) );
  NAND3_X1 U15936 ( .A1(n13959), .A2(n13958), .A3(n13957), .ZN(P1_U3250) );
  INV_X1 U15937 ( .A(n13960), .ZN(n13965) );
  NOR3_X1 U15938 ( .A1(n13963), .A2(n13962), .A3(n13961), .ZN(n13964) );
  OAI21_X1 U15939 ( .B1(n13965), .B2(n13964), .A(n14011), .ZN(n13977) );
  OAI21_X1 U15940 ( .B1(n14596), .B2(n6951), .A(n13966), .ZN(n13967) );
  AOI21_X1 U15941 ( .B1(n13968), .B2(n13984), .A(n13967), .ZN(n13976) );
  MUX2_X1 U15942 ( .A(n11273), .B(P1_REG2_REG_9__SCAN_IN), .S(n13968), .Z(
        n13971) );
  INV_X1 U15943 ( .A(n13969), .ZN(n13970) );
  NAND2_X1 U15944 ( .A1(n13971), .A2(n13970), .ZN(n13973) );
  OAI211_X1 U15945 ( .C1(n13974), .C2(n13973), .A(n13972), .B(n14012), .ZN(
        n13975) );
  NAND3_X1 U15946 ( .A1(n13977), .A2(n13976), .A3(n13975), .ZN(P1_U3252) );
  OAI21_X1 U15947 ( .B1(n13980), .B2(n13979), .A(n13978), .ZN(n13981) );
  NAND2_X1 U15948 ( .A1(n13981), .A2(n14011), .ZN(n13993) );
  OAI21_X1 U15949 ( .B1(n14596), .B2(n15351), .A(n13982), .ZN(n13983) );
  AOI21_X1 U15950 ( .B1(n13985), .B2(n13984), .A(n13983), .ZN(n13992) );
  OR3_X1 U15951 ( .A1(n13988), .A2(n13987), .A3(n13986), .ZN(n13989) );
  NAND3_X1 U15952 ( .A1(n13990), .A2(n14012), .A3(n13989), .ZN(n13991) );
  NAND3_X1 U15953 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(P1_U3254) );
  NAND2_X1 U15954 ( .A1(n13995), .A2(n13994), .ZN(n13996) );
  XNOR2_X1 U15955 ( .A(n14591), .B(n13996), .ZN(n14586) );
  NAND2_X1 U15956 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14586), .ZN(n14585) );
  NAND2_X1 U15957 ( .A1(n14005), .A2(n13996), .ZN(n13997) );
  NAND2_X1 U15958 ( .A1(n14585), .A2(n13997), .ZN(n13998) );
  XOR2_X1 U15959 ( .A(n13998), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14013) );
  INV_X1 U15960 ( .A(n14013), .ZN(n14009) );
  INV_X1 U15961 ( .A(n13999), .ZN(n14003) );
  INV_X1 U15962 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14000) );
  OAI22_X1 U15963 ( .A1(n14003), .A2(n14002), .B1(n14001), .B2(n14000), .ZN(
        n14004) );
  XNOR2_X1 U15964 ( .A(n14591), .B(n14004), .ZN(n14584) );
  NAND2_X1 U15965 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14584), .ZN(n14583) );
  NAND2_X1 U15966 ( .A1(n14005), .A2(n14004), .ZN(n14006) );
  NAND2_X1 U15967 ( .A1(n14583), .A2(n14006), .ZN(n14007) );
  INV_X1 U15968 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15413) );
  XNOR2_X1 U15969 ( .A(n14007), .B(n15413), .ZN(n14010) );
  OAI21_X1 U15970 ( .B1(n14010), .B2(n14590), .A(n14592), .ZN(n14008) );
  AOI21_X1 U15971 ( .B1(n14012), .B2(n14009), .A(n14008), .ZN(n14016) );
  AOI22_X1 U15972 ( .A1(n14013), .A2(n14012), .B1(n14011), .B2(n14010), .ZN(
        n14015) );
  MUX2_X1 U15973 ( .A(n14016), .B(n14015), .S(n14014), .Z(n14019) );
  INV_X1 U15974 ( .A(n14017), .ZN(n14018) );
  OAI211_X1 U15975 ( .C1(n7813), .C2(n14596), .A(n14019), .B(n14018), .ZN(
        P1_U3262) );
  NAND2_X1 U15976 ( .A1(n14257), .A2(n14026), .ZN(n14025) );
  XNOR2_X1 U15977 ( .A(n14254), .B(n14025), .ZN(n14020) );
  NAND2_X1 U15978 ( .A1(n14020), .A2(n14622), .ZN(n14253) );
  NAND2_X1 U15979 ( .A1(n14022), .A2(n14021), .ZN(n14255) );
  NOR2_X1 U15980 ( .A1(n14642), .A2(n14255), .ZN(n14028) );
  NOR2_X1 U15981 ( .A1(n14254), .A2(n14616), .ZN(n14023) );
  AOI211_X1 U15982 ( .C1(n14642), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14028), 
        .B(n14023), .ZN(n14024) );
  OAI21_X1 U15983 ( .B1(n14253), .B2(n14196), .A(n14024), .ZN(P1_U3263) );
  OAI211_X1 U15984 ( .C1(n14257), .C2(n14026), .A(n14622), .B(n14025), .ZN(
        n14256) );
  AND2_X1 U15985 ( .A1(n14642), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14027) );
  NOR2_X1 U15986 ( .A1(n14028), .A2(n14027), .ZN(n14031) );
  NAND2_X1 U15987 ( .A1(n14029), .A2(n14512), .ZN(n14030) );
  OAI211_X1 U15988 ( .C1(n14256), .C2(n14196), .A(n14031), .B(n14030), .ZN(
        P1_U3264) );
  XNOR2_X1 U15989 ( .A(n14032), .B(n7325), .ZN(n14035) );
  AOI222_X1 U15990 ( .A1(n14611), .A2(n14035), .B1(n14034), .B2(n14207), .C1(
        n14033), .C2(n14209), .ZN(n14272) );
  INV_X1 U15991 ( .A(n14051), .ZN(n14038) );
  INV_X1 U15992 ( .A(n14036), .ZN(n14037) );
  AOI211_X1 U15993 ( .C1(n14270), .C2(n14038), .A(n14242), .B(n14037), .ZN(
        n14269) );
  AOI22_X1 U15994 ( .A1(n14642), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14039), 
        .B2(n14599), .ZN(n14040) );
  OAI21_X1 U15995 ( .B1(n14041), .B2(n14616), .A(n14040), .ZN(n14045) );
  INV_X1 U15996 ( .A(n14042), .ZN(n14043) );
  AOI21_X1 U15997 ( .B1(n7328), .B2(n14044), .A(n14043), .ZN(n14273) );
  OAI21_X1 U15998 ( .B1(n14272), .B2(n14642), .A(n14046), .ZN(P1_U3266) );
  XNOR2_X1 U15999 ( .A(n14048), .B(n14047), .ZN(n14050) );
  AOI21_X1 U16000 ( .B1(n14050), .B2(n14611), .A(n14049), .ZN(n14277) );
  AOI211_X1 U16001 ( .C1(n14275), .C2(n6598), .A(n14242), .B(n14051), .ZN(
        n14274) );
  INV_X1 U16002 ( .A(n14275), .ZN(n14055) );
  INV_X1 U16003 ( .A(n14052), .ZN(n14053) );
  AOI22_X1 U16004 ( .A1(n14642), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14053), 
        .B2(n14599), .ZN(n14054) );
  OAI21_X1 U16005 ( .B1(n14055), .B2(n14616), .A(n14054), .ZN(n14061) );
  OR2_X1 U16006 ( .A1(n14057), .A2(n14056), .ZN(n14058) );
  NAND2_X1 U16007 ( .A1(n14059), .A2(n14058), .ZN(n14278) );
  NOR2_X1 U16008 ( .A1(n14278), .A2(n14249), .ZN(n14060) );
  AOI211_X1 U16009 ( .C1(n14274), .C2(n14626), .A(n14061), .B(n14060), .ZN(
        n14062) );
  OAI21_X1 U16010 ( .B1(n14642), .B2(n14277), .A(n14062), .ZN(P1_U3267) );
  NAND2_X1 U16011 ( .A1(n14064), .A2(n14063), .ZN(n14065) );
  NAND2_X1 U16012 ( .A1(n14066), .A2(n14065), .ZN(n14067) );
  NAND2_X1 U16013 ( .A1(n14067), .A2(n14611), .ZN(n14070) );
  INV_X1 U16014 ( .A(n14068), .ZN(n14069) );
  NAND2_X1 U16015 ( .A1(n14070), .A2(n14069), .ZN(n14284) );
  AOI21_X1 U16016 ( .B1(n14082), .B2(n14077), .A(n14242), .ZN(n14071) );
  NAND2_X1 U16017 ( .A1(n14071), .A2(n6598), .ZN(n14280) );
  NAND2_X1 U16018 ( .A1(n6675), .A2(n14072), .ZN(n14279) );
  NAND3_X1 U16019 ( .A1(n14279), .A2(n14627), .A3(n14073), .ZN(n14079) );
  NAND2_X1 U16020 ( .A1(n14642), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14074) );
  OAI21_X1 U16021 ( .B1(n14637), .B2(n14075), .A(n14074), .ZN(n14076) );
  AOI21_X1 U16022 ( .B1(n14077), .B2(n14512), .A(n14076), .ZN(n14078) );
  OAI211_X1 U16023 ( .C1(n14280), .C2(n14196), .A(n14079), .B(n14078), .ZN(
        n14080) );
  AOI21_X1 U16024 ( .B1(n14284), .B2(n14226), .A(n14080), .ZN(n14081) );
  INV_X1 U16025 ( .A(n14081), .ZN(P1_U3268) );
  OAI211_X1 U16026 ( .C1(n14104), .C2(n14288), .A(n14622), .B(n14082), .ZN(
        n14286) );
  INV_X1 U16027 ( .A(n14083), .ZN(n14084) );
  AOI21_X1 U16028 ( .B1(n14084), .B2(n7344), .A(n14234), .ZN(n14093) );
  INV_X1 U16029 ( .A(n14100), .ZN(n14087) );
  OAI21_X1 U16030 ( .B1(n14087), .B2(n14086), .A(n14085), .ZN(n14089) );
  AOI21_X1 U16031 ( .B1(n14089), .B2(n14088), .A(n14404), .ZN(n14090) );
  AOI211_X1 U16032 ( .C1(n14093), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14287) );
  OR2_X1 U16033 ( .A1(n14287), .A2(n14642), .ZN(n14099) );
  NAND2_X1 U16034 ( .A1(n14642), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n14094) );
  OAI21_X1 U16035 ( .B1(n14637), .B2(n14095), .A(n14094), .ZN(n14096) );
  AOI21_X1 U16036 ( .B1(n14097), .B2(n14512), .A(n14096), .ZN(n14098) );
  OAI211_X1 U16037 ( .C1(n14286), .C2(n14196), .A(n14099), .B(n14098), .ZN(
        P1_U3269) );
  INV_X1 U16038 ( .A(n14105), .ZN(n14101) );
  OAI21_X1 U16039 ( .B1(n7701), .B2(n14101), .A(n14100), .ZN(n14294) );
  NAND2_X1 U16040 ( .A1(n14125), .A2(n14291), .ZN(n14102) );
  NAND2_X1 U16041 ( .A1(n14102), .A2(n14622), .ZN(n14103) );
  NOR2_X1 U16042 ( .A1(n14104), .A2(n14103), .ZN(n14289) );
  INV_X1 U16043 ( .A(n14289), .ZN(n14111) );
  XNOR2_X1 U16044 ( .A(n14106), .B(n14105), .ZN(n14107) );
  NAND2_X1 U16045 ( .A1(n14107), .A2(n14611), .ZN(n14293) );
  INV_X1 U16046 ( .A(n14108), .ZN(n14109) );
  AOI21_X1 U16047 ( .B1(n14109), .B2(n14599), .A(n14290), .ZN(n14110) );
  OAI211_X1 U16048 ( .C1(n14143), .C2(n14111), .A(n14293), .B(n14110), .ZN(
        n14112) );
  NAND2_X1 U16049 ( .A1(n14112), .A2(n14226), .ZN(n14114) );
  AOI22_X1 U16050 ( .A1(n14291), .A2(n14512), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n14642), .ZN(n14113) );
  OAI211_X1 U16051 ( .C1(n14294), .C2(n14249), .A(n14114), .B(n14113), .ZN(
        P1_U3270) );
  INV_X1 U16052 ( .A(n14115), .ZN(n14116) );
  NAND2_X1 U16053 ( .A1(n14116), .A2(n14707), .ZN(n14120) );
  AOI22_X1 U16054 ( .A1(n14117), .A2(n14611), .B1(n14115), .B2(n14707), .ZN(
        n14119) );
  MUX2_X1 U16055 ( .A(n14120), .B(n14119), .S(n14118), .Z(n14123) );
  AOI22_X1 U16056 ( .A1(n14152), .A2(n14209), .B1(n14207), .B2(n14121), .ZN(
        n14122) );
  OAI211_X1 U16057 ( .C1(n14234), .C2(n14124), .A(n14123), .B(n14122), .ZN(
        n14295) );
  AOI21_X1 U16058 ( .B1(n14128), .B2(n14133), .A(n14242), .ZN(n14126) );
  NAND2_X1 U16059 ( .A1(n14126), .A2(n14125), .ZN(n14296) );
  AOI22_X1 U16060 ( .A1(n14642), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14127), 
        .B2(n14599), .ZN(n14130) );
  NAND2_X1 U16061 ( .A1(n14128), .A2(n14512), .ZN(n14129) );
  OAI211_X1 U16062 ( .C1(n14296), .C2(n14196), .A(n14130), .B(n14129), .ZN(
        n14131) );
  AOI21_X1 U16063 ( .B1(n14295), .B2(n14226), .A(n14131), .ZN(n14132) );
  INV_X1 U16064 ( .A(n14132), .ZN(P1_U3271) );
  OAI211_X1 U16065 ( .C1(n14149), .C2(n6714), .A(n14622), .B(n14133), .ZN(
        n14301) );
  OAI21_X1 U16066 ( .B1(n14136), .B2(n9554), .A(n14135), .ZN(n14138) );
  AOI21_X1 U16067 ( .B1(n14138), .B2(n14707), .A(n14137), .ZN(n14302) );
  NAND3_X1 U16068 ( .A1(n14139), .A2(n9554), .A3(n14140), .ZN(n14141) );
  NAND3_X1 U16069 ( .A1(n14142), .A2(n14611), .A3(n14141), .ZN(n14303) );
  OAI211_X1 U16070 ( .C1(n14143), .C2(n14301), .A(n14302), .B(n14303), .ZN(
        n14144) );
  NAND2_X1 U16071 ( .A1(n14144), .A2(n14226), .ZN(n14148) );
  INV_X1 U16072 ( .A(n14145), .ZN(n14146) );
  AOI22_X1 U16073 ( .A1(n14642), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14146), 
        .B2(n14599), .ZN(n14147) );
  OAI211_X1 U16074 ( .C1(n14149), .C2(n14616), .A(n14148), .B(n14147), .ZN(
        P1_U3272) );
  OAI211_X1 U16075 ( .C1(n14150), .C2(n14161), .A(n14139), .B(n14611), .ZN(
        n14154) );
  AOI22_X1 U16076 ( .A1(n14152), .A2(n14207), .B1(n14209), .B2(n14151), .ZN(
        n14153) );
  AND2_X1 U16077 ( .A1(n14154), .A2(n14153), .ZN(n14310) );
  NAND2_X1 U16078 ( .A1(n14304), .A2(n14166), .ZN(n14155) );
  NAND2_X1 U16079 ( .A1(n14155), .A2(n14622), .ZN(n14156) );
  OR2_X1 U16080 ( .A1(n6714), .A2(n14156), .ZN(n14307) );
  AOI22_X1 U16081 ( .A1(n14642), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14157), 
        .B2(n14599), .ZN(n14159) );
  NAND2_X1 U16082 ( .A1(n14304), .A2(n14512), .ZN(n14158) );
  OAI211_X1 U16083 ( .C1(n14307), .C2(n14196), .A(n14159), .B(n14158), .ZN(
        n14160) );
  INV_X1 U16084 ( .A(n14160), .ZN(n14164) );
  NAND2_X1 U16085 ( .A1(n14162), .A2(n14161), .ZN(n14305) );
  NAND3_X1 U16086 ( .A1(n14306), .A2(n14305), .A3(n14627), .ZN(n14163) );
  OAI211_X1 U16087 ( .C1(n14310), .C2(n14642), .A(n14164), .B(n14163), .ZN(
        P1_U3273) );
  XNOR2_X1 U16088 ( .A(n14165), .B(n14174), .ZN(n14316) );
  AOI21_X1 U16089 ( .B1(n14313), .B2(n14181), .A(n14242), .ZN(n14167) );
  AND2_X1 U16090 ( .A1(n14167), .A2(n14166), .ZN(n14311) );
  NAND2_X1 U16091 ( .A1(n14313), .A2(n14512), .ZN(n14171) );
  NOR2_X1 U16092 ( .A1(n14637), .A2(n14168), .ZN(n14169) );
  AOI21_X1 U16093 ( .B1(n14642), .B2(P1_REG2_REG_19__SCAN_IN), .A(n14169), 
        .ZN(n14170) );
  NAND2_X1 U16094 ( .A1(n14171), .A2(n14170), .ZN(n14179) );
  INV_X1 U16095 ( .A(n14172), .ZN(n14175) );
  OAI21_X1 U16096 ( .B1(n14175), .B2(n14174), .A(n14173), .ZN(n14176) );
  NAND2_X1 U16097 ( .A1(n14176), .A2(n14611), .ZN(n14315) );
  INV_X1 U16098 ( .A(n14312), .ZN(n14177) );
  AOI21_X1 U16099 ( .B1(n14315), .B2(n14177), .A(n14642), .ZN(n14178) );
  AOI211_X1 U16100 ( .C1(n14311), .C2(n14626), .A(n14179), .B(n14178), .ZN(
        n14180) );
  OAI21_X1 U16101 ( .B1(n14316), .B2(n14249), .A(n14180), .ZN(P1_U3274) );
  OAI211_X1 U16102 ( .C1(n14198), .C2(n14318), .A(n14622), .B(n14181), .ZN(
        n14317) );
  XNOR2_X1 U16103 ( .A(n14182), .B(n14185), .ZN(n14183) );
  NAND2_X1 U16104 ( .A1(n14183), .A2(n14707), .ZN(n14189) );
  OAI211_X1 U16105 ( .C1(n14186), .C2(n14185), .A(n14184), .B(n14611), .ZN(
        n14188) );
  NAND3_X1 U16106 ( .A1(n14189), .A2(n14188), .A3(n14187), .ZN(n14320) );
  NAND2_X1 U16107 ( .A1(n14320), .A2(n14226), .ZN(n14195) );
  OAI22_X1 U16108 ( .A1(n14226), .A2(n14191), .B1(n14190), .B2(n14637), .ZN(
        n14192) );
  AOI21_X1 U16109 ( .B1(n14193), .B2(n14512), .A(n14192), .ZN(n14194) );
  OAI211_X1 U16110 ( .C1(n14317), .C2(n14196), .A(n14195), .B(n14194), .ZN(
        P1_U3275) );
  XOR2_X1 U16111 ( .A(n14197), .B(n14203), .Z(n14327) );
  OAI21_X1 U16112 ( .B1(n14225), .B2(n14202), .A(n14622), .ZN(n14199) );
  NOR2_X1 U16113 ( .A1(n14199), .A2(n14198), .ZN(n14323) );
  AOI22_X1 U16114 ( .A1(n14642), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14200), 
        .B2(n14599), .ZN(n14201) );
  OAI21_X1 U16115 ( .B1(n14202), .B2(n14616), .A(n14201), .ZN(n14214) );
  INV_X1 U16116 ( .A(n14203), .ZN(n14205) );
  OAI211_X1 U16117 ( .C1(n6723), .C2(n14205), .A(n14611), .B(n14204), .ZN(
        n14325) );
  NAND2_X1 U16118 ( .A1(n14207), .A2(n14206), .ZN(n14211) );
  NAND2_X1 U16119 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  NAND2_X1 U16120 ( .A1(n14211), .A2(n14210), .ZN(n14324) );
  INV_X1 U16121 ( .A(n14324), .ZN(n14212) );
  AOI21_X1 U16122 ( .B1(n14325), .B2(n14212), .A(n14642), .ZN(n14213) );
  AOI211_X1 U16123 ( .C1(n14323), .C2(n14626), .A(n14214), .B(n14213), .ZN(
        n14215) );
  OAI21_X1 U16124 ( .B1(n14249), .B2(n14327), .A(n14215), .ZN(P1_U3276) );
  XOR2_X1 U16125 ( .A(n14216), .B(n14228), .Z(n14219) );
  OAI222_X1 U16126 ( .A1(n14221), .A2(n14220), .B1(n14219), .B2(n14234), .C1(
        n14218), .C2(n14217), .ZN(n14328) );
  AOI21_X1 U16127 ( .B1(n14222), .B2(n14599), .A(n14328), .ZN(n14233) );
  NAND2_X1 U16128 ( .A1(n14240), .A2(n14330), .ZN(n14223) );
  NAND2_X1 U16129 ( .A1(n14223), .A2(n14622), .ZN(n14224) );
  NOR2_X1 U16130 ( .A1(n14225), .A2(n14224), .ZN(n14329) );
  OAI22_X1 U16131 ( .A1(n14227), .A2(n14616), .B1(n11317), .B2(n14226), .ZN(
        n14231) );
  XOR2_X1 U16132 ( .A(n14229), .B(n14228), .Z(n14332) );
  NOR2_X1 U16133 ( .A1(n14332), .A2(n14249), .ZN(n14230) );
  AOI211_X1 U16134 ( .C1(n14329), .C2(n14626), .A(n14231), .B(n14230), .ZN(
        n14232) );
  OAI21_X1 U16135 ( .B1(n14642), .B2(n14233), .A(n14232), .ZN(P1_U3277) );
  AOI21_X1 U16136 ( .B1(n14236), .B2(n14235), .A(n14234), .ZN(n14239) );
  AOI21_X1 U16137 ( .B1(n14239), .B2(n14238), .A(n14237), .ZN(n14336) );
  INV_X1 U16138 ( .A(n14240), .ZN(n14241) );
  AOI211_X1 U16139 ( .C1(n14334), .C2(n14519), .A(n14242), .B(n14241), .ZN(
        n14333) );
  INV_X1 U16140 ( .A(n14243), .ZN(n14244) );
  AOI22_X1 U16141 ( .A1(n14642), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14244), 
        .B2(n14599), .ZN(n14245) );
  OAI21_X1 U16142 ( .B1(n14246), .B2(n14616), .A(n14245), .ZN(n14251) );
  AOI21_X1 U16143 ( .B1(n14248), .B2(n14247), .A(n6720), .ZN(n14337) );
  NOR2_X1 U16144 ( .A1(n14337), .A2(n14249), .ZN(n14250) );
  AOI211_X1 U16145 ( .C1(n14333), .C2(n14626), .A(n14251), .B(n14250), .ZN(
        n14252) );
  OAI21_X1 U16146 ( .B1(n14642), .B2(n14336), .A(n14252), .ZN(P1_U3278) );
  OAI211_X1 U16147 ( .C1(n14254), .C2(n14702), .A(n14253), .B(n14255), .ZN(
        n14338) );
  MUX2_X1 U16148 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14338), .S(n14720), .Z(
        P1_U3559) );
  OAI211_X1 U16149 ( .C1(n14257), .C2(n14702), .A(n14256), .B(n14255), .ZN(
        n14339) );
  MUX2_X1 U16150 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14339), .S(n14720), .Z(
        P1_U3558) );
  AOI21_X1 U16151 ( .B1(n14697), .B2(n14265), .A(n14264), .ZN(n14266) );
  OAI211_X1 U16152 ( .C1(n14404), .C2(n14268), .A(n14267), .B(n14266), .ZN(
        n14341) );
  MUX2_X1 U16153 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14341), .S(n14720), .Z(
        P1_U3556) );
  AOI21_X1 U16154 ( .B1(n14697), .B2(n14270), .A(n14269), .ZN(n14271) );
  OAI211_X1 U16155 ( .C1(n14273), .C2(n14404), .A(n14272), .B(n14271), .ZN(
        n14342) );
  MUX2_X1 U16156 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14342), .S(n14720), .Z(
        P1_U3555) );
  AOI21_X1 U16157 ( .B1(n14697), .B2(n14275), .A(n14274), .ZN(n14276) );
  OAI211_X1 U16158 ( .C1(n14404), .C2(n14278), .A(n14277), .B(n14276), .ZN(
        n14343) );
  MUX2_X1 U16159 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14343), .S(n14720), .Z(
        P1_U3554) );
  INV_X1 U16160 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15323) );
  NAND3_X1 U16161 ( .A1(n14279), .A2(n14707), .A3(n14073), .ZN(n14281) );
  OAI211_X1 U16162 ( .C1(n14282), .C2(n14702), .A(n14281), .B(n14280), .ZN(
        n14283) );
  NOR2_X1 U16163 ( .A1(n14284), .A2(n14283), .ZN(n14344) );
  MUX2_X1 U16164 ( .A(n15323), .B(n14344), .S(n14720), .Z(n14285) );
  INV_X1 U16165 ( .A(n14285), .ZN(P1_U3553) );
  OAI211_X1 U16166 ( .C1(n14288), .C2(n14702), .A(n14287), .B(n14286), .ZN(
        n14347) );
  MUX2_X1 U16167 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14347), .S(n14720), .Z(
        P1_U3552) );
  AOI211_X1 U16168 ( .C1(n14697), .C2(n14291), .A(n14290), .B(n14289), .ZN(
        n14292) );
  OAI211_X1 U16169 ( .C1(n14404), .C2(n14294), .A(n14293), .B(n14292), .ZN(
        n14348) );
  MUX2_X1 U16170 ( .A(n14348), .B(P1_REG1_REG_23__SCAN_IN), .S(n14718), .Z(
        P1_U3551) );
  INV_X1 U16171 ( .A(n14295), .ZN(n14297) );
  OAI211_X1 U16172 ( .C1(n14702), .C2(n14298), .A(n14297), .B(n14296), .ZN(
        n14349) );
  MUX2_X1 U16173 ( .A(n14349), .B(P1_REG1_REG_22__SCAN_IN), .S(n14718), .Z(
        P1_U3550) );
  NAND2_X1 U16174 ( .A1(n14299), .A2(n14697), .ZN(n14300) );
  NAND4_X1 U16175 ( .A1(n14303), .A2(n14302), .A3(n14301), .A4(n14300), .ZN(
        n14350) );
  MUX2_X1 U16176 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14350), .S(n14720), .Z(
        P1_U3549) );
  NAND2_X1 U16177 ( .A1(n14304), .A2(n14697), .ZN(n14309) );
  NAND3_X1 U16178 ( .A1(n14306), .A2(n14305), .A3(n14707), .ZN(n14308) );
  NAND4_X1 U16179 ( .A1(n14310), .A2(n14309), .A3(n14308), .A4(n14307), .ZN(
        n14351) );
  MUX2_X1 U16180 ( .A(n14351), .B(P1_REG1_REG_20__SCAN_IN), .S(n14718), .Z(
        P1_U3548) );
  AOI211_X1 U16181 ( .C1(n14697), .C2(n14313), .A(n14312), .B(n14311), .ZN(
        n14314) );
  OAI211_X1 U16182 ( .C1(n14316), .C2(n14404), .A(n14315), .B(n14314), .ZN(
        n14352) );
  MUX2_X1 U16183 ( .A(n14352), .B(P1_REG1_REG_19__SCAN_IN), .S(n14718), .Z(
        P1_U3547) );
  OAI21_X1 U16184 ( .B1(n14318), .B2(n14702), .A(n14317), .ZN(n14319) );
  NOR2_X1 U16185 ( .A1(n14320), .A2(n14319), .ZN(n14353) );
  MUX2_X1 U16186 ( .A(n14321), .B(n14353), .S(n14720), .Z(n14322) );
  INV_X1 U16187 ( .A(n14322), .ZN(P1_U3546) );
  AOI211_X1 U16188 ( .C1(n14697), .C2(n12204), .A(n14324), .B(n14323), .ZN(
        n14326) );
  OAI211_X1 U16189 ( .C1(n14327), .C2(n14404), .A(n14326), .B(n14325), .ZN(
        n14355) );
  MUX2_X1 U16190 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14355), .S(n14720), .Z(
        P1_U3545) );
  AOI211_X1 U16191 ( .C1(n14697), .C2(n14330), .A(n14329), .B(n14328), .ZN(
        n14331) );
  OAI21_X1 U16192 ( .B1(n14404), .B2(n14332), .A(n14331), .ZN(n14356) );
  MUX2_X1 U16193 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14356), .S(n14720), .Z(
        P1_U3544) );
  AOI21_X1 U16194 ( .B1(n14697), .B2(n14334), .A(n14333), .ZN(n14335) );
  OAI211_X1 U16195 ( .C1(n14337), .C2(n14404), .A(n14336), .B(n14335), .ZN(
        n14357) );
  MUX2_X1 U16196 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14357), .S(n14720), .Z(
        P1_U3543) );
  MUX2_X1 U16197 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14338), .S(n14710), .Z(
        P1_U3527) );
  MUX2_X1 U16198 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14339), .S(n14710), .Z(
        P1_U3526) );
  MUX2_X1 U16199 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14341), .S(n14710), .Z(
        P1_U3524) );
  MUX2_X1 U16200 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14342), .S(n14710), .Z(
        P1_U3523) );
  MUX2_X1 U16201 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14343), .S(n14710), .Z(
        P1_U3522) );
  INV_X1 U16202 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n14345) );
  MUX2_X1 U16203 ( .A(n14345), .B(n14344), .S(n14710), .Z(n14346) );
  INV_X1 U16204 ( .A(n14346), .ZN(P1_U3521) );
  MUX2_X1 U16205 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14347), .S(n14710), .Z(
        P1_U3520) );
  MUX2_X1 U16206 ( .A(n14348), .B(P1_REG0_REG_23__SCAN_IN), .S(n14708), .Z(
        P1_U3519) );
  MUX2_X1 U16207 ( .A(n14349), .B(P1_REG0_REG_22__SCAN_IN), .S(n14708), .Z(
        P1_U3518) );
  MUX2_X1 U16208 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14350), .S(n14710), .Z(
        P1_U3517) );
  MUX2_X1 U16209 ( .A(n14351), .B(P1_REG0_REG_20__SCAN_IN), .S(n14708), .Z(
        P1_U3516) );
  MUX2_X1 U16210 ( .A(n14352), .B(P1_REG0_REG_19__SCAN_IN), .S(n14708), .Z(
        P1_U3515) );
  MUX2_X1 U16211 ( .A(n15270), .B(n14353), .S(n14710), .Z(n14354) );
  INV_X1 U16212 ( .A(n14354), .ZN(P1_U3513) );
  MUX2_X1 U16213 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14355), .S(n14710), .Z(
        P1_U3510) );
  MUX2_X1 U16214 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14356), .S(n14710), .Z(
        P1_U3507) );
  MUX2_X1 U16215 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14357), .S(n14710), .Z(
        P1_U3504) );
  NOR4_X1 U16216 ( .A1(n14358), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9287), .A4(
        P1_U3086), .ZN(n14359) );
  AOI21_X1 U16217 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14360), .A(n14359), 
        .ZN(n14361) );
  OAI21_X1 U16218 ( .B1(n14362), .B2(n14369), .A(n14361), .ZN(P1_U3324) );
  OAI222_X1 U16219 ( .A1(n14369), .A2(n14365), .B1(n14364), .B2(P1_U3086), 
        .C1(n14363), .C2(n14366), .ZN(P1_U3326) );
  OAI222_X1 U16220 ( .A1(P1_U3086), .A2(n14370), .B1(n14369), .B2(n14368), 
        .C1(n14367), .C2(n14366), .ZN(P1_U3328) );
  MUX2_X1 U16221 ( .A(n14372), .B(n14371), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16222 ( .A(n14373), .B(n14566), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  XNOR2_X1 U16223 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14374), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16224 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14375) );
  OAI21_X1 U16225 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n14375), 
        .ZN(U28) );
  AOI21_X1 U16226 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14376) );
  OAI21_X1 U16227 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14376), 
        .ZN(U29) );
  NOR2_X1 U16228 ( .A1(n14378), .A2(n14377), .ZN(n14379) );
  XOR2_X1 U16229 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n14379), .Z(SUB_1596_U61) );
  INV_X1 U16230 ( .A(SI_9_), .ZN(n14380) );
  OAI22_X1 U16231 ( .A1(n14381), .A2(n15458), .B1(n14380), .B2(n15456), .ZN(
        n14382) );
  INV_X1 U16232 ( .A(n14382), .ZN(n14383) );
  OAI21_X1 U16233 ( .B1(P3_U3151), .B2(n14384), .A(n14383), .ZN(P3_U3286) );
  INV_X1 U16234 ( .A(n14385), .ZN(n14388) );
  AOI22_X1 U16235 ( .A1(n14388), .A2(n14387), .B1(SI_12_), .B2(n14386), .ZN(
        n14389) );
  OAI21_X1 U16236 ( .B1(P3_U3151), .B2(n14390), .A(n14389), .ZN(P3_U3283) );
  XOR2_X1 U16237 ( .A(n14392), .B(n14391), .Z(SUB_1596_U57) );
  XNOR2_X1 U16238 ( .A(n14393), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  AOI21_X1 U16239 ( .B1(n14396), .B2(n14395), .A(n14394), .ZN(n14397) );
  XOR2_X1 U16240 ( .A(n14397), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  NOR2_X1 U16241 ( .A1(n14399), .A2(n14398), .ZN(n14400) );
  XOR2_X1 U16242 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14400), .Z(SUB_1596_U70)
         );
  NAND2_X1 U16243 ( .A1(n14401), .A2(n14697), .ZN(n14402) );
  AND2_X1 U16244 ( .A1(n14403), .A2(n14402), .ZN(n14407) );
  OR2_X1 U16245 ( .A1(n14405), .A2(n14404), .ZN(n14406) );
  INV_X1 U16246 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U16247 ( .A1(n14710), .A2(n14410), .B1(n14409), .B2(n14708), .ZN(
        P1_U3495) );
  AOI22_X1 U16248 ( .A1(n14720), .A2(n14410), .B1(n10304), .B2(n14718), .ZN(
        P1_U3540) );
  NOR2_X1 U16249 ( .A1(n14412), .A2(n14411), .ZN(n14413) );
  XOR2_X1 U16250 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14413), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16251 ( .B1(n14416), .B2(n14415), .A(n14414), .ZN(n14417) );
  OAI21_X1 U16252 ( .B1(n14419), .B2(n14418), .A(n14417), .ZN(n14431) );
  OR2_X1 U16253 ( .A1(n14421), .A2(n14420), .ZN(n14424) );
  NAND2_X1 U16254 ( .A1(n14424), .A2(n14422), .ZN(n14429) );
  NAND2_X1 U16255 ( .A1(n14424), .A2(n14423), .ZN(n14426) );
  NAND2_X1 U16256 ( .A1(n14426), .A2(n14425), .ZN(n14428) );
  AOI21_X1 U16257 ( .B1(n14429), .B2(n14428), .A(n14427), .ZN(n14430) );
  AOI211_X1 U16258 ( .C1(n14441), .C2(n14481), .A(n14431), .B(n14430), .ZN(
        n14432) );
  OAI21_X1 U16259 ( .B1(n14434), .B2(n14433), .A(n14432), .ZN(P3_U3155) );
  NAND2_X1 U16260 ( .A1(n14436), .A2(n14435), .ZN(n14437) );
  NAND2_X1 U16261 ( .A1(n14438), .A2(n14437), .ZN(n14440) );
  AOI222_X1 U16262 ( .A1(n14444), .A2(n14443), .B1(n14442), .B2(n14441), .C1(
        n14440), .C2(n14439), .ZN(n14445) );
  NAND2_X1 U16263 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14463)
         );
  OAI211_X1 U16264 ( .C1(n14447), .C2(n14446), .A(n14445), .B(n14463), .ZN(
        P3_U3166) );
  AOI22_X1 U16265 ( .A1(n15021), .A2(n14448), .B1(n14990), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14465) );
  OAI21_X1 U16266 ( .B1(n14451), .B2(n14450), .A(n14449), .ZN(n14458) );
  INV_X1 U16267 ( .A(n14452), .ZN(n14454) );
  NAND2_X1 U16268 ( .A1(n14454), .A2(n14453), .ZN(n14455) );
  XNOR2_X1 U16269 ( .A(n14456), .B(n14455), .ZN(n14457) );
  AOI22_X1 U16270 ( .A1(n14458), .A2(n15023), .B1(n15031), .B2(n14457), .ZN(
        n14464) );
  OAI221_X1 U16271 ( .B1(n14461), .B2(n14460), .C1(n14461), .C2(n14459), .A(
        n14474), .ZN(n14462) );
  NAND4_X1 U16272 ( .A1(n14465), .A2(n14464), .A3(n14463), .A4(n14462), .ZN(
        P3_U3198) );
  AOI22_X1 U16273 ( .A1(n15021), .A2(n14466), .B1(n14990), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14480) );
  XNOR2_X1 U16274 ( .A(n14467), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n14472) );
  AOI211_X1 U16275 ( .C1(n14470), .C2(n14469), .A(n15010), .B(n14468), .ZN(
        n14471) );
  AOI21_X1 U16276 ( .B1(n14472), .B2(n15023), .A(n14471), .ZN(n14479) );
  NAND2_X1 U16277 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14478)
         );
  OAI221_X1 U16278 ( .B1(n14473), .B2(n14476), .C1(n14473), .C2(n14475), .A(
        n14474), .ZN(n14477) );
  NAND4_X1 U16279 ( .A1(n14480), .A2(n14479), .A3(n14478), .A4(n14477), .ZN(
        P3_U3199) );
  INV_X1 U16280 ( .A(n14481), .ZN(n14482) );
  OAI22_X1 U16281 ( .A1(n14483), .A2(n14498), .B1(n14482), .B2(n15124), .ZN(
        n14484) );
  NOR2_X1 U16282 ( .A1(n14485), .A2(n14484), .ZN(n14503) );
  INV_X1 U16283 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U16284 ( .A1(n15144), .A2(n14503), .B1(n14486), .B2(n15141), .ZN(
        P3_U3473) );
  NOR2_X1 U16285 ( .A1(n14487), .A2(n14498), .ZN(n14489) );
  AOI211_X1 U16286 ( .C1(n14490), .C2(n15105), .A(n14489), .B(n14488), .ZN(
        n14504) );
  INV_X1 U16287 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U16288 ( .A1(n15144), .A2(n14504), .B1(n14491), .B2(n15141), .ZN(
        P3_U3472) );
  OAI22_X1 U16289 ( .A1(n14493), .A2(n14498), .B1(n15124), .B2(n14492), .ZN(
        n14494) );
  NOR2_X1 U16290 ( .A1(n14495), .A2(n14494), .ZN(n14505) );
  AOI22_X1 U16291 ( .A1(n15144), .A2(n14505), .B1(n14496), .B2(n15141), .ZN(
        P3_U3471) );
  OAI22_X1 U16292 ( .A1(n14499), .A2(n14498), .B1(n14497), .B2(n15124), .ZN(
        n14500) );
  NOR2_X1 U16293 ( .A1(n14501), .A2(n14500), .ZN(n14506) );
  INV_X1 U16294 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U16295 ( .A1(n15144), .A2(n14506), .B1(n14502), .B2(n15141), .ZN(
        P3_U3470) );
  AOI22_X1 U16296 ( .A1(n15130), .A2(n14503), .B1(n8027), .B2(n8319), .ZN(
        P3_U3432) );
  AOI22_X1 U16297 ( .A1(n15130), .A2(n14504), .B1(n8014), .B2(n8319), .ZN(
        P3_U3429) );
  AOI22_X1 U16298 ( .A1(n15130), .A2(n14505), .B1(n8001), .B2(n8319), .ZN(
        P3_U3426) );
  AOI22_X1 U16299 ( .A1(n15130), .A2(n14506), .B1(n7981), .B2(n8319), .ZN(
        P3_U3423) );
  XNOR2_X1 U16300 ( .A(n14507), .B(n9475), .ZN(n14509) );
  AOI21_X1 U16301 ( .B1(n14509), .B2(n14611), .A(n14508), .ZN(n14526) );
  INV_X1 U16302 ( .A(n14510), .ZN(n14511) );
  AOI222_X1 U16303 ( .A1(n14513), .A2(n14512), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n14642), .C1(n14599), .C2(n14511), .ZN(n14523) );
  INV_X1 U16304 ( .A(n14514), .ZN(n14515) );
  AOI21_X1 U16305 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n14529) );
  INV_X1 U16306 ( .A(n14518), .ZN(n14520) );
  OAI211_X1 U16307 ( .C1(n14525), .C2(n14520), .A(n14622), .B(n14519), .ZN(
        n14524) );
  INV_X1 U16308 ( .A(n14524), .ZN(n14521) );
  AOI22_X1 U16309 ( .A1(n14529), .A2(n14627), .B1(n14626), .B2(n14521), .ZN(
        n14522) );
  OAI211_X1 U16310 ( .C1(n14642), .C2(n14526), .A(n14523), .B(n14522), .ZN(
        P1_U3279) );
  OAI21_X1 U16311 ( .B1(n14525), .B2(n14702), .A(n14524), .ZN(n14528) );
  INV_X1 U16312 ( .A(n14526), .ZN(n14527) );
  AOI211_X1 U16313 ( .C1(n14707), .C2(n14529), .A(n14528), .B(n14527), .ZN(
        n14538) );
  AOI22_X1 U16314 ( .A1(n14720), .A2(n14538), .B1(n9467), .B2(n14718), .ZN(
        P1_U3542) );
  OR2_X1 U16315 ( .A1(n14530), .A2(n14702), .ZN(n14531) );
  AND2_X1 U16316 ( .A1(n14532), .A2(n14531), .ZN(n14535) );
  NAND2_X1 U16317 ( .A1(n14533), .A2(n14707), .ZN(n14534) );
  AND3_X1 U16318 ( .A1(n14536), .A2(n14535), .A3(n14534), .ZN(n14540) );
  AOI22_X1 U16319 ( .A1(n14720), .A2(n14540), .B1(n9423), .B2(n14718), .ZN(
        P1_U3539) );
  INV_X1 U16320 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14537) );
  AOI22_X1 U16321 ( .A1(n14710), .A2(n14538), .B1(n14537), .B2(n14708), .ZN(
        P1_U3501) );
  INV_X1 U16322 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14539) );
  AOI22_X1 U16323 ( .A1(n14710), .A2(n14540), .B1(n14539), .B2(n14708), .ZN(
        P1_U3492) );
  AOI21_X1 U16324 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(n14545) );
  XNOR2_X1 U16325 ( .A(n14545), .B(n14544), .ZN(SUB_1596_U69) );
  AOI21_X1 U16326 ( .B1(n14548), .B2(n14547), .A(n14546), .ZN(n14549) );
  XNOR2_X1 U16327 ( .A(n14549), .B(n14768), .ZN(SUB_1596_U68) );
  NOR2_X1 U16328 ( .A1(n14551), .A2(n14550), .ZN(n14552) );
  XOR2_X1 U16329 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14552), .Z(SUB_1596_U67)
         );
  NOR2_X1 U16330 ( .A1(n14554), .A2(n14553), .ZN(n14555) );
  XOR2_X1 U16331 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14555), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16332 ( .B1(n14558), .B2(n14557), .A(n14556), .ZN(n14559) );
  XNOR2_X1 U16333 ( .A(n14559), .B(n15321), .ZN(SUB_1596_U65) );
  NOR2_X1 U16334 ( .A1(n14561), .A2(n14560), .ZN(n14562) );
  XOR2_X1 U16335 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14562), .Z(SUB_1596_U64)
         );
  OAI21_X1 U16336 ( .B1(n14564), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14563), .ZN(
        n14565) );
  XOR2_X1 U16337 ( .A(n14566), .B(n14565), .Z(n14571) );
  AOI22_X1 U16338 ( .A1(n14568), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14569) );
  OAI21_X1 U16339 ( .B1(n14571), .B2(n14570), .A(n14569), .ZN(P1_U3243) );
  AOI21_X1 U16340 ( .B1(n14573), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14572), 
        .ZN(n14577) );
  AOI21_X1 U16341 ( .B1(n14575), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14574), 
        .ZN(n14576) );
  OAI222_X1 U16342 ( .A1(n14592), .A2(n14578), .B1(n14590), .B2(n14577), .C1(
        n14588), .C2(n14576), .ZN(n14579) );
  INV_X1 U16343 ( .A(n14579), .ZN(n14581) );
  OAI211_X1 U16344 ( .C1(n14582), .C2(n14596), .A(n14581), .B(n14580), .ZN(
        P1_U3258) );
  OAI21_X1 U16345 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n14584), .A(n14583), 
        .ZN(n14589) );
  OAI21_X1 U16346 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n14586), .A(n14585), 
        .ZN(n14587) );
  OAI222_X1 U16347 ( .A1(n14592), .A2(n14591), .B1(n14590), .B2(n14589), .C1(
        n14588), .C2(n14587), .ZN(n14593) );
  INV_X1 U16348 ( .A(n14593), .ZN(n14595) );
  OAI211_X1 U16349 ( .C1(n14597), .C2(n14596), .A(n14595), .B(n14594), .ZN(
        P1_U3261) );
  NAND2_X1 U16350 ( .A1(n14598), .A2(n14626), .ZN(n14602) );
  AOI22_X1 U16351 ( .A1(n14642), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n14600), 
        .B2(n14599), .ZN(n14601) );
  OAI211_X1 U16352 ( .C1(n14603), .C2(n14616), .A(n14602), .B(n14601), .ZN(
        n14604) );
  AOI21_X1 U16353 ( .B1(n14605), .B2(n14627), .A(n14604), .ZN(n14606) );
  OAI21_X1 U16354 ( .B1(n14642), .B2(n14607), .A(n14606), .ZN(P1_U3283) );
  XNOR2_X1 U16355 ( .A(n14608), .B(n14618), .ZN(n14612) );
  INV_X1 U16356 ( .A(n14609), .ZN(n14610) );
  AOI21_X1 U16357 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14685) );
  NOR2_X1 U16358 ( .A1(n14637), .A2(n14613), .ZN(n14614) );
  AOI21_X1 U16359 ( .B1(n14642), .B2(P1_REG2_REG_4__SCAN_IN), .A(n14614), .ZN(
        n14615) );
  OAI21_X1 U16360 ( .B1(n14616), .B2(n14684), .A(n14615), .ZN(n14617) );
  INV_X1 U16361 ( .A(n14617), .ZN(n14629) );
  XOR2_X1 U16362 ( .A(n14619), .B(n14618), .Z(n14688) );
  INV_X1 U16363 ( .A(n14620), .ZN(n14624) );
  INV_X1 U16364 ( .A(n14621), .ZN(n14623) );
  OAI211_X1 U16365 ( .C1(n14684), .C2(n14624), .A(n14623), .B(n14622), .ZN(
        n14683) );
  INV_X1 U16366 ( .A(n14683), .ZN(n14625) );
  AOI22_X1 U16367 ( .A1(n14688), .A2(n14627), .B1(n14626), .B2(n14625), .ZN(
        n14628) );
  OAI211_X1 U16368 ( .C1(n14642), .C2(n14685), .A(n14629), .B(n14628), .ZN(
        P1_U3289) );
  NAND2_X1 U16369 ( .A1(n14631), .A2(n14630), .ZN(n14633) );
  NAND2_X1 U16370 ( .A1(n14633), .A2(n14632), .ZN(n14634) );
  OAI211_X1 U16371 ( .C1(n14637), .C2(n14636), .A(n14635), .B(n14634), .ZN(
        n14638) );
  INV_X1 U16372 ( .A(n14638), .ZN(n14641) );
  NOR2_X1 U16373 ( .A1(n14642), .A2(n14639), .ZN(n14640) );
  AOI22_X1 U16374 ( .A1(n9297), .A2(n14642), .B1(n14641), .B2(n14640), .ZN(
        P1_U3293) );
  INV_X1 U16375 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14643) );
  NOR2_X1 U16376 ( .A1(n14669), .A2(n14643), .ZN(P1_U3294) );
  INV_X1 U16377 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14644) );
  NOR2_X1 U16378 ( .A1(n14669), .A2(n14644), .ZN(P1_U3295) );
  INV_X1 U16379 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14645) );
  NOR2_X1 U16380 ( .A1(n14669), .A2(n14645), .ZN(P1_U3296) );
  INV_X1 U16381 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14646) );
  NOR2_X1 U16382 ( .A1(n14669), .A2(n14646), .ZN(P1_U3297) );
  INV_X1 U16383 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14647) );
  NOR2_X1 U16384 ( .A1(n14669), .A2(n14647), .ZN(P1_U3298) );
  INV_X1 U16385 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14648) );
  NOR2_X1 U16386 ( .A1(n14669), .A2(n14648), .ZN(P1_U3299) );
  NOR2_X1 U16387 ( .A1(n14669), .A2(n15372), .ZN(P1_U3300) );
  INV_X1 U16388 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14649) );
  NOR2_X1 U16389 ( .A1(n14669), .A2(n14649), .ZN(P1_U3301) );
  INV_X1 U16390 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14650) );
  NOR2_X1 U16391 ( .A1(n14669), .A2(n14650), .ZN(P1_U3302) );
  INV_X1 U16392 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14651) );
  NOR2_X1 U16393 ( .A1(n14669), .A2(n14651), .ZN(P1_U3303) );
  INV_X1 U16394 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14652) );
  NOR2_X1 U16395 ( .A1(n14669), .A2(n14652), .ZN(P1_U3304) );
  INV_X1 U16396 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14653) );
  NOR2_X1 U16397 ( .A1(n14669), .A2(n14653), .ZN(P1_U3305) );
  INV_X1 U16398 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14654) );
  NOR2_X1 U16399 ( .A1(n14669), .A2(n14654), .ZN(P1_U3306) );
  INV_X1 U16400 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14655) );
  NOR2_X1 U16401 ( .A1(n14669), .A2(n14655), .ZN(P1_U3307) );
  INV_X1 U16402 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14656) );
  NOR2_X1 U16403 ( .A1(n14669), .A2(n14656), .ZN(P1_U3308) );
  INV_X1 U16404 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14657) );
  NOR2_X1 U16405 ( .A1(n14669), .A2(n14657), .ZN(P1_U3309) );
  NOR2_X1 U16406 ( .A1(n14669), .A2(n15229), .ZN(P1_U3310) );
  NOR2_X1 U16407 ( .A1(n14669), .A2(n15310), .ZN(P1_U3311) );
  INV_X1 U16408 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14658) );
  NOR2_X1 U16409 ( .A1(n14669), .A2(n14658), .ZN(P1_U3312) );
  INV_X1 U16410 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14659) );
  NOR2_X1 U16411 ( .A1(n14669), .A2(n14659), .ZN(P1_U3313) );
  INV_X1 U16412 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14660) );
  NOR2_X1 U16413 ( .A1(n14669), .A2(n14660), .ZN(P1_U3314) );
  INV_X1 U16414 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14661) );
  NOR2_X1 U16415 ( .A1(n14669), .A2(n14661), .ZN(P1_U3315) );
  NOR2_X1 U16416 ( .A1(n14669), .A2(n15418), .ZN(P1_U3316) );
  INV_X1 U16417 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14662) );
  NOR2_X1 U16418 ( .A1(n14669), .A2(n14662), .ZN(P1_U3317) );
  INV_X1 U16419 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14663) );
  NOR2_X1 U16420 ( .A1(n14669), .A2(n14663), .ZN(P1_U3318) );
  INV_X1 U16421 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14664) );
  NOR2_X1 U16422 ( .A1(n14669), .A2(n14664), .ZN(P1_U3319) );
  INV_X1 U16423 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14665) );
  NOR2_X1 U16424 ( .A1(n14669), .A2(n14665), .ZN(P1_U3320) );
  INV_X1 U16425 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14666) );
  NOR2_X1 U16426 ( .A1(n14669), .A2(n14666), .ZN(P1_U3321) );
  INV_X1 U16427 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14667) );
  NOR2_X1 U16428 ( .A1(n14669), .A2(n14667), .ZN(P1_U3322) );
  INV_X1 U16429 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14668) );
  NOR2_X1 U16430 ( .A1(n14669), .A2(n14668), .ZN(P1_U3323) );
  INV_X1 U16431 ( .A(n14670), .ZN(n14671) );
  OAI21_X1 U16432 ( .B1(n14672), .B2(n14702), .A(n14671), .ZN(n14674) );
  AOI211_X1 U16433 ( .C1(n14707), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14711) );
  INV_X1 U16434 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15434) );
  AOI22_X1 U16435 ( .A1(n14710), .A2(n14711), .B1(n15434), .B2(n14708), .ZN(
        P1_U3462) );
  INV_X1 U16436 ( .A(n14676), .ZN(n14681) );
  OAI21_X1 U16437 ( .B1(n7439), .B2(n14702), .A(n14677), .ZN(n14680) );
  INV_X1 U16438 ( .A(n14678), .ZN(n14679) );
  AOI211_X1 U16439 ( .C1(n14707), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        n14712) );
  INV_X1 U16440 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14682) );
  AOI22_X1 U16441 ( .A1(n14710), .A2(n14712), .B1(n14682), .B2(n14708), .ZN(
        P1_U3468) );
  OAI21_X1 U16442 ( .B1(n14684), .B2(n14702), .A(n14683), .ZN(n14687) );
  INV_X1 U16443 ( .A(n14685), .ZN(n14686) );
  AOI211_X1 U16444 ( .C1(n14707), .C2(n14688), .A(n14687), .B(n14686), .ZN(
        n14713) );
  INV_X1 U16445 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14689) );
  AOI22_X1 U16446 ( .A1(n14710), .A2(n14713), .B1(n14689), .B2(n14708), .ZN(
        P1_U3471) );
  AOI211_X1 U16447 ( .C1(n14697), .C2(n14692), .A(n14691), .B(n14690), .ZN(
        n14715) );
  INV_X1 U16448 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14693) );
  AOI22_X1 U16449 ( .A1(n14710), .A2(n14715), .B1(n14693), .B2(n14708), .ZN(
        P1_U3474) );
  AOI211_X1 U16450 ( .C1(n14697), .C2(n14696), .A(n14695), .B(n14694), .ZN(
        n14717) );
  INV_X1 U16451 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U16452 ( .A1(n14710), .A2(n14717), .B1(n14698), .B2(n14708), .ZN(
        P1_U3477) );
  INV_X1 U16453 ( .A(n14699), .ZN(n14701) );
  OAI211_X1 U16454 ( .C1(n14703), .C2(n14702), .A(n14701), .B(n14700), .ZN(
        n14705) );
  AOI211_X1 U16455 ( .C1(n14707), .C2(n14706), .A(n14705), .B(n14704), .ZN(
        n14719) );
  INV_X1 U16456 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14709) );
  AOI22_X1 U16457 ( .A1(n14710), .A2(n14719), .B1(n14709), .B2(n14708), .ZN(
        P1_U3483) );
  AOI22_X1 U16458 ( .A1(n14720), .A2(n14711), .B1(n10084), .B2(n14718), .ZN(
        P1_U3529) );
  AOI22_X1 U16459 ( .A1(n14720), .A2(n14712), .B1(n10089), .B2(n14718), .ZN(
        P1_U3531) );
  AOI22_X1 U16460 ( .A1(n14720), .A2(n14713), .B1(n9330), .B2(n14718), .ZN(
        P1_U3532) );
  AOI22_X1 U16461 ( .A1(n14720), .A2(n14715), .B1(n14714), .B2(n14718), .ZN(
        P1_U3533) );
  AOI22_X1 U16462 ( .A1(n14720), .A2(n14717), .B1(n14716), .B2(n14718), .ZN(
        P1_U3534) );
  AOI22_X1 U16463 ( .A1(n14720), .A2(n14719), .B1(n10117), .B2(n14718), .ZN(
        P1_U3536) );
  NOR2_X1 U16464 ( .A1(n14788), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16465 ( .A(n14721), .ZN(n14722) );
  OAI21_X1 U16466 ( .B1(n14795), .B2(n14723), .A(n14722), .ZN(n14724) );
  AOI21_X1 U16467 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(n14788), .A(n14724), .ZN(
        n14734) );
  AOI211_X1 U16468 ( .C1(n14727), .C2(n14726), .A(n14744), .B(n14725), .ZN(
        n14728) );
  INV_X1 U16469 ( .A(n14728), .ZN(n14733) );
  OAI211_X1 U16470 ( .C1(n14731), .C2(n14730), .A(n14782), .B(n14729), .ZN(
        n14732) );
  NAND3_X1 U16471 ( .A1(n14734), .A2(n14733), .A3(n14732), .ZN(P2_U3220) );
  NAND2_X1 U16472 ( .A1(n14788), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n14737) );
  INV_X1 U16473 ( .A(n14735), .ZN(n14736) );
  OAI211_X1 U16474 ( .C1(n14795), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        n14739) );
  INV_X1 U16475 ( .A(n14739), .ZN(n14750) );
  OAI211_X1 U16476 ( .C1(n14742), .C2(n14741), .A(n14782), .B(n14740), .ZN(
        n14749) );
  AOI211_X1 U16477 ( .C1(n14746), .C2(n14745), .A(n14744), .B(n14743), .ZN(
        n14747) );
  INV_X1 U16478 ( .A(n14747), .ZN(n14748) );
  NAND3_X1 U16479 ( .A1(n14750), .A2(n14749), .A3(n14748), .ZN(P2_U3222) );
  NOR3_X1 U16480 ( .A1(n14753), .A2(n14752), .A3(n14751), .ZN(n14755) );
  OAI21_X1 U16481 ( .B1(n14755), .B2(n14754), .A(n14790), .ZN(n14762) );
  AOI21_X1 U16482 ( .B1(n14758), .B2(n14757), .A(n14756), .ZN(n14760) );
  OAI21_X1 U16483 ( .B1(n14760), .B2(n14759), .A(n14782), .ZN(n14761) );
  OAI211_X1 U16484 ( .C1(n14795), .C2(n14763), .A(n14762), .B(n14761), .ZN(
        n14764) );
  INV_X1 U16485 ( .A(n14764), .ZN(n14766) );
  OAI211_X1 U16486 ( .C1(n14768), .C2(n14767), .A(n14766), .B(n14765), .ZN(
        P2_U3226) );
  OAI211_X1 U16487 ( .C1(n14771), .C2(n14770), .A(n14769), .B(n14782), .ZN(
        n14772) );
  NAND2_X1 U16488 ( .A1(n14773), .A2(n14772), .ZN(n14774) );
  AOI21_X1 U16489 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n14788), .A(n14774), 
        .ZN(n14779) );
  OAI211_X1 U16490 ( .C1(n14777), .C2(n14776), .A(n14775), .B(n14790), .ZN(
        n14778) );
  OAI211_X1 U16491 ( .C1(n14795), .C2(n14780), .A(n14779), .B(n14778), .ZN(
        P2_U3227) );
  OAI211_X1 U16492 ( .C1(n14784), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        n14785) );
  NAND2_X1 U16493 ( .A1(n14786), .A2(n14785), .ZN(n14787) );
  AOI21_X1 U16494 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n14788), .A(n14787), 
        .ZN(n14793) );
  OAI211_X1 U16495 ( .C1(n14791), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14790), 
        .B(n14789), .ZN(n14792) );
  OAI211_X1 U16496 ( .C1(n14795), .C2(n14794), .A(n14793), .B(n14792), .ZN(
        P2_U3228) );
  NAND2_X1 U16497 ( .A1(n14798), .A2(n14797), .ZN(n14802) );
  AOI22_X1 U16498 ( .A1(n13469), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14800), 
        .B2(n14799), .ZN(n14801) );
  OAI211_X1 U16499 ( .C1(n7124), .C2(n14803), .A(n14802), .B(n14801), .ZN(
        n14804) );
  AOI21_X1 U16500 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14807) );
  OAI21_X1 U16501 ( .B1(n14809), .B2(n14808), .A(n14807), .ZN(P2_U3258) );
  AND2_X1 U16502 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14811), .ZN(P2_U3266) );
  AND2_X1 U16503 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14811), .ZN(P2_U3267) );
  AND2_X1 U16504 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14811), .ZN(P2_U3268) );
  NOR2_X1 U16505 ( .A1(n14814), .A2(n15341), .ZN(P2_U3269) );
  AND2_X1 U16506 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14811), .ZN(P2_U3270) );
  AND2_X1 U16507 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14811), .ZN(P2_U3271) );
  AND2_X1 U16508 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14811), .ZN(P2_U3272) );
  AND2_X1 U16509 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14811), .ZN(P2_U3273) );
  AND2_X1 U16510 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14811), .ZN(P2_U3274) );
  AND2_X1 U16511 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14811), .ZN(P2_U3275) );
  AND2_X1 U16512 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14811), .ZN(P2_U3276) );
  AND2_X1 U16513 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14811), .ZN(P2_U3277) );
  AND2_X1 U16514 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14811), .ZN(P2_U3278) );
  AND2_X1 U16515 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14811), .ZN(P2_U3279) );
  AND2_X1 U16516 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14811), .ZN(P2_U3280) );
  AND2_X1 U16517 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14811), .ZN(P2_U3281) );
  AND2_X1 U16518 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14811), .ZN(P2_U3282) );
  NOR2_X1 U16519 ( .A1(n14814), .A2(n15304), .ZN(P2_U3283) );
  AND2_X1 U16520 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14811), .ZN(P2_U3284) );
  AND2_X1 U16521 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14811), .ZN(P2_U3285) );
  AND2_X1 U16522 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14811), .ZN(P2_U3286) );
  AND2_X1 U16523 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14811), .ZN(P2_U3287) );
  AND2_X1 U16524 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14811), .ZN(P2_U3288) );
  AND2_X1 U16525 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14811), .ZN(P2_U3289) );
  AND2_X1 U16526 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14811), .ZN(P2_U3290) );
  AND2_X1 U16527 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14811), .ZN(P2_U3291) );
  AND2_X1 U16528 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14811), .ZN(P2_U3292) );
  NOR2_X1 U16529 ( .A1(n14814), .A2(n15397), .ZN(P2_U3293) );
  NOR2_X1 U16530 ( .A1(n14814), .A2(n15371), .ZN(P2_U3294) );
  AND2_X1 U16531 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14811), .ZN(P2_U3295) );
  AOI22_X1 U16532 ( .A1(n14814), .A2(n14813), .B1(n14812), .B2(n14811), .ZN(
        P2_U3416) );
  AOI22_X1 U16533 ( .A1(n14818), .A2(n14817), .B1(n14816), .B2(n14815), .ZN(
        P2_U3417) );
  AOI211_X1 U16534 ( .C1(n14821), .C2(n14877), .A(n14820), .B(n14819), .ZN(
        n14881) );
  INV_X1 U16535 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14822) );
  AOI22_X1 U16536 ( .A1(n14880), .A2(n14881), .B1(n14822), .B2(n14878), .ZN(
        P2_U3430) );
  AOI21_X1 U16537 ( .B1(n14847), .B2(n6560), .A(n14823), .ZN(n14824) );
  OAI211_X1 U16538 ( .C1(n14827), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        n14828) );
  INV_X1 U16539 ( .A(n14828), .ZN(n14882) );
  INV_X1 U16540 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14829) );
  AOI22_X1 U16541 ( .A1(n14880), .A2(n14882), .B1(n14829), .B2(n14878), .ZN(
        P2_U3433) );
  AOI21_X1 U16542 ( .B1(n14847), .B2(n14831), .A(n14830), .ZN(n14832) );
  OAI211_X1 U16543 ( .C1(n14840), .C2(n14834), .A(n14833), .B(n14832), .ZN(
        n14835) );
  INV_X1 U16544 ( .A(n14835), .ZN(n14883) );
  INV_X1 U16545 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14836) );
  AOI22_X1 U16546 ( .A1(n14880), .A2(n14883), .B1(n14836), .B2(n14878), .ZN(
        P2_U3436) );
  AND2_X1 U16547 ( .A1(n14837), .A2(n14847), .ZN(n14838) );
  NOR2_X1 U16548 ( .A1(n14839), .A2(n14838), .ZN(n14843) );
  OR2_X1 U16549 ( .A1(n14841), .A2(n14840), .ZN(n14842) );
  AND3_X1 U16550 ( .A1(n14844), .A2(n14843), .A3(n14842), .ZN(n14884) );
  INV_X1 U16551 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14845) );
  AOI22_X1 U16552 ( .A1(n14880), .A2(n14884), .B1(n14845), .B2(n14878), .ZN(
        P2_U3439) );
  NAND2_X1 U16553 ( .A1(n14846), .A2(n14877), .ZN(n14853) );
  NAND2_X1 U16554 ( .A1(n14846), .A2(n14862), .ZN(n14852) );
  NAND2_X1 U16555 ( .A1(n14848), .A2(n14847), .ZN(n14849) );
  AND2_X1 U16556 ( .A1(n14850), .A2(n14849), .ZN(n14851) );
  INV_X1 U16557 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14855) );
  AOI22_X1 U16558 ( .A1(n14880), .A2(n14885), .B1(n14855), .B2(n14878), .ZN(
        P2_U3442) );
  NAND2_X1 U16559 ( .A1(n14861), .A2(n14877), .ZN(n14857) );
  OAI211_X1 U16560 ( .C1(n14858), .C2(n14872), .A(n14857), .B(n14856), .ZN(
        n14859) );
  AOI211_X1 U16561 ( .C1(n14862), .C2(n14861), .A(n14860), .B(n14859), .ZN(
        n14886) );
  INV_X1 U16562 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14863) );
  AOI22_X1 U16563 ( .A1(n14880), .A2(n14886), .B1(n14863), .B2(n14878), .ZN(
        P2_U3445) );
  OAI21_X1 U16564 ( .B1(n14865), .B2(n14872), .A(n14864), .ZN(n14867) );
  AOI211_X1 U16565 ( .C1(n14877), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14887) );
  INV_X1 U16566 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U16567 ( .A1(n14880), .A2(n14887), .B1(n14869), .B2(n14878), .ZN(
        P2_U3454) );
  INV_X1 U16568 ( .A(n14870), .ZN(n14876) );
  OAI21_X1 U16569 ( .B1(n14873), .B2(n14872), .A(n14871), .ZN(n14875) );
  AOI211_X1 U16570 ( .C1(n14877), .C2(n14876), .A(n14875), .B(n14874), .ZN(
        n14890) );
  INV_X1 U16571 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14879) );
  AOI22_X1 U16572 ( .A1(n14880), .A2(n14890), .B1(n14879), .B2(n14878), .ZN(
        P2_U3460) );
  AOI22_X1 U16573 ( .A1(n14891), .A2(n14881), .B1(n8381), .B2(n14888), .ZN(
        P2_U3499) );
  AOI22_X1 U16574 ( .A1(n14891), .A2(n14882), .B1(n10148), .B2(n14888), .ZN(
        P2_U3500) );
  AOI22_X1 U16575 ( .A1(n14891), .A2(n14883), .B1(n10150), .B2(n14888), .ZN(
        P2_U3501) );
  AOI22_X1 U16576 ( .A1(n14891), .A2(n14884), .B1(n10153), .B2(n14888), .ZN(
        P2_U3502) );
  AOI22_X1 U16577 ( .A1(n14891), .A2(n14885), .B1(n10157), .B2(n14888), .ZN(
        P2_U3503) );
  AOI22_X1 U16578 ( .A1(n14891), .A2(n14886), .B1(n10158), .B2(n14888), .ZN(
        P2_U3504) );
  AOI22_X1 U16579 ( .A1(n14891), .A2(n14887), .B1(n10267), .B2(n14888), .ZN(
        P2_U3507) );
  AOI22_X1 U16580 ( .A1(n14891), .A2(n14890), .B1(n14889), .B2(n14888), .ZN(
        P2_U3509) );
  NOR2_X1 U16581 ( .A1(P3_U3897), .A2(n14990), .ZN(P3_U3150) );
  NOR2_X1 U16582 ( .A1(n14892), .A2(n6922), .ZN(n14894) );
  NAND3_X1 U16583 ( .A1(n15036), .A2(n14908), .A3(n15010), .ZN(n14893) );
  OAI21_X1 U16584 ( .B1(n14895), .B2(n14894), .A(n14893), .ZN(n14898) );
  AOI22_X1 U16585 ( .A1(n15021), .A2(n6922), .B1(P3_REG3_REG_0__SCAN_IN), .B2(
        P3_U3151), .ZN(n14897) );
  OAI211_X1 U16586 ( .C1(n14899), .C2(n15041), .A(n14898), .B(n14897), .ZN(
        P3_U3182) );
  INV_X1 U16587 ( .A(n14900), .ZN(n14901) );
  NAND3_X1 U16588 ( .A1(n14903), .A2(n14902), .A3(n14901), .ZN(n14904) );
  AOI21_X1 U16589 ( .B1(n14920), .B2(n14904), .A(n15010), .ZN(n14912) );
  AOI21_X1 U16590 ( .B1(n11037), .B2(n14906), .A(n14905), .ZN(n14910) );
  XNOR2_X1 U16591 ( .A(n14907), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n14909) );
  OAI22_X1 U16592 ( .A1(n15036), .A2(n14910), .B1(n14909), .B2(n14908), .ZN(
        n14911) );
  AOI211_X1 U16593 ( .C1(n15021), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        n14915) );
  NAND2_X1 U16594 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n14914) );
  OAI211_X1 U16595 ( .C1(n14916), .C2(n15041), .A(n14915), .B(n14914), .ZN(
        P3_U3185) );
  INV_X1 U16596 ( .A(n14917), .ZN(n14918) );
  NAND3_X1 U16597 ( .A1(n14920), .A2(n14919), .A3(n14918), .ZN(n14921) );
  AOI21_X1 U16598 ( .B1(n14940), .B2(n14921), .A(n15010), .ZN(n14932) );
  AOI21_X1 U16599 ( .B1(n14924), .B2(n14923), .A(n14922), .ZN(n14930) );
  OAI21_X1 U16600 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14928) );
  NAND2_X1 U16601 ( .A1(n15023), .A2(n14928), .ZN(n14929) );
  OAI21_X1 U16602 ( .B1(n15036), .B2(n14930), .A(n14929), .ZN(n14931) );
  AOI211_X1 U16603 ( .C1(n15021), .C2(n14933), .A(n14932), .B(n14931), .ZN(
        n14935) );
  NAND2_X1 U16604 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n14934) );
  OAI211_X1 U16605 ( .C1(n14936), .C2(n15041), .A(n14935), .B(n14934), .ZN(
        P3_U3186) );
  INV_X1 U16606 ( .A(n14937), .ZN(n14938) );
  NAND3_X1 U16607 ( .A1(n14940), .A2(n14939), .A3(n14938), .ZN(n14941) );
  AOI21_X1 U16608 ( .B1(n14968), .B2(n14941), .A(n15010), .ZN(n14950) );
  AOI21_X1 U16609 ( .B1(n14943), .B2(n11051), .A(n14942), .ZN(n14948) );
  OAI21_X1 U16610 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14945), .A(n14944), .ZN(
        n14946) );
  NAND2_X1 U16611 ( .A1(n15023), .A2(n14946), .ZN(n14947) );
  OAI21_X1 U16612 ( .B1(n15036), .B2(n14948), .A(n14947), .ZN(n14949) );
  AOI211_X1 U16613 ( .C1(n15021), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14953) );
  NAND2_X1 U16614 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n14952) );
  OAI211_X1 U16615 ( .C1(n14954), .C2(n15041), .A(n14953), .B(n14952), .ZN(
        P3_U3187) );
  INV_X1 U16616 ( .A(n14955), .ZN(n14956) );
  AOI21_X1 U16617 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(n14964) );
  OAI21_X1 U16618 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14962) );
  NAND2_X1 U16619 ( .A1(n15023), .A2(n14962), .ZN(n14963) );
  OAI21_X1 U16620 ( .B1(n15036), .B2(n14964), .A(n14963), .ZN(n14971) );
  INV_X1 U16621 ( .A(n14965), .ZN(n14966) );
  NAND3_X1 U16622 ( .A1(n14968), .A2(n14967), .A3(n14966), .ZN(n14969) );
  AOI21_X1 U16623 ( .B1(n14983), .B2(n14969), .A(n15010), .ZN(n14970) );
  AOI211_X1 U16624 ( .C1(n15021), .C2(n14972), .A(n14971), .B(n14970), .ZN(
        n14974) );
  NAND2_X1 U16625 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14973) );
  OAI211_X1 U16626 ( .C1(n14975), .C2(n15041), .A(n14974), .B(n14973), .ZN(
        P3_U3188) );
  AOI21_X1 U16627 ( .B1(n11117), .B2(n14977), .A(n14976), .ZN(n14996) );
  NOR2_X1 U16628 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14978), .ZN(n14989) );
  INV_X1 U16629 ( .A(n14979), .ZN(n14980) );
  NOR2_X1 U16630 ( .A1(n14981), .A2(n14980), .ZN(n14984) );
  INV_X1 U16631 ( .A(n15009), .ZN(n14982) );
  AOI21_X1 U16632 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n14987) );
  OAI22_X1 U16633 ( .A1(n14987), .A2(n15010), .B1(n14986), .B2(n14985), .ZN(
        n14988) );
  AOI211_X1 U16634 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14990), .A(n14989), .B(
        n14988), .ZN(n14995) );
  OAI21_X1 U16635 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14992), .A(n14991), .ZN(
        n14993) );
  NAND2_X1 U16636 ( .A1(n14993), .A2(n15023), .ZN(n14994) );
  OAI211_X1 U16637 ( .C1(n14996), .C2(n15036), .A(n14995), .B(n14994), .ZN(
        P3_U3189) );
  AOI21_X1 U16638 ( .B1(n14998), .B2(n14997), .A(n6615), .ZN(n15005) );
  OAI21_X1 U16639 ( .B1(n15001), .B2(n15000), .A(n14999), .ZN(n15003) );
  AOI22_X1 U16640 ( .A1(n15003), .A2(n15023), .B1(n15021), .B2(n15002), .ZN(
        n15004) );
  OAI21_X1 U16641 ( .B1(n15005), .B2(n15036), .A(n15004), .ZN(n15013) );
  INV_X1 U16642 ( .A(n15006), .ZN(n15007) );
  NAND3_X1 U16643 ( .A1(n15009), .A2(n15008), .A3(n15007), .ZN(n15011) );
  AOI21_X1 U16644 ( .B1(n15025), .B2(n15011), .A(n15010), .ZN(n15012) );
  NOR2_X1 U16645 ( .A1(n15013), .A2(n15012), .ZN(n15015) );
  NAND2_X1 U16646 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15014) );
  OAI211_X1 U16647 ( .C1(n15016), .C2(n15041), .A(n15015), .B(n15014), .ZN(
        P3_U3190) );
  AOI21_X1 U16648 ( .B1(n15018), .B2(n11077), .A(n15017), .ZN(n15037) );
  OAI21_X1 U16649 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15020), .A(n15019), .ZN(
        n15024) );
  AOI22_X1 U16650 ( .A1(n15024), .A2(n15023), .B1(n15022), .B2(n15021), .ZN(
        n15035) );
  INV_X1 U16651 ( .A(n15025), .ZN(n15029) );
  INV_X1 U16652 ( .A(n15026), .ZN(n15028) );
  NOR3_X1 U16653 ( .A1(n15029), .A2(n15028), .A3(n15027), .ZN(n15033) );
  INV_X1 U16654 ( .A(n15030), .ZN(n15032) );
  OAI21_X1 U16655 ( .B1(n15033), .B2(n15032), .A(n15031), .ZN(n15034) );
  OAI211_X1 U16656 ( .C1(n15037), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15038) );
  INV_X1 U16657 ( .A(n15038), .ZN(n15040) );
  NAND2_X1 U16658 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15039) );
  OAI211_X1 U16659 ( .C1(n15234), .C2(n15041), .A(n15040), .B(n15039), .ZN(
        P3_U3191) );
  XNOR2_X1 U16660 ( .A(n15047), .B(n15042), .ZN(n15055) );
  INV_X1 U16661 ( .A(n15055), .ZN(n15086) );
  NOR2_X1 U16662 ( .A1(n15043), .A2(n15124), .ZN(n15085) );
  INV_X1 U16663 ( .A(n15085), .ZN(n15044) );
  OAI22_X1 U16664 ( .A1(n15072), .A2(n15046), .B1(n15045), .B2(n15044), .ZN(
        n15056) );
  XNOR2_X1 U16665 ( .A(n15048), .B(n15047), .ZN(n15053) );
  OAI22_X1 U16666 ( .A1(n15051), .A2(n15050), .B1(n7838), .B2(n15049), .ZN(
        n15052) );
  AOI21_X1 U16667 ( .B1(n15053), .B2(n15067), .A(n15052), .ZN(n15054) );
  OAI21_X1 U16668 ( .B1(n15108), .B2(n15055), .A(n15054), .ZN(n15084) );
  AOI211_X1 U16669 ( .C1(n15057), .C2(n15086), .A(n15056), .B(n15084), .ZN(
        n15058) );
  AOI22_X1 U16670 ( .A1(n15079), .A2(n10669), .B1(n15058), .B2(n15077), .ZN(
        P3_U3231) );
  NOR2_X1 U16671 ( .A1(n15059), .A2(n15124), .ZN(n15082) );
  XNOR2_X1 U16672 ( .A(n15060), .B(n15066), .ZN(n15080) );
  AOI22_X1 U16673 ( .A1(n15064), .A2(n15063), .B1(n15062), .B2(n15061), .ZN(
        n15070) );
  XNOR2_X1 U16674 ( .A(n15066), .B(n15065), .ZN(n15068) );
  NAND2_X1 U16675 ( .A1(n15068), .A2(n15067), .ZN(n15069) );
  OAI211_X1 U16676 ( .C1(n15080), .C2(n15108), .A(n15070), .B(n15069), .ZN(
        n15081) );
  AOI21_X1 U16677 ( .B1(n15082), .B2(n15071), .A(n15081), .ZN(n15078) );
  OAI22_X1 U16678 ( .A1(n15074), .A2(n15080), .B1(n15073), .B2(n15072), .ZN(
        n15075) );
  INV_X1 U16679 ( .A(n15075), .ZN(n15076) );
  OAI221_X1 U16680 ( .B1(n15079), .B2(n15078), .C1(n15077), .C2(n10544), .A(
        n15076), .ZN(P3_U3232) );
  INV_X1 U16681 ( .A(n15080), .ZN(n15083) );
  AOI211_X1 U16682 ( .C1(n15129), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15131) );
  AOI22_X1 U16683 ( .A1(n15130), .A2(n15131), .B1(n7825), .B2(n8319), .ZN(
        P3_U3393) );
  AOI211_X1 U16684 ( .C1(n15086), .C2(n15129), .A(n15085), .B(n15084), .ZN(
        n15132) );
  AOI22_X1 U16685 ( .A1(n15130), .A2(n15132), .B1(n7843), .B2(n8319), .ZN(
        P3_U3396) );
  NAND2_X1 U16686 ( .A1(n15091), .A2(n15129), .ZN(n15087) );
  OAI211_X1 U16687 ( .C1(n15089), .C2(n15124), .A(n15088), .B(n15087), .ZN(
        n15090) );
  AOI21_X1 U16688 ( .B1(n15091), .B2(n15118), .A(n15090), .ZN(n15133) );
  AOI22_X1 U16689 ( .A1(n15130), .A2(n15133), .B1(n7855), .B2(n8319), .ZN(
        P3_U3399) );
  INV_X1 U16690 ( .A(n15129), .ZN(n15114) );
  AOI21_X1 U16691 ( .B1(n15108), .B2(n15114), .A(n15092), .ZN(n15095) );
  INV_X1 U16692 ( .A(n15093), .ZN(n15094) );
  AOI211_X1 U16693 ( .C1(n15105), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        n15134) );
  AOI22_X1 U16694 ( .A1(n15130), .A2(n15134), .B1(n7870), .B2(n8319), .ZN(
        P3_U3402) );
  NOR2_X1 U16695 ( .A1(n15097), .A2(n15124), .ZN(n15099) );
  AOI211_X1 U16696 ( .C1(n15100), .C2(n15129), .A(n15099), .B(n15098), .ZN(
        n15135) );
  AOI22_X1 U16697 ( .A1(n15130), .A2(n15135), .B1(n7888), .B2(n8319), .ZN(
        P3_U3405) );
  AOI21_X1 U16698 ( .B1(n15108), .B2(n15114), .A(n15101), .ZN(n15103) );
  AOI211_X1 U16699 ( .C1(n15105), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n15136) );
  AOI22_X1 U16700 ( .A1(n15130), .A2(n15136), .B1(n7906), .B2(n8319), .ZN(
        P3_U3408) );
  OAI22_X1 U16701 ( .A1(n15109), .A2(n15114), .B1(n15124), .B2(n15106), .ZN(
        n15107) );
  INV_X1 U16702 ( .A(n15107), .ZN(n15111) );
  OR2_X1 U16703 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  AOI22_X1 U16704 ( .A1(n15130), .A2(n15137), .B1(n7920), .B2(n8319), .ZN(
        P3_U3411) );
  INV_X1 U16705 ( .A(n15115), .ZN(n15119) );
  OAI22_X1 U16706 ( .A1(n15115), .A2(n15114), .B1(n15113), .B2(n15124), .ZN(
        n15117) );
  AOI211_X1 U16707 ( .C1(n15119), .C2(n15118), .A(n15117), .B(n15116), .ZN(
        n15139) );
  AOI22_X1 U16708 ( .A1(n15130), .A2(n15139), .B1(n7936), .B2(n8319), .ZN(
        P3_U3414) );
  NOR2_X1 U16709 ( .A1(n15120), .A2(n15124), .ZN(n15122) );
  AOI211_X1 U16710 ( .C1(n15123), .C2(n15129), .A(n15122), .B(n15121), .ZN(
        n15140) );
  AOI22_X1 U16711 ( .A1(n15130), .A2(n15140), .B1(n7950), .B2(n8319), .ZN(
        P3_U3417) );
  NOR2_X1 U16712 ( .A1(n15125), .A2(n15124), .ZN(n15127) );
  AOI211_X1 U16713 ( .C1(n15129), .C2(n15128), .A(n15127), .B(n15126), .ZN(
        n15143) );
  AOI22_X1 U16714 ( .A1(n15130), .A2(n15143), .B1(n7965), .B2(n8319), .ZN(
        P3_U3420) );
  AOI22_X1 U16715 ( .A1(n15144), .A2(n15131), .B1(n10543), .B2(n15141), .ZN(
        P3_U3460) );
  AOI22_X1 U16716 ( .A1(n15144), .A2(n15132), .B1(n10668), .B2(n15141), .ZN(
        P3_U3461) );
  AOI22_X1 U16717 ( .A1(n15144), .A2(n15133), .B1(n11036), .B2(n15141), .ZN(
        P3_U3462) );
  AOI22_X1 U16718 ( .A1(n15144), .A2(n15134), .B1(n11043), .B2(n15141), .ZN(
        P3_U3463) );
  AOI22_X1 U16719 ( .A1(n15144), .A2(n15135), .B1(n11050), .B2(n15141), .ZN(
        P3_U3464) );
  AOI22_X1 U16720 ( .A1(n15144), .A2(n15136), .B1(n11057), .B2(n15141), .ZN(
        P3_U3465) );
  AOI22_X1 U16721 ( .A1(n15144), .A2(n15137), .B1(n11064), .B2(n15141), .ZN(
        P3_U3466) );
  AOI22_X1 U16722 ( .A1(n15144), .A2(n15139), .B1(n15138), .B2(n15141), .ZN(
        P3_U3467) );
  AOI22_X1 U16723 ( .A1(n15144), .A2(n15140), .B1(n11076), .B2(n15141), .ZN(
        P3_U3468) );
  AOI22_X1 U16724 ( .A1(n15144), .A2(n15143), .B1(n15142), .B2(n15141), .ZN(
        P3_U3469) );
  NAND2_X1 U16725 ( .A1(keyinput31), .A2(keyinput39), .ZN(n15145) );
  NOR3_X1 U16726 ( .A1(keyinput57), .A2(keyinput4), .A3(n15145), .ZN(n15146)
         );
  NAND3_X1 U16727 ( .A1(keyinput121), .A2(keyinput66), .A3(n15146), .ZN(n15159) );
  NAND2_X1 U16728 ( .A1(keyinput10), .A2(keyinput126), .ZN(n15147) );
  NOR3_X1 U16729 ( .A1(keyinput0), .A2(keyinput23), .A3(n15147), .ZN(n15157)
         );
  NOR4_X1 U16730 ( .A1(keyinput46), .A2(keyinput8), .A3(keyinput108), .A4(
        keyinput98), .ZN(n15156) );
  NOR2_X1 U16731 ( .A1(keyinput28), .A2(keyinput109), .ZN(n15148) );
  NAND3_X1 U16732 ( .A1(keyinput20), .A2(keyinput63), .A3(n15148), .ZN(n15154)
         );
  NOR2_X1 U16733 ( .A1(keyinput16), .A2(keyinput97), .ZN(n15149) );
  NAND3_X1 U16734 ( .A1(keyinput52), .A2(keyinput17), .A3(n15149), .ZN(n15153)
         );
  NOR2_X1 U16735 ( .A1(keyinput49), .A2(keyinput45), .ZN(n15150) );
  NAND3_X1 U16736 ( .A1(keyinput5), .A2(keyinput48), .A3(n15150), .ZN(n15152)
         );
  NAND4_X1 U16737 ( .A1(keyinput18), .A2(keyinput115), .A3(keyinput106), .A4(
        keyinput83), .ZN(n15151) );
  NOR4_X1 U16738 ( .A1(n15154), .A2(n15153), .A3(n15152), .A4(n15151), .ZN(
        n15155) );
  NAND3_X1 U16739 ( .A1(n15157), .A2(n15156), .A3(n15155), .ZN(n15158) );
  NOR4_X1 U16740 ( .A1(keyinput14), .A2(keyinput111), .A3(n15159), .A4(n15158), 
        .ZN(n15208) );
  INV_X1 U16741 ( .A(keyinput87), .ZN(n15162) );
  INV_X1 U16742 ( .A(keyinput71), .ZN(n15160) );
  NAND4_X1 U16743 ( .A1(keyinput100), .A2(keyinput55), .A3(keyinput35), .A4(
        n15160), .ZN(n15161) );
  NOR4_X1 U16744 ( .A1(keyinput34), .A2(keyinput102), .A3(n15162), .A4(n15161), 
        .ZN(n15174) );
  NOR4_X1 U16745 ( .A1(keyinput101), .A2(keyinput90), .A3(keyinput47), .A4(
        keyinput36), .ZN(n15173) );
  NAND3_X1 U16746 ( .A1(keyinput15), .A2(keyinput62), .A3(keyinput93), .ZN(
        n15163) );
  NOR2_X1 U16747 ( .A1(keyinput94), .A2(n15163), .ZN(n15172) );
  NAND4_X1 U16748 ( .A1(keyinput77), .A2(keyinput68), .A3(keyinput103), .A4(
        keyinput107), .ZN(n15170) );
  NOR2_X1 U16749 ( .A1(keyinput38), .A2(keyinput105), .ZN(n15164) );
  NAND3_X1 U16750 ( .A1(keyinput82), .A2(keyinput41), .A3(n15164), .ZN(n15169)
         );
  INV_X1 U16751 ( .A(keyinput67), .ZN(n15165) );
  NAND4_X1 U16752 ( .A1(keyinput79), .A2(keyinput19), .A3(keyinput104), .A4(
        n15165), .ZN(n15168) );
  NOR3_X1 U16753 ( .A1(keyinput56), .A2(keyinput6), .A3(keyinput78), .ZN(
        n15166) );
  NAND2_X1 U16754 ( .A1(keyinput26), .A2(n15166), .ZN(n15167) );
  NOR4_X1 U16755 ( .A1(n15170), .A2(n15169), .A3(n15168), .A4(n15167), .ZN(
        n15171) );
  NAND4_X1 U16756 ( .A1(n15174), .A2(n15173), .A3(n15172), .A4(n15171), .ZN(
        n15206) );
  NOR4_X1 U16757 ( .A1(keyinput3), .A2(keyinput58), .A3(keyinput70), .A4(
        keyinput54), .ZN(n15180) );
  NAND2_X1 U16758 ( .A1(keyinput37), .A2(keyinput88), .ZN(n15175) );
  NOR3_X1 U16759 ( .A1(keyinput81), .A2(keyinput9), .A3(n15175), .ZN(n15179)
         );
  AND4_X1 U16760 ( .A1(keyinput13), .A2(keyinput91), .A3(keyinput86), .A4(
        keyinput24), .ZN(n15178) );
  INV_X1 U16761 ( .A(keyinput11), .ZN(n15176) );
  NOR4_X1 U16762 ( .A1(keyinput75), .A2(keyinput120), .A3(keyinput72), .A4(
        n15176), .ZN(n15177) );
  NAND4_X1 U16763 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        n15205) );
  AND4_X1 U16764 ( .A1(keyinput112), .A2(keyinput42), .A3(keyinput25), .A4(
        keyinput117), .ZN(n15185) );
  INV_X1 U16765 ( .A(keyinput123), .ZN(n15181) );
  NOR4_X1 U16766 ( .A1(keyinput74), .A2(keyinput85), .A3(keyinput44), .A4(
        n15181), .ZN(n15184) );
  AND4_X1 U16767 ( .A1(keyinput89), .A2(keyinput114), .A3(keyinput116), .A4(
        keyinput92), .ZN(n15183) );
  NOR4_X1 U16768 ( .A1(keyinput80), .A2(keyinput124), .A3(keyinput60), .A4(
        keyinput125), .ZN(n15182) );
  NAND4_X1 U16769 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15204) );
  NAND2_X1 U16770 ( .A1(keyinput40), .A2(keyinput118), .ZN(n15186) );
  NOR3_X1 U16771 ( .A1(keyinput33), .A2(keyinput2), .A3(n15186), .ZN(n15202)
         );
  INV_X1 U16772 ( .A(keyinput53), .ZN(n15187) );
  NOR4_X1 U16773 ( .A1(keyinput119), .A2(keyinput122), .A3(keyinput61), .A4(
        n15187), .ZN(n15201) );
  INV_X1 U16774 ( .A(keyinput99), .ZN(n15188) );
  NAND2_X1 U16775 ( .A1(keyinput51), .A2(n15188), .ZN(n15190) );
  NAND4_X1 U16776 ( .A1(keyinput84), .A2(keyinput64), .A3(keyinput1), .A4(
        keyinput30), .ZN(n15189) );
  NOR4_X1 U16777 ( .A1(keyinput12), .A2(keyinput96), .A3(n15190), .A4(n15189), 
        .ZN(n15200) );
  INV_X1 U16778 ( .A(keyinput95), .ZN(n15191) );
  NAND4_X1 U16779 ( .A1(keyinput76), .A2(keyinput113), .A3(keyinput65), .A4(
        n15191), .ZN(n15198) );
  NOR2_X1 U16780 ( .A1(keyinput21), .A2(keyinput69), .ZN(n15192) );
  NAND3_X1 U16781 ( .A1(keyinput29), .A2(keyinput27), .A3(n15192), .ZN(n15197)
         );
  INV_X1 U16782 ( .A(keyinput73), .ZN(n15193) );
  NAND4_X1 U16783 ( .A1(keyinput7), .A2(keyinput50), .A3(keyinput43), .A4(
        n15193), .ZN(n15196) );
  NOR2_X1 U16784 ( .A1(keyinput32), .A2(keyinput22), .ZN(n15194) );
  NAND3_X1 U16785 ( .A1(keyinput59), .A2(keyinput110), .A3(n15194), .ZN(n15195) );
  NOR4_X1 U16786 ( .A1(n15198), .A2(n15197), .A3(n15196), .A4(n15195), .ZN(
        n15199) );
  NAND4_X1 U16787 ( .A1(n15202), .A2(n15201), .A3(n15200), .A4(n15199), .ZN(
        n15203) );
  NOR4_X1 U16788 ( .A1(n15206), .A2(n15205), .A3(n15204), .A4(n15203), .ZN(
        n15207) );
  AOI21_X1 U16789 ( .B1(n15208), .B2(n15207), .A(keyinput127), .ZN(n15452) );
  AOI22_X1 U16790 ( .A1(n15211), .A2(keyinput111), .B1(keyinput46), .B2(n15210), .ZN(n15209) );
  OAI221_X1 U16791 ( .B1(n15211), .B2(keyinput111), .C1(n15210), .C2(
        keyinput46), .A(n15209), .ZN(n15219) );
  AOI22_X1 U16792 ( .A1(n10552), .A2(keyinput66), .B1(n7982), .B2(keyinput31), 
        .ZN(n15212) );
  OAI221_X1 U16793 ( .B1(n10552), .B2(keyinput66), .C1(n7982), .C2(keyinput31), 
        .A(n15212), .ZN(n15218) );
  XOR2_X1 U16794 ( .A(n8485), .B(keyinput121), .Z(n15216) );
  XNOR2_X1 U16795 ( .A(SI_2_), .B(keyinput57), .ZN(n15215) );
  XNOR2_X1 U16796 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput4), .ZN(n15214) );
  XNOR2_X1 U16797 ( .A(P3_REG0_REG_16__SCAN_IN), .B(keyinput14), .ZN(n15213)
         );
  NAND4_X1 U16798 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15217) );
  NOR3_X1 U16799 ( .A1(n15219), .A2(n15218), .A3(n15217), .ZN(n15264) );
  XOR2_X1 U16800 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput0), .Z(n15223) );
  XOR2_X1 U16801 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput8), .Z(n15222) );
  XNOR2_X1 U16802 ( .A(n15220), .B(keyinput52), .ZN(n15221) );
  NOR3_X1 U16803 ( .A1(n15223), .A2(n15222), .A3(n15221), .ZN(n15226) );
  XNOR2_X1 U16804 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput126), .ZN(n15225)
         );
  XNOR2_X1 U16805 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput10), .ZN(n15224) );
  NAND3_X1 U16806 ( .A1(n15226), .A2(n15225), .A3(n15224), .ZN(n15232) );
  AOI22_X1 U16807 ( .A1(n15228), .A2(keyinput23), .B1(n8027), .B2(keyinput108), 
        .ZN(n15227) );
  OAI221_X1 U16808 ( .B1(n15228), .B2(keyinput23), .C1(n8027), .C2(keyinput108), .A(n15227), .ZN(n15231) );
  XNOR2_X1 U16809 ( .A(n15229), .B(keyinput98), .ZN(n15230) );
  NOR3_X1 U16810 ( .A1(n15232), .A2(n15231), .A3(n15230), .ZN(n15263) );
  AOI22_X1 U16811 ( .A1(n15235), .A2(keyinput97), .B1(keyinput16), .B2(n15234), 
        .ZN(n15233) );
  OAI221_X1 U16812 ( .B1(n15235), .B2(keyinput97), .C1(n15234), .C2(keyinput16), .A(n15233), .ZN(n15245) );
  INV_X1 U16813 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n15237) );
  AOI22_X1 U16814 ( .A1(n15238), .A2(keyinput28), .B1(keyinput63), .B2(n15237), 
        .ZN(n15236) );
  OAI221_X1 U16815 ( .B1(n15238), .B2(keyinput28), .C1(n15237), .C2(keyinput63), .A(n15236), .ZN(n15244) );
  XNOR2_X1 U16816 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput20), .ZN(n15242) );
  XNOR2_X1 U16817 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput18), .ZN(n15241)
         );
  XNOR2_X1 U16818 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput109), .ZN(n15240) );
  XNOR2_X1 U16819 ( .A(keyinput17), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n15239)
         );
  NAND4_X1 U16820 ( .A1(n15242), .A2(n15241), .A3(n15240), .A4(n15239), .ZN(
        n15243) );
  NOR3_X1 U16821 ( .A1(n15245), .A2(n15244), .A3(n15243), .ZN(n15262) );
  AOI22_X1 U16822 ( .A1(n15248), .A2(keyinput115), .B1(n15247), .B2(keyinput5), 
        .ZN(n15246) );
  OAI221_X1 U16823 ( .B1(n15248), .B2(keyinput115), .C1(n15247), .C2(keyinput5), .A(n15246), .ZN(n15260) );
  INV_X1 U16824 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n15251) );
  AOI22_X1 U16825 ( .A1(n15251), .A2(keyinput49), .B1(n15250), .B2(keyinput48), 
        .ZN(n15249) );
  OAI221_X1 U16826 ( .B1(n15251), .B2(keyinput49), .C1(n15250), .C2(keyinput48), .A(n15249), .ZN(n15259) );
  INV_X1 U16827 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15253) );
  AOI22_X1 U16828 ( .A1(n15254), .A2(keyinput45), .B1(keyinput106), .B2(n15253), .ZN(n15252) );
  OAI221_X1 U16829 ( .B1(n15254), .B2(keyinput45), .C1(n15253), .C2(
        keyinput106), .A(n15252), .ZN(n15258) );
  AOI22_X1 U16830 ( .A1(n11076), .A2(keyinput83), .B1(keyinput29), .B2(n15256), 
        .ZN(n15255) );
  OAI221_X1 U16831 ( .B1(n11076), .B2(keyinput83), .C1(n15256), .C2(keyinput29), .A(n15255), .ZN(n15257) );
  NOR4_X1 U16832 ( .A1(n15260), .A2(n15259), .A3(n15258), .A4(n15257), .ZN(
        n15261) );
  NAND4_X1 U16833 ( .A1(n15264), .A2(n15263), .A3(n15262), .A4(n15261), .ZN(
        n15450) );
  AOI22_X1 U16834 ( .A1(n15266), .A2(keyinput65), .B1(n10304), .B2(keyinput59), 
        .ZN(n15265) );
  OAI221_X1 U16835 ( .B1(n15266), .B2(keyinput65), .C1(n10304), .C2(keyinput59), .A(n15265), .ZN(n15277) );
  AOI22_X1 U16836 ( .A1(n11117), .A2(keyinput69), .B1(keyinput95), .B2(n15268), 
        .ZN(n15267) );
  OAI221_X1 U16837 ( .B1(n11117), .B2(keyinput69), .C1(n15268), .C2(keyinput95), .A(n15267), .ZN(n15276) );
  AOI22_X1 U16838 ( .A1(n15271), .A2(keyinput76), .B1(keyinput113), .B2(n15270), .ZN(n15269) );
  OAI221_X1 U16839 ( .B1(n15271), .B2(keyinput76), .C1(n15270), .C2(
        keyinput113), .A(n15269), .ZN(n15275) );
  XNOR2_X1 U16840 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput27), .ZN(n15273)
         );
  XNOR2_X1 U16841 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput21), .ZN(n15272) );
  NAND2_X1 U16842 ( .A1(n15273), .A2(n15272), .ZN(n15274) );
  NOR4_X1 U16843 ( .A1(n15277), .A2(n15276), .A3(n15275), .A4(n15274), .ZN(
        n15318) );
  AOI22_X1 U16844 ( .A1(n15279), .A2(keyinput22), .B1(keyinput50), .B2(n7981), 
        .ZN(n15278) );
  OAI221_X1 U16845 ( .B1(n15279), .B2(keyinput22), .C1(n7981), .C2(keyinput50), 
        .A(n15278), .ZN(n15289) );
  AOI22_X1 U16846 ( .A1(n15281), .A2(keyinput7), .B1(n7906), .B2(keyinput73), 
        .ZN(n15280) );
  OAI221_X1 U16847 ( .B1(n15281), .B2(keyinput7), .C1(n7906), .C2(keyinput73), 
        .A(n15280), .ZN(n15288) );
  XNOR2_X1 U16848 ( .A(SI_5_), .B(keyinput119), .ZN(n15284) );
  XNOR2_X1 U16849 ( .A(P1_REG1_REG_23__SCAN_IN), .B(keyinput110), .ZN(n15283)
         );
  XNOR2_X1 U16850 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput32), .ZN(n15282)
         );
  NAND3_X1 U16851 ( .A1(n15284), .A2(n15283), .A3(n15282), .ZN(n15287) );
  XNOR2_X1 U16852 ( .A(n15285), .B(keyinput43), .ZN(n15286) );
  NOR4_X1 U16853 ( .A1(n15289), .A2(n15288), .A3(n15287), .A4(n15286), .ZN(
        n15317) );
  AOI22_X1 U16854 ( .A1(n15291), .A2(keyinput40), .B1(keyinput99), .B2(n10163), 
        .ZN(n15290) );
  OAI221_X1 U16855 ( .B1(n15291), .B2(keyinput40), .C1(n10163), .C2(keyinput99), .A(n15290), .ZN(n15301) );
  AOI22_X1 U16856 ( .A1(n15294), .A2(keyinput61), .B1(n15293), .B2(keyinput118), .ZN(n15292) );
  OAI221_X1 U16857 ( .B1(n15294), .B2(keyinput61), .C1(n15293), .C2(
        keyinput118), .A(n15292), .ZN(n15300) );
  XNOR2_X1 U16858 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput122), .ZN(n15298)
         );
  XNOR2_X1 U16859 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput53), .ZN(n15297) );
  XNOR2_X1 U16860 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput2), .ZN(n15296) );
  XNOR2_X1 U16861 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput33), .ZN(n15295) );
  NAND4_X1 U16862 ( .A1(n15298), .A2(n15297), .A3(n15296), .A4(n15295), .ZN(
        n15299) );
  NOR3_X1 U16863 ( .A1(n15301), .A2(n15300), .A3(n15299), .ZN(n15316) );
  AOI22_X1 U16864 ( .A1(n15304), .A2(keyinput51), .B1(keyinput84), .B2(n15303), 
        .ZN(n15302) );
  OAI221_X1 U16865 ( .B1(n15304), .B2(keyinput51), .C1(n15303), .C2(keyinput84), .A(n15302), .ZN(n15314) );
  AOI22_X1 U16866 ( .A1(n9263), .A2(keyinput64), .B1(n10150), .B2(keyinput96), 
        .ZN(n15305) );
  OAI221_X1 U16867 ( .B1(n9263), .B2(keyinput64), .C1(n10150), .C2(keyinput96), 
        .A(n15305), .ZN(n15313) );
  AOI22_X1 U16868 ( .A1(n6810), .A2(keyinput12), .B1(n15307), .B2(keyinput1), 
        .ZN(n15306) );
  OAI221_X1 U16869 ( .B1(n6810), .B2(keyinput12), .C1(n15307), .C2(keyinput1), 
        .A(n15306), .ZN(n15312) );
  AOI22_X1 U16870 ( .A1(n15310), .A2(keyinput34), .B1(keyinput30), .B2(n15309), 
        .ZN(n15308) );
  OAI221_X1 U16871 ( .B1(n15310), .B2(keyinput34), .C1(n15309), .C2(keyinput30), .A(n15308), .ZN(n15311) );
  NOR4_X1 U16872 ( .A1(n15314), .A2(n15313), .A3(n15312), .A4(n15311), .ZN(
        n15315) );
  NAND4_X1 U16873 ( .A1(n15318), .A2(n15317), .A3(n15316), .A4(n15315), .ZN(
        n15449) );
  INV_X1 U16874 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15320) );
  AOI22_X1 U16875 ( .A1(n15321), .A2(keyinput114), .B1(n15320), .B2(
        keyinput116), .ZN(n15319) );
  OAI221_X1 U16876 ( .B1(n15321), .B2(keyinput114), .C1(n15320), .C2(
        keyinput116), .A(n15319), .ZN(n15332) );
  AOI22_X1 U16877 ( .A1(n15324), .A2(keyinput92), .B1(n15323), .B2(keyinput81), 
        .ZN(n15322) );
  OAI221_X1 U16878 ( .B1(n15324), .B2(keyinput92), .C1(n15323), .C2(keyinput81), .A(n15322), .ZN(n15331) );
  INV_X1 U16879 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15326) );
  AOI22_X1 U16880 ( .A1(n7720), .A2(keyinput124), .B1(keyinput60), .B2(n15326), 
        .ZN(n15325) );
  OAI221_X1 U16881 ( .B1(n7720), .B2(keyinput124), .C1(n15326), .C2(keyinput60), .A(n15325), .ZN(n15330) );
  XOR2_X1 U16882 ( .A(n9267), .B(keyinput89), .Z(n15328) );
  XNOR2_X1 U16883 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput125), .ZN(n15327) );
  NAND2_X1 U16884 ( .A1(n15328), .A2(n15327), .ZN(n15329) );
  NOR4_X1 U16885 ( .A1(n15332), .A2(n15331), .A3(n15330), .A4(n15329), .ZN(
        n15380) );
  INV_X1 U16886 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15335) );
  INV_X1 U16887 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n15334) );
  AOI22_X1 U16888 ( .A1(n15335), .A2(keyinput42), .B1(keyinput25), .B2(n15334), 
        .ZN(n15333) );
  OAI221_X1 U16889 ( .B1(n15335), .B2(keyinput42), .C1(n15334), .C2(keyinput25), .A(n15333), .ZN(n15346) );
  AOI22_X1 U16890 ( .A1(n15337), .A2(keyinput123), .B1(n8807), .B2(keyinput112), .ZN(n15336) );
  OAI221_X1 U16891 ( .B1(n15337), .B2(keyinput123), .C1(n8807), .C2(
        keyinput112), .A(n15336), .ZN(n15345) );
  INV_X1 U16892 ( .A(keyinput80), .ZN(n15339) );
  AOI22_X1 U16893 ( .A1(n7825), .A2(keyinput44), .B1(P1_WR_REG_SCAN_IN), .B2(
        n15339), .ZN(n15338) );
  OAI221_X1 U16894 ( .B1(n7825), .B2(keyinput44), .C1(n15339), .C2(
        P1_WR_REG_SCAN_IN), .A(n15338), .ZN(n15344) );
  INV_X1 U16895 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U16896 ( .A1(n15342), .A2(keyinput117), .B1(n15341), .B2(keyinput85), .ZN(n15340) );
  OAI221_X1 U16897 ( .B1(n15342), .B2(keyinput117), .C1(n15341), .C2(
        keyinput85), .A(n15340), .ZN(n15343) );
  NOR4_X1 U16898 ( .A1(n15346), .A2(n15345), .A3(n15344), .A4(n15343), .ZN(
        n15379) );
  AOI22_X1 U16899 ( .A1(n15349), .A2(keyinput91), .B1(n15348), .B2(keyinput75), 
        .ZN(n15347) );
  OAI221_X1 U16900 ( .B1(n15349), .B2(keyinput91), .C1(n15348), .C2(keyinput75), .A(n15347), .ZN(n15361) );
  AOI22_X1 U16901 ( .A1(n15351), .A2(keyinput120), .B1(n8740), .B2(keyinput13), 
        .ZN(n15350) );
  OAI221_X1 U16902 ( .B1(n15351), .B2(keyinput120), .C1(n8740), .C2(keyinput13), .A(n15350), .ZN(n15360) );
  AOI22_X1 U16903 ( .A1(n15354), .A2(keyinput24), .B1(keyinput39), .B2(n15353), 
        .ZN(n15352) );
  OAI221_X1 U16904 ( .B1(n15354), .B2(keyinput24), .C1(n15353), .C2(keyinput39), .A(n15352), .ZN(n15359) );
  AOI22_X1 U16905 ( .A1(n15357), .A2(keyinput72), .B1(keyinput86), .B2(n15356), 
        .ZN(n15355) );
  OAI221_X1 U16906 ( .B1(n15357), .B2(keyinput72), .C1(n15356), .C2(keyinput86), .A(n15355), .ZN(n15358) );
  NOR4_X1 U16907 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        n15378) );
  AOI22_X1 U16908 ( .A1(n15364), .A2(keyinput58), .B1(keyinput70), .B2(n15363), 
        .ZN(n15362) );
  OAI221_X1 U16909 ( .B1(n15364), .B2(keyinput58), .C1(n15363), .C2(keyinput70), .A(n15362), .ZN(n15376) );
  INV_X1 U16910 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U16911 ( .A1(n15367), .A2(keyinput88), .B1(keyinput3), .B2(n15366), 
        .ZN(n15365) );
  OAI221_X1 U16912 ( .B1(n15367), .B2(keyinput88), .C1(n15366), .C2(keyinput3), 
        .A(n15365), .ZN(n15375) );
  AOI22_X1 U16913 ( .A1(n15369), .A2(keyinput37), .B1(keyinput11), .B2(n9297), 
        .ZN(n15368) );
  OAI221_X1 U16914 ( .B1(n15369), .B2(keyinput37), .C1(n9297), .C2(keyinput11), 
        .A(n15368), .ZN(n15374) );
  AOI22_X1 U16915 ( .A1(n15372), .A2(keyinput54), .B1(n15371), .B2(keyinput9), 
        .ZN(n15370) );
  OAI221_X1 U16916 ( .B1(n15372), .B2(keyinput54), .C1(n15371), .C2(keyinput9), 
        .A(n15370), .ZN(n15373) );
  NOR4_X1 U16917 ( .A1(n15376), .A2(n15375), .A3(n15374), .A4(n15373), .ZN(
        n15377) );
  NAND4_X1 U16918 ( .A1(n15380), .A2(n15379), .A3(n15378), .A4(n15377), .ZN(
        n15448) );
  AOI22_X1 U16919 ( .A1(n15383), .A2(keyinput107), .B1(keyinput38), .B2(n15382), .ZN(n15381) );
  OAI221_X1 U16920 ( .B1(n15383), .B2(keyinput107), .C1(n15382), .C2(
        keyinput38), .A(n15381), .ZN(n15395) );
  INV_X1 U16921 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n15386) );
  AOI22_X1 U16922 ( .A1(n15386), .A2(keyinput41), .B1(keyinput26), .B2(n15385), 
        .ZN(n15384) );
  OAI221_X1 U16923 ( .B1(n15386), .B2(keyinput41), .C1(n15385), .C2(keyinput26), .A(n15384), .ZN(n15394) );
  INV_X1 U16924 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n15389) );
  INV_X1 U16925 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15388) );
  AOI22_X1 U16926 ( .A1(n15389), .A2(keyinput105), .B1(keyinput77), .B2(n15388), .ZN(n15387) );
  OAI221_X1 U16927 ( .B1(n15389), .B2(keyinput105), .C1(n15388), .C2(
        keyinput77), .A(n15387), .ZN(n15393) );
  XNOR2_X1 U16928 ( .A(P2_REG0_REG_30__SCAN_IN), .B(keyinput68), .ZN(n15391)
         );
  XNOR2_X1 U16929 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput103), .ZN(n15390) );
  NAND2_X1 U16930 ( .A1(n15391), .A2(n15390), .ZN(n15392) );
  NOR4_X1 U16931 ( .A1(n15395), .A2(n15394), .A3(n15393), .A4(n15392), .ZN(
        n15446) );
  INV_X1 U16932 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n15398) );
  AOI22_X1 U16933 ( .A1(n15398), .A2(keyinput100), .B1(n15397), .B2(keyinput55), .ZN(n15396) );
  OAI221_X1 U16934 ( .B1(n15398), .B2(keyinput100), .C1(n15397), .C2(
        keyinput55), .A(n15396), .ZN(n15411) );
  INV_X1 U16935 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n15405) );
  XNOR2_X1 U16936 ( .A(n15399), .B(keyinput71), .ZN(n15402) );
  XNOR2_X1 U16937 ( .A(n15400), .B(keyinput35), .ZN(n15401) );
  NOR2_X1 U16938 ( .A1(n15402), .A2(n15401), .ZN(n15404) );
  XNOR2_X1 U16939 ( .A(P2_REG1_REG_28__SCAN_IN), .B(keyinput102), .ZN(n15403)
         );
  OAI211_X1 U16940 ( .C1(keyinput127), .C2(n15405), .A(n15404), .B(n15403), 
        .ZN(n15410) );
  XNOR2_X1 U16941 ( .A(n15406), .B(keyinput87), .ZN(n15409) );
  XNOR2_X1 U16942 ( .A(keyinput82), .B(n15407), .ZN(n15408) );
  NOR4_X1 U16943 ( .A1(n15411), .A2(n15410), .A3(n15409), .A4(n15408), .ZN(
        n15445) );
  AOI22_X1 U16944 ( .A1(n12265), .A2(keyinput90), .B1(n15413), .B2(keyinput47), 
        .ZN(n15412) );
  OAI221_X1 U16945 ( .B1(n12265), .B2(keyinput90), .C1(n15413), .C2(keyinput47), .A(n15412), .ZN(n15426) );
  AOI22_X1 U16946 ( .A1(n15416), .A2(keyinput94), .B1(n15415), .B2(keyinput101), .ZN(n15414) );
  OAI221_X1 U16947 ( .B1(n15416), .B2(keyinput94), .C1(n15415), .C2(
        keyinput101), .A(n15414), .ZN(n15425) );
  AOI22_X1 U16948 ( .A1(n15419), .A2(keyinput15), .B1(n15418), .B2(keyinput74), 
        .ZN(n15417) );
  OAI221_X1 U16949 ( .B1(n15419), .B2(keyinput15), .C1(n15418), .C2(keyinput74), .A(n15417), .ZN(n15424) );
  INV_X1 U16950 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U16951 ( .A1(n15422), .A2(keyinput36), .B1(n15421), .B2(keyinput62), 
        .ZN(n15420) );
  OAI221_X1 U16952 ( .B1(n15422), .B2(keyinput36), .C1(n15421), .C2(keyinput62), .A(n15420), .ZN(n15423) );
  NOR4_X1 U16953 ( .A1(n15426), .A2(n15425), .A3(n15424), .A4(n15423), .ZN(
        n15444) );
  AOI22_X1 U16954 ( .A1(n15429), .A2(keyinput6), .B1(n15428), .B2(keyinput67), 
        .ZN(n15427) );
  OAI221_X1 U16955 ( .B1(n15429), .B2(keyinput6), .C1(n15428), .C2(keyinput67), 
        .A(n15427), .ZN(n15442) );
  INV_X1 U16956 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U16957 ( .A1(n15432), .A2(keyinput78), .B1(keyinput56), .B2(n15431), 
        .ZN(n15430) );
  OAI221_X1 U16958 ( .B1(n15432), .B2(keyinput78), .C1(n15431), .C2(keyinput56), .A(n15430), .ZN(n15441) );
  AOI22_X1 U16959 ( .A1(n15435), .A2(keyinput104), .B1(keyinput93), .B2(n15434), .ZN(n15433) );
  OAI221_X1 U16960 ( .B1(n15435), .B2(keyinput104), .C1(n15434), .C2(
        keyinput93), .A(n15433), .ZN(n15440) );
  AOI22_X1 U16961 ( .A1(n15438), .A2(keyinput79), .B1(n15437), .B2(keyinput19), 
        .ZN(n15436) );
  OAI221_X1 U16962 ( .B1(n15438), .B2(keyinput79), .C1(n15437), .C2(keyinput19), .A(n15436), .ZN(n15439) );
  NOR4_X1 U16963 ( .A1(n15442), .A2(n15441), .A3(n15440), .A4(n15439), .ZN(
        n15443) );
  NAND4_X1 U16964 ( .A1(n15446), .A2(n15445), .A3(n15444), .A4(n15443), .ZN(
        n15447) );
  NOR4_X1 U16965 ( .A1(n15450), .A2(n15449), .A3(n15448), .A4(n15447), .ZN(
        n15451) );
  OAI21_X1 U16966 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(n15452), .A(n15451), 
        .ZN(n15460) );
  INV_X1 U16967 ( .A(n15453), .ZN(n15457) );
  OAI222_X1 U16968 ( .A1(n15458), .A2(n15457), .B1(n15456), .B2(n15455), .C1(
        n15454), .C2(P3_U3151), .ZN(n15459) );
  XNOR2_X1 U16969 ( .A(n15460), .B(n15459), .ZN(P3_U3284) );
  XOR2_X1 U16970 ( .A(n15462), .B(n15461), .Z(SUB_1596_U59) );
  XNOR2_X1 U16971 ( .A(n15463), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16972 ( .B1(n15465), .B2(n15464), .A(n15473), .ZN(SUB_1596_U53) );
  XOR2_X1 U16973 ( .A(n15466), .B(n15467), .Z(SUB_1596_U56) );
  OAI21_X1 U16974 ( .B1(n15470), .B2(n15469), .A(n15468), .ZN(n15471) );
  XNOR2_X1 U16975 ( .A(n15471), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16976 ( .A(n15472), .B(n15473), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7361 ( .A(n12464), .Z(n6962) );
  NOR4_X1 U7370 ( .A1(n12345), .A2(n12344), .A3(n12343), .A4(n12342), .ZN(
        n12350) );
endmodule

