

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669;

  INV_X1 U7145 ( .A(n14978), .ZN(n14903) );
  MUX2_X1 U7146 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13860), .S(n15454), .Z(
        n13749) );
  INV_X1 U7147 ( .A(n15262), .ZN(n14971) );
  INV_X4 U7148 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7149 ( .A1(n14911), .A2(n14912), .ZN(n14910) );
  NAND2_X1 U7150 ( .A1(n14766), .A2(n14788), .ZN(n15025) );
  INV_X2 U7151 ( .A(n15260), .ZN(n14798) );
  NOR2_X2 U7152 ( .A1(n14841), .A2(n7871), .ZN(n14766) );
  NAND2_X1 U7153 ( .A1(n9786), .A2(n9785), .ZN(n13880) );
  CLKBUF_X1 U7154 ( .A(n9256), .Z(n15071) );
  NAND2_X1 U7155 ( .A1(n11238), .A2(n11242), .ZN(n11237) );
  AND2_X1 U7156 ( .A1(n9230), .A2(n8758), .ZN(n10783) );
  INV_X1 U7157 ( .A(n14466), .ZN(n9063) );
  INV_X1 U7158 ( .A(n8382), .ZN(n8218) );
  NAND4_X2 U7160 ( .A1(n8735), .A2(n8733), .A3(n8734), .A4(n7014), .ZN(n14581)
         );
  INV_X4 U7162 ( .A(n7960), .ZN(n8386) );
  INV_X2 U7163 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13905) );
  INV_X1 U7164 ( .A(n13277), .ZN(n13224) );
  AND2_X1 U7165 ( .A1(n13674), .A2(n7342), .ZN(n7346) );
  NAND2_X1 U7166 ( .A1(n6933), .A2(n6932), .ZN(n8453) );
  INV_X2 U7167 ( .A(n6425), .ZN(n12214) );
  NOR2_X1 U7168 ( .A1(n13674), .A2(n7518), .ZN(n7517) );
  INV_X4 U7169 ( .A(n14011), .ZN(n10284) );
  AND2_X1 U7170 ( .A1(n10284), .A2(n10283), .ZN(n14108) );
  INV_X1 U7171 ( .A(n14108), .ZN(n14052) );
  INV_X1 U7172 ( .A(n8755), .ZN(n9062) );
  INV_X1 U7174 ( .A(n12695), .ZN(n12419) );
  INV_X2 U7175 ( .A(n8390), .ZN(n7997) );
  NAND2_X1 U7176 ( .A1(n10633), .A2(n7378), .ZN(n7377) );
  NAND2_X1 U7177 ( .A1(n6479), .A2(n12658), .ZN(n12657) );
  INV_X1 U7178 ( .A(n7918), .ZN(n8217) );
  NAND2_X1 U7179 ( .A1(n11966), .A2(n11777), .ZN(n8475) );
  INV_X2 U7180 ( .A(n10126), .ZN(n9385) );
  AND3_X1 U7181 ( .A1(n7996), .A2(n7995), .A3(n7994), .ZN(n11121) );
  NAND2_X1 U7182 ( .A1(n8428), .A2(n8421), .ZN(n9326) );
  INV_X1 U7183 ( .A(n9510), .ZN(n12277) );
  AND2_X1 U7184 ( .A1(n14007), .A2(n14006), .ZN(n14246) );
  INV_X1 U7185 ( .A(n12290), .ZN(n7789) );
  NAND2_X1 U7187 ( .A1(n9280), .A2(n9279), .ZN(n14111) );
  AND2_X1 U7188 ( .A1(n8832), .A2(n8831), .ZN(n15298) );
  XNOR2_X1 U7189 ( .A(n7377), .B(n10635), .ZN(n10875) );
  INV_X2 U7190 ( .A(n8171), .ZN(n8381) );
  NOR2_X1 U7191 ( .A1(n13480), .A2(n9821), .ZN(n13493) );
  MUX2_X1 U7192 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13860), .S(n15448), .Z(
        n13861) );
  NAND2_X1 U7193 ( .A1(n9601), .A2(n9600), .ZN(n13145) );
  NAND2_X1 U7195 ( .A1(n9101), .A2(n9100), .ZN(n15030) );
  AOI211_X1 U7196 ( .C1(n7040), .C2(n14601), .A(n14600), .B(n14599), .ZN(
        n15223) );
  AND2_X2 U7197 ( .A1(n14395), .A2(n14872), .ZN(n14912) );
  OR2_X1 U7198 ( .A1(n10300), .A2(n10297), .ZN(n15236) );
  INV_X1 U7199 ( .A(n10283), .ZN(n15240) );
  AOI211_X1 U7200 ( .C1(n15006), .C2(n15315), .A(n15005), .B(n15004), .ZN(
        n15007) );
  NAND2_X1 U7201 ( .A1(n15134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8630) );
  OR2_X1 U7202 ( .A1(n8856), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U7203 ( .A1(n7236), .A2(n7234), .ZN(n7895) );
  NAND4_X2 U7204 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n13353)
         );
  INV_X1 U7206 ( .A(n14798), .ZN(n15269) );
  INV_X1 U7207 ( .A(n13264), .ZN(n9556) );
  NAND2_X2 U7208 ( .A1(n9372), .A2(n9371), .ZN(n10622) );
  AND2_X2 U7209 ( .A1(n7731), .A2(n7730), .ZN(n6479) );
  OR2_X2 U7210 ( .A1(n8964), .A2(n6857), .ZN(n6716) );
  NAND2_X2 U7211 ( .A1(n8680), .A2(n8679), .ZN(n8964) );
  NOR2_X2 U7212 ( .A1(n10985), .A2(n13119), .ZN(n10748) );
  OAI211_X2 U7213 ( .C1(n9536), .C2(n9967), .A(n9535), .B(n9534), .ZN(n13119)
         );
  NOR2_X2 U7214 ( .A1(n7364), .A2(n7771), .ZN(n7021) );
  INV_X4 U7215 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7039) );
  INV_X4 U7216 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7040) );
  XNOR2_X2 U7217 ( .A(n12248), .B(n12247), .ZN(n13051) );
  NAND2_X2 U7218 ( .A1(n8454), .A2(n8453), .ZN(n11164) );
  NOR2_X2 U7219 ( .A1(n6411), .A2(n14927), .ZN(n7022) );
  AND2_X2 U7220 ( .A1(n7499), .A2(n7495), .ZN(n9858) );
  NAND2_X1 U7221 ( .A1(n9286), .A2(n9290), .ZN(n6397) );
  NAND2_X2 U7222 ( .A1(n9286), .A2(n9290), .ZN(n8755) );
  AOI21_X2 U7223 ( .B1(n13571), .B2(n9784), .A(n6453), .ZN(n7532) );
  XNOR2_X1 U7224 ( .A(n9443), .B(n9446), .ZN(n13325) );
  XNOR2_X2 U7225 ( .A(n13828), .B(n9843), .ZN(n13674) );
  XNOR2_X2 U7226 ( .A(n6761), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9481) );
  OAI21_X2 U7227 ( .B1(n7210), .B2(n6450), .A(n6655), .ZN(n12746) );
  CLKBUF_X2 U7228 ( .A(n10402), .Z(n6399) );
  XNOR2_X1 U7229 ( .A(n6750), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10402) );
  CLKBUF_X3 U7230 ( .A(n9556), .Z(n6400) );
  NAND2_X1 U7231 ( .A1(n10089), .A2(n9464), .ZN(n13264) );
  OAI21_X2 U7232 ( .B1(n15211), .B2(n10193), .A(n10192), .ZN(n10191) );
  OR2_X2 U7233 ( .A1(n13471), .A2(n13472), .ZN(n13474) );
  XNOR2_X2 U7234 ( .A(n9477), .B(n9476), .ZN(n9480) );
  NAND2_X2 U7235 ( .A1(n6605), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9477) );
  AOI21_X1 U7236 ( .B1(n13326), .B2(n6398), .A(n13324), .ZN(n13327) );
  AND2_X1 U7237 ( .A1(n7787), .A2(n7786), .ZN(n14734) );
  NAND2_X1 U7238 ( .A1(n12370), .A2(n12317), .ZN(n12437) );
  AOI21_X1 U7239 ( .B1(n12331), .B2(n12330), .A(n12332), .ZN(n12418) );
  NAND2_X1 U7240 ( .A1(n7762), .A2(n7761), .ZN(n12823) );
  INV_X1 U7241 ( .A(n13515), .ZN(n6401) );
  NAND2_X1 U7242 ( .A1(n12271), .A2(n12270), .ZN(n13765) );
  AND2_X2 U7243 ( .A1(n14777), .A2(n14214), .ZN(n14747) );
  NAND2_X1 U7244 ( .A1(n9737), .A2(n9736), .ZN(n13809) );
  OR2_X1 U7245 ( .A1(n15078), .A2(n15082), .ZN(n14390) );
  CLKBUF_X1 U7246 ( .A(n15102), .Z(n7165) );
  XNOR2_X1 U7247 ( .A(n8982), .B(n8981), .ZN(n10825) );
  XNOR2_X1 U7248 ( .A(n9072), .B(SI_20_), .ZN(n9099) );
  NAND2_X1 U7249 ( .A1(n8954), .A2(n8953), .ZN(n15086) );
  INV_X2 U7250 ( .A(n13687), .ZN(n6402) );
  CLKBUF_X2 U7251 ( .A(P2_U3947), .Z(n6404) );
  INV_X1 U7252 ( .A(n15246), .ZN(n15285) );
  INV_X2 U7253 ( .A(n10805), .ZN(n7152) );
  NAND4_X1 U7254 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n14579)
         );
  NAND4_X1 U7255 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .ZN(n15250)
         );
  INV_X1 U7256 ( .A(n12457), .ZN(n6933) );
  INV_X1 U7257 ( .A(n11419), .ZN(n6932) );
  INV_X1 U7258 ( .A(n12454), .ZN(n11777) );
  NAND2_X1 U7259 ( .A1(n10836), .A2(n11412), .ZN(n8555) );
  NAND4_X1 U7261 ( .A1(n9541), .A2(n9540), .A3(n9539), .A4(n9538), .ZN(n13352)
         );
  INV_X1 U7262 ( .A(n15458), .ZN(n10587) );
  XNOR2_X1 U7263 ( .A(n10406), .B(n10455), .ZN(n10448) );
  BUF_X1 U7265 ( .A(n9510), .Z(n13100) );
  BUF_X1 U7266 ( .A(n9290), .Z(n6410) );
  CLKBUF_X2 U7267 ( .A(n9509), .Z(n9479) );
  INV_X2 U7268 ( .A(n10089), .ZN(n9735) );
  NAND2_X2 U7269 ( .A1(n6670), .A2(n6669), .ZN(n13328) );
  AND2_X1 U7270 ( .A1(n6675), .A2(n6531), .ZN(n6669) );
  INV_X4 U7271 ( .A(n8659), .ZN(n9464) );
  NAND3_X1 U7272 ( .A1(n7318), .A2(n6898), .A3(n6899), .ZN(n8073) );
  AND3_X1 U7273 ( .A1(n7684), .A2(n7683), .A3(n7682), .ZN(n7681) );
  NOR2_X1 U7274 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8624) );
  NOR2_X1 U7275 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8623) );
  NOR2_X1 U7276 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9435) );
  NOR2_X1 U7277 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n9434) );
  NOR2_X1 U7278 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7683) );
  NOR2_X1 U7279 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7684) );
  NOR2_X1 U7280 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n9458) );
  NOR2_X1 U7281 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n9456) );
  AND2_X1 U7282 ( .A1(n7755), .A2(n7753), .ZN(n12849) );
  NOR2_X1 U7283 ( .A1(n12138), .A2(n12129), .ZN(n14712) );
  AND2_X1 U7284 ( .A1(n7137), .A2(n7122), .ZN(n14991) );
  NOR2_X1 U7285 ( .A1(n15015), .A2(n7066), .ZN(n7065) );
  AND2_X1 U7286 ( .A1(n7373), .A2(n15308), .ZN(n14992) );
  OR2_X1 U7287 ( .A1(n15014), .A2(n15013), .ZN(n15120) );
  OAI21_X1 U7288 ( .B1(n14732), .B2(n14733), .A(n14731), .ZN(n14995) );
  OR3_X1 U7289 ( .A1(n15024), .A2(n15023), .A3(n15022), .ZN(n15122) );
  AOI21_X1 U7290 ( .B1(n12134), .B2(n15308), .A(n12133), .ZN(n14716) );
  AOI21_X1 U7291 ( .B1(n14794), .B2(n14793), .A(n14792), .ZN(n14797) );
  NAND2_X1 U7292 ( .A1(n14677), .A2(n15240), .ZN(n14979) );
  NAND2_X1 U7293 ( .A1(n7534), .A2(n7533), .ZN(n13794) );
  NAND2_X1 U7294 ( .A1(n14811), .A2(n14815), .ZN(n14810) );
  OR2_X1 U7295 ( .A1(n13445), .A2(n13444), .ZN(n13748) );
  NAND2_X1 U7296 ( .A1(n12150), .A2(n14545), .ZN(n12149) );
  OR2_X1 U7297 ( .A1(n13594), .A2(n13608), .ZN(n13595) );
  NAND2_X1 U7298 ( .A1(n6678), .A2(n6447), .ZN(n6677) );
  NOR2_X1 U7299 ( .A1(n14993), .A2(n7372), .ZN(n7371) );
  NAND2_X1 U7300 ( .A1(n6680), .A2(n6447), .ZN(n6679) );
  NAND2_X1 U7301 ( .A1(n7810), .A2(n7809), .ZN(n14765) );
  NAND2_X1 U7302 ( .A1(n6929), .A2(n7513), .ZN(n13594) );
  NAND2_X1 U7303 ( .A1(n14747), .A2(n7448), .ZN(n12140) );
  NOR2_X1 U7304 ( .A1(n13517), .A2(n7694), .ZN(n13480) );
  OR2_X1 U7305 ( .A1(n7337), .A2(n6431), .ZN(n7333) );
  OR2_X1 U7306 ( .A1(n6799), .A2(n14074), .ZN(n6798) );
  NAND2_X1 U7307 ( .A1(n7068), .A2(n7067), .ZN(n7066) );
  NAND2_X1 U7308 ( .A1(n12693), .A2(n12692), .ZN(n12691) );
  NAND2_X1 U7309 ( .A1(n14931), .A2(n14930), .ZN(n14929) );
  NAND2_X1 U7310 ( .A1(n13661), .A2(n9845), .ZN(n13640) );
  CLKBUF_X1 U7311 ( .A(n12041), .Z(n12044) );
  AND2_X1 U7312 ( .A1(n7455), .A2(n7454), .ZN(n14074) );
  AND2_X1 U7313 ( .A1(n13657), .A2(n13895), .ZN(n13658) );
  NAND2_X1 U7314 ( .A1(n9796), .A2(n9795), .ZN(n13535) );
  NAND2_X1 U7315 ( .A1(n9630), .A2(n9629), .ZN(n11860) );
  NAND2_X1 U7316 ( .A1(n9761), .A2(n9760), .ZN(n13587) );
  INV_X1 U7317 ( .A(n14962), .ZN(n7444) );
  NAND2_X1 U7318 ( .A1(n9748), .A2(n9747), .ZN(n13804) );
  XNOR2_X1 U7319 ( .A(n9077), .B(n9076), .ZN(n11497) );
  NAND2_X2 U7320 ( .A1(n9689), .A2(n9688), .ZN(n13828) );
  NAND2_X1 U7321 ( .A1(n9676), .A2(n9675), .ZN(n13707) );
  NAND2_X1 U7322 ( .A1(n9043), .A2(n9042), .ZN(n15045) );
  XNOR2_X1 U7323 ( .A(n15102), .B(n15092), .ZN(n14539) );
  NAND2_X1 U7324 ( .A1(n9020), .A2(n9019), .ZN(n15064) );
  NAND2_X1 U7325 ( .A1(n8979), .A2(n8968), .ZN(n10570) );
  INV_X1 U7326 ( .A(n9072), .ZN(n7429) );
  INV_X1 U7327 ( .A(n14359), .ZN(n15108) );
  NAND2_X1 U7328 ( .A1(n11660), .A2(n11659), .ZN(n11661) );
  OR2_X1 U7329 ( .A1(n8967), .A2(n8966), .ZN(n8979) );
  NAND2_X1 U7330 ( .A1(n6852), .A2(n8696), .ZN(n9072) );
  OAI21_X2 U7331 ( .B1(n10256), .B2(n13091), .A(n9619), .ZN(n13152) );
  OAI22_X1 U7332 ( .A1(n11213), .A2(n6992), .B1(n6994), .B2(n6991), .ZN(n11397) );
  XNOR2_X1 U7333 ( .A(n8913), .B(n8912), .ZN(n10422) );
  OR2_X1 U7334 ( .A1(n8964), .A2(n10271), .ZN(n7351) );
  NAND2_X1 U7335 ( .A1(n8911), .A2(n8891), .ZN(n10256) );
  AOI21_X1 U7336 ( .B1(n11801), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11800), .ZN(
        n11802) );
  NAND2_X1 U7337 ( .A1(n10923), .A2(n10924), .ZN(n11213) );
  NAND2_X1 U7338 ( .A1(n6620), .A2(n11462), .ZN(n11577) );
  OR2_X1 U7339 ( .A1(n8890), .A2(n9973), .ZN(n8911) );
  NAND2_X1 U7340 ( .A1(n9589), .A2(n9588), .ZN(n13148) );
  AND3_X1 U7341 ( .A1(n10562), .A2(n10560), .A3(n10561), .ZN(n10762) );
  NAND2_X1 U7342 ( .A1(n8879), .A2(n8878), .ZN(n14355) );
  NAND2_X1 U7343 ( .A1(n7220), .A2(n7218), .ZN(n10951) );
  NAND3_X1 U7344 ( .A1(n10462), .A2(n10461), .A3(n10460), .ZN(n10562) );
  INV_X1 U7345 ( .A(n14348), .ZN(n15303) );
  NAND2_X1 U7346 ( .A1(n9577), .A2(n9576), .ZN(n13136) );
  NAND2_X1 U7347 ( .A1(n10821), .A2(n13683), .ZN(n13087) );
  NAND2_X1 U7348 ( .A1(n10313), .A2(n10314), .ZN(n10462) );
  INV_X1 U7349 ( .A(n15292), .ZN(n6406) );
  AOI21_X1 U7350 ( .B1(n10309), .B2(n10308), .A(n10307), .ZN(n10467) );
  INV_X2 U7351 ( .A(n15323), .ZN(n6403) );
  NAND2_X1 U7352 ( .A1(n9561), .A2(n9560), .ZN(n13129) );
  INV_X2 U7353 ( .A(n11174), .ZN(n12293) );
  AND2_X2 U7355 ( .A1(n14468), .A2(n14310), .ZN(n14448) );
  NAND2_X1 U7356 ( .A1(n7099), .A2(n6773), .ZN(n10976) );
  INV_X1 U7357 ( .A(n11204), .ZN(n14131) );
  NAND2_X1 U7358 ( .A1(n8824), .A2(n7352), .ZN(n8827) );
  NAND3_X2 U7359 ( .A1(n8745), .A2(n8744), .A3(n8743), .ZN(n14580) );
  AND3_X1 U7360 ( .A1(n8775), .A2(n8774), .A3(n8773), .ZN(n15275) );
  OR2_X1 U7361 ( .A1(n10168), .A2(n10167), .ZN(n10346) );
  NAND2_X1 U7362 ( .A1(n8806), .A2(n8662), .ZN(n8824) );
  NAND4_X2 U7363 ( .A1(n7986), .A2(n7985), .A3(n7984), .A4(n7983), .ZN(n12458)
         );
  NAND3_X1 U7364 ( .A1(n7899), .A2(n6420), .A3(n7898), .ZN(n15481) );
  AND2_X1 U7365 ( .A1(n8675), .A2(n7422), .ZN(n7421) );
  NAND4_X1 U7366 ( .A1(n9584), .A2(n9583), .A3(n9582), .A4(n9581), .ZN(n13349)
         );
  CLKBUF_X1 U7367 ( .A(n6449), .Z(n10010) );
  INV_X1 U7368 ( .A(n7415), .ZN(n7414) );
  OR2_X1 U7369 ( .A1(n8759), .A2(n11207), .ZN(n8723) );
  NAND4_X1 U7370 ( .A1(n9572), .A2(n9571), .A3(n9570), .A4(n9569), .ZN(n13350)
         );
  AND3_X1 U7371 ( .A1(n7906), .A2(n7905), .A3(n7904), .ZN(n15476) );
  AND2_X1 U7372 ( .A1(n8852), .A2(n7112), .ZN(n7519) );
  OAI21_X1 U7373 ( .B1(n7417), .B2(n7416), .A(n8687), .ZN(n7415) );
  OR2_X1 U7374 ( .A1(n9510), .A2(n9496), .ZN(n6905) );
  AND2_X1 U7375 ( .A1(n8666), .A2(n6614), .ZN(n8852) );
  AND2_X1 U7376 ( .A1(n9859), .A2(n13433), .ZN(n13111) );
  NAND2_X1 U7378 ( .A1(n7298), .A2(n7896), .ZN(n7982) );
  AOI21_X1 U7379 ( .B1(n8674), .B2(n8931), .A(n8673), .ZN(n8675) );
  NAND2_X2 U7380 ( .A1(n11264), .A2(n11081), .ZN(n10126) );
  NAND2_X1 U7381 ( .A1(n9227), .A2(n9226), .ZN(n11375) );
  MUX2_X1 U7382 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9225), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9226) );
  XNOR2_X1 U7383 ( .A(n9221), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14304) );
  NAND2_X2 U7384 ( .A1(n7895), .A2(n7896), .ZN(n8372) );
  XNOR2_X1 U7385 ( .A(n9440), .B(n9876), .ZN(n9859) );
  NAND2_X1 U7386 ( .A1(n9481), .A2(n9478), .ZN(n9751) );
  OR2_X1 U7387 ( .A1(n8835), .A2(n7520), .ZN(n7112) );
  INV_X2 U7388 ( .A(n11473), .ZN(n12937) );
  INV_X1 U7389 ( .A(n12933), .ZN(n7896) );
  XNOR2_X1 U7390 ( .A(n8417), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11264) );
  XNOR2_X1 U7391 ( .A(n8396), .B(n8582), .ZN(n11564) );
  NAND2_X1 U7392 ( .A1(n13325), .A2(n10800), .ZN(n13284) );
  OR2_X1 U7393 ( .A1(n9481), .A2(n9480), .ZN(n9509) );
  NAND2_X1 U7394 ( .A1(n8716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U7395 ( .A1(n8599), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U7396 ( .A1(n7463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8632) );
  INV_X1 U7397 ( .A(n7368), .ZN(n8835) );
  INV_X1 U7398 ( .A(n13666), .ZN(n13433) );
  CLKBUF_X1 U7399 ( .A(n10800), .Z(n13323) );
  NAND2_X1 U7400 ( .A1(n9875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9440) );
  XNOR2_X1 U7401 ( .A(n9819), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10800) );
  INV_X1 U7402 ( .A(n8966), .ZN(n8681) );
  OAI21_X1 U7403 ( .B1(n7434), .B2(n7094), .A(n7093), .ZN(n8665) );
  NAND2_X1 U7404 ( .A1(n13906), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6761) );
  NAND2_X2 U7405 ( .A1(n7434), .A2(P2_U3088), .ZN(n13913) );
  NAND2_X1 U7406 ( .A1(n9463), .A2(n6608), .ZN(n6670) );
  OAI21_X1 U7407 ( .B1(n9880), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9443) );
  AND2_X1 U7408 ( .A1(n7811), .A2(n8631), .ZN(n7464) );
  NAND2_X1 U7409 ( .A1(n7819), .A2(n7817), .ZN(n6930) );
  AND2_X1 U7410 ( .A1(n8619), .A2(n7788), .ZN(n8627) );
  NAND2_X1 U7411 ( .A1(n6644), .A2(n9515), .ZN(n13362) );
  OR2_X1 U7412 ( .A1(n8073), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7816) );
  AND2_X1 U7413 ( .A1(n7813), .A2(n8715), .ZN(n7811) );
  AND2_X1 U7414 ( .A1(n7331), .A2(n6533), .ZN(n7512) );
  NOR2_X1 U7415 ( .A1(n7814), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U7416 ( .A1(n8732), .A2(n8746), .ZN(n14586) );
  INV_X1 U7417 ( .A(n7318), .ZN(n7931) );
  NOR2_X1 U7418 ( .A1(n9296), .A2(n8856), .ZN(n8626) );
  AND2_X1 U7419 ( .A1(n6662), .A2(n7381), .ZN(n7318) );
  NAND4_X1 U7420 ( .A1(n8985), .A2(n8624), .A3(n8623), .A4(n8984), .ZN(n9038)
         );
  NAND4_X1 U7421 ( .A1(n7901), .A2(n13436), .A3(n7537), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7536) );
  NAND3_X1 U7422 ( .A1(n9457), .A2(n9458), .A3(n9456), .ZN(n9881) );
  NAND4_X1 U7423 ( .A1(n7886), .A2(n8039), .A3(n8011), .A4(n8013), .ZN(n8056)
         );
  NAND4_X1 U7424 ( .A1(n7277), .A2(n7276), .A3(n8132), .A4(n8184), .ZN(n8215)
         );
  NAND3_X1 U7425 ( .A1(n9003), .A2(n7008), .A3(n7007), .ZN(n9037) );
  INV_X1 U7426 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9685) );
  NOR2_X1 U7427 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7886) );
  INV_X1 U7428 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8184) );
  INV_X4 U7429 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7430 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7277) );
  INV_X1 U7431 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8013) );
  INV_X1 U7432 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13436) );
  INV_X1 U7433 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7901) );
  NOR2_X2 U7434 ( .A1(n13479), .A2(n13478), .ZN(n13767) );
  NAND4_X2 U7435 ( .A1(n7444), .A2(n14921), .A3(n7443), .A4(n7447), .ZN(n14892) );
  OR2_X2 U7436 ( .A1(n11642), .A2(n14535), .ZN(n11644) );
  AOI21_X1 U7437 ( .B1(n10557), .B2(n10556), .A(n10555), .ZN(n10767) );
  NOR2_X1 U7438 ( .A1(n11064), .A2(n13129), .ZN(n11249) );
  NAND2_X1 U7439 ( .A1(n10748), .A2(n7686), .ZN(n11064) );
  INV_X1 U7440 ( .A(n7406), .ZN(n7405) );
  INV_X1 U7441 ( .A(n14463), .ZN(n14450) );
  OR2_X1 U7442 ( .A1(n9136), .A2(n14582), .ZN(n8721) );
  NAND2_X4 U7443 ( .A1(n8633), .A2(n7789), .ZN(n9136) );
  OAI21_X2 U7444 ( .B1(n12381), .B2(n7880), .A(n7649), .ZN(n7648) );
  INV_X4 U7445 ( .A(n14455), .ZN(n9209) );
  OAI21_X2 U7446 ( .B1(n9244), .B2(n7043), .A(n7041), .ZN(n11756) );
  OAI211_X1 U7447 ( .C1(n14466), .C2(n9981), .A(n8814), .B(n8813), .ZN(n15292)
         );
  INV_X1 U7448 ( .A(n14463), .ZN(n6408) );
  INV_X1 U7449 ( .A(n14463), .ZN(n6409) );
  NAND2_X2 U7450 ( .A1(n6397), .A2(n9464), .ZN(n14463) );
  OAI21_X2 U7451 ( .B1(n9250), .B2(n7047), .A(n7044), .ZN(n14907) );
  OAI222_X1 U7452 ( .A1(n9286), .A2(P1_U3086), .B1(n15147), .B2(n13914), .C1(
        n12205), .C2(n15144), .ZN(P1_U3327) );
  XNOR2_X1 U7453 ( .A(n8718), .B(n8717), .ZN(n9290) );
  INV_X4 U7454 ( .A(n13091), .ZN(n13262) );
  XNOR2_X2 U7455 ( .A(n7392), .B(n8715), .ZN(n9286) );
  OR2_X2 U7456 ( .A1(n10001), .A2(n10288), .ZN(n14600) );
  NAND2_X1 U7457 ( .A1(n7718), .A2(n13164), .ZN(n7717) );
  OR2_X1 U7458 ( .A1(n12848), .A2(n12451), .ZN(n8414) );
  NAND2_X1 U7459 ( .A1(n10639), .A2(n10640), .ZN(n7273) );
  OR2_X1 U7460 ( .A1(n12850), .A2(n12355), .ZN(n8544) );
  NOR2_X1 U7461 ( .A1(n7736), .A2(n7189), .ZN(n7188) );
  INV_X1 U7462 ( .A(n7193), .ZN(n7189) );
  OR2_X1 U7463 ( .A1(n12340), .A2(n12682), .ZN(n8285) );
  XNOR2_X1 U7464 ( .A(n6652), .B(n7903), .ZN(n8602) );
  NAND2_X1 U7465 ( .A1(n6653), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6652) );
  AND2_X1 U7466 ( .A1(n8216), .A2(n7820), .ZN(n6654) );
  AOI21_X1 U7467 ( .B1(n6828), .B2(n6830), .A(n6589), .ZN(n6826) );
  NAND2_X1 U7468 ( .A1(n6675), .A2(n6674), .ZN(n6673) );
  NOR2_X1 U7469 ( .A1(n9462), .A2(n13905), .ZN(n6674) );
  INV_X1 U7470 ( .A(n6541), .ZN(n7473) );
  INV_X1 U7471 ( .A(n14048), .ZN(n7474) );
  INV_X2 U7472 ( .A(n14111), .ZN(n14051) );
  NAND2_X1 U7473 ( .A1(n14439), .A2(n14438), .ZN(n14445) );
  OR2_X1 U7474 ( .A1(n9193), .A2(n9192), .ZN(n9208) );
  INV_X1 U7475 ( .A(n14572), .ZN(n14010) );
  AND2_X2 U7476 ( .A1(n9285), .A2(n11375), .ZN(n14479) );
  AND2_X1 U7477 ( .A1(n7742), .A2(n7200), .ZN(n7199) );
  INV_X1 U7478 ( .A(n7749), .ZN(n7742) );
  NAND2_X1 U7479 ( .A1(n12647), .A2(n8524), .ZN(n7200) );
  OR2_X1 U7480 ( .A1(n10126), .A2(n9360), .ZN(n15469) );
  AND2_X1 U7481 ( .A1(n9385), .A2(n9360), .ZN(n12704) );
  NAND2_X1 U7482 ( .A1(n13331), .A2(n13323), .ZN(n10812) );
  OR3_X1 U7483 ( .A1(n15415), .A2(n10811), .A3(n10972), .ZN(n10819) );
  AND2_X1 U7484 ( .A1(n7529), .A2(n6459), .ZN(n7339) );
  NAND2_X1 U7485 ( .A1(n6864), .A2(n6459), .ZN(n7338) );
  INV_X1 U7486 ( .A(n14280), .ZN(n7475) );
  NAND2_X1 U7487 ( .A1(n7806), .A2(n9271), .ZN(n7061) );
  NAND2_X1 U7488 ( .A1(n14765), .A2(n9268), .ZN(n12146) );
  INV_X1 U7489 ( .A(n8759), .ZN(n9210) );
  NAND2_X1 U7490 ( .A1(n14359), .A2(n14574), .ZN(n8909) );
  NAND2_X1 U7491 ( .A1(n7040), .A2(n7039), .ZN(n8746) );
  OR2_X1 U7492 ( .A1(n13277), .A2(n13113), .ZN(n7705) );
  NAND2_X1 U7493 ( .A1(n7086), .A2(n7085), .ZN(n13115) );
  NAND2_X1 U7494 ( .A1(n13277), .A2(n13113), .ZN(n7085) );
  OR2_X1 U7495 ( .A1(n6602), .A2(n13277), .ZN(n7086) );
  NAND2_X1 U7496 ( .A1(n13146), .A2(n7715), .ZN(n7714) );
  NAND2_X1 U7497 ( .A1(n6776), .A2(n13171), .ZN(n6775) );
  NAND2_X1 U7498 ( .A1(n14309), .A2(n14307), .ZN(n14472) );
  AOI21_X1 U7499 ( .B1(n8536), .B2(n7305), .A(n6507), .ZN(n7304) );
  INV_X1 U7500 ( .A(n8533), .ZN(n7305) );
  NAND2_X1 U7501 ( .A1(n8537), .A2(n9391), .ZN(n8538) );
  OR2_X1 U7502 ( .A1(n12867), .A2(n12644), .ZN(n7870) );
  NOR2_X2 U7503 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n9457) );
  NOR2_X1 U7504 ( .A1(n6871), .A2(n8706), .ZN(n6870) );
  INV_X1 U7505 ( .A(n6872), .ZN(n6871) );
  NOR2_X1 U7506 ( .A1(n9075), .A2(SI_21_), .ZN(n8698) );
  AOI21_X1 U7507 ( .B1(n7414), .B2(n6856), .A(n6510), .ZN(n6855) );
  NOR2_X1 U7508 ( .A1(n7413), .A2(n8689), .ZN(n6856) );
  NAND2_X1 U7509 ( .A1(n7414), .A2(n6858), .ZN(n6857) );
  INV_X1 U7510 ( .A(n8689), .ZN(n6858) );
  OAI21_X1 U7511 ( .B1(n7434), .B2(P2_DATAO_REG_15__SCAN_IN), .A(n6613), .ZN(
        n8684) );
  NAND2_X1 U7512 ( .A1(n7434), .A2(n10827), .ZN(n6613) );
  NAND2_X1 U7513 ( .A1(n6877), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U7514 ( .A1(n12614), .A2(n9426), .ZN(n8537) );
  OR2_X1 U7515 ( .A1(n12614), .A2(n9426), .ZN(n8539) );
  NAND2_X1 U7516 ( .A1(n6461), .A2(n9334), .ZN(n7221) );
  OR2_X1 U7517 ( .A1(n12893), .A2(n12732), .ZN(n8553) );
  AND2_X1 U7518 ( .A1(n8418), .A2(n8498), .ZN(n12711) );
  AND2_X1 U7519 ( .A1(n7852), .A2(n6514), .ZN(n7214) );
  NAND2_X1 U7520 ( .A1(n11966), .A2(n12454), .ZN(n7859) );
  INV_X1 U7521 ( .A(n7562), .ZN(n7561) );
  OAI21_X1 U7522 ( .B1(n8168), .B2(n7563), .A(n8196), .ZN(n7562) );
  NOR2_X1 U7523 ( .A1(n7554), .A2(n7550), .ZN(n7549) );
  INV_X1 U7524 ( .A(n8008), .ZN(n7550) );
  INV_X1 U7525 ( .A(n8027), .ZN(n7554) );
  OR2_X1 U7526 ( .A1(n7916), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n7968) );
  INV_X1 U7527 ( .A(n12230), .ZN(n7596) );
  NOR2_X1 U7528 ( .A1(n12990), .A2(n12238), .ZN(n7604) );
  INV_X1 U7529 ( .A(n7333), .ZN(n6680) );
  AOI21_X1 U7530 ( .B1(n7514), .B2(n6519), .A(n6430), .ZN(n7513) );
  NAND2_X1 U7531 ( .A1(n6683), .A2(n6685), .ZN(n6681) );
  XNOR2_X1 U7532 ( .A(n13113), .B(n10801), .ZN(n7099) );
  NAND2_X1 U7533 ( .A1(n7483), .A2(n6473), .ZN(n12177) );
  NAND2_X1 U7534 ( .A1(n11939), .A2(n7485), .ZN(n7483) );
  AND2_X1 U7535 ( .A1(n14139), .A2(n6468), .ZN(n7461) );
  AND2_X1 U7536 ( .A1(n11443), .A2(n14177), .ZN(n6814) );
  NAND2_X1 U7537 ( .A1(n7411), .A2(n7410), .ZN(n14513) );
  NAND2_X1 U7538 ( .A1(n14461), .A2(n14460), .ZN(n7410) );
  AND2_X1 U7539 ( .A1(n7780), .A2(n6555), .ZN(n7024) );
  AND2_X1 U7540 ( .A1(n7063), .A2(n14733), .ZN(n7062) );
  OR2_X1 U7541 ( .A1(n7802), .A2(n7064), .ZN(n7063) );
  NOR2_X1 U7542 ( .A1(n14746), .A2(n7785), .ZN(n7784) );
  INV_X1 U7543 ( .A(n9143), .ZN(n7785) );
  INV_X1 U7544 ( .A(n14535), .ZN(n7043) );
  NAND2_X1 U7545 ( .A1(n14131), .A2(n7111), .ZN(n14317) );
  OAI21_X1 U7546 ( .B1(n9204), .B2(n9203), .A(n9205), .ZN(n12197) );
  XNOR2_X1 U7547 ( .A(n8671), .B(SI_11_), .ZN(n8912) );
  OR2_X1 U7548 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  OAI21_X1 U7549 ( .B1(n12402), .B2(n12372), .A(n12371), .ZN(n12370) );
  INV_X1 U7550 ( .A(n8372), .ZN(n8385) );
  NAND2_X1 U7551 ( .A1(n10520), .A2(n8421), .ZN(n10581) );
  NAND2_X1 U7552 ( .A1(n12297), .A2(n12770), .ZN(n7649) );
  AND4_X1 U7553 ( .A1(n6484), .A2(n7861), .A3(n7543), .A4(n6524), .ZN(n8572)
         );
  AND4_X1 U7555 ( .A1(n8049), .A2(n8048), .A3(n8047), .A4(n8046), .ZN(n11431)
         );
  OR2_X1 U7556 ( .A1(n10640), .A2(n10401), .ZN(n7378) );
  NAND2_X1 U7557 ( .A1(n6419), .A2(n10878), .ZN(n7665) );
  OR2_X1 U7558 ( .A1(n7666), .A2(n10635), .ZN(n7664) );
  NAND2_X1 U7559 ( .A1(n7270), .A2(n7273), .ZN(n7269) );
  AOI21_X1 U7560 ( .B1(n10549), .B2(n7274), .A(n7272), .ZN(n7271) );
  NAND2_X1 U7561 ( .A1(n7377), .A2(n10878), .ZN(n6748) );
  NAND2_X1 U7562 ( .A1(n10875), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U7563 ( .A1(n6940), .A2(n6941), .ZN(n6939) );
  AND2_X1 U7564 ( .A1(n6943), .A2(n6535), .ZN(n6940) );
  NAND2_X1 U7565 ( .A1(n11536), .A2(n6942), .ZN(n6938) );
  NAND2_X1 U7566 ( .A1(n7746), .A2(n12647), .ZN(n7198) );
  NAND2_X1 U7567 ( .A1(n8334), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8335) );
  AOI21_X1 U7568 ( .B1(n8516), .B2(n8508), .A(n8519), .ZN(n7730) );
  INV_X1 U7569 ( .A(n12596), .ZN(n12593) );
  OR2_X1 U7570 ( .A1(n8382), .A2(n9931), .ZN(n7905) );
  NOR2_X1 U7571 ( .A1(n12355), .A2(n15469), .ZN(n9361) );
  NAND2_X1 U7572 ( .A1(n8332), .A2(n8331), .ZN(n12793) );
  OR2_X1 U7573 ( .A1(n12884), .A2(n12718), .ZN(n7740) );
  XNOR2_X1 U7574 ( .A(n12884), .B(n12718), .ZN(n12702) );
  NAND2_X1 U7575 ( .A1(n7192), .A2(n8553), .ZN(n12701) );
  NAND2_X1 U7576 ( .A1(n12823), .A2(n7193), .ZN(n7192) );
  OR2_X1 U7577 ( .A1(n12738), .A2(n12749), .ZN(n8418) );
  INV_X1 U7578 ( .A(n7851), .ZN(n7210) );
  NAND2_X1 U7579 ( .A1(n7851), .A2(n7214), .ZN(n7212) );
  AND2_X1 U7580 ( .A1(n9401), .A2(n11564), .ZN(n12829) );
  AND2_X1 U7581 ( .A1(n12922), .A2(n10233), .ZN(n10252) );
  NOR2_X1 U7582 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n6898) );
  NOR2_X1 U7583 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n6899) );
  OAI211_X1 U7584 ( .C1(n7577), .C2(n6840), .A(n6586), .B(n6836), .ZN(n8352)
         );
  INV_X1 U7585 ( .A(n6842), .ZN(n6840) );
  NAND2_X1 U7586 ( .A1(n6837), .A2(n6443), .ZN(n6836) );
  OAI211_X1 U7587 ( .C1(n8300), .C2(n7579), .A(n7577), .B(n8316), .ZN(n8329)
         );
  NAND2_X1 U7588 ( .A1(n8258), .A2(n8257), .ZN(n7557) );
  OAI21_X1 U7589 ( .B1(P1_DATAO_REG_20__SCAN_IN), .B2(n11374), .A(n8259), .ZN(
        n8256) );
  AND2_X1 U7590 ( .A1(n8231), .A2(n8214), .ZN(n8229) );
  OR2_X1 U7591 ( .A1(n8113), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U7592 ( .A1(n8110), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8127) );
  NOR2_X2 U7593 ( .A1(n8073), .A2(n8056), .ZN(n8591) );
  OAI21_X1 U7594 ( .B1(n12982), .B2(n7004), .A(n7001), .ZN(n12971) );
  AOI21_X1 U7595 ( .B1(n7003), .B2(n7601), .A(n7002), .ZN(n7001) );
  INV_X1 U7596 ( .A(n7601), .ZN(n7004) );
  INV_X1 U7597 ( .A(n12247), .ZN(n7002) );
  NAND2_X1 U7598 ( .A1(n12982), .A2(n12235), .ZN(n13040) );
  XNOR2_X1 U7599 ( .A(n10805), .B(n6425), .ZN(n10808) );
  NAND2_X1 U7600 ( .A1(n6723), .A2(n6421), .ZN(n13319) );
  INV_X1 U7601 ( .A(n9479), .ZN(n12278) );
  OR2_X1 U7602 ( .A1(n9510), .A2(n6895), .ZN(n9506) );
  NAND2_X1 U7603 ( .A1(n9503), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9504) );
  OR2_X1 U7604 ( .A1(n9509), .A2(n10142), .ZN(n9505) );
  OR2_X1 U7605 ( .A1(n9659), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9684) );
  NOR2_X1 U7606 ( .A1(n13765), .A2(n7691), .ZN(n7690) );
  NAND2_X1 U7607 ( .A1(n13762), .A2(n7692), .ZN(n7691) );
  INV_X1 U7608 ( .A(n9784), .ZN(n7530) );
  AOI21_X1 U7609 ( .B1(n6921), .B2(n9853), .A(n6503), .ZN(n6922) );
  NAND2_X1 U7610 ( .A1(n13627), .A2(n6924), .ZN(n6923) );
  NAND2_X1 U7611 ( .A1(n6666), .A2(n6665), .ZN(n13704) );
  AND2_X1 U7612 ( .A1(n7524), .A2(n9673), .ZN(n6666) );
  AND2_X1 U7613 ( .A1(n13703), .A2(n9839), .ZN(n9840) );
  XNOR2_X1 U7614 ( .A(n7105), .B(n13345), .ZN(n13315) );
  NAND2_X1 U7615 ( .A1(n10705), .A2(n9508), .ZN(n10980) );
  NOR2_X1 U7616 ( .A1(n10811), .A2(n9906), .ZN(n10712) );
  NAND2_X1 U7617 ( .A1(n13266), .A2(n13265), .ZN(n13437) );
  NAND2_X1 U7618 ( .A1(n9909), .A2(n9908), .ZN(n10972) );
  NOR2_X1 U7619 ( .A1(n13905), .A2(n7151), .ZN(n6608) );
  NAND2_X1 U7620 ( .A1(n9877), .A2(n9876), .ZN(n9910) );
  OR2_X1 U7621 ( .A1(n9532), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9543) );
  AOI21_X1 U7622 ( .B1(n7472), .B2(n7475), .A(n7469), .ZN(n7468) );
  INV_X1 U7623 ( .A(n14058), .ZN(n7469) );
  NAND2_X1 U7624 ( .A1(n6782), .A2(n10894), .ZN(n7477) );
  AND2_X1 U7625 ( .A1(n14048), .A2(n14046), .ZN(n14156) );
  XNOR2_X1 U7626 ( .A(n6783), .B(n14111), .ZN(n10654) );
  NAND2_X1 U7627 ( .A1(n10649), .A2(n6784), .ZN(n6783) );
  NAND2_X1 U7628 ( .A1(n9228), .A2(n10286), .ZN(n6784) );
  AND2_X1 U7629 ( .A1(n6541), .A2(n6708), .ZN(n14280) );
  NAND2_X1 U7630 ( .A1(n14057), .A2(n14056), .ZN(n6708) );
  AOI21_X1 U7631 ( .B1(n14700), .B2(n9216), .A(n9215), .ZN(n14484) );
  AND2_X1 U7632 ( .A1(n8639), .A2(n8638), .ZN(n14042) );
  NAND2_X2 U7633 ( .A1(n12203), .A2(n7789), .ZN(n14455) );
  NAND3_X1 U7634 ( .A1(n9308), .A2(n9311), .A3(n9309), .ZN(n10288) );
  NOR2_X1 U7635 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  NOR2_X1 U7636 ( .A1(n7449), .A2(n14449), .ZN(n7448) );
  INV_X1 U7637 ( .A(n7450), .ZN(n7449) );
  NAND2_X1 U7638 ( .A1(n12128), .A2(n12127), .ZN(n14547) );
  XNOR2_X1 U7639 ( .A(n14985), .B(n14567), .ZN(n14718) );
  OR2_X1 U7640 ( .A1(n15006), .A2(n14160), .ZN(n9143) );
  NAND2_X1 U7641 ( .A1(n12149), .A2(n7784), .ZN(n7787) );
  NAND2_X1 U7642 ( .A1(n14825), .A2(n7354), .ZN(n7810) );
  NOR2_X1 U7643 ( .A1(n9265), .A2(n7355), .ZN(n7354) );
  INV_X1 U7644 ( .A(n9264), .ZN(n7355) );
  NOR2_X1 U7645 ( .A1(n14790), .A2(n7440), .ZN(n7439) );
  INV_X1 U7646 ( .A(n7441), .ZN(n7440) );
  AND2_X1 U7647 ( .A1(n9033), .A2(n7365), .ZN(n7364) );
  NAND2_X1 U7648 ( .A1(n14912), .A2(n7366), .ZN(n7365) );
  NOR2_X1 U7649 ( .A1(n8851), .A2(n7776), .ZN(n7775) );
  INV_X1 U7650 ( .A(n8833), .ZN(n7776) );
  AOI21_X1 U7651 ( .B1(n14719), .B2(n14718), .A(n9180), .ZN(n12130) );
  AND2_X1 U7652 ( .A1(n14985), .A2(n14311), .ZN(n9180) );
  NAND2_X1 U7653 ( .A1(n8720), .A2(n8719), .ZN(n14998) );
  NAND2_X1 U7654 ( .A1(n9006), .A2(n9005), .ZN(n15057) );
  NAND2_X1 U7655 ( .A1(n9284), .A2(n11201), .ZN(n15315) );
  OAI211_X1 U7656 ( .C1(n11998), .C2(P1_B_REG_SCAN_IN), .A(n9311), .B(n9310), 
        .ZN(n10278) );
  INV_X1 U7657 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8715) );
  INV_X1 U7658 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U7659 ( .A1(n10607), .A2(n10606), .ZN(n10690) );
  AND2_X1 U7660 ( .A1(n10604), .A2(n10605), .ZN(n10607) );
  NAND2_X1 U7661 ( .A1(n6749), .A2(n6748), .ZN(n6747) );
  NAND2_X1 U7662 ( .A1(n7202), .A2(n9428), .ZN(n12186) );
  NAND2_X1 U7663 ( .A1(n7203), .A2(n12784), .ZN(n7202) );
  NOR2_X1 U7664 ( .A1(n12186), .A2(n15509), .ZN(n7754) );
  OR3_X1 U7665 ( .A1(n11997), .A2(n11949), .A3(n13918), .ZN(n10093) );
  OAI211_X1 U7666 ( .C1(n13362), .C2(n10100), .A(n13361), .B(n6609), .ZN(
        n13359) );
  NAND2_X1 U7667 ( .A1(n13362), .A2(n10100), .ZN(n6609) );
  OAI21_X1 U7668 ( .B1(n10256), .B2(n14463), .A(n8899), .ZN(n7374) );
  OAI21_X1 U7669 ( .B1(n6715), .B2(n9136), .A(n9162), .ZN(n14568) );
  NAND2_X1 U7670 ( .A1(n14586), .A2(n10158), .ZN(n7143) );
  OR2_X1 U7671 ( .A1(n14586), .A2(n10158), .ZN(n7144) );
  XNOR2_X1 U7672 ( .A(n6886), .B(n15181), .ZN(n15183) );
  NAND2_X1 U7673 ( .A1(n7708), .A2(n13127), .ZN(n7707) );
  NAND2_X1 U7674 ( .A1(n7084), .A2(n7083), .ZN(n13124) );
  OR2_X1 U7675 ( .A1(n7625), .A2(n14349), .ZN(n7623) );
  NAND2_X1 U7676 ( .A1(n7625), .A2(n14349), .ZN(n7624) );
  INV_X1 U7677 ( .A(n14351), .ZN(n7397) );
  INV_X1 U7678 ( .A(n8452), .ZN(n7285) );
  INV_X1 U7679 ( .A(n8451), .ZN(n7280) );
  AND2_X1 U7680 ( .A1(n8447), .A2(n10833), .ZN(n7287) );
  NOR2_X1 U7681 ( .A1(n8452), .A2(n7283), .ZN(n7282) );
  OAI21_X1 U7682 ( .B1(n7294), .B2(n8476), .A(n6492), .ZN(n7292) );
  AOI21_X1 U7683 ( .B1(n6433), .B2(n8472), .A(n7295), .ZN(n7294) );
  INV_X1 U7684 ( .A(n8474), .ZN(n7295) );
  OR2_X1 U7685 ( .A1(n13151), .A2(n13150), .ZN(n6763) );
  OR2_X1 U7686 ( .A1(n14393), .A2(n7119), .ZN(n7118) );
  INV_X1 U7687 ( .A(n14392), .ZN(n7121) );
  NOR2_X1 U7688 ( .A1(n7403), .A2(n7404), .ZN(n7402) );
  OAI21_X1 U7689 ( .B1(n14416), .B2(n14415), .A(n14414), .ZN(n14418) );
  NAND2_X1 U7690 ( .A1(n7311), .A2(n7309), .ZN(n7308) );
  NOR2_X1 U7691 ( .A1(n12702), .A2(n7310), .ZN(n7309) );
  OAI21_X1 U7692 ( .B1(n8503), .B2(n12739), .A(n8502), .ZN(n7311) );
  INV_X1 U7693 ( .A(n8504), .ZN(n7310) );
  NAND2_X1 U7694 ( .A1(n6597), .A2(n6596), .ZN(n14429) );
  NAND2_X1 U7695 ( .A1(n14424), .A2(n14426), .ZN(n6596) );
  NAND2_X1 U7696 ( .A1(n7389), .A2(n6598), .ZN(n6597) );
  AND2_X1 U7697 ( .A1(n14306), .A2(n14305), .ZN(n14309) );
  INV_X1 U7698 ( .A(n8669), .ZN(n7423) );
  NAND2_X1 U7699 ( .A1(n12304), .A2(n12694), .ZN(n7647) );
  NAND2_X1 U7700 ( .A1(n7314), .A2(n12658), .ZN(n7313) );
  NAND2_X1 U7701 ( .A1(n7316), .A2(n7315), .ZN(n7314) );
  OR2_X1 U7702 ( .A1(n8518), .A2(n10126), .ZN(n7315) );
  NAND2_X1 U7703 ( .A1(n6824), .A2(n9385), .ZN(n6823) );
  NAND2_X1 U7704 ( .A1(n8539), .A2(n8538), .ZN(n6824) );
  NOR2_X1 U7705 ( .A1(n6741), .A2(n12541), .ZN(n6738) );
  AND2_X1 U7706 ( .A1(n6584), .A2(n6697), .ZN(n6696) );
  INV_X1 U7707 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n6697) );
  AOI21_X1 U7708 ( .B1(n7230), .B2(n7228), .A(n6523), .ZN(n7227) );
  INV_X1 U7709 ( .A(n9349), .ZN(n7228) );
  INV_X1 U7710 ( .A(n9351), .ZN(n7821) );
  INV_X1 U7711 ( .A(n13190), .ZN(n6771) );
  NAND2_X1 U7712 ( .A1(n13184), .A2(n7720), .ZN(n7719) );
  NOR2_X1 U7713 ( .A1(n13608), .A2(n6721), .ZN(n6720) );
  OR2_X1 U7714 ( .A1(n13626), .A2(n6457), .ZN(n6721) );
  NOR2_X1 U7715 ( .A1(n13044), .A2(n6692), .ZN(n6691) );
  AOI21_X1 U7716 ( .B1(n6802), .B2(n6458), .A(n6801), .ZN(n6800) );
  NAND2_X1 U7717 ( .A1(n13970), .A2(n14191), .ZN(n6801) );
  AND3_X1 U7718 ( .A1(n7412), .A2(n14512), .A3(n14513), .ZN(n14505) );
  INV_X1 U7719 ( .A(n8691), .ZN(n6853) );
  INV_X1 U7720 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9003) );
  OR2_X1 U7721 ( .A1(n7640), .A2(n7636), .ZN(n7635) );
  INV_X1 U7722 ( .A(n7647), .ZN(n7636) );
  AND2_X1 U7723 ( .A1(n12409), .A2(n7641), .ZN(n7640) );
  NAND2_X1 U7724 ( .A1(n7642), .A2(n7645), .ZN(n7641) );
  NAND2_X1 U7725 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  AND2_X1 U7726 ( .A1(n12389), .A2(n7329), .ZN(n6908) );
  INV_X1 U7727 ( .A(n7637), .ZN(n6909) );
  NAND2_X1 U7728 ( .A1(n7647), .A2(n7642), .ZN(n7637) );
  NAND2_X1 U7729 ( .A1(n8546), .A2(n9385), .ZN(n7542) );
  NAND2_X1 U7730 ( .A1(n11480), .A2(n11529), .ZN(n6943) );
  NAND3_X1 U7731 ( .A1(n6939), .A2(n6938), .A3(n6569), .ZN(n7663) );
  NAND2_X1 U7732 ( .A1(n6753), .A2(n6751), .ZN(n12497) );
  OR2_X1 U7733 ( .A1(n6573), .A2(n6752), .ZN(n6751) );
  NAND2_X1 U7734 ( .A1(n12000), .A2(n6754), .ZN(n6753) );
  INV_X1 U7735 ( .A(n6760), .ZN(n6752) );
  INV_X1 U7736 ( .A(n6563), .ZN(n7250) );
  NAND2_X1 U7737 ( .A1(n7255), .A2(n7253), .ZN(n7252) );
  INV_X1 U7738 ( .A(n12592), .ZN(n6732) );
  NOR2_X1 U7739 ( .A1(n6474), .A2(n8538), .ZN(n7745) );
  AND2_X1 U7740 ( .A1(n12666), .A2(n7232), .ZN(n7230) );
  INV_X1 U7741 ( .A(n8018), .ZN(n6705) );
  INV_X1 U7742 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7166) );
  AND2_X1 U7743 ( .A1(n7224), .A2(n7223), .ZN(n9334) );
  NAND2_X1 U7744 ( .A1(n9333), .A2(n10830), .ZN(n7224) );
  OR2_X1 U7745 ( .A1(n12461), .A2(n15476), .ZN(n8428) );
  NOR2_X1 U7746 ( .A1(n7837), .A2(n7833), .ZN(n7832) );
  INV_X1 U7747 ( .A(n7873), .ZN(n7833) );
  INV_X1 U7748 ( .A(n7838), .ZN(n7837) );
  NAND2_X1 U7749 ( .A1(n8536), .A2(n6445), .ZN(n7838) );
  NAND2_X1 U7750 ( .A1(n7870), .A2(n7824), .ZN(n7823) );
  INV_X1 U7751 ( .A(n7879), .ZN(n7824) );
  NAND2_X1 U7752 ( .A1(n7227), .A2(n7229), .ZN(n7226) );
  INV_X1 U7753 ( .A(n7230), .ZN(n7229) );
  NOR2_X1 U7754 ( .A1(n7848), .A2(n7847), .ZN(n7846) );
  NOR2_X1 U7755 ( .A1(n12778), .A2(n7175), .ZN(n7174) );
  INV_X1 U7756 ( .A(n8124), .ZN(n7175) );
  INV_X1 U7757 ( .A(n8125), .ZN(n7178) );
  AND2_X1 U7758 ( .A1(n7757), .A2(n7184), .ZN(n7183) );
  NAND2_X1 U7759 ( .A1(n7185), .A2(n8050), .ZN(n7184) );
  NOR2_X1 U7760 ( .A1(n7760), .A2(n7758), .ZN(n7757) );
  INV_X1 U7761 ( .A(n8459), .ZN(n7185) );
  INV_X1 U7762 ( .A(n8050), .ZN(n7186) );
  AOI21_X1 U7763 ( .B1(n6842), .B2(n8328), .A(n6588), .ZN(n6841) );
  NAND2_X1 U7764 ( .A1(n6842), .A2(n6839), .ZN(n6838) );
  INV_X1 U7765 ( .A(n8316), .ZN(n6839) );
  NOR2_X1 U7766 ( .A1(n7579), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7578) );
  NOR2_X1 U7767 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8590) );
  NOR2_X1 U7768 ( .A1(n8593), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n7321) );
  INV_X1 U7769 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8588) );
  INV_X1 U7770 ( .A(n8180), .ZN(n7563) );
  AOI21_X1 U7771 ( .B1(n7583), .B2(n7585), .A(n7582), .ZN(n7581) );
  INV_X1 U7772 ( .A(n8106), .ZN(n7582) );
  INV_X1 U7773 ( .A(n7588), .ZN(n7583) );
  NOR2_X1 U7774 ( .A1(n7584), .A2(n6851), .ZN(n6850) );
  INV_X1 U7775 ( .A(n8068), .ZN(n6851) );
  INV_X1 U7776 ( .A(n7585), .ZN(n7584) );
  INV_X1 U7777 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8132) );
  NOR2_X1 U7778 ( .A1(n8090), .A2(n7589), .ZN(n7588) );
  AND2_X1 U7779 ( .A1(n10423), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8090) );
  INV_X1 U7780 ( .A(n8070), .ZN(n7589) );
  AND2_X1 U7781 ( .A1(n6547), .A2(n6845), .ZN(n6844) );
  NAND2_X1 U7782 ( .A1(n6848), .A2(n7549), .ZN(n6845) );
  INV_X1 U7783 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8011) );
  INV_X1 U7784 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6662) );
  INV_X1 U7785 ( .A(n9738), .ZN(n9471) );
  OAI21_X1 U7786 ( .B1(n6997), .B2(n6996), .A(n11392), .ZN(n6995) );
  NAND2_X1 U7787 ( .A1(n11391), .A2(n11390), .ZN(n6998) );
  INV_X1 U7788 ( .A(n7605), .ZN(n6980) );
  NAND2_X1 U7789 ( .A1(n6979), .A2(n7605), .ZN(n6978) );
  INV_X1 U7790 ( .A(n12083), .ZN(n6979) );
  INV_X1 U7791 ( .A(n9637), .ZN(n6686) );
  NAND2_X1 U7792 ( .A1(n11603), .A2(n11602), .ZN(n11604) );
  OR2_X1 U7793 ( .A1(n13413), .A2(n13422), .ZN(n13425) );
  AND2_X1 U7794 ( .A1(n7498), .A2(n7496), .ZN(n7495) );
  INV_X1 U7795 ( .A(n7497), .ZN(n7496) );
  OR2_X1 U7796 ( .A1(n9810), .A2(n15516), .ZN(n9490) );
  NAND2_X1 U7797 ( .A1(n13551), .A2(n9855), .ZN(n7494) );
  AND2_X1 U7798 ( .A1(n13526), .A2(n7506), .ZN(n7505) );
  NAND2_X1 U7799 ( .A1(n9856), .A2(n9855), .ZN(n7506) );
  NOR2_X1 U7800 ( .A1(n9850), .A2(n7515), .ZN(n7514) );
  INV_X1 U7801 ( .A(n9849), .ZN(n7515) );
  NAND2_X1 U7802 ( .A1(n9698), .A2(n7345), .ZN(n7344) );
  NOR2_X1 U7803 ( .A1(n7344), .A2(n7341), .ZN(n7340) );
  INV_X1 U7804 ( .A(n9683), .ZN(n7341) );
  INV_X1 U7805 ( .A(n9842), .ZN(n7518) );
  INV_X1 U7806 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U7807 ( .A1(n6906), .A2(n11051), .ZN(n13108) );
  INV_X1 U7808 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U7809 ( .A1(n7700), .A2(n9461), .ZN(n6675) );
  INV_X1 U7810 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9884) );
  INV_X1 U7811 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9586) );
  NOR2_X2 U7812 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9499) );
  OR2_X1 U7813 ( .A1(n14479), .A2(n10282), .ZN(n14011) );
  NAND2_X1 U7814 ( .A1(n10825), .A2(n6409), .ZN(n7358) );
  NAND2_X1 U7815 ( .A1(n14505), .A2(n14504), .ZN(n14491) );
  AND2_X1 U7816 ( .A1(n8857), .A2(n7788), .ZN(n9040) );
  NOR2_X1 U7817 ( .A1(n7027), .A2(n7031), .ZN(n7026) );
  INV_X1 U7818 ( .A(n7781), .ZN(n7780) );
  OAI21_X1 U7819 ( .B1(n7784), .B2(n7783), .A(n7782), .ZN(n7781) );
  INV_X1 U7820 ( .A(n7786), .ZN(n7783) );
  OR2_X1 U7821 ( .A1(n9129), .A2(n7114), .ZN(n7028) );
  NAND2_X1 U7822 ( .A1(n8612), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9089) );
  INV_X1 U7823 ( .A(n9045), .ZN(n8612) );
  OR2_X1 U7824 ( .A1(n15045), .A2(n15054), .ZN(n14405) );
  OR2_X1 U7825 ( .A1(n9027), .A2(n9007), .ZN(n9045) );
  AND2_X1 U7826 ( .A1(n14932), .A2(n7446), .ZN(n7443) );
  NAND2_X1 U7827 ( .A1(n9256), .A2(n15074), .ZN(n14395) );
  NOR2_X1 U7829 ( .A1(n15074), .A2(n7357), .ZN(n7356) );
  INV_X1 U7830 ( .A(n8989), .ZN(n7357) );
  INV_X1 U7831 ( .A(n7791), .ZN(n7045) );
  AOI21_X1 U7832 ( .B1(n9253), .B2(n7792), .A(n6500), .ZN(n7791) );
  INV_X1 U7833 ( .A(n9252), .ZN(n7792) );
  INV_X1 U7834 ( .A(n9249), .ZN(n7046) );
  AND2_X1 U7835 ( .A1(n9242), .A2(n15303), .ZN(n7438) );
  INV_X1 U7836 ( .A(n14326), .ZN(n7763) );
  INV_X1 U7837 ( .A(n14934), .ZN(n14672) );
  OR2_X1 U7838 ( .A1(n14579), .A2(n15275), .ZN(n14327) );
  NAND2_X1 U7839 ( .A1(n8628), .A2(n7815), .ZN(n7814) );
  INV_X1 U7840 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U7841 ( .A1(n9166), .A2(n9165), .ZN(n9184) );
  OAI21_X1 U7842 ( .B1(n9164), .B2(n12942), .A(n9163), .ZN(n9166) );
  NAND2_X1 U7843 ( .A1(n6869), .A2(n6867), .ZN(n9146) );
  AOI21_X1 U7844 ( .B1(n6868), .B2(n6872), .A(n6511), .ZN(n6867) );
  NOR2_X1 U7845 ( .A1(n8697), .A2(n8698), .ZN(n7428) );
  AOI21_X1 U7846 ( .B1(n6412), .B2(n8683), .A(n6505), .ZN(n7417) );
  NAND2_X1 U7847 ( .A1(n7097), .A2(n6876), .ZN(n8888) );
  NAND2_X1 U7848 ( .A1(n7434), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7097) );
  OAI21_X1 U7849 ( .B1(n7369), .B2(SI_7_), .A(n8664), .ZN(n7368) );
  NAND2_X1 U7850 ( .A1(n8827), .A2(n8663), .ZN(n8836) );
  NAND2_X1 U7851 ( .A1(n7426), .A2(n8658), .ZN(n8803) );
  AOI21_X1 U7852 ( .B1(n8657), .B2(n8784), .A(n8656), .ZN(n8658) );
  OR2_X1 U7853 ( .A1(n9941), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n9942) );
  OR2_X1 U7854 ( .A1(n9989), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n9990) );
  AND2_X1 U7855 ( .A1(n6968), .A2(n6967), .ZN(n10491) );
  NAND2_X1 U7856 ( .A1(n10480), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6967) );
  INV_X1 U7857 ( .A(n10478), .ZN(n6969) );
  INV_X1 U7858 ( .A(n6964), .ZN(n6963) );
  OAI21_X1 U7859 ( .B1(n11558), .B2(n6965), .A(n11712), .ZN(n6964) );
  INV_X1 U7860 ( .A(n11560), .ZN(n6965) );
  INV_X1 U7861 ( .A(n6971), .ZN(n15168) );
  OAI21_X1 U7862 ( .B1(n15163), .B2(n6591), .A(n15164), .ZN(n6971) );
  INV_X1 U7863 ( .A(n7634), .ZN(n7633) );
  OAI21_X1 U7864 ( .B1(n12438), .B2(n12319), .A(n12322), .ZN(n7634) );
  OR2_X1 U7865 ( .A1(n12397), .A2(n12309), .ZN(n7134) );
  NAND2_X1 U7866 ( .A1(n6624), .A2(n6623), .ZN(n7326) );
  INV_X1 U7867 ( .A(n12334), .ZN(n6623) );
  INV_X1 U7868 ( .A(n12335), .ZN(n6624) );
  INV_X1 U7869 ( .A(n12402), .ZN(n7327) );
  INV_X1 U7870 ( .A(n10695), .ZN(n6625) );
  AOI21_X1 U7871 ( .B1(n11307), .B2(n11191), .A(n6481), .ZN(n7651) );
  NAND2_X1 U7872 ( .A1(n11190), .A2(n11307), .ZN(n6897) );
  NAND2_X1 U7873 ( .A1(n12596), .A2(n11362), .ZN(n10515) );
  NAND2_X1 U7874 ( .A1(n7302), .A2(n7301), .ZN(n7303) );
  AND4_X1 U7875 ( .A1(n8086), .A2(n8085), .A3(n8084), .A4(n8083), .ZN(n11908)
         );
  BUF_X1 U7876 ( .A(n7982), .Z(n8080) );
  OR2_X1 U7877 ( .A1(n8080), .A2(n11405), .ZN(n7965) );
  OR2_X1 U7878 ( .A1(n7960), .A2(n6622), .ZN(n7196) );
  INV_X1 U7879 ( .A(n10321), .ZN(n10204) );
  INV_X1 U7880 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10336) );
  XNOR2_X1 U7881 ( .A(n7238), .B(n10321), .ZN(n10323) );
  NAND2_X1 U7882 ( .A1(n7667), .A2(n7669), .ZN(n7666) );
  NAND2_X1 U7883 ( .A1(n7668), .A2(n6419), .ZN(n6934) );
  NOR2_X1 U7884 ( .A1(n7275), .A2(n7268), .ZN(n7267) );
  INV_X1 U7885 ( .A(n7273), .ZN(n7268) );
  INV_X1 U7886 ( .A(n10880), .ZN(n7265) );
  NAND2_X1 U7887 ( .A1(n7259), .A2(n11471), .ZN(n7258) );
  INV_X1 U7888 ( .A(n7261), .ZN(n7259) );
  NAND2_X1 U7889 ( .A1(n11927), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U7890 ( .A1(n11915), .A2(n11914), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11917), .ZN(n12000) );
  INV_X1 U7891 ( .A(n12543), .ZN(n6741) );
  NAND2_X1 U7892 ( .A1(n12542), .A2(n6743), .ZN(n6740) );
  NOR2_X1 U7893 ( .A1(n12523), .A2(n12522), .ZN(n12532) );
  INV_X1 U7894 ( .A(n7252), .ZN(n7248) );
  AOI21_X1 U7895 ( .B1(n6418), .B2(n7256), .A(n6580), .ZN(n7255) );
  NAND4_X1 U7896 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(
        P3_REG2_REG_17__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U7897 ( .A1(n6953), .A2(n12576), .ZN(n12573) );
  NAND2_X1 U7898 ( .A1(n6954), .A2(n7678), .ZN(n6953) );
  OR2_X1 U7899 ( .A1(n9423), .A2(n9426), .ZN(n7876) );
  NAND2_X1 U7900 ( .A1(n7168), .A2(n8333), .ZN(n8345) );
  INV_X1 U7901 ( .A(n8334), .ZN(n7168) );
  OR2_X1 U7902 ( .A1(n8345), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U7903 ( .A1(n8531), .A2(n8415), .ZN(n7748) );
  NAND2_X1 U7904 ( .A1(n7841), .A2(n9356), .ZN(n12618) );
  OR2_X1 U7905 ( .A1(n12793), .A2(n12357), .ZN(n8339) );
  NAND2_X1 U7906 ( .A1(n12619), .A2(n15479), .ZN(n12622) );
  AND2_X1 U7907 ( .A1(n8521), .A2(n8520), .ZN(n12658) );
  AND2_X1 U7908 ( .A1(n7737), .A2(n7733), .ZN(n7732) );
  NAND2_X1 U7909 ( .A1(n12679), .A2(n9349), .ZN(n7231) );
  NAND2_X1 U7910 ( .A1(n7231), .A2(n7230), .ZN(n12665) );
  INV_X1 U7911 ( .A(n6656), .ZN(n6655) );
  AND2_X1 U7912 ( .A1(n9339), .A2(n8457), .ZN(n11349) );
  AOI21_X1 U7913 ( .B1(n7828), .B2(n7830), .A(n6471), .ZN(n7826) );
  NAND2_X1 U7914 ( .A1(n7999), .A2(n7998), .ZN(n8018) );
  INV_X1 U7915 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n7998) );
  INV_X1 U7916 ( .A(n8000), .ZN(n7999) );
  OR2_X1 U7917 ( .A1(n12460), .A2(n11406), .ZN(n11082) );
  NAND2_X1 U7918 ( .A1(n10626), .A2(n10625), .ZN(n11288) );
  NAND2_X1 U7919 ( .A1(n12648), .A2(n12647), .ZN(n12646) );
  OR2_X1 U7920 ( .A1(n8415), .A2(n8530), .ZN(n12633) );
  NAND2_X1 U7921 ( .A1(n8304), .A2(n8303), .ZN(n12313) );
  NAND2_X1 U7922 ( .A1(n12691), .A2(n6649), .ZN(n12679) );
  NAND2_X1 U7923 ( .A1(n6650), .A2(n12681), .ZN(n6649) );
  NAND2_X1 U7924 ( .A1(n7738), .A2(n8509), .ZN(n7737) );
  NAND2_X1 U7925 ( .A1(n7728), .A2(n8510), .ZN(n7738) );
  NAND2_X1 U7926 ( .A1(n12702), .A2(n7740), .ZN(n7728) );
  OR2_X1 U7927 ( .A1(n8508), .A2(n8513), .ZN(n12676) );
  AND2_X1 U7928 ( .A1(n6651), .A2(n6534), .ZN(n12693) );
  AND2_X1 U7929 ( .A1(n8211), .A2(n8210), .ZN(n12749) );
  AND2_X1 U7930 ( .A1(n8241), .A2(n8240), .ZN(n12718) );
  AND2_X1 U7931 ( .A1(n8486), .A2(n8491), .ZN(n12767) );
  NAND2_X1 U7932 ( .A1(n7853), .A2(n7859), .ZN(n7852) );
  NAND2_X1 U7933 ( .A1(n9342), .A2(n6478), .ZN(n7851) );
  AOI21_X1 U7934 ( .B1(n11951), .B2(n7726), .A(n7725), .ZN(n7724) );
  INV_X1 U7935 ( .A(n8470), .ZN(n7726) );
  NAND2_X1 U7936 ( .A1(n9342), .A2(n7857), .ZN(n7856) );
  OR2_X1 U7937 ( .A1(n11787), .A2(n11955), .ZN(n8470) );
  AND2_X1 U7938 ( .A1(n8474), .A2(n8475), .ZN(n11951) );
  NAND2_X1 U7939 ( .A1(n11364), .A2(n9340), .ZN(n9342) );
  NAND2_X1 U7940 ( .A1(n8088), .A2(n8087), .ZN(n11598) );
  INV_X1 U7941 ( .A(n15469), .ZN(n15479) );
  NAND2_X1 U7942 ( .A1(n7574), .A2(n8378), .ZN(n7573) );
  NAND2_X1 U7943 ( .A1(n7570), .A2(n8380), .ZN(n7569) );
  INV_X1 U7944 ( .A(n8378), .ZN(n7570) );
  NOR2_X1 U7945 ( .A1(n7572), .A2(n7574), .ZN(n7571) );
  INV_X1 U7946 ( .A(n7575), .ZN(n7572) );
  NOR2_X1 U7947 ( .A1(n8368), .A2(n7576), .ZN(n7575) );
  INV_X1 U7948 ( .A(n8365), .ZN(n7576) );
  NAND2_X1 U7949 ( .A1(n8288), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8300) );
  NOR2_X1 U7950 ( .A1(n8273), .A2(n7556), .ZN(n7555) );
  INV_X1 U7951 ( .A(n8262), .ZN(n7556) );
  AOI21_X1 U7952 ( .B1(n6834), .B2(n6566), .A(n6833), .ZN(n6832) );
  OR2_X1 U7953 ( .A1(n8397), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8416) );
  INV_X1 U7954 ( .A(n6835), .ZN(n6834) );
  OAI21_X1 U7955 ( .B1(n7558), .B2(n6566), .A(n8213), .ZN(n6835) );
  INV_X1 U7956 ( .A(n8397), .ZN(n7655) );
  NOR2_X1 U7957 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7654) );
  AOI21_X1 U7958 ( .B1(n7561), .B2(n7563), .A(n7559), .ZN(n7558) );
  INV_X1 U7959 ( .A(n8198), .ZN(n7559) );
  AND2_X1 U7960 ( .A1(n8180), .A2(n8167), .ZN(n8168) );
  NAND2_X1 U7961 ( .A1(n8169), .A2(n8168), .ZN(n8181) );
  AND2_X1 U7962 ( .A1(n8109), .A2(n8126), .ZN(n8110) );
  NAND2_X1 U7963 ( .A1(n8071), .A2(n7588), .ZN(n7587) );
  NOR2_X1 U7964 ( .A1(n8093), .A2(n7586), .ZN(n7585) );
  INV_X1 U7965 ( .A(n8089), .ZN(n7586) );
  INV_X1 U7966 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8076) );
  INV_X1 U7967 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8039) );
  XNOR2_X1 U7968 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8025) );
  NAND2_X1 U7969 ( .A1(n8009), .A2(n8008), .ZN(n8026) );
  NAND2_X1 U7970 ( .A1(n7991), .A2(n6847), .ZN(n8009) );
  XNOR2_X1 U7971 ( .A(n7993), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10640) );
  XNOR2_X1 U7972 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7987) );
  INV_X1 U7973 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7953) );
  AND2_X1 U7974 ( .A1(n7924), .A2(n7922), .ZN(n7545) );
  XNOR2_X1 U7975 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7972) );
  NOR2_X1 U7976 ( .A1(n11220), .A2(n11211), .ZN(n6997) );
  NOR2_X1 U7977 ( .A1(n12210), .A2(n12114), .ZN(n7605) );
  OR2_X1 U7978 ( .A1(n12963), .A2(n12964), .ZN(n13007) );
  NAND2_X1 U7979 ( .A1(n11397), .A2(n11396), .ZN(n11660) );
  INV_X1 U7980 ( .A(n13344), .ZN(n13695) );
  NAND2_X1 U7981 ( .A1(n7160), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9810) );
  INV_X1 U7982 ( .A(n9808), .ZN(n7160) );
  INV_X1 U7983 ( .A(n13642), .ZN(n13294) );
  NAND2_X1 U7984 ( .A1(n9472), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9797) );
  INV_X1 U7985 ( .A(n9788), .ZN(n9472) );
  NAND2_X1 U7986 ( .A1(n13040), .A2(n13041), .ZN(n13039) );
  NOR2_X1 U7987 ( .A1(n7603), .A2(n7006), .ZN(n7005) );
  INV_X1 U7988 ( .A(n12235), .ZN(n7006) );
  INV_X1 U7989 ( .A(n7604), .ZN(n7603) );
  AOI21_X1 U7990 ( .B1(n7604), .B2(n7602), .A(n6475), .ZN(n7601) );
  INV_X1 U7991 ( .A(n13041), .ZN(n7602) );
  AND2_X1 U7992 ( .A1(n7594), .A2(n7592), .ZN(n7591) );
  INV_X1 U7993 ( .A(n12984), .ZN(n7592) );
  NAND2_X1 U7994 ( .A1(n10801), .A2(n12272), .ZN(n10802) );
  INV_X1 U7995 ( .A(n6398), .ZN(n13298) );
  AND2_X1 U7996 ( .A1(n13463), .A2(n9864), .ZN(n12276) );
  INV_X1 U7997 ( .A(n15361), .ZN(n6632) );
  AOI21_X1 U7998 ( .B1(n15361), .B2(n6631), .A(n6460), .ZN(n6630) );
  INV_X1 U7999 ( .A(n10084), .ZN(n6631) );
  NAND2_X1 U8000 ( .A1(n15386), .A2(n10371), .ZN(n10373) );
  OR2_X1 U8001 ( .A1(n10373), .A2(n10372), .ZN(n10593) );
  NAND2_X1 U8002 ( .A1(n15380), .A2(n15379), .ZN(n6642) );
  OR2_X1 U8003 ( .A1(n11144), .A2(n11143), .ZN(n11603) );
  XNOR2_X1 U8004 ( .A(n11604), .B(n11609), .ZN(n11678) );
  XNOR2_X1 U8005 ( .A(n13465), .B(n13336), .ZN(n13755) );
  NAND2_X1 U8006 ( .A1(n13453), .A2(n13290), .ZN(n13475) );
  OR2_X1 U8007 ( .A1(n9863), .A2(n9862), .ZN(n13463) );
  AND2_X1 U8008 ( .A1(n9858), .A2(n13450), .ZN(n9861) );
  OR2_X1 U8009 ( .A1(n13289), .A2(n13678), .ZN(n9872) );
  AOI21_X1 U8010 ( .B1(n7338), .B2(n7336), .A(n6501), .ZN(n7335) );
  INV_X1 U8011 ( .A(n7339), .ZN(n7336) );
  INV_X1 U8012 ( .A(n7338), .ZN(n7337) );
  NAND2_X1 U8013 ( .A1(n7494), .A2(n7505), .ZN(n7511) );
  OR2_X1 U8014 ( .A1(n13551), .A2(n9856), .ZN(n7504) );
  INV_X1 U8015 ( .A(n7159), .ZN(n9777) );
  NOR2_X1 U8016 ( .A1(n13630), .A2(n13809), .ZN(n13615) );
  NAND2_X1 U8017 ( .A1(n13645), .A2(n6457), .ZN(n13644) );
  NAND2_X1 U8018 ( .A1(n6451), .A2(n9683), .ZN(n7342) );
  AND2_X1 U8019 ( .A1(n9643), .A2(n6413), .ZN(n7528) );
  NAND2_X1 U8020 ( .A1(n7523), .A2(n12043), .ZN(n7526) );
  NAND2_X1 U8021 ( .A1(n9644), .A2(n9643), .ZN(n7523) );
  NAND2_X1 U8022 ( .A1(n6682), .A2(n6494), .ZN(n9630) );
  INV_X1 U8023 ( .A(n6448), .ZN(n7490) );
  NAND2_X1 U8024 ( .A1(n9828), .A2(n13305), .ZN(n11244) );
  NAND2_X1 U8025 ( .A1(n11058), .A2(n11241), .ZN(n9828) );
  NAND2_X1 U8026 ( .A1(n10746), .A2(n9537), .ZN(n10993) );
  NAND2_X1 U8027 ( .A1(n7350), .A2(n10803), .ZN(n10705) );
  INV_X1 U8028 ( .A(n13108), .ZN(n6773) );
  NAND2_X1 U8029 ( .A1(n9652), .A2(n9651), .ZN(n13846) );
  NAND2_X1 U8030 ( .A1(n10422), .A2(n13262), .ZN(n9635) );
  OR2_X1 U8031 ( .A1(n9536), .A2(n9968), .ZN(n7701) );
  AND2_X1 U8032 ( .A1(n10712), .A2(n10711), .ZN(n10974) );
  NAND2_X1 U8033 ( .A1(n13666), .A2(n9455), .ZN(n15422) );
  INV_X1 U8034 ( .A(n9881), .ZN(n9882) );
  XNOR2_X1 U8035 ( .A(n9911), .B(n15527), .ZN(n11491) );
  OAI21_X1 U8036 ( .B1(n9880), .B2(n6417), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9819) );
  INV_X1 U8037 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9446) );
  AND2_X1 U8038 ( .A1(n9533), .A2(n9543), .ZN(n13389) );
  INV_X1 U8039 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6646) );
  INV_X1 U8040 ( .A(n9499), .ZN(n9515) );
  AOI21_X1 U8041 ( .B1(n11815), .B2(n11814), .A(n7860), .ZN(n11939) );
  OAI211_X1 U8042 ( .C1(n12177), .C2(n13932), .A(n13957), .B(n6786), .ZN(n6785) );
  OR2_X1 U8043 ( .A1(n12176), .A2(n13932), .ZN(n6786) );
  AND2_X1 U8044 ( .A1(n7456), .A2(n6792), .ZN(n6791) );
  NAND2_X1 U8045 ( .A1(n7458), .A2(n13994), .ZN(n6792) );
  INV_X1 U8046 ( .A(n14245), .ZN(n7457) );
  AOI21_X1 U8047 ( .B1(n14270), .B2(n13980), .A(n6502), .ZN(n7481) );
  NAND2_X1 U8048 ( .A1(n6798), .A2(n6795), .ZN(n7480) );
  NOR2_X1 U8049 ( .A1(n6796), .A2(n7482), .ZN(n6795) );
  INV_X1 U8050 ( .A(n14270), .ZN(n7482) );
  NAND2_X1 U8051 ( .A1(n14226), .A2(n14225), .ZN(n7462) );
  INV_X1 U8052 ( .A(n14568), .ZN(n14161) );
  INV_X1 U8053 ( .A(n6707), .ZN(n9133) );
  NAND2_X1 U8054 ( .A1(n6707), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9135) );
  INV_X1 U8055 ( .A(n14479), .ZN(n9279) );
  NAND2_X1 U8056 ( .A1(n9080), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9106) );
  OR2_X1 U8057 ( .A1(n9106), .A2(n14254), .ZN(n9123) );
  INV_X1 U8058 ( .A(n6796), .ZN(n6794) );
  NAND2_X1 U8059 ( .A1(n11443), .A2(n11444), .ZN(n6811) );
  NAND2_X1 U8060 ( .A1(n6808), .A2(n6810), .ZN(n6807) );
  INV_X1 U8061 ( .A(n6814), .ZN(n6810) );
  AND2_X1 U8062 ( .A1(n6816), .A2(n14178), .ZN(n6815) );
  OR2_X1 U8063 ( .A1(n11443), .A2(n14177), .ZN(n6816) );
  AND2_X1 U8064 ( .A1(n6814), .A2(n11444), .ZN(n6813) );
  NAND2_X1 U8065 ( .A1(n7394), .A2(n7617), .ZN(n7616) );
  AND4_X1 U8066 ( .A1(n8870), .A2(n8869), .A3(n8868), .A4(n8867), .ZN(n11933)
         );
  INV_X1 U8067 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14602) );
  OR2_X1 U8068 ( .A1(n8859), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U8069 ( .A1(n11793), .A2(n7073), .ZN(n11794) );
  OR2_X1 U8070 ( .A1(n11801), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U8071 ( .A1(n14452), .A2(n14451), .ZN(n14681) );
  NAND2_X1 U8072 ( .A1(n9207), .A2(n9206), .ZN(n14486) );
  AOI21_X1 U8073 ( .B1(n7806), .B2(n7782), .A(n12136), .ZN(n7805) );
  NAND2_X1 U8074 ( .A1(n14998), .A2(n14042), .ZN(n7786) );
  AND2_X1 U8075 ( .A1(n9267), .A2(n14542), .ZN(n7809) );
  AND2_X1 U8076 ( .A1(n14856), .A2(n6529), .ZN(n14799) );
  AND2_X1 U8077 ( .A1(n7053), .A2(n9262), .ZN(n7052) );
  AND2_X1 U8078 ( .A1(n14880), .A2(n14855), .ZN(n14856) );
  INV_X1 U8079 ( .A(n7016), .ZN(n7015) );
  AND2_X1 U8080 ( .A1(n6525), .A2(n9260), .ZN(n7058) );
  NOR2_X2 U8081 ( .A1(n14892), .A2(n15057), .ZN(n14880) );
  NAND2_X1 U8082 ( .A1(n14929), .A2(n14390), .ZN(n14911) );
  NAND2_X1 U8083 ( .A1(n8937), .A2(n8936), .ZN(n14972) );
  NAND2_X1 U8084 ( .A1(n11756), .A2(n11757), .ZN(n9247) );
  NAND2_X1 U8085 ( .A1(n7363), .A2(n8908), .ZN(n7766) );
  AND2_X1 U8086 ( .A1(n8909), .A2(n8887), .ZN(n7363) );
  INV_X1 U8087 ( .A(n11757), .ZN(n14538) );
  NAND2_X1 U8088 ( .A1(n14348), .A2(n15313), .ZN(n7777) );
  NOR2_X1 U8089 ( .A1(n6489), .A2(n7011), .ZN(n7010) );
  INV_X1 U8090 ( .A(n8815), .ZN(n7011) );
  NAND2_X1 U8091 ( .A1(n7037), .A2(n9239), .ZN(n15230) );
  NAND2_X1 U8092 ( .A1(n11337), .A2(n14530), .ZN(n7037) );
  NAND2_X1 U8093 ( .A1(n11200), .A2(n11199), .ZN(n14693) );
  NAND2_X1 U8094 ( .A1(n14527), .A2(n14321), .ZN(n10786) );
  INV_X1 U8095 ( .A(n14581), .ZN(n7013) );
  INV_X1 U8096 ( .A(n14984), .ZN(n14987) );
  INV_X1 U8097 ( .A(n15016), .ZN(n7068) );
  NAND2_X1 U8098 ( .A1(n9519), .A2(n6408), .ZN(n7407) );
  OAI22_X1 U8099 ( .A1(n14466), .A2(n9969), .B1(n8755), .B2(n14605), .ZN(n7406) );
  INV_X1 U8100 ( .A(n15310), .ZN(n15090) );
  AOI21_X1 U8101 ( .B1(n12197), .B2(n12196), .A(n12195), .ZN(n12200) );
  INV_X1 U8102 ( .A(n7814), .ZN(n7812) );
  XNOR2_X1 U8103 ( .A(n9302), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9311) );
  AND2_X1 U8104 ( .A1(n9219), .A2(n9220), .ZN(n7628) );
  INV_X1 U8105 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9220) );
  INV_X1 U8106 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9059) );
  XNOR2_X1 U8107 ( .A(n6727), .B(n9057), .ZN(n9734) );
  OAI21_X1 U8108 ( .B1(n9052), .B2(n8690), .A(n9054), .ZN(n6727) );
  NAND2_X1 U8109 ( .A1(n6854), .A2(n7414), .ZN(n9001) );
  NAND2_X1 U8110 ( .A1(n8964), .A2(n7413), .ZN(n6854) );
  NAND2_X1 U8111 ( .A1(n8897), .A2(n8896), .ZN(n8987) );
  NAND2_X1 U8112 ( .A1(n8836), .A2(n8835), .ZN(n8838) );
  NAND2_X1 U8113 ( .A1(n6616), .A2(n6615), .ZN(n6614) );
  INV_X1 U8114 ( .A(n8665), .ZN(n6616) );
  NAND2_X1 U8115 ( .A1(n10499), .A2(n10498), .ZN(n10931) );
  OAI22_X1 U8116 ( .A1(n15158), .A2(n6894), .B1(n6893), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n10940) );
  INV_X1 U8117 ( .A(n15156), .ZN(n6893) );
  NOR2_X1 U8118 ( .A1(n15156), .A2(n7095), .ZN(n6894) );
  NAND2_X1 U8119 ( .A1(n11553), .A2(n11552), .ZN(n11559) );
  NAND2_X1 U8120 ( .A1(n12093), .A2(n12092), .ZN(n6892) );
  XNOR2_X1 U8121 ( .A(n15168), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n15169) );
  INV_X1 U8122 ( .A(n6966), .ZN(n15192) );
  AND2_X1 U8123 ( .A1(n8326), .A2(n8325), .ZN(n12645) );
  NAND2_X1 U8124 ( .A1(n8276), .A2(n8275), .ZN(n12340) );
  AOI21_X1 U8125 ( .B1(n12426), .B2(n12425), .A(n7868), .ZN(n12344) );
  AND2_X1 U8126 ( .A1(n8098), .A2(n8097), .ZN(n11909) );
  INV_X1 U8127 ( .A(n12668), .ZN(n12644) );
  AND2_X1 U8128 ( .A1(n12295), .A2(n12383), .ZN(n7650) );
  NAND2_X1 U8129 ( .A1(n8188), .A2(n8187), .ZN(n12392) );
  NAND2_X1 U8130 ( .A1(n7652), .A2(n11188), .ZN(n11308) );
  INV_X1 U8131 ( .A(n6621), .ZN(n7652) );
  INV_X1 U8132 ( .A(n7638), .ZN(n12410) );
  AOI21_X1 U8133 ( .B1(n12426), .B2(n7639), .A(n7643), .ZN(n7638) );
  INV_X1 U8134 ( .A(n7645), .ZN(n7639) );
  NAND2_X1 U8135 ( .A1(n10582), .A2(n10583), .ZN(n10606) );
  NAND2_X1 U8136 ( .A1(n10249), .A2(n15460), .ZN(n12414) );
  AND2_X1 U8137 ( .A1(n8313), .A2(n8312), .ZN(n12656) );
  NAND2_X1 U8138 ( .A1(n10609), .A2(n11517), .ZN(n12441) );
  NAND2_X1 U8139 ( .A1(n8271), .A2(n8270), .ZN(n12695) );
  OAI211_X1 U8140 ( .C1(n8372), .C2(n12832), .A(n8178), .B(n8177), .ZN(n12770)
         );
  NAND4_X1 U8141 ( .A1(n8105), .A2(n8104), .A3(n8103), .A4(n8102), .ZN(n12454)
         );
  INV_X1 U8142 ( .A(n11908), .ZN(n11955) );
  INV_X1 U8143 ( .A(n11431), .ZN(n11365) );
  NAND4_X2 U8144 ( .A1(n7915), .A2(n7914), .A3(n7913), .A4(n7912), .ZN(n10836)
         );
  OAI22_X1 U8145 ( .A1(n10322), .A2(n10323), .B1(n10321), .B2(n7238), .ZN(
        n10383) );
  NAND2_X1 U8146 ( .A1(n7658), .A2(n7659), .ZN(n11478) );
  INV_X1 U8147 ( .A(n10877), .ZN(n6746) );
  OAI22_X1 U8148 ( .A1(n11528), .A2(n11568), .B1(n7375), .B2(n11529), .ZN(
        n11915) );
  INV_X1 U8149 ( .A(n7376), .ZN(n7375) );
  NAND2_X1 U8150 ( .A1(n6939), .A2(n6938), .ZN(n11916) );
  NAND2_X1 U8151 ( .A1(n6944), .A2(n6945), .ZN(n12536) );
  INV_X1 U8152 ( .A(n6946), .ZN(n6945) );
  NAND2_X1 U8153 ( .A1(n6949), .A2(n6429), .ZN(n6944) );
  OAI21_X1 U8154 ( .B1(n12493), .B2(n6947), .A(n12531), .ZN(n6946) );
  NAND2_X1 U8155 ( .A1(n7674), .A2(n12590), .ZN(n7672) );
  NAND2_X1 U8156 ( .A1(n6590), .A2(n7675), .ZN(n7674) );
  XNOR2_X1 U8157 ( .A(n7243), .B(n12603), .ZN(n7242) );
  AOI21_X1 U8158 ( .B1(n12574), .B2(n12573), .A(n12572), .ZN(n12589) );
  NOR2_X1 U8159 ( .A1(n7673), .A2(n12566), .ZN(n7671) );
  AND2_X1 U8160 ( .A1(n7675), .A2(n12601), .ZN(n7673) );
  INV_X1 U8161 ( .A(n12606), .ZN(n7245) );
  XNOR2_X1 U8162 ( .A(n9393), .B(n7301), .ZN(n12617) );
  NAND2_X1 U8163 ( .A1(n8344), .A2(n8343), .ZN(n12614) );
  NAND2_X1 U8164 ( .A1(n8264), .A2(n8263), .ZN(n12686) );
  NOR2_X1 U8165 ( .A1(n12739), .A2(n8497), .ZN(n7761) );
  NAND2_X1 U8166 ( .A1(n8204), .A2(n8203), .ZN(n12738) );
  AND2_X1 U8167 ( .A1(n12593), .A2(n11362), .ZN(n15462) );
  INV_X1 U8168 ( .A(n15460), .ZN(n15488) );
  NAND2_X1 U8169 ( .A1(n10248), .A2(n15462), .ZN(n15460) );
  NAND2_X1 U8170 ( .A1(n7756), .A2(n15501), .ZN(n7755) );
  INV_X1 U8171 ( .A(n12186), .ZN(n7753) );
  NAND2_X1 U8172 ( .A1(n15514), .A2(n12829), .ZN(n12821) );
  AND2_X1 U8173 ( .A1(n8384), .A2(n8383), .ZN(n8548) );
  NAND2_X1 U8174 ( .A1(n8354), .A2(n8353), .ZN(n12850) );
  AOI21_X1 U8175 ( .B1(n7754), .B2(n12797), .A(n6440), .ZN(n7751) );
  NOR2_X1 U8176 ( .A1(n6565), .A2(n9361), .ZN(n9362) );
  NAND2_X1 U8177 ( .A1(n8220), .A2(n8219), .ZN(n12893) );
  AND2_X1 U8178 ( .A1(n8137), .A2(n8136), .ZN(n12916) );
  NAND2_X1 U8179 ( .A1(n8116), .A2(n8115), .ZN(n12110) );
  AND2_X1 U8180 ( .A1(n15510), .A2(n12829), .ZN(n12915) );
  OAI21_X1 U8181 ( .B1(n9412), .B2(n10250), .A(n9411), .ZN(n9413) );
  OR2_X1 U8182 ( .A1(n10247), .A2(n9410), .ZN(n9411) );
  NAND2_X1 U8183 ( .A1(n11213), .A2(n6997), .ZN(n6993) );
  INV_X1 U8184 ( .A(n13456), .ZN(n13289) );
  NAND2_X1 U8185 ( .A1(n7135), .A2(n13262), .ZN(n9676) );
  OAI21_X1 U8186 ( .B1(n7600), .B2(n6985), .A(n6981), .ZN(n6987) );
  NAND2_X1 U8187 ( .A1(n6986), .A2(n12265), .ZN(n6985) );
  AOI21_X1 U8188 ( .B1(n6986), .B2(n6983), .A(n6982), .ZN(n6981) );
  INV_X1 U8189 ( .A(n12953), .ZN(n6986) );
  INV_X1 U8190 ( .A(n13341), .ZN(n13581) );
  NAND2_X1 U8191 ( .A1(n9702), .A2(n9701), .ZN(n13180) );
  NAND2_X1 U8192 ( .A1(n9662), .A2(n9661), .ZN(n13839) );
  INV_X1 U8193 ( .A(n13074), .ZN(n13061) );
  NOR2_X1 U8194 ( .A1(n13074), .A2(n13676), .ZN(n13083) );
  NOR2_X1 U8195 ( .A1(n10810), .A2(n10809), .ZN(n10861) );
  OR2_X1 U8196 ( .A1(n10819), .A2(n10813), .ZN(n13089) );
  NOR2_X2 U8197 ( .A1(n13282), .A2(n13281), .ZN(n13326) );
  NAND2_X1 U8198 ( .A1(n9486), .A2(n9485), .ZN(n13449) );
  OR2_X1 U8199 ( .A1(n13489), .A2(n9811), .ZN(n9486) );
  NAND2_X1 U8200 ( .A1(n9804), .A2(n9803), .ZN(n13339) );
  NAND2_X1 U8201 ( .A1(n9783), .A2(n9782), .ZN(n13340) );
  NAND2_X1 U8202 ( .A1(n10103), .A2(n13374), .ZN(n13385) );
  AND2_X1 U8203 ( .A1(n10099), .A2(n10098), .ZN(n15405) );
  OR2_X1 U8204 ( .A1(n15399), .A2(n13436), .ZN(n6635) );
  OAI21_X1 U8205 ( .B1(n13431), .B2(n13430), .A(n6637), .ZN(n6636) );
  AOI21_X1 U8206 ( .B1(n13432), .B2(n15405), .A(n6638), .ZN(n6637) );
  OR2_X1 U8207 ( .A1(n13768), .A2(n13738), .ZN(n7091) );
  INV_X1 U8208 ( .A(n13738), .ZN(n13714) );
  OR2_X1 U8209 ( .A1(n10089), .A2(n13372), .ZN(n9523) );
  OR2_X1 U8210 ( .A1(n13264), .A2(n9927), .ZN(n9521) );
  NAND2_X1 U8211 ( .A1(n13093), .A2(n13092), .ZN(n13862) );
  NAND2_X1 U8212 ( .A1(n6863), .A2(n6859), .ZN(n13864) );
  AOI21_X1 U8213 ( .B1(n13759), .B2(n6860), .A(n13763), .ZN(n6859) );
  INV_X1 U8214 ( .A(n13760), .ZN(n6863) );
  AOI22_X1 U8215 ( .A1(n7468), .A2(n7471), .B1(n7470), .B2(n7475), .ZN(n7467)
         );
  NAND2_X1 U8216 ( .A1(n7468), .A2(n6714), .ZN(n6713) );
  NAND2_X1 U8217 ( .A1(n7476), .A2(n7477), .ZN(n14092) );
  AND2_X1 U8218 ( .A1(n10902), .A2(n10898), .ZN(n7476) );
  NAND2_X1 U8219 ( .A1(n7480), .A2(n7478), .ZN(n14101) );
  NOR2_X1 U8220 ( .A1(n7479), .A2(n14099), .ZN(n7478) );
  INV_X1 U8221 ( .A(n7481), .ZN(n7479) );
  AND4_X1 U8222 ( .A1(n8886), .A2(n8885), .A3(n8884), .A4(n8883), .ZN(n15311)
         );
  AND2_X1 U8223 ( .A1(n10912), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14295) );
  AND2_X1 U8224 ( .A1(n10296), .A2(n10295), .ZN(n14281) );
  OAI21_X2 U8225 ( .B1(n10298), .B2(n11201), .A(n15236), .ZN(n14300) );
  NAND2_X1 U8226 ( .A1(n9200), .A2(n9199), .ZN(n14566) );
  INV_X1 U8227 ( .A(n15053), .ZN(n14884) );
  NAND2_X1 U8228 ( .A1(n14607), .A2(n10161), .ZN(n14619) );
  AND2_X1 U8229 ( .A1(n10170), .A2(n10169), .ZN(n15217) );
  OAI21_X1 U8230 ( .B1(n14464), .B2(n14463), .A(n14467), .ZN(n14689) );
  AND2_X1 U8231 ( .A1(n12140), .A2(n12139), .ZN(n14715) );
  NAND2_X1 U8232 ( .A1(n14717), .A2(n14718), .ZN(n7122) );
  NAND2_X1 U8233 ( .A1(n14731), .A2(n9272), .ZN(n14717) );
  NAND2_X1 U8234 ( .A1(n12148), .A2(n9270), .ZN(n14760) );
  NAND2_X1 U8235 ( .A1(n12149), .A2(n9143), .ZN(n14745) );
  INV_X1 U8236 ( .A(n7787), .ZN(n14744) );
  NAND2_X1 U8237 ( .A1(n11759), .A2(n8909), .ZN(n12028) );
  NAND2_X1 U8238 ( .A1(n6452), .A2(n9968), .ZN(n7431) );
  INV_X1 U8239 ( .A(n14974), .ZN(n15266) );
  INV_X1 U8240 ( .A(n7869), .ZN(n7798) );
  INV_X1 U8241 ( .A(n12132), .ZN(n12133) );
  AOI21_X1 U8242 ( .B1(n14567), .B2(n15107), .A(n12131), .ZN(n12132) );
  NAND2_X1 U8243 ( .A1(n7125), .A2(n7124), .ZN(n15117) );
  INV_X1 U8244 ( .A(n14992), .ZN(n7124) );
  INV_X1 U8245 ( .A(n7370), .ZN(n7125) );
  OAI21_X1 U8246 ( .B1(n14995), .B2(n15289), .A(n7371), .ZN(n7370) );
  NAND2_X1 U8247 ( .A1(n10506), .A2(n10504), .ZN(n15158) );
  OAI22_X1 U8248 ( .A1(n15183), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(n15182), 
        .B2(n6885), .ZN(n15188) );
  INV_X1 U8249 ( .A(n6886), .ZN(n6885) );
  OAI21_X1 U8250 ( .B1(n7706), .B2(n7703), .A(n7132), .ZN(n13123) );
  INV_X1 U8251 ( .A(n13123), .ZN(n7084) );
  INV_X1 U8252 ( .A(n13122), .ZN(n7083) );
  NAND2_X1 U8253 ( .A1(n14335), .A2(n14338), .ZN(n7408) );
  NOR2_X1 U8254 ( .A1(n14338), .A2(n14335), .ZN(n7409) );
  INV_X1 U8255 ( .A(n8439), .ZN(n7283) );
  OAI21_X1 U8256 ( .B1(n14352), .B2(n7398), .A(n7396), .ZN(n14358) );
  NOR2_X1 U8257 ( .A1(n14351), .A2(n14354), .ZN(n7398) );
  OR2_X1 U8258 ( .A1(n7397), .A2(n14353), .ZN(n7396) );
  NOR2_X1 U8259 ( .A1(n11164), .A2(n7280), .ZN(n7279) );
  NAND2_X1 U8260 ( .A1(n6434), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U8261 ( .A1(n8446), .A2(n7285), .ZN(n7278) );
  INV_X1 U8262 ( .A(n14391), .ZN(n7120) );
  INV_X1 U8263 ( .A(n8472), .ZN(n7296) );
  INV_X1 U8264 ( .A(n7292), .ZN(n7291) );
  NOR2_X1 U8265 ( .A1(n7297), .A2(n7290), .ZN(n7289) );
  NAND2_X1 U8266 ( .A1(n12779), .A2(n12071), .ZN(n7297) );
  NOR2_X1 U8267 ( .A1(n7292), .A2(n7293), .ZN(n7290) );
  NOR2_X1 U8268 ( .A1(n7296), .A2(n8476), .ZN(n7293) );
  NAND2_X1 U8269 ( .A1(n13153), .A2(n13155), .ZN(n7710) );
  NOR2_X1 U8270 ( .A1(n7401), .A2(n7402), .ZN(n7400) );
  NOR2_X1 U8271 ( .A1(n14394), .A2(n7118), .ZN(n7399) );
  AND2_X1 U8272 ( .A1(n14396), .A2(n7611), .ZN(n7401) );
  NAND2_X1 U8273 ( .A1(n14422), .A2(n7391), .ZN(n7390) );
  INV_X1 U8274 ( .A(n13168), .ZN(n7163) );
  OR2_X1 U8275 ( .A1(n6776), .A2(n13171), .ZN(n6774) );
  AND2_X1 U8276 ( .A1(n7388), .A2(n6542), .ZN(n6598) );
  NAND2_X1 U8277 ( .A1(n14421), .A2(n14423), .ZN(n7388) );
  NAND2_X1 U8278 ( .A1(n7308), .A2(n7307), .ZN(n8512) );
  NOR2_X1 U8279 ( .A1(n12692), .A2(n8507), .ZN(n7307) );
  NAND2_X1 U8280 ( .A1(n13182), .A2(n6767), .ZN(n6766) );
  INV_X1 U8281 ( .A(n13181), .ZN(n6767) );
  NAND2_X1 U8282 ( .A1(n13183), .A2(n13181), .ZN(n6768) );
  INV_X1 U8283 ( .A(n13185), .ZN(n7720) );
  INV_X1 U8284 ( .A(n13292), .ZN(n7502) );
  INV_X1 U8285 ( .A(n8999), .ZN(n8688) );
  NAND2_X1 U8286 ( .A1(n12476), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6760) );
  AND2_X1 U8287 ( .A1(n6760), .A2(n6759), .ZN(n6754) );
  INV_X1 U8288 ( .A(n12477), .ZN(n6755) );
  INV_X1 U8289 ( .A(n8051), .ZN(n7758) );
  INV_X1 U8290 ( .A(n6829), .ZN(n6828) );
  OAI21_X1 U8291 ( .B1(n7555), .B2(n6830), .A(n8286), .ZN(n6829) );
  INV_X1 U8292 ( .A(n8274), .ZN(n6830) );
  NAND2_X1 U8293 ( .A1(n7553), .A2(n8027), .ZN(n7552) );
  INV_X1 U8294 ( .A(n8025), .ZN(n7553) );
  OAI21_X1 U8295 ( .B1(n7509), .B2(n7502), .A(n13291), .ZN(n7497) );
  NOR2_X1 U8296 ( .A1(n7503), .A2(n7502), .ZN(n7501) );
  OR2_X1 U8297 ( .A1(n7508), .A2(n7502), .ZN(n7498) );
  NOR2_X1 U8298 ( .A1(n7489), .A2(n6903), .ZN(n6900) );
  INV_X1 U8299 ( .A(n11241), .ZN(n6903) );
  NAND2_X1 U8300 ( .A1(n9462), .A2(n13905), .ZN(n6671) );
  NAND2_X1 U8301 ( .A1(n14435), .A2(n14437), .ZN(n7116) );
  INV_X1 U8302 ( .A(n7862), .ZN(n7361) );
  NOR2_X1 U8303 ( .A1(n8990), .A2(n6711), .ZN(n6710) );
  NAND2_X1 U8304 ( .A1(n8608), .A2(n6424), .ZN(n8881) );
  NAND2_X1 U8305 ( .A1(n7883), .A2(n9236), .ZN(n9237) );
  INV_X1 U8306 ( .A(n11316), .ZN(n9236) );
  NOR2_X1 U8307 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8617) );
  NOR2_X1 U8308 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8618) );
  INV_X1 U8309 ( .A(n9117), .ZN(n8707) );
  NOR2_X1 U8310 ( .A1(n8702), .A2(n8706), .ZN(n6868) );
  INV_X1 U8311 ( .A(SI_16_), .ZN(n8685) );
  NAND2_X1 U8312 ( .A1(n7424), .A2(n7423), .ZN(n7422) );
  OAI21_X1 U8313 ( .B1(n7434), .B2(n10151), .A(n7080), .ZN(n8676) );
  NAND2_X1 U8314 ( .A1(n7434), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7080) );
  AND2_X1 U8315 ( .A1(n8784), .A2(n8765), .ZN(n6619) );
  NAND2_X1 U8316 ( .A1(n8659), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U8317 ( .A1(n8659), .A2(n9927), .ZN(n7115) );
  INV_X1 U8318 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7537) );
  OR2_X1 U8319 ( .A1(n11176), .A2(n12458), .ZN(n6931) );
  NAND2_X1 U8320 ( .A1(n7304), .A2(n12625), .ZN(n7302) );
  NAND2_X1 U8321 ( .A1(n7313), .A2(n7312), .ZN(n8529) );
  NOR2_X1 U8322 ( .A1(n8525), .A2(n12643), .ZN(n7312) );
  NOR2_X1 U8323 ( .A1(n6497), .A2(n7300), .ZN(n7299) );
  NAND2_X1 U8324 ( .A1(n8539), .A2(n10126), .ZN(n6822) );
  INV_X1 U8325 ( .A(n8548), .ZN(n8542) );
  INV_X1 U8326 ( .A(n10885), .ZN(n7661) );
  INV_X1 U8327 ( .A(n12006), .ZN(n6937) );
  OAI21_X1 U8328 ( .B1(n12542), .B2(n6742), .A(n6508), .ZN(n7386) );
  NAND2_X1 U8329 ( .A1(n12543), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n6742) );
  OR2_X1 U8330 ( .A1(n12555), .A2(n12832), .ZN(n7387) );
  OR2_X1 U8331 ( .A1(n8530), .A2(n7750), .ZN(n7749) );
  INV_X1 U8332 ( .A(n8527), .ZN(n7750) );
  INV_X1 U8333 ( .A(n7870), .ZN(n7825) );
  NAND2_X1 U8334 ( .A1(n7169), .A2(n6444), .ZN(n8307) );
  INV_X1 U8335 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n6695) );
  AND2_X1 U8336 ( .A1(n7732), .A2(n8516), .ZN(n7195) );
  NAND2_X1 U8337 ( .A1(n7735), .A2(n7191), .ZN(n7190) );
  INV_X1 U8338 ( .A(n8553), .ZN(n7191) );
  INV_X1 U8339 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n6698) );
  INV_X1 U8340 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8250) );
  NOR2_X1 U8341 ( .A1(n8205), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8222) );
  NOR2_X1 U8342 ( .A1(n8235), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7169) );
  INV_X1 U8343 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n6703) );
  NOR2_X1 U8344 ( .A1(n8140), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7170) );
  NOR2_X1 U8345 ( .A1(n8081), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7167) );
  INV_X1 U8346 ( .A(n7829), .ZN(n7828) );
  OAI21_X1 U8347 ( .B1(n11164), .B2(n7830), .A(n9338), .ZN(n7829) );
  INV_X1 U8348 ( .A(n9337), .ZN(n7830) );
  NAND2_X1 U8349 ( .A1(n6705), .A2(n7166), .ZN(n8044) );
  AND2_X1 U8350 ( .A1(n8441), .A2(n8442), .ZN(n7975) );
  INV_X1 U8351 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7942) );
  INV_X1 U8352 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n7941) );
  NAND2_X1 U8353 ( .A1(n11082), .A2(n8442), .ZN(n9333) );
  NOR2_X1 U8354 ( .A1(n8228), .A2(n7194), .ZN(n7193) );
  INV_X1 U8355 ( .A(n8418), .ZN(n7194) );
  NOR2_X1 U8356 ( .A1(n7727), .A2(n11595), .ZN(n7723) );
  INV_X1 U8357 ( .A(n11951), .ZN(n7727) );
  INV_X1 U8358 ( .A(n8475), .ZN(n7725) );
  NAND2_X1 U8359 ( .A1(n10950), .A2(n9337), .ZN(n11283) );
  INV_X1 U8360 ( .A(n8380), .ZN(n7574) );
  INV_X1 U8361 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8580) );
  NOR2_X1 U8362 ( .A1(n8340), .A2(n6843), .ZN(n6842) );
  INV_X1 U8363 ( .A(n8327), .ZN(n6843) );
  INV_X1 U8364 ( .A(n8229), .ZN(n6833) );
  NAND2_X1 U8365 ( .A1(n6849), .A2(n6427), .ZN(n8109) );
  OR2_X1 U8366 ( .A1(n8057), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U8367 ( .A1(n6821), .A2(n7972), .ZN(n6820) );
  INV_X1 U8368 ( .A(n7951), .ZN(n6821) );
  INV_X1 U8369 ( .A(n7005), .ZN(n7003) );
  NOR2_X1 U8370 ( .A1(n9703), .A2(n6689), .ZN(n6688) );
  NOR2_X1 U8371 ( .A1(n13070), .A2(n7599), .ZN(n7598) );
  INV_X1 U8372 ( .A(n12262), .ZN(n7599) );
  INV_X1 U8373 ( .A(n9690), .ZN(n9470) );
  OAI21_X1 U8374 ( .B1(n13188), .B2(n13187), .A(n13195), .ZN(n6772) );
  NOR2_X1 U8375 ( .A1(n6722), .A2(n6719), .ZN(n6718) );
  NAND2_X1 U8376 ( .A1(n13318), .A2(n13576), .ZN(n6722) );
  INV_X1 U8377 ( .A(n7694), .ZN(n7692) );
  NAND2_X1 U8378 ( .A1(n13869), .A2(n13231), .ZN(n7694) );
  NAND2_X1 U8379 ( .A1(n13521), .A2(n13197), .ZN(n7509) );
  NAND2_X1 U8380 ( .A1(n6401), .A2(n9857), .ZN(n7508) );
  AND2_X1 U8381 ( .A1(n9471), .A2(n6572), .ZN(n7159) );
  AND2_X1 U8382 ( .A1(n13887), .A2(n7695), .ZN(n7698) );
  INV_X1 U8383 ( .A(n7699), .ZN(n7695) );
  INV_X1 U8384 ( .A(n9854), .ZN(n6928) );
  NAND2_X1 U8385 ( .A1(n9471), .A2(n6691), .ZN(n9762) );
  NAND2_X1 U8386 ( .A1(n13606), .A2(n7696), .ZN(n7699) );
  INV_X1 U8387 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U8388 ( .A1(n7526), .A2(n7522), .ZN(n7524) );
  AND2_X1 U8389 ( .A1(n6413), .A2(n9672), .ZN(n7522) );
  NAND2_X1 U8390 ( .A1(n6686), .A2(n6568), .ZN(n9677) );
  NOR2_X1 U8391 ( .A1(n9664), .A2(n10722), .ZN(n7158) );
  NOR2_X1 U8392 ( .A1(n7105), .A2(n13846), .ZN(n7689) );
  NAND2_X1 U8393 ( .A1(n10751), .A2(n6676), .ZN(n9822) );
  NAND2_X1 U8394 ( .A1(n7152), .A2(n10806), .ZN(n6676) );
  INV_X1 U8395 ( .A(n9822), .ZN(n13300) );
  AND2_X1 U8396 ( .A1(n15412), .A2(n9905), .ZN(n10811) );
  NOR3_X1 U8397 ( .A1(n13517), .A2(n13765), .A3(n7694), .ZN(n13481) );
  OAI21_X1 U8398 ( .B1(n10094), .B2(n13438), .A(n9500), .ZN(n9501) );
  INV_X1 U8399 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9459) );
  INV_X1 U8400 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n15527) );
  INV_X1 U8401 ( .A(n7461), .ZN(n7460) );
  INV_X1 U8402 ( .A(n14225), .ZN(n7459) );
  OR2_X1 U8403 ( .A1(n12174), .A2(n12173), .ZN(n7866) );
  NOR2_X1 U8404 ( .A1(n9123), .A2(n9122), .ZN(n6707) );
  AOI21_X1 U8405 ( .B1(n7485), .B2(n11938), .A(n12160), .ZN(n7484) );
  AND2_X1 U8406 ( .A1(n8614), .A2(n8613), .ZN(n9080) );
  NAND2_X1 U8407 ( .A1(n6797), .A2(n14192), .ZN(n6796) );
  XNOR2_X1 U8408 ( .A(n6709), .B(n14051), .ZN(n14055) );
  NAND2_X1 U8409 ( .A1(n14049), .A2(n14050), .ZN(n6709) );
  CLKBUF_X1 U8410 ( .A(n14448), .Z(n14460) );
  INV_X1 U8411 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7008) );
  INV_X1 U8412 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7007) );
  AND2_X1 U8413 ( .A1(n6466), .A2(n7451), .ZN(n7450) );
  INV_X1 U8414 ( .A(n9272), .ZN(n7807) );
  NOR2_X1 U8415 ( .A1(n14850), .A2(n15030), .ZN(n7441) );
  NOR2_X1 U8416 ( .A1(n7056), .A2(n7050), .ZN(n7049) );
  OR2_X1 U8417 ( .A1(n7361), .A2(n7057), .ZN(n7056) );
  INV_X1 U8418 ( .A(n9261), .ZN(n7057) );
  OR2_X1 U8419 ( .A1(n7361), .A2(n7054), .ZN(n7053) );
  NAND2_X1 U8420 ( .A1(n7055), .A2(n9261), .ZN(n7054) );
  INV_X1 U8421 ( .A(n7058), .ZN(n7055) );
  INV_X1 U8422 ( .A(n14390), .ZN(n7366) );
  NOR2_X1 U8423 ( .A1(n7021), .A2(n7019), .ZN(n7018) );
  INV_X1 U8424 ( .A(n8963), .ZN(n7019) );
  INV_X1 U8425 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9007) );
  AND2_X1 U8426 ( .A1(n7367), .A2(n9255), .ZN(n7150) );
  NAND2_X1 U8427 ( .A1(n8611), .A2(n6710), .ZN(n9025) );
  NAND2_X1 U8428 ( .A1(n8610), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8956) );
  INV_X1 U8429 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8955) );
  INV_X1 U8430 ( .A(n8973), .ZN(n8611) );
  NAND2_X1 U8431 ( .A1(n8609), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8938) );
  INV_X1 U8432 ( .A(n8919), .ZN(n8609) );
  INV_X1 U8433 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8900) );
  OR2_X1 U8434 ( .A1(n8901), .A2(n8900), .ZN(n8919) );
  NOR2_X1 U8435 ( .A1(n7038), .A2(n7883), .ZN(n7033) );
  NAND3_X1 U8436 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U8437 ( .A1(n9185), .A2(n7108), .ZN(n9204) );
  NAND2_X1 U8438 ( .A1(n7109), .A2(SI_27_), .ZN(n7108) );
  INV_X1 U8439 ( .A(n9184), .ZN(n7109) );
  AOI21_X1 U8440 ( .B1(n8695), .B2(n9056), .A(n8694), .ZN(n8696) );
  NAND2_X1 U8441 ( .A1(n9059), .A2(n9060), .ZN(n6806) );
  NAND2_X1 U8442 ( .A1(n6716), .A2(n6855), .ZN(n9053) );
  XNOR2_X1 U8443 ( .A(n9053), .B(SI_18_), .ZN(n9052) );
  AND2_X1 U8444 ( .A1(n6412), .A2(n9012), .ZN(n7413) );
  OR2_X1 U8445 ( .A1(n8987), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8935) );
  INV_X1 U8446 ( .A(n8888), .ZN(n8672) );
  AOI21_X1 U8447 ( .B1(n8888), .B2(SI_10_), .A(n8912), .ZN(n8929) );
  NAND2_X1 U8448 ( .A1(n7434), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U8449 ( .A1(n6729), .A2(n7521), .ZN(n6728) );
  NAND2_X1 U8450 ( .A1(n8659), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U8451 ( .A1(n6728), .A2(SI_6_), .ZN(n8663) );
  XNOR2_X1 U8452 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n9948) );
  INV_X1 U8453 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n6879) );
  NOR2_X1 U8454 ( .A1(n10935), .A2(n6974), .ZN(n6973) );
  NAND2_X1 U8455 ( .A1(n10932), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n7136) );
  NAND2_X1 U8456 ( .A1(n12098), .A2(n12097), .ZN(n15163) );
  NOR2_X1 U8457 ( .A1(n15172), .A2(n15171), .ZN(n15178) );
  XNOR2_X1 U8458 ( .A(n15178), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15179) );
  INV_X1 U8459 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10610) );
  AND2_X1 U8460 ( .A1(n10515), .A2(n10514), .ZN(n10516) );
  INV_X1 U8461 ( .A(n10512), .ZN(n7328) );
  OAI21_X1 U8462 ( .B1(n7648), .B2(n6512), .A(n6907), .ZN(n12363) );
  AND2_X1 U8463 ( .A1(n7635), .A2(n6910), .ZN(n6907) );
  XNOR2_X1 U8464 ( .A(n11412), .B(n11174), .ZN(n10687) );
  INV_X1 U8465 ( .A(n7868), .ZN(n7644) );
  OR2_X1 U8466 ( .A1(n12343), .A2(n7646), .ZN(n7645) );
  INV_X1 U8467 ( .A(n12425), .ZN(n7646) );
  NAND2_X1 U8468 ( .A1(n7170), .A2(n6701), .ZN(n8205) );
  AND2_X1 U8469 ( .A1(n6439), .A2(n6702), .ZN(n6701) );
  INV_X1 U8470 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n6702) );
  OAI21_X1 U8471 ( .B1(n8551), .B2(n8547), .A(n7540), .ZN(n8549) );
  NOR2_X1 U8472 ( .A1(n7541), .A2(n8545), .ZN(n7540) );
  NAND2_X1 U8473 ( .A1(n7543), .A2(n7542), .ZN(n7541) );
  AND2_X1 U8474 ( .A1(n10513), .A2(n11564), .ZN(n10512) );
  NAND2_X1 U8475 ( .A1(n7240), .A2(n7239), .ZN(n7238) );
  OR2_X1 U8476 ( .A1(n12937), .A2(n15491), .ZN(n7240) );
  NAND2_X1 U8477 ( .A1(n12937), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7239) );
  OR2_X1 U8478 ( .A1(n10405), .A2(n10390), .ZN(n6958) );
  NAND2_X1 U8479 ( .A1(n10394), .A2(n10547), .ZN(n10395) );
  OR2_X1 U8480 ( .A1(n10541), .A2(n11090), .ZN(n10543) );
  AOI21_X1 U8481 ( .B1(n7263), .B2(n7262), .A(n6515), .ZN(n7261) );
  INV_X1 U8482 ( .A(n7267), .ZN(n7262) );
  NAND2_X1 U8483 ( .A1(n10882), .A2(n7661), .ZN(n7659) );
  AND2_X1 U8484 ( .A1(n6941), .A2(n6943), .ZN(n11481) );
  NAND2_X1 U8485 ( .A1(n6570), .A2(n6941), .ZN(n11538) );
  OAI21_X1 U8486 ( .B1(n6749), .B2(n10877), .A(n6744), .ZN(n7376) );
  INV_X1 U8487 ( .A(n6745), .ZN(n6744) );
  OAI21_X1 U8488 ( .B1(n6748), .B2(n10877), .A(n6518), .ZN(n6745) );
  NOR2_X1 U8489 ( .A1(n7663), .A2(n11927), .ZN(n7662) );
  NAND2_X1 U8490 ( .A1(n11918), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U8491 ( .A1(n12003), .A2(n6937), .ZN(n6935) );
  XNOR2_X1 U8492 ( .A(n12497), .B(n12478), .ZN(n12479) );
  INV_X1 U8493 ( .A(n12536), .ZN(n12538) );
  NAND3_X1 U8494 ( .A1(n7679), .A2(n6442), .A3(n12536), .ZN(n7677) );
  NAND2_X1 U8495 ( .A1(n7677), .A2(n7680), .ZN(n6955) );
  NAND2_X1 U8496 ( .A1(n12538), .A2(n12537), .ZN(n7678) );
  NAND2_X1 U8497 ( .A1(n7252), .A2(n6563), .ZN(n7251) );
  NOR2_X1 U8498 ( .A1(n7250), .A2(n12558), .ZN(n7249) );
  NAND2_X1 U8499 ( .A1(n12588), .A2(n7676), .ZN(n7675) );
  NAND2_X1 U8500 ( .A1(n7383), .A2(n6732), .ZN(n6731) );
  AOI21_X1 U8501 ( .B1(n7745), .B2(n7197), .A(n7744), .ZN(n7743) );
  INV_X1 U8502 ( .A(n8539), .ZN(n7744) );
  NAND2_X1 U8503 ( .A1(n8306), .A2(n6699), .ZN(n8334) );
  AND2_X1 U8504 ( .A1(n8305), .A2(n6700), .ZN(n6699) );
  NAND2_X1 U8505 ( .A1(n8306), .A2(n8305), .ZN(n8320) );
  XNOR2_X1 U8506 ( .A(n6661), .B(n12643), .ZN(n6660) );
  AOI21_X1 U8507 ( .B1(n12654), .B2(n7879), .A(n7825), .ZN(n6661) );
  NAND2_X1 U8508 ( .A1(n12665), .A2(n9351), .ZN(n12654) );
  NAND2_X1 U8509 ( .A1(n7169), .A2(n6584), .ZN(n8277) );
  NAND2_X1 U8510 ( .A1(n7169), .A2(n8250), .ZN(n8265) );
  NAND2_X1 U8511 ( .A1(n8222), .A2(n8221), .ZN(n8235) );
  INV_X1 U8512 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8221) );
  INV_X1 U8513 ( .A(n7169), .ZN(n8251) );
  AOI21_X1 U8514 ( .B1(n12746), .B2(n12745), .A(n7842), .ZN(n12731) );
  INV_X1 U8515 ( .A(n7850), .ZN(n7842) );
  INV_X1 U8516 ( .A(n12770), .ZN(n12748) );
  NAND2_X1 U8517 ( .A1(n7170), .A2(n6439), .ZN(n8189) );
  NAND2_X1 U8518 ( .A1(n7170), .A2(n8157), .ZN(n8175) );
  INV_X1 U8519 ( .A(n7170), .ZN(n8158) );
  NAND2_X1 U8520 ( .A1(n6694), .A2(n8117), .ZN(n8140) );
  INV_X1 U8521 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8117) );
  INV_X1 U8522 ( .A(n8118), .ZN(n6694) );
  NAND2_X1 U8523 ( .A1(n7167), .A2(n8099), .ZN(n8118) );
  INV_X1 U8524 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8099) );
  INV_X1 U8525 ( .A(n7167), .ZN(n8100) );
  AND2_X1 U8526 ( .A1(n7166), .A2(n8043), .ZN(n6704) );
  INV_X1 U8527 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8043) );
  OR2_X1 U8528 ( .A1(n8062), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8081) );
  INV_X1 U8529 ( .A(n12456), .ZN(n11353) );
  AND2_X1 U8530 ( .A1(n7219), .A2(n9336), .ZN(n7218) );
  NAND2_X1 U8531 ( .A1(n10951), .A2(n11164), .ZN(n10950) );
  NAND4_X1 U8532 ( .A1(n7941), .A2(n10610), .A3(n6706), .A4(n7942), .ZN(n8000)
         );
  INV_X1 U8533 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U8534 ( .A1(n8450), .A2(n8449), .ZN(n10966) );
  NAND2_X1 U8535 ( .A1(n10610), .A2(n7941), .ZN(n7963) );
  OAI21_X1 U8536 ( .B1(n7936), .B2(n10736), .A(n8556), .ZN(n7937) );
  NAND2_X1 U8537 ( .A1(n10581), .A2(n8428), .ZN(n15457) );
  INV_X1 U8538 ( .A(n10520), .ZN(n8425) );
  AND2_X1 U8539 ( .A1(n10252), .A2(n12829), .ZN(n10248) );
  AND2_X1 U8540 ( .A1(n10235), .A2(n10619), .ZN(n10623) );
  AND2_X1 U8541 ( .A1(n12450), .A2(n12142), .ZN(n12844) );
  AOI21_X1 U8542 ( .B1(n12627), .B2(n8355), .A(n8338), .ZN(n12357) );
  AND2_X1 U8543 ( .A1(n7836), .A2(n12352), .ZN(n7835) );
  NAND2_X1 U8544 ( .A1(n7838), .A2(n7840), .ZN(n7836) );
  OR2_X1 U8545 ( .A1(n9358), .A2(n12352), .ZN(n9359) );
  NAND2_X1 U8546 ( .A1(n7834), .A2(n7838), .ZN(n9358) );
  NAND2_X1 U8547 ( .A1(n7841), .A2(n7839), .ZN(n7834) );
  AND2_X1 U8548 ( .A1(n7823), .A2(n12643), .ZN(n7822) );
  NAND2_X1 U8549 ( .A1(n7845), .A2(n7843), .ZN(n7201) );
  NAND2_X1 U8550 ( .A1(n7849), .A2(n7844), .ZN(n7843) );
  NAND2_X1 U8551 ( .A1(n9348), .A2(n7850), .ZN(n7844) );
  AOI21_X1 U8552 ( .B1(n7205), .B2(n7208), .A(n6521), .ZN(n7204) );
  NOR2_X1 U8553 ( .A1(n6416), .A2(n9345), .ZN(n7205) );
  NAND2_X1 U8554 ( .A1(n7173), .A2(n7176), .ZN(n12766) );
  AOI21_X1 U8555 ( .B1(n12779), .B2(n7178), .A(n7177), .ZN(n7176) );
  INV_X1 U8556 ( .A(n8480), .ZN(n7177) );
  NOR2_X1 U8557 ( .A1(n11951), .A2(n7855), .ZN(n7854) );
  INV_X1 U8558 ( .A(n9343), .ZN(n7855) );
  NAND2_X1 U8559 ( .A1(n7856), .A2(n9343), .ZN(n11952) );
  AOI21_X1 U8560 ( .B1(n7183), .B2(n7186), .A(n7182), .ZN(n7181) );
  INV_X1 U8561 ( .A(n8467), .ZN(n7182) );
  NAND2_X1 U8562 ( .A1(n11350), .A2(n11349), .ZN(n6648) );
  OR2_X1 U8563 ( .A1(n9406), .A2(n9405), .ZN(n10250) );
  OAI21_X1 U8564 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8362) );
  INV_X1 U8565 ( .A(n8073), .ZN(n7819) );
  AND2_X1 U8566 ( .A1(n7903), .A2(n7892), .ZN(n7817) );
  INV_X1 U8567 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7893) );
  INV_X1 U8568 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U8569 ( .A1(n8216), .A2(n7820), .ZN(n7818) );
  INV_X1 U8570 ( .A(n8602), .ZN(n11473) );
  XNOR2_X1 U8571 ( .A(n7319), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U8572 ( .A1(n7320), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7319) );
  AND2_X1 U8573 ( .A1(n8590), .A2(n8588), .ZN(n7133) );
  XNOR2_X1 U8574 ( .A(n8587), .B(n8588), .ZN(n10124) );
  OAI21_X1 U8575 ( .B1(n8586), .B2(n8585), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8587) );
  INV_X1 U8576 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8582) );
  OR2_X1 U8577 ( .A1(n8183), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8200) );
  OR2_X1 U8578 ( .A1(n8148), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8150) );
  XNOR2_X1 U8579 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8068) );
  OAI21_X1 U8580 ( .B1(n7991), .B2(n6846), .A(n6844), .ZN(n8037) );
  INV_X1 U8581 ( .A(n7549), .ZN(n6846) );
  XNOR2_X1 U8582 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8052) );
  OR2_X1 U8583 ( .A1(n8028), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8038) );
  INV_X1 U8584 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U8585 ( .A1(n7900), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7919) );
  INV_X1 U8586 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U8587 ( .A1(n6690), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9738) );
  INV_X1 U8588 ( .A(n9725), .ZN(n6690) );
  NAND2_X1 U8589 ( .A1(n9471), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9749) );
  AOI21_X1 U8590 ( .B1(n7595), .B2(n13025), .A(n6520), .ZN(n7594) );
  INV_X1 U8591 ( .A(n12232), .ZN(n7597) );
  NOR2_X1 U8592 ( .A1(n7598), .A2(n6984), .ZN(n6983) );
  INV_X1 U8593 ( .A(n12265), .ZN(n6984) );
  NOR2_X1 U8594 ( .A1(n12268), .A2(n12267), .ZN(n6982) );
  NAND2_X1 U8595 ( .A1(n9468), .A2(n6423), .ZN(n9604) );
  INV_X1 U8596 ( .A(n6998), .ZN(n6991) );
  NAND2_X1 U8597 ( .A1(n6999), .A2(n6998), .ZN(n6992) );
  INV_X1 U8598 ( .A(n6995), .ZN(n6994) );
  OR2_X1 U8599 ( .A1(n12214), .A2(n11051), .ZN(n10804) );
  NAND2_X1 U8600 ( .A1(n9470), .A2(n6687), .ZN(n9725) );
  AND2_X1 U8601 ( .A1(n6688), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6687) );
  AND2_X1 U8602 ( .A1(n6977), .A2(n6528), .ZN(n6976) );
  NAND2_X1 U8603 ( .A1(n6414), .A2(n6980), .ZN(n6977) );
  NOR2_X1 U8604 ( .A1(n12971), .A2(n12250), .ZN(n7146) );
  OR2_X1 U8605 ( .A1(n9797), .A2(n13034), .ZN(n9808) );
  NAND2_X1 U8606 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9550) );
  NAND2_X1 U8607 ( .A1(n9469), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9621) );
  INV_X1 U8608 ( .A(n9606), .ZN(n9469) );
  NAND2_X1 U8609 ( .A1(n11661), .A2(n11662), .ZN(n11740) );
  NAND2_X1 U8610 ( .A1(n7590), .A2(n12272), .ZN(n10956) );
  OR2_X1 U8611 ( .A1(n9621), .A2(n9620), .ZN(n9637) );
  NAND2_X1 U8612 ( .A1(n6686), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U8613 ( .A1(n7607), .A2(n7609), .ZN(n7606) );
  XNOR2_X1 U8614 ( .A(n6425), .B(n13113), .ZN(n6990) );
  NAND2_X1 U8615 ( .A1(n12229), .A2(n12228), .ZN(n13023) );
  INV_X1 U8616 ( .A(n13022), .ZN(n12229) );
  NAND2_X1 U8617 ( .A1(n9468), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U8618 ( .A1(n7157), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9690) );
  INV_X1 U8619 ( .A(n9677), .ZN(n7157) );
  NAND2_X1 U8620 ( .A1(n9470), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9704) );
  AND2_X1 U8621 ( .A1(n13275), .A2(n13276), .ZN(n7106) );
  AND2_X1 U8622 ( .A1(n6398), .A2(n13666), .ZN(n13286) );
  OR2_X1 U8623 ( .A1(n9814), .A2(n11004), .ZN(n9540) );
  AOI21_X1 U8624 ( .B1(n6630), .B2(n6632), .A(n6628), .ZN(n6627) );
  INV_X1 U8625 ( .A(n15374), .ZN(n6628) );
  OR2_X1 U8626 ( .A1(n15384), .A2(n15383), .ZN(n15386) );
  AOI21_X1 U8627 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n15380) );
  INV_X1 U8628 ( .A(n6642), .ZN(n15381) );
  AND2_X1 U8629 ( .A1(n10593), .A2(n10592), .ZN(n10596) );
  NAND2_X1 U8630 ( .A1(n10596), .A2(n10595), .ZN(n10728) );
  INV_X1 U8631 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10722) );
  XNOR2_X1 U8632 ( .A(n11886), .B(n11611), .ZN(n11888) );
  NAND2_X1 U8633 ( .A1(n11606), .A2(n11605), .ZN(n11883) );
  AOI22_X1 U8634 ( .A1(n11888), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n11886), 
        .B2(n11887), .ZN(n13400) );
  OAI22_X1 U8635 ( .A1(n13400), .A2(n13399), .B1(n13398), .B2(n15531), .ZN(
        n15401) );
  AOI21_X1 U8636 ( .B1(n15401), .B2(n15402), .A(n6643), .ZN(n13420) );
  AND2_X1 U8637 ( .A1(n13410), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6643) );
  XNOR2_X1 U8638 ( .A(n13428), .B(n13427), .ZN(n13432) );
  NAND2_X1 U8639 ( .A1(n13337), .A2(n13771), .ZN(n7087) );
  NAND2_X1 U8640 ( .A1(n13453), .A2(n13717), .ZN(n7078) );
  AND2_X1 U8641 ( .A1(n9490), .A2(n9489), .ZN(n13502) );
  NAND2_X1 U8642 ( .A1(n7505), .A2(n6401), .ZN(n7503) );
  AND2_X1 U8643 ( .A1(n7508), .A2(n7509), .ZN(n7507) );
  NAND2_X1 U8644 ( .A1(n7159), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U8645 ( .A1(n7697), .A2(n7698), .ZN(n13584) );
  AND2_X1 U8646 ( .A1(n6925), .A2(n9853), .ZN(n6924) );
  NAND2_X1 U8647 ( .A1(n6927), .A2(n6926), .ZN(n6925) );
  INV_X1 U8648 ( .A(n7514), .ZN(n6926) );
  INV_X1 U8649 ( .A(n13576), .ZN(n13582) );
  NAND2_X1 U8650 ( .A1(n13627), .A2(n7514), .ZN(n6929) );
  NAND2_X1 U8651 ( .A1(n6664), .A2(n6667), .ZN(n13645) );
  INV_X1 U8652 ( .A(n6668), .ZN(n6667) );
  NAND2_X1 U8653 ( .A1(n7340), .A2(n13704), .ZN(n6664) );
  NOR2_X1 U8654 ( .A1(n13705), .A2(n13828), .ZN(n13657) );
  NAND2_X1 U8655 ( .A1(n6607), .A2(n6606), .ZN(n13705) );
  AND3_X1 U8656 ( .A1(n11698), .A2(n11695), .A3(n7689), .ZN(n13727) );
  OR2_X1 U8657 ( .A1(n13152), .A2(n7687), .ZN(n12047) );
  NAND2_X1 U8658 ( .A1(n11695), .A2(n7688), .ZN(n7687) );
  AND2_X1 U8659 ( .A1(n13315), .A2(n9833), .ZN(n7127) );
  NAND2_X1 U8660 ( .A1(n11691), .A2(n13311), .ZN(n11690) );
  XNOR2_X1 U8661 ( .A(n13152), .B(n13346), .ZN(n13311) );
  INV_X1 U8662 ( .A(n9612), .ZN(n6685) );
  AND2_X1 U8663 ( .A1(n9616), .A2(n6684), .ZN(n6683) );
  NAND2_X1 U8664 ( .A1(n9612), .A2(n13306), .ZN(n6684) );
  NAND2_X1 U8665 ( .A1(n11695), .A2(n11698), .ZN(n11856) );
  XNOR2_X1 U8666 ( .A(n13348), .B(n13145), .ZN(n9830) );
  INV_X1 U8667 ( .A(n11296), .ZN(n6620) );
  NAND2_X1 U8668 ( .A1(n11294), .A2(n11297), .ZN(n11573) );
  NAND2_X1 U8669 ( .A1(n10978), .A2(n9525), .ZN(n10747) );
  NAND2_X1 U8670 ( .A1(n10747), .A2(n10752), .ZN(n10746) );
  CLKBUF_X1 U8671 ( .A(n9822), .Z(n10979) );
  NAND2_X1 U8672 ( .A1(n10979), .A2(n10980), .ZN(n10978) );
  NAND2_X1 U8673 ( .A1(n10974), .A2(n10973), .ZN(n10984) );
  INV_X1 U8674 ( .A(n10814), .ZN(n10820) );
  AND2_X1 U8675 ( .A1(n13242), .A2(n13241), .ZN(n13762) );
  NAND2_X1 U8676 ( .A1(n6862), .A2(n6861), .ZN(n6860) );
  NOR2_X1 U8677 ( .A1(n13755), .A2(n13470), .ZN(n6861) );
  INV_X1 U8678 ( .A(n13758), .ZN(n6862) );
  XNOR2_X1 U8679 ( .A(n13758), .B(n13470), .ZN(n13768) );
  NAND2_X1 U8680 ( .A1(n13771), .A2(n13851), .ZN(n7077) );
  NAND2_X1 U8681 ( .A1(n13696), .A2(n9842), .ZN(n13675) );
  INV_X1 U8682 ( .A(n12272), .ZN(n13840) );
  OR2_X1 U8683 ( .A1(n15421), .A2(n13286), .ZN(n15439) );
  INV_X1 U8684 ( .A(n15439), .ZN(n13851) );
  NAND2_X1 U8685 ( .A1(n13840), .A2(n13433), .ZN(n10814) );
  AND2_X1 U8686 ( .A1(n10093), .A2(n11491), .ZN(n10855) );
  INV_X1 U8687 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9476) );
  INV_X1 U8688 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9438) );
  NOR2_X1 U8689 ( .A1(n6417), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n7610) );
  INV_X1 U8690 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9876) );
  AND2_X1 U8691 ( .A1(n9660), .A2(n9684), .ZN(n11608) );
  OR2_X1 U8692 ( .A1(n9645), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n9647) );
  OR2_X1 U8693 ( .A1(n9617), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9712) );
  OR2_X1 U8694 ( .A1(n9558), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U8695 ( .A1(n8608), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8864) );
  NOR2_X1 U8696 ( .A1(n14058), .A2(n7471), .ZN(n7470) );
  INV_X1 U8697 ( .A(n7458), .ZN(n6793) );
  NAND2_X1 U8698 ( .A1(n12177), .A2(n12176), .ZN(n13934) );
  NAND2_X1 U8699 ( .A1(n7466), .A2(n7468), .ZN(n14121) );
  NOR2_X1 U8700 ( .A1(n11826), .A2(n7486), .ZN(n7485) );
  INV_X1 U8701 ( .A(n7488), .ZN(n7486) );
  NAND2_X1 U8702 ( .A1(n11820), .A2(n11819), .ZN(n7488) );
  OR2_X1 U8703 ( .A1(n11939), .A2(n11938), .ZN(n7487) );
  OAI21_X1 U8704 ( .B1(n11445), .B2(n11444), .A(n11443), .ZN(n11450) );
  AND2_X1 U8705 ( .A1(n14155), .A2(n14037), .ZN(n14203) );
  AND2_X1 U8706 ( .A1(n14081), .A2(n14019), .ZN(n14245) );
  XNOR2_X1 U8707 ( .A(n10661), .B(n14111), .ZN(n10895) );
  OR2_X1 U8708 ( .A1(n9156), .A2(n14285), .ZN(n9172) );
  NAND2_X1 U8709 ( .A1(n8615), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9156) );
  INV_X1 U8710 ( .A(n9135), .ZN(n8615) );
  NAND2_X1 U8711 ( .A1(n7358), .A2(n8989), .ZN(n9256) );
  NOR2_X1 U8712 ( .A1(n14491), .A2(n7615), .ZN(n7612) );
  INV_X1 U8713 ( .A(n6526), .ZN(n7615) );
  INV_X1 U8714 ( .A(n14518), .ZN(n7613) );
  AOI21_X1 U8715 ( .B1(n14778), .B2(n9216), .A(n9128), .ZN(n14251) );
  OR2_X1 U8716 ( .A1(n9136), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8761) );
  OAI21_X1 U8717 ( .B1(n10349), .B2(n10225), .A(n10224), .ZN(n10309) );
  OAI21_X1 U8718 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(n10557) );
  AOI21_X1 U8719 ( .B1(n10768), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10767), .ZN(
        n10772) );
  INV_X1 U8720 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8984) );
  NOR2_X2 U8721 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n8985) );
  XNOR2_X1 U8722 ( .A(n11794), .B(n7072), .ZN(n11972) );
  AOI21_X1 U8723 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n14643) );
  AOI21_X1 U8724 ( .B1(n14644), .B2(P1_REG2_REG_17__SCAN_IN), .A(n14643), .ZN(
        n14662) );
  XNOR2_X1 U8725 ( .A(n14660), .B(n7145), .ZN(n14659) );
  INV_X1 U8726 ( .A(n9208), .ZN(n14700) );
  AND2_X1 U8727 ( .A1(n9208), .A2(n9194), .ZN(n14708) );
  AOI21_X1 U8728 ( .B1(n7780), .B2(n7783), .A(n6522), .ZN(n7778) );
  NAND2_X1 U8729 ( .A1(n14758), .A2(n9271), .ZN(n14732) );
  NAND2_X1 U8730 ( .A1(n14747), .A2(n14755), .ZN(n14748) );
  NOR2_X1 U8731 ( .A1(n14759), .A2(n7803), .ZN(n7802) );
  INV_X1 U8732 ( .A(n9270), .ZN(n7803) );
  NAND2_X1 U8733 ( .A1(n7029), .A2(n7028), .ZN(n12150) );
  NAND2_X1 U8734 ( .A1(n14856), .A2(n15038), .ZN(n14829) );
  INV_X1 U8735 ( .A(n15064), .ZN(n7447) );
  INV_X1 U8736 ( .A(n7443), .ZN(n7445) );
  NAND2_X1 U8737 ( .A1(n7444), .A2(n6567), .ZN(n14916) );
  OR2_X1 U8738 ( .A1(n8956), .A2(n8955), .ZN(n8973) );
  NAND2_X1 U8739 ( .A1(n8611), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8991) );
  NAND2_X1 U8740 ( .A1(n15240), .A2(n14672), .ZN(n10300) );
  INV_X1 U8741 ( .A(n7790), .ZN(n7047) );
  AOI21_X1 U8742 ( .B1(n7046), .B2(n7790), .A(n7045), .ZN(n7044) );
  NOR2_X1 U8743 ( .A1(n14944), .A2(n14961), .ZN(n7790) );
  NOR2_X1 U8744 ( .A1(n14962), .A2(n15086), .ZN(n14954) );
  AND2_X1 U8745 ( .A1(n7765), .A2(n14539), .ZN(n7764) );
  NAND2_X1 U8746 ( .A1(n7766), .A2(n8909), .ZN(n7765) );
  INV_X1 U8747 ( .A(n7042), .ZN(n7041) );
  NAND2_X1 U8748 ( .A1(n15241), .A2(n6495), .ZN(n11760) );
  NAND2_X1 U8749 ( .A1(n15241), .A2(n7438), .ZN(n11646) );
  INV_X1 U8750 ( .A(n14696), .ZN(n14964) );
  AND2_X1 U8751 ( .A1(n15264), .A2(n15298), .ZN(n15241) );
  AND3_X1 U8752 ( .A1(n11506), .A2(n15246), .A3(n7435), .ZN(n15264) );
  AND2_X1 U8753 ( .A1(n6406), .A2(n15275), .ZN(n7435) );
  XNOR2_X1 U8754 ( .A(n14578), .B(n6407), .ZN(n15252) );
  NAND2_X1 U8755 ( .A1(n7436), .A2(n15246), .ZN(n15265) );
  INV_X1 U8756 ( .A(n11505), .ZN(n7436) );
  OAI21_X1 U8757 ( .B1(n7763), .B2(n14318), .A(n14327), .ZN(n7071) );
  NAND2_X1 U8758 ( .A1(n11506), .A2(n15275), .ZN(n11505) );
  NAND2_X1 U8759 ( .A1(n6452), .A2(n7434), .ZN(n7430) );
  NOR2_X1 U8760 ( .A1(n14484), .A2(n15310), .ZN(n12131) );
  AND2_X1 U8761 ( .A1(n14994), .A2(n15315), .ZN(n7372) );
  NAND2_X1 U8762 ( .A1(n15017), .A2(n15315), .ZN(n7067) );
  AND2_X1 U8763 ( .A1(n9087), .A2(n9086), .ZN(n15027) );
  OR2_X1 U8764 ( .A1(n14818), .A2(n9136), .ZN(n9087) );
  AND3_X1 U8765 ( .A1(n9030), .A2(n9029), .A3(n9028), .ZN(n15053) );
  INV_X1 U8766 ( .A(n15315), .ZN(n15302) );
  XNOR2_X1 U8767 ( .A(n12197), .B(n12196), .ZN(n13239) );
  XNOR2_X1 U8768 ( .A(n9204), .B(n9203), .ZN(n12269) );
  XNOR2_X1 U8769 ( .A(n9184), .B(n9167), .ZN(n12064) );
  XNOR2_X1 U8770 ( .A(n9303), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9309) );
  AND2_X1 U8771 ( .A1(n9300), .A2(n9299), .ZN(n9308) );
  AOI21_X1 U8772 ( .B1(n8702), .B2(n6873), .A(n6513), .ZN(n6872) );
  INV_X1 U8773 ( .A(n7428), .ZN(n6873) );
  XNOR2_X1 U8774 ( .A(n9306), .B(n9305), .ZN(n10041) );
  INV_X1 U8775 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9305) );
  OAI21_X1 U8776 ( .B1(n9304), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9306) );
  XNOR2_X1 U8777 ( .A(n9222), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U8778 ( .A1(n6805), .A2(n6804), .ZN(n9227) );
  NOR2_X1 U8779 ( .A1(n6806), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8780 ( .A1(n7418), .A2(n7417), .ZN(n9013) );
  NAND2_X1 U8781 ( .A1(n6412), .A2(n8964), .ZN(n7418) );
  AND2_X1 U8782 ( .A1(n9018), .A2(n9017), .ZN(n14636) );
  NAND2_X1 U8783 ( .A1(n8979), .A2(n7351), .ZN(n8982) );
  AND2_X1 U8784 ( .A1(n8969), .A2(n8952), .ZN(n11112) );
  NAND2_X1 U8785 ( .A1(n8911), .A2(n8910), .ZN(n8913) );
  OR2_X1 U8786 ( .A1(n8928), .A2(n8888), .ZN(n8889) );
  AND2_X1 U8787 ( .A1(n8860), .A2(n9002), .ZN(n10312) );
  OR2_X1 U8788 ( .A1(n8829), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8839) );
  OAI21_X1 U8789 ( .B1(SI_6_), .B2(n6728), .A(n8663), .ZN(n8825) );
  INV_X1 U8790 ( .A(n8803), .ZN(n8805) );
  INV_X1 U8791 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8809) );
  AND2_X1 U8792 ( .A1(n10069), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9949) );
  AND2_X1 U8793 ( .A1(n9939), .A2(n9938), .ZN(n9946) );
  OR2_X1 U8794 ( .A1(n10052), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10054) );
  XNOR2_X1 U8795 ( .A(n10491), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U8796 ( .A1(n6962), .A2(n11560), .ZN(n11713) );
  NAND2_X1 U8797 ( .A1(n11559), .A2(n11558), .ZN(n6962) );
  OAI22_X1 U8798 ( .A1(n15161), .A2(n6888), .B1(P2_ADDR_REG_11__SCAN_IN), .B2(
        n6887), .ZN(n11709) );
  NOR2_X1 U8799 ( .A1(n15159), .A2(n6889), .ZN(n6888) );
  INV_X1 U8800 ( .A(n15159), .ZN(n6887) );
  AOI21_X1 U8801 ( .B1(n6963), .B2(n6965), .A(n6961), .ZN(n6960) );
  INV_X1 U8802 ( .A(n11714), .ZN(n6961) );
  OR2_X1 U8803 ( .A1(n11848), .A2(n11847), .ZN(n12098) );
  XNOR2_X1 U8804 ( .A(n15192), .B(n15191), .ZN(n15190) );
  NAND2_X1 U8805 ( .A1(n15177), .A2(n15176), .ZN(n6886) );
  NAND2_X1 U8806 ( .A1(n12436), .A2(n12320), .ZN(n12321) );
  XNOR2_X1 U8807 ( .A(n10687), .B(n10836), .ZN(n10605) );
  AOI21_X1 U8808 ( .B1(n7633), .B2(n12319), .A(n12350), .ZN(n7632) );
  INV_X1 U8809 ( .A(n7648), .ZN(n12390) );
  AND2_X1 U8810 ( .A1(n7327), .A2(n12682), .ZN(n7324) );
  AOI21_X1 U8811 ( .B1(n7327), .B2(n12400), .A(n12434), .ZN(n7322) );
  NAND2_X1 U8812 ( .A1(n8292), .A2(n8291), .ZN(n12406) );
  CLKBUF_X1 U8813 ( .A(n11190), .Z(n6621) );
  OAI21_X1 U8814 ( .B1(n11772), .B2(n11721), .A(n11720), .ZN(n6896) );
  AND2_X1 U8815 ( .A1(n11771), .A2(n11955), .ZN(n11721) );
  NAND2_X1 U8816 ( .A1(n7648), .A2(n7330), .ZN(n6912) );
  AND2_X1 U8817 ( .A1(n8319), .A2(n8318), .ZN(n12449) );
  AND2_X1 U8818 ( .A1(n8393), .A2(n8360), .ZN(n12355) );
  INV_X1 U8819 ( .A(n12357), .ZN(n12637) );
  INV_X1 U8820 ( .A(n12656), .ZN(n9352) );
  INV_X1 U8821 ( .A(n12718), .ZN(n12694) );
  INV_X1 U8822 ( .A(n12430), .ZN(n12732) );
  NAND2_X1 U8823 ( .A1(n8386), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8005) );
  NAND4_X2 U8824 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n12460)
         );
  OR2_X1 U8825 ( .A1(n8390), .A2(n7959), .ZN(n7967) );
  OR2_X1 U8826 ( .A1(n8372), .A2(n7907), .ZN(n7910) );
  OR2_X1 U8827 ( .A1(n8372), .A2(n10536), .ZN(n7899) );
  OAI21_X1 U8828 ( .B1(n10548), .B2(n10549), .A(n7274), .ZN(n10642) );
  AOI21_X1 U8829 ( .B1(n6432), .B2(n10635), .A(n10882), .ZN(n10636) );
  NAND2_X1 U8830 ( .A1(n10636), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U8831 ( .A1(n7266), .A2(n7269), .ZN(n10881) );
  NAND2_X1 U8832 ( .A1(n10548), .A2(n7267), .ZN(n7266) );
  XNOR2_X1 U8833 ( .A(n7376), .B(n11486), .ZN(n11528) );
  NAND2_X1 U8834 ( .A1(n7263), .A2(n11471), .ZN(n7260) );
  XNOR2_X1 U8835 ( .A(n12000), .B(n12012), .ZN(n12002) );
  NAND2_X1 U8836 ( .A1(n6936), .A2(n6935), .ZN(n12462) );
  NAND2_X1 U8837 ( .A1(n12000), .A2(n6759), .ZN(n6756) );
  OAI21_X1 U8838 ( .B1(n12542), .B2(n12835), .A(n6743), .ZN(n12544) );
  NAND2_X1 U8839 ( .A1(n6740), .A2(n6739), .ZN(n12554) );
  AOI21_X1 U8840 ( .B1(n6743), .B2(n12835), .A(n6741), .ZN(n6739) );
  NOR2_X1 U8841 ( .A1(n12532), .A2(n6418), .ZN(n12559) );
  NAND2_X1 U8842 ( .A1(n6956), .A2(n7678), .ZN(n6952) );
  AND2_X1 U8843 ( .A1(n7677), .A2(n6957), .ZN(n6956) );
  AND2_X1 U8844 ( .A1(n7680), .A2(n7385), .ZN(n6957) );
  NAND2_X1 U8845 ( .A1(n6955), .A2(n12576), .ZN(n6951) );
  OR2_X1 U8846 ( .A1(n7678), .A2(n7385), .ZN(n6950) );
  NAND2_X1 U8847 ( .A1(n12532), .A2(n7256), .ZN(n7254) );
  NAND2_X1 U8848 ( .A1(n7747), .A2(n7748), .ZN(n12626) );
  AOI21_X1 U8849 ( .B1(n12624), .B2(n12784), .A(n12623), .ZN(n12795) );
  NAND2_X1 U8850 ( .A1(n12622), .A2(n12621), .ZN(n12623) );
  XNOR2_X1 U8851 ( .A(n12618), .B(n12625), .ZN(n12624) );
  NAND2_X1 U8852 ( .A1(n6659), .A2(n6657), .ZN(n12800) );
  INV_X1 U8853 ( .A(n6658), .ZN(n6657) );
  NAND2_X1 U8854 ( .A1(n6660), .A2(n12784), .ZN(n6659) );
  OAI22_X1 U8855 ( .A1(n12645), .A2(n15469), .B1(n12644), .B2(n15467), .ZN(
        n6658) );
  NAND2_X1 U8856 ( .A1(n7729), .A2(n8514), .ZN(n12664) );
  NAND2_X1 U8857 ( .A1(n7734), .A2(n7732), .ZN(n7729) );
  AND2_X1 U8858 ( .A1(n7231), .A2(n7232), .ZN(n12667) );
  NAND2_X1 U8859 ( .A1(n7762), .A2(n8420), .ZN(n12740) );
  AND3_X1 U8860 ( .A1(n7958), .A2(n7957), .A3(n7956), .ZN(n11093) );
  INV_X1 U8861 ( .A(n12790), .ZN(n12741) );
  INV_X1 U8862 ( .A(n15472), .ZN(n15493) );
  AOI21_X1 U8863 ( .B1(n12206), .B2(n8381), .A(n6583), .ZN(n12848) );
  INV_X1 U8864 ( .A(n12449), .ZN(n12856) );
  NAND2_X1 U8865 ( .A1(n12646), .A2(n8527), .ZN(n12634) );
  INV_X1 U8866 ( .A(n12406), .ZN(n12867) );
  NAND2_X1 U8867 ( .A1(n7734), .A2(n7737), .ZN(n12677) );
  NAND2_X1 U8868 ( .A1(n7739), .A2(n7740), .ZN(n12690) );
  OR2_X1 U8869 ( .A1(n12701), .A2(n12702), .ZN(n7739) );
  NAND2_X1 U8870 ( .A1(n8234), .A2(n8233), .ZN(n12884) );
  NAND2_X1 U8871 ( .A1(n12823), .A2(n8418), .ZN(n12723) );
  NAND2_X1 U8872 ( .A1(n8174), .A2(n8173), .ZN(n12902) );
  NAND2_X1 U8873 ( .A1(n7209), .A2(n7208), .ZN(n12768) );
  NAND2_X1 U8874 ( .A1(n7210), .A2(n6416), .ZN(n7209) );
  NAND2_X1 U8875 ( .A1(n7212), .A2(n7216), .ZN(n12780) );
  NAND2_X1 U8876 ( .A1(n12070), .A2(n8124), .ZN(n7179) );
  NAND2_X1 U8877 ( .A1(n7851), .A2(n7852), .ZN(n12068) );
  INV_X1 U8878 ( .A(n11909), .ZN(n11966) );
  NAND2_X1 U8879 ( .A1(n11598), .A2(n8470), .ZN(n11950) );
  NAND2_X1 U8880 ( .A1(n8079), .A2(n8078), .ZN(n11787) );
  NAND2_X1 U8881 ( .A1(n7759), .A2(n8051), .ZN(n11368) );
  NAND2_X1 U8882 ( .A1(n11348), .A2(n8050), .ZN(n7759) );
  AND2_X1 U8883 ( .A1(n10124), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12922) );
  INV_X1 U8884 ( .A(n7568), .ZN(n7567) );
  OAI21_X1 U8885 ( .B1(n7575), .B2(n7573), .A(n7569), .ZN(n7568) );
  XNOR2_X1 U8886 ( .A(n8352), .B(n8342), .ZN(n12123) );
  OAI21_X1 U8887 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(n8341) );
  INV_X1 U8888 ( .A(SI_26_), .ZN(n12942) );
  NAND2_X1 U8889 ( .A1(n7580), .A2(n8300), .ZN(n8315) );
  NAND2_X1 U8890 ( .A1(n8290), .A2(n15647), .ZN(n7580) );
  NAND2_X1 U8891 ( .A1(n6827), .A2(n8274), .ZN(n8287) );
  NAND2_X1 U8892 ( .A1(n7557), .A2(n7555), .ZN(n6827) );
  NAND2_X1 U8893 ( .A1(n7557), .A2(n8262), .ZN(n8272) );
  OAI21_X1 U8894 ( .B1(n8416), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8417) );
  INV_X1 U8895 ( .A(SI_20_), .ZN(n11363) );
  NAND2_X1 U8896 ( .A1(n8399), .A2(n8416), .ZN(n11362) );
  OAI21_X1 U8897 ( .B1(n7560), .B2(n6566), .A(n6834), .ZN(n8230) );
  NAND2_X1 U8898 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n7656) );
  NOR2_X1 U8899 ( .A1(n7655), .A2(n7654), .ZN(n7653) );
  NOR2_X1 U8900 ( .A1(n8586), .A2(n8215), .ZN(n7657) );
  INV_X1 U8901 ( .A(SI_18_), .ZN(n10844) );
  NAND2_X1 U8902 ( .A1(n7560), .A2(n7558), .ZN(n8212) );
  NAND2_X1 U8903 ( .A1(n8181), .A2(n8180), .ZN(n8197) );
  INV_X1 U8904 ( .A(SI_15_), .ZN(n10477) );
  INV_X1 U8905 ( .A(SI_14_), .ZN(n10271) );
  NAND2_X1 U8906 ( .A1(n8127), .A2(n8126), .ZN(n8130) );
  INV_X1 U8907 ( .A(SI_12_), .ZN(n9999) );
  NAND2_X1 U8908 ( .A1(n7587), .A2(n7585), .ZN(n8107) );
  NAND2_X1 U8909 ( .A1(n7587), .A2(n8089), .ZN(n8094) );
  INV_X1 U8910 ( .A(SI_11_), .ZN(n9991) );
  INV_X1 U8911 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U8912 ( .A1(n7551), .A2(n8027), .ZN(n8035) );
  NAND2_X1 U8913 ( .A1(n8026), .A2(n8025), .ZN(n7551) );
  NAND2_X1 U8914 ( .A1(n7991), .A2(n7990), .ZN(n8007) );
  NAND2_X1 U8915 ( .A1(n6819), .A2(n7951), .ZN(n7971) );
  NAND2_X1 U8916 ( .A1(n7932), .A2(n7933), .ZN(n7548) );
  NAND2_X1 U8917 ( .A1(n7931), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6750) );
  NOR2_X1 U8918 ( .A1(n7434), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12929) );
  AOI22_X1 U8919 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n7382), .B1(n7381), .B2(
        n7380), .ZN(n7379) );
  AND2_X1 U8920 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7382) );
  INV_X1 U8921 ( .A(n11491), .ZN(n10092) );
  NAND2_X1 U8922 ( .A1(n13068), .A2(n12265), .ZN(n12952) );
  NAND2_X1 U8923 ( .A1(n12116), .A2(n7605), .ZN(n12961) );
  AND2_X1 U8924 ( .A1(n11740), .A2(n11739), .ZN(n11983) );
  NAND2_X1 U8925 ( .A1(n7593), .A2(n7594), .ZN(n12985) );
  NAND2_X1 U8926 ( .A1(n9734), .A2(n13262), .ZN(n9737) );
  NAND2_X1 U8927 ( .A1(n13039), .A2(n12239), .ZN(n12991) );
  AND2_X1 U8928 ( .A1(n11026), .A2(n10859), .ZN(n6989) );
  INV_X1 U8929 ( .A(n12272), .ZN(n10917) );
  INV_X1 U8930 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U8931 ( .A1(n12116), .A2(n12115), .ZN(n12209) );
  NAND2_X1 U8932 ( .A1(n13023), .A2(n12230), .ZN(n13059) );
  NAND2_X1 U8933 ( .A1(n11213), .A2(n11212), .ZN(n11221) );
  INV_X1 U8934 ( .A(n13089), .ZN(n13042) );
  NAND2_X1 U8935 ( .A1(n6725), .A2(n6724), .ZN(n13324) );
  NOR2_X1 U8936 ( .A1(n13334), .A2(n13323), .ZN(n6724) );
  XNOR2_X1 U8937 ( .A(n6726), .B(n13433), .ZN(n6725) );
  INV_X1 U8938 ( .A(n9859), .ZN(n13331) );
  NAND2_X1 U8939 ( .A1(n9869), .A2(n9868), .ZN(n13456) );
  NAND2_X1 U8940 ( .A1(n9794), .A2(n9793), .ZN(n13561) );
  NAND2_X1 U8941 ( .A1(n9769), .A2(n9768), .ZN(n13599) );
  NAND2_X1 U8942 ( .A1(n9503), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6904) );
  CLKBUF_X1 U8943 ( .A(n13355), .Z(n7148) );
  NAND2_X1 U8944 ( .A1(n13385), .A2(n13384), .ZN(n10106) );
  NAND2_X1 U8945 ( .A1(n15345), .A2(n15346), .ZN(n15344) );
  NAND2_X1 U8946 ( .A1(n10262), .A2(n10084), .ZN(n15360) );
  NAND2_X1 U8947 ( .A1(n15360), .A2(n15361), .ZN(n15359) );
  NAND2_X1 U8948 ( .A1(n6629), .A2(n6630), .ZN(n15373) );
  OR2_X1 U8949 ( .A1(n10262), .A2(n6632), .ZN(n6629) );
  NAND2_X1 U8950 ( .A1(n15371), .A2(n15372), .ZN(n15370) );
  NAND2_X1 U8951 ( .A1(n10591), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U8952 ( .A1(n11140), .A2(n11139), .ZN(n11144) );
  NAND2_X1 U8953 ( .A1(n13409), .A2(n13408), .ZN(n15408) );
  INV_X1 U8954 ( .A(n13755), .ZN(n13752) );
  AND2_X1 U8955 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  OR2_X1 U8956 ( .A1(n13232), .A2(n13676), .ZN(n9871) );
  OAI21_X1 U8957 ( .B1(n13572), .B2(n7333), .A(n7332), .ZN(n13501) );
  NAND2_X1 U8958 ( .A1(n7334), .A2(n7338), .ZN(n13516) );
  NAND2_X1 U8959 ( .A1(n13572), .A2(n7339), .ZN(n7334) );
  AND2_X1 U8960 ( .A1(n7511), .A2(n7510), .ZN(n13512) );
  NAND2_X1 U8961 ( .A1(n7504), .A2(n9855), .ZN(n13525) );
  INV_X1 U8962 ( .A(n13571), .ZN(n7533) );
  INV_X1 U8963 ( .A(n13572), .ZN(n7534) );
  NAND2_X1 U8964 ( .A1(n7516), .A2(n9849), .ZN(n13612) );
  OR2_X1 U8965 ( .A1(n13627), .A2(n6519), .ZN(n7516) );
  NAND2_X1 U8966 ( .A1(n9715), .A2(n9714), .ZN(n13819) );
  NAND2_X1 U8967 ( .A1(n7343), .A2(n9698), .ZN(n13668) );
  NAND2_X1 U8968 ( .A1(n7347), .A2(n7346), .ZN(n7343) );
  NAND2_X1 U8969 ( .A1(n13704), .A2(n9683), .ZN(n7347) );
  OAI21_X1 U8970 ( .B1(n13704), .B2(n6451), .A(n9683), .ZN(n13673) );
  NAND2_X1 U8971 ( .A1(n7527), .A2(n7525), .ZN(n13737) );
  NAND2_X1 U8972 ( .A1(n7526), .A2(n6413), .ZN(n7525) );
  OAI21_X1 U8973 ( .B1(n11860), .B2(n9644), .A(n9643), .ZN(n12050) );
  NAND2_X1 U8974 ( .A1(n11244), .A2(n7490), .ZN(n11298) );
  AOI21_X1 U8975 ( .B1(n13262), .B2(n9971), .A(n7104), .ZN(n7103) );
  OAI21_X1 U8976 ( .B1(n7079), .B2(n6773), .A(n10976), .ZN(n10708) );
  NAND2_X2 U8977 ( .A1(n10984), .A2(n13683), .ZN(n13687) );
  OR2_X1 U8978 ( .A1(n10984), .A2(n13433), .ZN(n13549) );
  AND2_X1 U8979 ( .A1(n13687), .A2(n10990), .ZN(n13649) );
  AND2_X1 U8980 ( .A1(n7171), .A2(n11045), .ZN(n11046) );
  INV_X1 U8981 ( .A(n13437), .ZN(n13859) );
  NAND2_X1 U8982 ( .A1(n7075), .A2(n7074), .ZN(n13870) );
  INV_X1 U8983 ( .A(n13770), .ZN(n7074) );
  NOR2_X1 U8984 ( .A1(n13769), .A2(n7076), .ZN(n7075) );
  OAI21_X1 U8985 ( .B1(n13772), .B2(n13855), .A(n7077), .ZN(n7076) );
  NAND2_X1 U8986 ( .A1(n6618), .A2(n6485), .ZN(n13878) );
  NAND2_X1 U8987 ( .A1(n13784), .A2(n13835), .ZN(n6618) );
  AND2_X1 U8988 ( .A1(n13785), .A2(n13787), .ZN(n6617) );
  INV_X1 U8989 ( .A(n13180), .ZN(n13895) );
  INV_X1 U8990 ( .A(n13900), .ZN(n13881) );
  OAI21_X1 U8991 ( .B1(n9895), .B2(n9907), .A(n9894), .ZN(n15415) );
  AND2_X1 U8992 ( .A1(n10855), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15416) );
  INV_X1 U8993 ( .A(n9481), .ZN(n12204) );
  INV_X1 U8994 ( .A(n9907), .ZN(n11949) );
  NAND2_X1 U8995 ( .A1(n9891), .A2(n9890), .ZN(n13918) );
  XNOR2_X1 U8996 ( .A(n9879), .B(n9878), .ZN(n11997) );
  INV_X1 U8997 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9878) );
  OAI21_X1 U8998 ( .B1(n9910), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9879) );
  INV_X1 U8999 ( .A(n10800), .ZN(n13104) );
  INV_X1 U9000 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n15584) );
  INV_X1 U9001 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10760) );
  INV_X1 U9002 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10618) );
  INV_X1 U9003 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10827) );
  INV_X1 U9004 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n15618) );
  INV_X1 U9005 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9975) );
  NOR2_X1 U9006 ( .A1(n7434), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13910) );
  INV_X1 U9007 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9977) );
  INV_X1 U9008 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9927) );
  NAND2_X1 U9009 ( .A1(n9518), .A2(n9532), .ZN(n13372) );
  AND2_X1 U9010 ( .A1(n6647), .A2(n6645), .ZN(n6644) );
  NAND2_X1 U9011 ( .A1(n13905), .A2(n6646), .ZN(n6645) );
  AND4_X1 U9012 ( .A1(n8998), .A2(n8997), .A3(n8996), .A4(n8995), .ZN(n15074)
         );
  INV_X1 U9013 ( .A(n14072), .ZN(n7454) );
  NAND2_X1 U9014 ( .A1(n6785), .A2(n6483), .ZN(n7455) );
  NAND2_X1 U9015 ( .A1(n6790), .A2(n6791), .ZN(n14248) );
  OR2_X1 U9016 ( .A1(n14101), .A2(n6793), .ZN(n6790) );
  NAND2_X1 U9017 ( .A1(n9121), .A2(n9120), .ZN(n15009) );
  NAND2_X1 U9018 ( .A1(n7477), .A2(n10898), .ZN(n14091) );
  AND2_X1 U9019 ( .A1(n9097), .A2(n9096), .ZN(n14848) );
  NAND2_X1 U9020 ( .A1(n7480), .A2(n7481), .ZN(n14100) );
  AND2_X1 U9021 ( .A1(n13925), .A2(n13924), .ZN(n14122) );
  AND2_X1 U9022 ( .A1(n7487), .A2(n7485), .ZN(n12161) );
  NAND2_X1 U9023 ( .A1(n7487), .A2(n7488), .ZN(n11827) );
  AND2_X1 U9024 ( .A1(n7462), .A2(n6468), .ZN(n14140) );
  AND3_X1 U9025 ( .A1(n9049), .A2(n9048), .A3(n9047), .ZN(n15054) );
  NAND2_X1 U9026 ( .A1(n14101), .A2(n13995), .ZN(n14226) );
  NAND2_X1 U9027 ( .A1(n10658), .A2(n10657), .ZN(n6782) );
  AND2_X1 U9028 ( .A1(n9070), .A2(n9069), .ZN(n15043) );
  NAND2_X1 U9029 ( .A1(n14269), .A2(n14270), .ZN(n14268) );
  NAND2_X1 U9030 ( .A1(n14195), .A2(n13981), .ZN(n14269) );
  AOI21_X1 U9031 ( .B1(n6815), .B2(n6817), .A(n6813), .ZN(n6812) );
  NAND2_X1 U9032 ( .A1(n11445), .A2(n6807), .ZN(n6809) );
  NAND2_X1 U9033 ( .A1(n6811), .A2(n11449), .ZN(n6817) );
  NAND2_X1 U9034 ( .A1(n14158), .A2(n14048), .ZN(n14279) );
  INV_X1 U9035 ( .A(n14281), .ZN(n14302) );
  NAND2_X1 U9036 ( .A1(n7395), .A2(n7618), .ZN(n14523) );
  AND2_X1 U9037 ( .A1(n14307), .A2(n14476), .ZN(n14554) );
  OR2_X1 U9038 ( .A1(n10301), .A2(P1_U3086), .ZN(n14558) );
  NAND2_X1 U9039 ( .A1(n9179), .A2(n9178), .ZN(n14567) );
  NAND2_X1 U9040 ( .A1(n9142), .A2(n9141), .ZN(n14570) );
  NAND2_X1 U9041 ( .A1(n9112), .A2(n9111), .ZN(n14572) );
  INV_X1 U9042 ( .A(n15027), .ZN(n14573) );
  INV_X1 U9043 ( .A(n14848), .ZN(n15035) );
  INV_X1 U9044 ( .A(n15054), .ZN(n15034) );
  AND4_X1 U9045 ( .A1(n8978), .A2(n8977), .A3(n8976), .A4(n8975), .ZN(n15082)
         );
  INV_X1 U9046 ( .A(n11933), .ZN(n14575) );
  NAND2_X1 U9047 ( .A1(n14453), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U9048 ( .A1(n9209), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8735) );
  OR2_X1 U9049 ( .A1(n8759), .A2(n11328), .ZN(n8734) );
  INV_X1 U9050 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U9051 ( .A1(n14671), .A2(n15217), .ZN(n7142) );
  OR2_X1 U9052 ( .A1(n12137), .A2(n7864), .ZN(n9278) );
  XNOR2_X1 U9053 ( .A(n14734), .B(n14733), .ZN(n7373) );
  NAND2_X1 U9054 ( .A1(n9132), .A2(n9131), .ZN(n15006) );
  NAND2_X1 U9055 ( .A1(n7810), .A2(n9267), .ZN(n14763) );
  NAND2_X1 U9056 ( .A1(n14856), .A2(n7439), .ZN(n14800) );
  INV_X1 U9057 ( .A(n7020), .ZN(n14867) );
  AOI21_X1 U9058 ( .B1(n14931), .B2(n7022), .A(n7021), .ZN(n7020) );
  NAND2_X1 U9059 ( .A1(n7051), .A2(n9261), .ZN(n14854) );
  NAND2_X1 U9060 ( .A1(n7059), .A2(n7058), .ZN(n7051) );
  NAND2_X1 U9061 ( .A1(n7059), .A2(n9260), .ZN(n14871) );
  AND3_X1 U9062 ( .A1(n9011), .A2(n9010), .A3(n9009), .ZN(n15061) );
  NAND2_X1 U9063 ( .A1(n14959), .A2(n9251), .ZN(n7793) );
  INV_X1 U9064 ( .A(n7766), .ZN(n7768) );
  NOR2_X1 U9065 ( .A1(n7770), .A2(n7769), .ZN(n11758) );
  INV_X1 U9066 ( .A(n8887), .ZN(n7769) );
  INV_X1 U9067 ( .A(n11644), .ZN(n7770) );
  NOR2_X1 U9068 ( .A1(n14524), .A2(n7773), .ZN(n7772) );
  INV_X1 U9069 ( .A(n7777), .ZN(n7773) );
  NAND2_X1 U9070 ( .A1(n7774), .A2(n7777), .ZN(n11378) );
  NAND2_X1 U9071 ( .A1(n8834), .A2(n8833), .ZN(n15228) );
  OR2_X1 U9072 ( .A1(n15269), .A2(n15277), .ZN(n14906) );
  OR2_X1 U9073 ( .A1(n14693), .A2(n14672), .ZN(n14974) );
  INV_X1 U9074 ( .A(n11317), .ZN(n11503) );
  NAND2_X1 U9075 ( .A1(n10786), .A2(n14318), .ZN(n11501) );
  NOR2_X1 U9076 ( .A1(n14989), .A2(n14988), .ZN(n14990) );
  NAND2_X1 U9077 ( .A1(n14987), .A2(n14986), .ZN(n14988) );
  NAND2_X1 U9078 ( .A1(n14985), .A2(n15315), .ZN(n14986) );
  NAND2_X1 U9079 ( .A1(n10000), .A2(n10278), .ZN(n15270) );
  INV_X1 U9080 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15135) );
  XNOR2_X1 U9081 ( .A(n13261), .B(n13260), .ZN(n15140) );
  NAND2_X1 U9082 ( .A1(n7427), .A2(n13258), .ZN(n14464) );
  NAND2_X1 U9083 ( .A1(n12202), .A2(n12201), .ZN(n7427) );
  INV_X1 U9084 ( .A(n7813), .ZN(n7393) );
  NAND2_X1 U9085 ( .A1(n8629), .A2(n7812), .ZN(n8716) );
  INV_X1 U9086 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11945) );
  INV_X1 U9087 ( .A(n9309), .ZN(n15149) );
  INV_X1 U9088 ( .A(n9308), .ZN(n11998) );
  OR2_X1 U9089 ( .A1(n9773), .A2(n7434), .ZN(n9105) );
  NAND2_X1 U9090 ( .A1(n9304), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9221) );
  INV_X1 U9091 ( .A(n9285), .ZN(n14307) );
  INV_X1 U9092 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11374) );
  NAND2_X1 U9093 ( .A1(n6805), .A2(n9059), .ZN(n9218) );
  INV_X1 U9094 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n15608) );
  INV_X1 U9095 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10569) );
  INV_X1 U9096 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10539) );
  XNOR2_X1 U9097 ( .A(n8970), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11801) );
  AND2_X1 U9098 ( .A1(n8898), .A2(n8987), .ZN(n10559) );
  INV_X1 U9099 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U9100 ( .A1(n8838), .A2(n8664), .ZN(n8853) );
  INV_X1 U9101 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9994) );
  NAND2_X2 U9102 ( .A1(n8748), .A2(n8856), .ZN(n14605) );
  NAND2_X1 U9103 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8731) );
  CLKBUF_X1 U9104 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n7069) );
  NAND2_X1 U9105 ( .A1(n6884), .A2(n6882), .ZN(n10503) );
  NOR2_X1 U9106 ( .A1(n6883), .A2(n10501), .ZN(n6882) );
  INV_X1 U9107 ( .A(n10487), .ZN(n6883) );
  NAND2_X1 U9108 ( .A1(n6884), .A2(n10487), .ZN(n10502) );
  AND2_X1 U9109 ( .A1(n10931), .A2(n10930), .ZN(n10937) );
  NAND2_X1 U9110 ( .A1(n10940), .A2(n10941), .ZN(n11547) );
  INV_X1 U9111 ( .A(n10940), .ZN(n10938) );
  XNOR2_X1 U9112 ( .A(n11709), .B(n11707), .ZN(n11706) );
  NAND2_X1 U9113 ( .A1(n12103), .A2(n12102), .ZN(n15166) );
  NAND2_X1 U9114 ( .A1(n6892), .A2(n6890), .ZN(n12103) );
  NOR2_X1 U9115 ( .A1(n12100), .A2(n6891), .ZN(n6890) );
  INV_X1 U9116 ( .A(n12096), .ZN(n6891) );
  NAND2_X1 U9117 ( .A1(n15166), .A2(n15165), .ZN(n15175) );
  NAND2_X1 U9118 ( .A1(n11308), .A2(n11307), .ZN(n11718) );
  NAND2_X1 U9119 ( .A1(n10690), .A2(n10689), .ZN(n10696) );
  INV_X1 U9120 ( .A(n6747), .ZN(n10876) );
  NAND2_X1 U9121 ( .A1(n7679), .A2(n12536), .ZN(n12514) );
  NAND2_X1 U9122 ( .A1(n7242), .A2(n12491), .ZN(n7241) );
  OR2_X1 U9123 ( .A1(n12589), .A2(n7672), .ZN(n7246) );
  MUX2_X1 U9124 ( .A(n12612), .B(n12611), .S(n15472), .Z(n12616) );
  OAI22_X1 U9125 ( .A1(n12187), .A2(n12821), .B1(n15514), .B2(n9430), .ZN(
        n9431) );
  INV_X1 U9126 ( .A(n7754), .ZN(n7752) );
  NAND2_X1 U9127 ( .A1(n6993), .A2(n6999), .ZN(n11393) );
  NOR2_X1 U9128 ( .A1(n10861), .A2(n10860), .ZN(n11027) );
  XNOR2_X1 U9129 ( .A(n6987), .B(n12275), .ZN(n12288) );
  AOI21_X1 U9130 ( .B1(n6636), .B2(n13433), .A(n6634), .ZN(n6633) );
  NAND2_X1 U9131 ( .A1(n6635), .A2(n13435), .ZN(n6634) );
  INV_X1 U9132 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U9133 ( .A1(n15452), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7348) );
  INV_X1 U9134 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U9135 ( .A1(n6712), .A2(n14281), .ZN(n14063) );
  OAI21_X1 U9136 ( .B1(n14716), .B2(n15260), .A(n7156), .ZN(n7155) );
  AOI21_X1 U9137 ( .B1(n14715), .B2(n15266), .A(n14714), .ZN(n7156) );
  NOR2_X1 U9138 ( .A1(n15327), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7799) );
  AND2_X1 U9139 ( .A1(n14716), .A2(n6476), .ZN(n7795) );
  NOR2_X1 U9140 ( .A1(n6403), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7796) );
  AND2_X1 U9141 ( .A1(n14716), .A2(n7797), .ZN(n7794) );
  NOR2_X1 U9142 ( .A1(n7798), .A2(n15323), .ZN(n7797) );
  NAND2_X1 U9143 ( .A1(n7123), .A2(n6581), .ZN(P1_U3522) );
  NAND2_X1 U9144 ( .A1(n15117), .A2(n6403), .ZN(n7123) );
  NAND2_X1 U9145 ( .A1(n7131), .A2(n6582), .ZN(P1_U3518) );
  INV_X1 U9146 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n7130) );
  AOI21_X1 U9147 ( .B1(n15188), .B2(n15189), .A(n6516), .ZN(n15198) );
  AND2_X2 U9148 ( .A1(n13284), .A2(n15422), .ZN(n6425) );
  OR2_X1 U9149 ( .A1(n7367), .A2(n7771), .ZN(n6411) );
  INV_X2 U9150 ( .A(n10518), .ZN(n11174) );
  INV_X2 U9151 ( .A(n13099), .ZN(n9814) );
  AND2_X1 U9152 ( .A1(n8980), .A2(n8682), .ZN(n6412) );
  OR2_X1 U9153 ( .A1(n13846), .A2(n13721), .ZN(n6413) );
  AND2_X1 U9154 ( .A1(n12203), .A2(n12290), .ZN(n8794) );
  NAND2_X1 U9155 ( .A1(n6454), .A2(n12541), .ZN(n7679) );
  INV_X1 U9156 ( .A(n7697), .ZN(n13630) );
  INV_X1 U9157 ( .A(n13667), .ZN(n7345) );
  NAND2_X1 U9158 ( .A1(n6912), .A2(n7329), .ZN(n12426) );
  AND2_X1 U9159 ( .A1(n6517), .A2(n6978), .ZN(n6414) );
  NAND3_X1 U9160 ( .A1(n6936), .A2(n6579), .A3(n6935), .ZN(n6415) );
  NOR2_X1 U9161 ( .A1(n7217), .A2(n7211), .ZN(n6416) );
  NAND2_X1 U9162 ( .A1(n8548), .A2(n12450), .ZN(n7543) );
  NAND2_X1 U9163 ( .A1(n9446), .A2(n9441), .ZN(n6417) );
  XNOR2_X1 U9164 ( .A(n15006), .B(n14570), .ZN(n14545) );
  INV_X1 U9165 ( .A(n14545), .ZN(n7027) );
  AND2_X1 U9166 ( .A1(n12533), .A2(n12541), .ZN(n6418) );
  AND2_X1 U9167 ( .A1(n7669), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6419) );
  AND2_X1 U9168 ( .A1(n7897), .A2(n7196), .ZN(n6420) );
  AND3_X1 U9169 ( .A1(n13526), .A2(n6718), .A3(n6717), .ZN(n6421) );
  INV_X1 U9170 ( .A(n12463), .ZN(n12494) );
  AND2_X1 U9171 ( .A1(n7384), .A2(n6733), .ZN(n6422) );
  AND2_X1 U9172 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n6423) );
  AND2_X1 U9173 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n6424) );
  AND3_X1 U9174 ( .A1(n7679), .A2(n12536), .A3(P3_REG2_REG_15__SCAN_IN), .ZN(
        n6426) );
  NAND2_X1 U9175 ( .A1(n9169), .A2(n9168), .ZN(n14985) );
  INV_X1 U9176 ( .A(n14985), .ZN(n7451) );
  INV_X1 U9177 ( .A(n12782), .ZN(n12383) );
  INV_X1 U9178 ( .A(n9036), .ZN(n7771) );
  OR2_X1 U9179 ( .A1(n12856), .A2(n12645), .ZN(n8532) );
  AND2_X1 U9180 ( .A1(n7581), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6427) );
  OR2_X1 U9181 ( .A1(n10640), .A2(n11096), .ZN(n6428) );
  AND2_X1 U9182 ( .A1(n12463), .A2(n12518), .ZN(n6429) );
  NOR2_X1 U9183 ( .A1(n13809), .A2(n13192), .ZN(n6430) );
  AND2_X1 U9184 ( .A1(n6693), .A2(n13197), .ZN(n6431) );
  AND2_X1 U9185 ( .A1(n6552), .A2(n6934), .ZN(n6432) );
  NAND2_X1 U9186 ( .A1(n7269), .A2(n7265), .ZN(n7264) );
  INV_X1 U9187 ( .A(n7264), .ZN(n7263) );
  NAND2_X1 U9188 ( .A1(n8087), .A2(n8468), .ZN(n6433) );
  AND2_X1 U9189 ( .A1(n7286), .A2(n8447), .ZN(n6434) );
  AND2_X1 U9190 ( .A1(n7660), .A2(n11486), .ZN(n11536) );
  INV_X1 U9191 ( .A(n14424), .ZN(n7621) );
  NOR2_X1 U9192 ( .A1(n12902), .A2(n12770), .ZN(n6435) );
  OR2_X1 U9193 ( .A1(n13765), .A2(n13289), .ZN(n13453) );
  INV_X1 U9194 ( .A(n12389), .ZN(n7330) );
  NOR2_X1 U9195 ( .A1(n9275), .A2(n9273), .ZN(n6436) );
  INV_X1 U9196 ( .A(n10629), .ZN(n10946) );
  AND2_X1 U9197 ( .A1(n7528), .A2(n9672), .ZN(n6437) );
  AND2_X1 U9198 ( .A1(n8677), .A2(n9999), .ZN(n6438) );
  INV_X1 U9199 ( .A(n13707), .ZN(n6606) );
  AND2_X1 U9200 ( .A1(n8157), .A2(n6703), .ZN(n6439) );
  INV_X1 U9201 ( .A(n12681), .ZN(n12705) );
  AOI21_X1 U9202 ( .B1(n12698), .B2(n8355), .A(n8255), .ZN(n12681) );
  NOR2_X1 U9203 ( .A1(n15510), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6440) );
  AND2_X1 U9204 ( .A1(n6756), .A2(n6758), .ZN(n6441) );
  AND2_X1 U9205 ( .A1(n12537), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6442) );
  INV_X1 U9206 ( .A(n8314), .ZN(n7579) );
  AND2_X1 U9207 ( .A1(n6842), .A2(n8314), .ZN(n6443) );
  AND2_X1 U9208 ( .A1(n6696), .A2(n6695), .ZN(n6444) );
  INV_X2 U9209 ( .A(n8794), .ZN(n9213) );
  CLKBUF_X3 U9210 ( .A(n9503), .Z(n13099) );
  OR2_X1 U9211 ( .A1(n12793), .A2(n12637), .ZN(n6445) );
  XNOR2_X1 U9212 ( .A(n12540), .B(n12531), .ZN(n12542) );
  NAND2_X1 U9213 ( .A1(n14943), .A2(n8963), .ZN(n14931) );
  NAND2_X1 U9214 ( .A1(n12701), .A2(n7735), .ZN(n7734) );
  INV_X1 U9215 ( .A(n12745), .ZN(n7847) );
  INV_X1 U9216 ( .A(n14902), .ZN(n7050) );
  OR3_X1 U9217 ( .A1(n14712), .A2(n14711), .A3(n15289), .ZN(n6446) );
  INV_X1 U9218 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9818) );
  XNOR2_X1 U9219 ( .A(n14850), .B(n15043), .ZN(n14399) );
  NAND2_X1 U9220 ( .A1(n9391), .A2(n8339), .ZN(n12625) );
  XNOR2_X1 U9221 ( .A(n14994), .B(n14161), .ZN(n14733) );
  INV_X1 U9222 ( .A(n14733), .ZN(n7782) );
  NAND2_X1 U9223 ( .A1(n7462), .A2(n7461), .ZN(n14138) );
  NAND2_X1 U9224 ( .A1(n13934), .A2(n13933), .ZN(n14064) );
  INV_X1 U9225 ( .A(n12055), .ZN(n6920) );
  OR2_X1 U9226 ( .A1(n13337), .A2(n13771), .ZN(n6447) );
  AND2_X1 U9227 ( .A1(n11056), .A2(n13133), .ZN(n6448) );
  AND2_X1 U9228 ( .A1(n9365), .A2(n9367), .ZN(n6449) );
  OAI22_X1 U9229 ( .A1(n12343), .A2(n7644), .B1(n12302), .B2(n12430), .ZN(
        n7643) );
  NAND2_X1 U9230 ( .A1(n14825), .A2(n9264), .ZN(n14785) );
  OR2_X1 U9231 ( .A1(n7206), .A2(n6435), .ZN(n6450) );
  AND2_X1 U9232 ( .A1(n13707), .A2(n13724), .ZN(n6451) );
  INV_X1 U9233 ( .A(n13550), .ZN(n6717) );
  OR2_X1 U9234 ( .A1(n9464), .A2(n7139), .ZN(n6452) );
  AOI21_X1 U9235 ( .B1(n14280), .B2(n7474), .A(n7473), .ZN(n7472) );
  INV_X1 U9236 ( .A(n7472), .ZN(n7471) );
  NOR2_X1 U9237 ( .A1(n13880), .A2(n13561), .ZN(n6453) );
  AND2_X1 U9238 ( .A1(n12513), .A2(n12518), .ZN(n6454) );
  AND2_X1 U9239 ( .A1(n6672), .A2(n6671), .ZN(n6455) );
  AND2_X1 U9240 ( .A1(n13449), .A2(n13491), .ZN(n6456) );
  AND2_X1 U9241 ( .A1(n7663), .A2(n11927), .ZN(n12003) );
  XOR2_X1 U9242 ( .A(n13819), .B(n13342), .Z(n6457) );
  AND2_X1 U9243 ( .A1(n13959), .A2(n13958), .ZN(n6458) );
  NAND2_X1 U9244 ( .A1(n13535), .A2(n13339), .ZN(n6459) );
  AND2_X1 U9245 ( .A1(n10111), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6460) );
  INV_X1 U9246 ( .A(n12352), .ZN(n7301) );
  NAND2_X1 U9247 ( .A1(n7923), .A2(n7922), .ZN(n7932) );
  INV_X1 U9248 ( .A(n13809), .ZN(n7696) );
  NAND2_X1 U9249 ( .A1(n9488), .A2(n9487), .ZN(n13771) );
  NOR2_X1 U9250 ( .A1(n14718), .A2(n7807), .ZN(n7806) );
  INV_X1 U9251 ( .A(n7806), .ZN(n7060) );
  INV_X1 U9252 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9462) );
  INV_X1 U9253 ( .A(n14355), .ZN(n7437) );
  NAND2_X1 U9254 ( .A1(n9332), .A2(n9333), .ZN(n6461) );
  NAND2_X1 U9255 ( .A1(n14856), .A2(n7441), .ZN(n7442) );
  OR2_X1 U9256 ( .A1(n15018), .A2(n15289), .ZN(n6462) );
  INV_X1 U9257 ( .A(n11486), .ZN(n11529) );
  NAND2_X1 U9258 ( .A1(n9155), .A2(n9154), .ZN(n14994) );
  INV_X1 U9259 ( .A(n14994), .ZN(n7452) );
  XNOR2_X1 U9260 ( .A(n8029), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11470) );
  AND2_X1 U9261 ( .A1(n6641), .A2(n6640), .ZN(n6463) );
  NAND2_X1 U9262 ( .A1(n9547), .A2(n7103), .ZN(n13126) );
  INV_X1 U9263 ( .A(n13126), .ZN(n7686) );
  INV_X1 U9264 ( .A(n14542), .ZN(n14771) );
  INV_X1 U9265 ( .A(n9058), .ZN(n6805) );
  OR2_X1 U9266 ( .A1(n14217), .A2(n12172), .ZN(n6464) );
  BUF_X1 U9267 ( .A(n9298), .Z(n9299) );
  NAND2_X1 U9268 ( .A1(n7600), .A2(n12262), .ZN(n13067) );
  OR3_X1 U9269 ( .A1(n13473), .A2(n13752), .A3(n7078), .ZN(n6465) );
  AND2_X1 U9270 ( .A1(n14755), .A2(n7452), .ZN(n6466) );
  AND2_X1 U9271 ( .A1(n13880), .A2(n13561), .ZN(n6467) );
  INV_X1 U9272 ( .A(n13147), .ZN(n7715) );
  INV_X1 U9273 ( .A(n7217), .ZN(n7216) );
  NAND2_X1 U9274 ( .A1(n14000), .A2(n14001), .ZN(n6468) );
  NAND2_X1 U9275 ( .A1(n12419), .A2(n12873), .ZN(n7232) );
  INV_X1 U9276 ( .A(n13306), .ZN(n11297) );
  OR2_X1 U9277 ( .A1(n12686), .A2(n12419), .ZN(n8514) );
  AND2_X1 U9278 ( .A1(n9234), .A2(n6406), .ZN(n6469) );
  AND2_X1 U9279 ( .A1(n7609), .A2(n11662), .ZN(n6470) );
  AND2_X1 U9280 ( .A1(n11436), .A2(n12456), .ZN(n6471) );
  NAND2_X1 U9281 ( .A1(n15150), .A2(n8755), .ZN(n14804) );
  AND2_X1 U9282 ( .A1(n6855), .A2(n6853), .ZN(n6472) );
  NAND2_X1 U9283 ( .A1(n8862), .A2(n8861), .ZN(n15316) );
  AND2_X1 U9284 ( .A1(n7484), .A2(n6464), .ZN(n6473) );
  AND3_X1 U9285 ( .A1(n7748), .A2(n8536), .A3(n7749), .ZN(n6474) );
  AND2_X1 U9286 ( .A1(n12242), .A2(n12241), .ZN(n6475) );
  INV_X1 U9287 ( .A(n14850), .ZN(n15038) );
  NAND2_X1 U9288 ( .A1(n9065), .A2(n9064), .ZN(n14850) );
  INV_X1 U9289 ( .A(n15313), .ZN(n14576) );
  AND4_X1 U9290 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n15313)
         );
  AND2_X1 U9291 ( .A1(n7869), .A2(n15327), .ZN(n6476) );
  AND2_X1 U9292 ( .A1(n13425), .A2(n13414), .ZN(n6477) );
  AND2_X1 U9293 ( .A1(n7859), .A2(n7857), .ZN(n6478) );
  NAND2_X1 U9294 ( .A1(n8629), .A2(n8628), .ZN(n9301) );
  OR2_X1 U9295 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15178), .ZN(n6480) );
  AND2_X1 U9296 ( .A1(n11717), .A2(n12455), .ZN(n6481) );
  NOR2_X1 U9297 ( .A1(n10364), .A2(n10365), .ZN(n6482) );
  NOR2_X1 U9298 ( .A1(n13956), .A2(n13955), .ZN(n6483) );
  INV_X1 U9299 ( .A(n13500), .ZN(n6723) );
  OR2_X1 U9300 ( .A1(n8548), .A2(n12450), .ZN(n6484) );
  AND2_X1 U9301 ( .A1(n13786), .A2(n6617), .ZN(n6485) );
  INV_X1 U9302 ( .A(n8909), .ZN(n7767) );
  INV_X1 U9303 ( .A(n9271), .ZN(n7064) );
  NAND2_X1 U9304 ( .A1(n7712), .A2(n13135), .ZN(n6486) );
  AND2_X1 U9305 ( .A1(n13167), .A2(n13166), .ZN(n6487) );
  INV_X1 U9306 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8595) );
  AND2_X1 U9307 ( .A1(n13174), .A2(n13173), .ZN(n6488) );
  NOR2_X1 U9308 ( .A1(n14577), .A2(n15298), .ZN(n6489) );
  INV_X1 U9309 ( .A(SI_10_), .ZN(n9973) );
  INV_X1 U9310 ( .A(n13165), .ZN(n7718) );
  INV_X1 U9311 ( .A(n14158), .ZN(n6714) );
  INV_X1 U9312 ( .A(n14419), .ZN(n7627) );
  INV_X1 U9313 ( .A(n14449), .ZN(n14710) );
  NAND2_X1 U9314 ( .A1(n9191), .A2(n9190), .ZN(n14449) );
  NAND2_X1 U9315 ( .A1(n7678), .A2(n7677), .ZN(n6490) );
  AND2_X1 U9316 ( .A1(n10802), .A2(n6990), .ZN(n6491) );
  INV_X1 U9317 ( .A(n14912), .ZN(n7367) );
  OR2_X1 U9318 ( .A1(n8475), .A2(n10126), .ZN(n6492) );
  INV_X1 U9319 ( .A(n7275), .ZN(n7274) );
  NOR2_X1 U9320 ( .A1(n10387), .A2(n10547), .ZN(n7275) );
  NAND2_X1 U9321 ( .A1(n9470), .A2(n6688), .ZN(n6493) );
  INV_X1 U9322 ( .A(n8664), .ZN(n7520) );
  NAND2_X1 U9323 ( .A1(n7369), .A2(SI_7_), .ZN(n8664) );
  AND2_X1 U9324 ( .A1(n9628), .A2(n6681), .ZN(n6494) );
  AND2_X1 U9325 ( .A1(n7438), .A2(n7437), .ZN(n6495) );
  INV_X1 U9326 ( .A(n11595), .ZN(n8087) );
  AND2_X1 U9327 ( .A1(n7248), .A2(n7254), .ZN(n6496) );
  INV_X1 U9328 ( .A(n9345), .ZN(n7207) );
  AND2_X1 U9329 ( .A1(n6823), .A2(n6822), .ZN(n6497) );
  NAND2_X1 U9330 ( .A1(n14747), .A2(n7450), .ZN(n7453) );
  NAND2_X1 U9331 ( .A1(n7627), .A2(n14420), .ZN(n6498) );
  NAND2_X1 U9332 ( .A1(n7169), .A2(n6696), .ZN(n6499) );
  NOR2_X1 U9333 ( .A1(n15086), .A2(n15091), .ZN(n6500) );
  INV_X1 U9334 ( .A(n7643), .ZN(n7642) );
  AND2_X1 U9335 ( .A1(n13521), .A2(n13338), .ZN(n6501) );
  INV_X1 U9336 ( .A(n9857), .ZN(n7510) );
  INV_X1 U9337 ( .A(n7736), .ZN(n7735) );
  NAND2_X1 U9338 ( .A1(n8509), .A2(n7740), .ZN(n7736) );
  NOR2_X1 U9339 ( .A1(n13986), .A2(n13985), .ZN(n6502) );
  NOR2_X1 U9340 ( .A1(n13792), .A2(n13580), .ZN(n6503) );
  AND2_X1 U9341 ( .A1(n10864), .A2(n10863), .ZN(n6504) );
  INV_X1 U9342 ( .A(n7840), .ZN(n7839) );
  NAND2_X1 U9343 ( .A1(n6445), .A2(n9356), .ZN(n7840) );
  AND2_X1 U9344 ( .A1(n8684), .A2(n10477), .ZN(n6505) );
  INV_X1 U9345 ( .A(n10396), .ZN(n7669) );
  INV_X1 U9346 ( .A(n8702), .ZN(n6874) );
  AND2_X1 U9347 ( .A1(n9102), .A2(n8701), .ZN(n8702) );
  INV_X1 U9348 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9603) );
  INV_X1 U9349 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8880) );
  OR2_X1 U9350 ( .A1(n14491), .A2(n14521), .ZN(n6506) );
  AND2_X1 U9351 ( .A1(n8535), .A2(n12629), .ZN(n6507) );
  INV_X1 U9352 ( .A(n7031), .ZN(n7030) );
  OR2_X1 U9353 ( .A1(n14074), .A2(n6458), .ZN(n6803) );
  AND2_X1 U9354 ( .A1(n9231), .A2(n9232), .ZN(n7883) );
  AND2_X1 U9355 ( .A1(n6737), .A2(n7387), .ZN(n6508) );
  INV_X1 U9356 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8717) );
  AND2_X1 U9357 ( .A1(n7513), .A2(n6928), .ZN(n6927) );
  INV_X1 U9358 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9219) );
  INV_X1 U9359 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U9360 ( .A1(n8156), .A2(n8155), .ZN(n12908) );
  AND3_X1 U9361 ( .A1(n13218), .A2(n13216), .A3(n13217), .ZN(n6509) );
  AND2_X1 U9362 ( .A1(n8688), .A2(SI_17_), .ZN(n6510) );
  AND2_X1 U9363 ( .A1(n8707), .A2(SI_23_), .ZN(n6511) );
  OR2_X1 U9364 ( .A1(n7637), .A2(n6911), .ZN(n6512) );
  AND2_X1 U9365 ( .A1(n8704), .A2(n8703), .ZN(n6513) );
  OR2_X1 U9366 ( .A1(n12110), .A2(n12781), .ZN(n6514) );
  NOR2_X1 U9367 ( .A1(n10879), .A2(n10878), .ZN(n6515) );
  AND2_X1 U9368 ( .A1(n15187), .A2(n15186), .ZN(n6516) );
  INV_X1 U9369 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10826) );
  INV_X1 U9370 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7380) );
  AND2_X1 U9371 ( .A1(n12959), .A2(n12960), .ZN(n6517) );
  OR2_X1 U9372 ( .A1(n11470), .A2(n8020), .ZN(n6518) );
  NOR2_X1 U9373 ( .A1(n13814), .A2(n13294), .ZN(n6519) );
  AND2_X1 U9374 ( .A1(n12231), .A2(n7597), .ZN(n6520) );
  AND2_X1 U9375 ( .A1(n12908), .A2(n12782), .ZN(n6521) );
  NOR2_X1 U9376 ( .A1(n7452), .A2(n14568), .ZN(n6522) );
  OR2_X1 U9377 ( .A1(n7825), .A2(n7821), .ZN(n6523) );
  INV_X1 U9378 ( .A(n14435), .ZN(n7620) );
  INV_X1 U9379 ( .A(n7849), .ZN(n7848) );
  INV_X1 U9380 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7094) );
  INV_X1 U9381 ( .A(n6999), .ZN(n6996) );
  OR2_X1 U9382 ( .A1(n11218), .A2(n11219), .ZN(n6999) );
  AND2_X1 U9383 ( .A1(n8544), .A2(n8543), .ZN(n6524) );
  INV_X1 U9384 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7900) );
  INV_X1 U9385 ( .A(n6848), .ZN(n6847) );
  NAND2_X1 U9386 ( .A1(n6560), .A2(n7990), .ZN(n6848) );
  INV_X1 U9387 ( .A(n9012), .ZN(n7416) );
  OR2_X1 U9388 ( .A1(n15057), .A2(n14858), .ZN(n6525) );
  NAND2_X1 U9389 ( .A1(n14488), .A2(n14487), .ZN(n6526) );
  AND2_X1 U9390 ( .A1(n9943), .A2(n6879), .ZN(n6527) );
  AND2_X1 U9391 ( .A1(n12220), .A2(n13006), .ZN(n6528) );
  AND2_X1 U9392 ( .A1(n7439), .A2(n14804), .ZN(n6529) );
  AND2_X1 U9393 ( .A1(n12856), .A2(n12645), .ZN(n8530) );
  NAND2_X1 U9394 ( .A1(n14449), .A2(n15315), .ZN(n6530) );
  OR2_X1 U9395 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n6531) );
  INV_X1 U9396 ( .A(n13971), .ZN(n6802) );
  AND2_X1 U9397 ( .A1(n7091), .A2(n13486), .ZN(n6532) );
  AND2_X1 U9398 ( .A1(n7748), .A2(n8536), .ZN(n7746) );
  INV_X1 U9399 ( .A(n7746), .ZN(n7197) );
  AND2_X1 U9400 ( .A1(n7151), .A2(n9462), .ZN(n6533) );
  NAND2_X1 U9401 ( .A1(n12884), .A2(n12694), .ZN(n6534) );
  AND2_X1 U9402 ( .A1(n12686), .A2(n12419), .ZN(n8513) );
  INV_X1 U9403 ( .A(n8513), .ZN(n7733) );
  AND2_X1 U9404 ( .A1(n6942), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6535) );
  AND2_X1 U9405 ( .A1(n8663), .A2(n8664), .ZN(n6536) );
  NAND2_X1 U9406 ( .A1(n12296), .A2(n12782), .ZN(n6537) );
  NAND2_X1 U9407 ( .A1(n11469), .A2(n11470), .ZN(n6538) );
  OR2_X1 U9408 ( .A1(n7627), .A2(n14420), .ZN(n6539) );
  OR2_X1 U9409 ( .A1(n12384), .A2(n12748), .ZN(n6540) );
  INV_X1 U9410 ( .A(n9844), .ZN(n6915) );
  INV_X1 U9411 ( .A(n7329), .ZN(n6911) );
  NAND2_X1 U9412 ( .A1(n12298), .A2(n12759), .ZN(n7329) );
  NAND2_X1 U9413 ( .A1(n14055), .A2(n14054), .ZN(n6541) );
  NAND2_X1 U9414 ( .A1(n14425), .A2(n7621), .ZN(n6542) );
  OR2_X1 U9415 ( .A1(n7718), .A2(n13164), .ZN(n6543) );
  AND2_X1 U9416 ( .A1(n7244), .A2(n7245), .ZN(n6544) );
  OR2_X1 U9417 ( .A1(n13155), .A2(n13153), .ZN(n6545) );
  INV_X1 U9418 ( .A(n7877), .ZN(n7493) );
  AND2_X1 U9419 ( .A1(n7698), .A2(n13566), .ZN(n6546) );
  AND2_X1 U9420 ( .A1(n8034), .A2(n7552), .ZN(n6547) );
  AND2_X1 U9421 ( .A1(n7661), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6548) );
  OR2_X1 U9422 ( .A1(n7715), .A2(n13146), .ZN(n6549) );
  NAND2_X1 U9423 ( .A1(n13273), .A2(n13322), .ZN(n6550) );
  AND2_X1 U9424 ( .A1(n7817), .A2(n7893), .ZN(n6551) );
  AND2_X1 U9425 ( .A1(n7666), .A2(n6428), .ZN(n6552) );
  INV_X1 U9426 ( .A(n7425), .ZN(n7424) );
  AND2_X1 U9427 ( .A1(n6423), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6553) );
  AND2_X1 U9428 ( .A1(n6424), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6554) );
  OR2_X1 U9429 ( .A1(n7028), .A2(n7027), .ZN(n6555) );
  INV_X1 U9430 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8631) );
  AND2_X1 U9431 ( .A1(n6820), .A2(n7952), .ZN(n6556) );
  AND2_X1 U9432 ( .A1(n7390), .A2(n6498), .ZN(n6557) );
  INV_X1 U9433 ( .A(n13172), .ZN(n6776) );
  INV_X1 U9434 ( .A(n14350), .ZN(n7625) );
  AND2_X1 U9435 ( .A1(n7195), .A2(n7190), .ZN(n6558) );
  INV_X1 U9436 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7381) );
  INV_X1 U9437 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9441) );
  INV_X1 U9438 ( .A(n7384), .ZN(n7383) );
  OR2_X1 U9439 ( .A1(n10635), .A2(n6428), .ZN(n6559) );
  INV_X1 U9440 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7903) );
  INV_X1 U9441 ( .A(n7215), .ZN(n7211) );
  NAND2_X1 U9442 ( .A1(n12916), .A2(n12769), .ZN(n7215) );
  INV_X1 U9443 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9979) );
  INV_X1 U9444 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10423) );
  NAND2_X1 U9445 ( .A1(n9975), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6560) );
  OR2_X1 U9446 ( .A1(n11470), .A2(n10883), .ZN(n6561) );
  NAND2_X1 U9447 ( .A1(n14436), .A2(n7620), .ZN(n6562) );
  INV_X1 U9448 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7098) );
  INV_X1 U9449 ( .A(n7362), .ZN(n7114) );
  NAND2_X1 U9450 ( .A1(n15009), .A2(n14251), .ZN(n7362) );
  INV_X1 U9451 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10425) );
  INV_X1 U9452 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7090) );
  INV_X1 U9453 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7151) );
  CLKBUF_X3 U9454 ( .A(n12214), .Z(n7171) );
  NAND2_X1 U9455 ( .A1(n12576), .A2(n12568), .ZN(n6563) );
  INV_X1 U9456 ( .A(n11976), .ZN(n7072) );
  NAND2_X1 U9457 ( .A1(n9250), .A2(n9249), .ZN(n14959) );
  INV_X1 U9458 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U9459 ( .A1(n12082), .A2(n12083), .ZN(n12116) );
  INV_X1 U9460 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U9461 ( .A1(n11644), .A2(n7768), .ZN(n11759) );
  NAND2_X1 U9462 ( .A1(n7483), .A2(n7484), .ZN(n6564) );
  INV_X1 U9463 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n7317) );
  NOR2_X1 U9464 ( .A1(n12357), .A2(n15467), .ZN(n6565) );
  INV_X1 U9465 ( .A(n13728), .ZN(n6607) );
  INV_X1 U9466 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7089) );
  INV_X1 U9467 ( .A(n7105), .ZN(n7688) );
  NAND2_X1 U9468 ( .A1(n7179), .A2(n8125), .ZN(n12777) );
  NAND2_X1 U9469 ( .A1(n7722), .A2(n7724), .ZN(n12070) );
  NAND2_X1 U9470 ( .A1(n8032), .A2(n8459), .ZN(n11348) );
  NAND2_X1 U9471 ( .A1(n6648), .A2(n9339), .ZN(n11364) );
  NAND2_X1 U9472 ( .A1(n7827), .A2(n7826), .ZN(n11350) );
  NAND2_X1 U9473 ( .A1(n9247), .A2(n9246), .ZN(n12026) );
  NAND2_X1 U9474 ( .A1(n7012), .A2(n8815), .ZN(n11338) );
  NAND2_X1 U9475 ( .A1(n9244), .A2(n9243), .ZN(n11645) );
  NAND2_X1 U9476 ( .A1(n7793), .A2(n9252), .ZN(n14942) );
  NAND2_X1 U9477 ( .A1(n8213), .A2(n8199), .ZN(n6566) );
  AND2_X1 U9478 ( .A1(n9699), .A2(n9687), .ZN(n11887) );
  INV_X1 U9479 ( .A(n14081), .ZN(n6788) );
  NAND2_X1 U9480 ( .A1(n9817), .A2(n9816), .ZN(n13338) );
  INV_X1 U9481 ( .A(n13338), .ZN(n13197) );
  NOR2_X1 U9482 ( .A1(n14962), .A2(n7445), .ZN(n14915) );
  AND2_X1 U9483 ( .A1(n8284), .A2(n8283), .ZN(n12682) );
  NAND2_X1 U9484 ( .A1(n8249), .A2(n8248), .ZN(n12879) );
  INV_X1 U9485 ( .A(n12879), .ZN(n6650) );
  INV_X1 U9486 ( .A(n12058), .ZN(n12769) );
  AND3_X1 U9487 ( .A1(n8144), .A2(n8143), .A3(n8142), .ZN(n12058) );
  NAND2_X1 U9488 ( .A1(n8195), .A2(n8194), .ZN(n12759) );
  INV_X1 U9489 ( .A(n6715), .ZN(n14739) );
  NAND2_X1 U9490 ( .A1(n9172), .A2(n9157), .ZN(n6715) );
  NAND2_X1 U9491 ( .A1(n9466), .A2(n9465), .ZN(n13491) );
  AND2_X1 U9492 ( .A1(n14921), .A2(n7443), .ZN(n6567) );
  INV_X1 U9493 ( .A(n10498), .ZN(n6974) );
  AND2_X1 U9494 ( .A1(n7158), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U9495 ( .A1(n11917), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6569) );
  INV_X1 U9496 ( .A(n9136), .ZN(n9216) );
  INV_X1 U9497 ( .A(n11537), .ZN(n6942) );
  INV_X1 U9498 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n15539) );
  INV_X1 U9499 ( .A(n13337), .ZN(n13232) );
  NAND2_X1 U9500 ( .A1(n9495), .A2(n9494), .ZN(n13337) );
  AND2_X1 U9501 ( .A1(n6943), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6570) );
  INV_X1 U9502 ( .A(n13184), .ZN(n7721) );
  NOR2_X1 U9503 ( .A1(n12592), .A2(n12830), .ZN(n6571) );
  AND2_X1 U9504 ( .A1(n6691), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6572) );
  NOR2_X1 U9505 ( .A1(n6755), .A2(n6757), .ZN(n6573) );
  AND2_X1 U9506 ( .A1(n6710), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6574) );
  AND2_X1 U9507 ( .A1(n7856), .A2(n7854), .ZN(n6575) );
  AND2_X1 U9508 ( .A1(n11690), .A2(n9833), .ZN(n6576) );
  AND2_X1 U9509 ( .A1(n6937), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6577) );
  OAI21_X1 U9510 ( .B1(n10935), .B2(n10930), .A(n7136), .ZN(n6972) );
  AND2_X1 U9511 ( .A1(n7721), .A2(n13185), .ZN(n6578) );
  OR2_X1 U9512 ( .A1(n12021), .A2(n12004), .ZN(n6579) );
  INV_X1 U9513 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10274) );
  AND2_X1 U9514 ( .A1(n8145), .A2(n8128), .ZN(n8129) );
  INV_X1 U9515 ( .A(n15395), .ZN(n6638) );
  XNOR2_X1 U9516 ( .A(n8185), .B(n8184), .ZN(n12576) );
  INV_X1 U9517 ( .A(n15484), .ZN(n12784) );
  NAND2_X1 U9518 ( .A1(n15241), .A2(n15303), .ZN(n11382) );
  BUF_X1 U9519 ( .A(n10806), .Z(n13354) );
  INV_X1 U9520 ( .A(n13355), .ZN(n6906) );
  INV_X1 U9521 ( .A(n10801), .ZN(n6602) );
  AND2_X1 U9522 ( .A1(n12555), .A2(n12534), .ZN(n6580) );
  AND3_X2 U9523 ( .A1(n9912), .A2(n10712), .A3(n15417), .ZN(n15454) );
  AND2_X1 U9524 ( .A1(n10132), .A2(n10131), .ZN(n12590) );
  INV_X1 U9525 ( .A(n12434), .ZN(n12439) );
  OR2_X1 U9526 ( .A1(n6403), .A2(n9160), .ZN(n6581) );
  OR2_X1 U9527 ( .A1(n6403), .A2(n7130), .ZN(n6582) );
  NOR2_X1 U9528 ( .A1(n6612), .A2(n12208), .ZN(n6583) );
  INV_X1 U9529 ( .A(n15086), .ZN(n7446) );
  AND2_X1 U9530 ( .A1(n8250), .A2(n6698), .ZN(n6584) );
  NAND2_X1 U9531 ( .A1(n7070), .A2(n7023), .ZN(n11318) );
  NAND2_X1 U9532 ( .A1(n9328), .A2(n9327), .ZN(n15463) );
  INV_X1 U9533 ( .A(n15481), .ZN(n7172) );
  OR2_X1 U9534 ( .A1(n15448), .A2(n7081), .ZN(n6585) );
  AND2_X1 U9535 ( .A1(n9283), .A2(n14307), .ZN(n9293) );
  INV_X1 U9536 ( .A(n12558), .ZN(n7256) );
  INV_X1 U9537 ( .A(n12518), .ZN(n6947) );
  INV_X1 U9538 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6711) );
  INV_X1 U9539 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6689) );
  INV_X1 U9540 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6692) );
  AND2_X1 U9541 ( .A1(n6841), .A2(n6838), .ZN(n6586) );
  AND2_X1 U9542 ( .A1(n8448), .A2(n8441), .ZN(n11086) );
  INV_X1 U9543 ( .A(n11086), .ZN(n7286) );
  AND2_X1 U9544 ( .A1(n6934), .A2(n7666), .ZN(n6587) );
  AND2_X1 U9545 ( .A1(n15143), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6588) );
  AND2_X1 U9546 ( .A1(n8705), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6589) );
  OR2_X1 U9547 ( .A1(n12588), .A2(n7676), .ZN(n6590) );
  AND2_X1 U9548 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15162), .ZN(n6591) );
  NAND2_X1 U9549 ( .A1(n6642), .A2(n6482), .ZN(n6641) );
  OR2_X1 U9550 ( .A1(n14645), .A2(n14646), .ZN(n6592) );
  AND2_X1 U9551 ( .A1(n6747), .A2(n6746), .ZN(n6593) );
  INV_X1 U9552 ( .A(n14664), .ZN(n7145) );
  INV_X1 U9553 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n6700) );
  AND2_X1 U9554 ( .A1(n6958), .A2(n10430), .ZN(n6594) );
  AND2_X1 U9555 ( .A1(n7804), .A2(n8724), .ZN(n7111) );
  INV_X1 U9556 ( .A(n6758), .ZN(n6757) );
  NAND2_X1 U9557 ( .A1(n12012), .A2(n12001), .ZN(n6758) );
  INV_X1 U9558 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n6622) );
  INV_X1 U9559 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7095) );
  INV_X1 U9560 ( .A(SI_8_), .ZN(n6615) );
  INV_X1 U9561 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6895) );
  INV_X1 U9562 ( .A(n12576), .ZN(n7385) );
  NAND2_X1 U9563 ( .A1(n7386), .A2(n12576), .ZN(n7384) );
  NAND2_X1 U9564 ( .A1(n8874), .A2(n8873), .ZN(n8876) );
  INV_X1 U9565 ( .A(n9295), .ZN(n7113) );
  NAND2_X1 U9566 ( .A1(n14824), .A2(n14827), .ZN(n14825) );
  NAND3_X1 U9567 ( .A1(n8649), .A2(n8648), .A3(n8751), .ZN(n8769) );
  NOR2_X2 U9568 ( .A1(n14840), .A2(n14399), .ZN(n14841) );
  INV_X1 U9569 ( .A(n7071), .ZN(n7070) );
  NAND2_X1 U9570 ( .A1(n11377), .A2(n8872), .ZN(n11642) );
  INV_X2 U9571 ( .A(n10781), .ZN(n8756) );
  NAND2_X1 U9572 ( .A1(n12027), .A2(n8926), .ZN(n7009) );
  NAND2_X1 U9573 ( .A1(n15245), .A2(n15252), .ZN(n7012) );
  NAND2_X1 U9574 ( .A1(n14943), .A2(n7018), .ZN(n7017) );
  NAND2_X1 U9575 ( .A1(n11318), .A2(n8791), .ZN(n8793) );
  NAND2_X1 U9576 ( .A1(n6462), .A2(n7065), .ZN(n15121) );
  NAND2_X1 U9577 ( .A1(n11860), .A2(n6437), .ZN(n6665) );
  OR2_X1 U9578 ( .A1(n13768), .A2(n13855), .ZN(n7161) );
  NAND2_X2 U9579 ( .A1(n9635), .A2(n9634), .ZN(n7105) );
  NAND2_X1 U9580 ( .A1(n6663), .A2(n9759), .ZN(n13583) );
  NAND2_X1 U9581 ( .A1(n9746), .A2(n13297), .ZN(n13607) );
  NAND2_X1 U9582 ( .A1(n6595), .A2(n7872), .ZN(n14413) );
  OAI22_X1 U9583 ( .A1(n7400), .A2(n7399), .B1(n7404), .B2(n14398), .ZN(n6595)
         );
  NAND2_X1 U9584 ( .A1(n7351), .A2(n8965), .ZN(n8967) );
  OAI21_X2 U9585 ( .B1(n10570), .B2(n14463), .A(n8971), .ZN(n15078) );
  NAND2_X1 U9586 ( .A1(n7017), .A2(n7015), .ZN(n14866) );
  OAI21_X1 U9587 ( .B1(n7022), .B2(n7021), .A(n9050), .ZN(n7016) );
  AOI21_X1 U9588 ( .B1(n6791), .B2(n6793), .A(n6788), .ZN(n6787) );
  AOI21_X2 U9589 ( .B1(n7461), .B2(n7459), .A(n14246), .ZN(n7458) );
  NAND3_X1 U9590 ( .A1(n6958), .A2(n10430), .A3(P3_REG2_REG_3__SCAN_IN), .ZN(
        n10449) );
  NOR2_X2 U9591 ( .A1(n9858), .A2(n13450), .ZN(n13471) );
  NOR2_X1 U9592 ( .A1(n12003), .A2(n7662), .ZN(n11918) );
  INV_X1 U9593 ( .A(n12492), .ZN(n6949) );
  AOI21_X1 U9594 ( .B1(n6914), .B2(n9844), .A(n7345), .ZN(n6913) );
  NAND2_X1 U9595 ( .A1(n6948), .A2(n12493), .ZN(n12513) );
  NAND3_X1 U9596 ( .A1(n7512), .A2(n9461), .A3(n9476), .ZN(n13906) );
  AND2_X4 U9597 ( .A1(n6599), .A2(n9585), .ZN(n9461) );
  NAND2_X1 U9598 ( .A1(n7713), .A2(n7714), .ZN(n13151) );
  NAND2_X1 U9599 ( .A1(n7705), .A2(n6601), .ZN(n7704) );
  OAI21_X1 U9600 ( .B1(n6487), .B2(n6603), .A(n6775), .ZN(n13175) );
  NAND2_X1 U9601 ( .A1(n6780), .A2(n7711), .ZN(n13139) );
  NAND2_X1 U9602 ( .A1(n13151), .A2(n13150), .ZN(n6765) );
  NOR2_X2 U9603 ( .A1(n9711), .A2(n9439), .ZN(n6599) );
  NAND2_X1 U9604 ( .A1(n6600), .A2(n7707), .ZN(n13131) );
  NAND3_X1 U9605 ( .A1(n13125), .A2(n7709), .A3(n13124), .ZN(n6600) );
  NAND2_X1 U9606 ( .A1(n9883), .A2(n7610), .ZN(n9875) );
  OAI21_X1 U9607 ( .B1(n13186), .B2(n6578), .A(n7719), .ZN(n13188) );
  OAI21_X1 U9608 ( .B1(n6772), .B2(n6770), .A(n6509), .ZN(n6769) );
  NAND2_X1 U9609 ( .A1(n6602), .A2(n13277), .ZN(n6601) );
  AND2_X4 U9610 ( .A1(n13111), .A2(n13094), .ZN(n13277) );
  NOR3_X2 U9611 ( .A1(n13471), .A2(n13472), .A3(n13475), .ZN(n13473) );
  NAND2_X1 U9612 ( .A1(n11628), .A2(n9832), .ZN(n11691) );
  NAND2_X1 U9613 ( .A1(n11584), .A2(n9831), .ZN(n11629) );
  NAND2_X2 U9614 ( .A1(n6455), .A2(n6673), .ZN(n9870) );
  NAND2_X2 U9615 ( .A1(n9848), .A2(n9847), .ZN(n13627) );
  NAND2_X1 U9616 ( .A1(n11583), .A2(n9830), .ZN(n11584) );
  NAND2_X1 U9617 ( .A1(n13170), .A2(n6774), .ZN(n6603) );
  OAI21_X1 U9618 ( .B1(n6488), .B2(n6604), .A(n6768), .ZN(n13186) );
  NAND2_X1 U9619 ( .A1(n13179), .A2(n6766), .ZN(n6604) );
  INV_X1 U9620 ( .A(n13169), .ZN(n7164) );
  NAND2_X1 U9621 ( .A1(n6477), .A2(n13415), .ZN(n13426) );
  OR2_X1 U9622 ( .A1(n13434), .A2(n13433), .ZN(n6639) );
  NAND2_X1 U9623 ( .A1(n6762), .A2(n7710), .ZN(n13158) );
  NAND2_X1 U9624 ( .A1(n7490), .A2(n7493), .ZN(n7489) );
  NAND2_X1 U9625 ( .A1(n7512), .A2(n9461), .ZN(n6605) );
  AOI21_X1 U9626 ( .B1(n13188), .B2(n13187), .A(n6771), .ZN(n6770) );
  NAND2_X1 U9627 ( .A1(n13238), .A2(n6769), .ZN(n13274) );
  NAND2_X1 U9628 ( .A1(n13274), .A2(n7878), .ZN(n7107) );
  AOI21_X2 U9629 ( .B1(n13881), .B2(n13862), .A(n13861), .ZN(n13863) );
  NAND2_X2 U9630 ( .A1(n13532), .A2(n6693), .ZN(n13517) );
  NAND2_X1 U9631 ( .A1(n7693), .A2(n7690), .ZN(n13461) );
  NAND2_X1 U9632 ( .A1(n7697), .A2(n6546), .ZN(n13564) );
  NAND2_X2 U9633 ( .A1(n13022), .A2(n7595), .ZN(n7593) );
  NAND2_X2 U9634 ( .A1(n7593), .A2(n7591), .ZN(n12982) );
  NAND2_X2 U9635 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  NAND2_X1 U9636 ( .A1(n10868), .A2(n10867), .ZN(n10922) );
  INV_X1 U9637 ( .A(n10861), .ZN(n6988) );
  NAND2_X1 U9638 ( .A1(n6639), .A2(n6633), .ZN(P2_U3233) );
  NOR2_X1 U9639 ( .A1(n11010), .A2(n6491), .ZN(n10810) );
  NAND2_X1 U9640 ( .A1(n11669), .A2(n13262), .ZN(n9775) );
  NAND2_X1 U9641 ( .A1(n7529), .A2(n7531), .ZN(n6865) );
  NAND2_X1 U9642 ( .A1(n6866), .A2(n6865), .ZN(n6864) );
  INV_X1 U9643 ( .A(n7332), .ZN(n6678) );
  NAND2_X1 U9644 ( .A1(n6897), .A2(n7651), .ZN(n11772) );
  NAND2_X1 U9645 ( .A1(n7208), .A2(n7207), .ZN(n7206) );
  NAND2_X1 U9646 ( .A1(n12746), .A2(n7846), .ZN(n7845) );
  NAND2_X1 U9647 ( .A1(n7201), .A2(n12702), .ZN(n6651) );
  NAND2_X1 U9648 ( .A1(n11187), .A2(n11186), .ZN(n11190) );
  XNOR2_X1 U9649 ( .A(n9425), .B(n6524), .ZN(n7203) );
  OAI21_X1 U9650 ( .B1(n7214), .B2(n7217), .A(n12778), .ZN(n7213) );
  INV_X1 U9651 ( .A(n7854), .ZN(n7853) );
  NAND2_X1 U9652 ( .A1(n7831), .A2(n7835), .ZN(n9424) );
  XNOR2_X2 U9653 ( .A(n6611), .B(n7892), .ZN(n12125) );
  OAI21_X2 U9654 ( .B1(n7818), .B2(n7816), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n6611) );
  OAI21_X1 U9655 ( .B1(n7756), .B2(n7752), .A(n7751), .ZN(n12852) );
  NAND2_X1 U9656 ( .A1(n12054), .A2(n6919), .ZN(n6918) );
  AOI21_X1 U9657 ( .B1(n7458), .B2(n7460), .A(n7457), .ZN(n7456) );
  NAND2_X1 U9658 ( .A1(n6789), .A2(n6787), .ZN(n14028) );
  NAND2_X2 U9659 ( .A1(n14047), .A2(n14156), .ZN(n14158) );
  NOR2_X1 U9660 ( .A1(n10350), .A2(n10351), .ZN(n10349) );
  OAI21_X1 U9661 ( .B1(n7346), .B2(n7344), .A(n9710), .ZN(n6668) );
  NAND2_X1 U9662 ( .A1(n13794), .A2(n9784), .ZN(n13541) );
  NAND2_X2 U9663 ( .A1(n9771), .A2(n9770), .ZN(n13572) );
  NAND3_X1 U9664 ( .A1(n14445), .A2(n14446), .A3(n14444), .ZN(n7618) );
  NAND2_X1 U9665 ( .A1(n8769), .A2(n6619), .ZN(n7426) );
  NAND2_X1 U9666 ( .A1(n7121), .A2(n7120), .ZN(n7119) );
  MUX2_X1 U9667 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13919), .S(n10089), .Z(n11051)
         );
  NOR2_X2 U9668 ( .A1(n11577), .A2(n13145), .ZN(n11624) );
  NAND2_X1 U9669 ( .A1(n7819), .A2(n6654), .ZN(n6653) );
  INV_X1 U9670 ( .A(n7271), .ZN(n7270) );
  INV_X1 U9671 ( .A(n10641), .ZN(n7272) );
  INV_X1 U9672 ( .A(n7257), .ZN(n11533) );
  INV_X1 U9673 ( .A(n12604), .ZN(n7243) );
  NAND4_X1 U9674 ( .A1(n7241), .A2(n7246), .A3(n7670), .A4(n6544), .ZN(
        P3_U3201) );
  NAND2_X1 U9675 ( .A1(n7142), .A2(n14672), .ZN(n7141) );
  NAND2_X1 U9676 ( .A1(n7000), .A2(n7601), .ZN(n12248) );
  NOR2_X1 U9677 ( .A1(n13058), .A2(n7596), .ZN(n7595) );
  XNOR2_X1 U9678 ( .A(n14666), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n14667) );
  INV_X1 U9679 ( .A(n14667), .ZN(n14671) );
  OAI21_X2 U9680 ( .B1(n6930), .B2(n7818), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7894) );
  AOI21_X2 U9681 ( .B1(n9350), .B2(n12336), .A(n12401), .ZN(n12342) );
  NAND2_X1 U9682 ( .A1(n6918), .A2(n6917), .ZN(n12294) );
  AOI22_X1 U9683 ( .A1(n11868), .A2(n11867), .B1(n11866), .B2(n12781), .ZN(
        n12054) );
  NAND2_X1 U9684 ( .A1(n10846), .A2(n10845), .ZN(n10847) );
  INV_X1 U9685 ( .A(n10575), .ZN(n15477) );
  INV_X1 U9686 ( .A(n6916), .ZN(n12381) );
  AND3_X2 U9687 ( .A1(n7326), .A2(n12398), .A3(n12682), .ZN(n12401) );
  NAND3_X1 U9688 ( .A1(n10690), .A2(n6625), .A3(n10689), .ZN(n10846) );
  OAI21_X1 U9689 ( .B1(n12294), .B2(n7650), .A(n6537), .ZN(n6916) );
  NAND2_X1 U9690 ( .A1(n6896), .A2(n11901), .ZN(n11868) );
  NAND2_X1 U9691 ( .A1(n8591), .A2(n8216), .ZN(n8397) );
  NOR2_X2 U9692 ( .A1(n8215), .A2(n7891), .ZN(n8216) );
  NAND2_X1 U9693 ( .A1(n12363), .A2(n12364), .ZN(n12362) );
  NAND2_X1 U9694 ( .A1(n7117), .A2(n7116), .ZN(n14440) );
  NOR2_X1 U9695 ( .A1(n7619), .A2(n14519), .ZN(n14557) );
  NAND2_X1 U9696 ( .A1(n6627), .A2(n6626), .ZN(n10087) );
  NAND2_X1 U9697 ( .A1(n10262), .A2(n6630), .ZN(n6626) );
  MUX2_X1 U9698 ( .A(n10072), .B(P2_REG1_REG_1__SCAN_IN), .S(n13362), .Z(
        n10074) );
  NAND3_X1 U9699 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n6647) );
  OAI21_X1 U9700 ( .B1(n7204), .B2(n6435), .A(n6540), .ZN(n6656) );
  OAI21_X1 U9701 ( .B1(n7210), .B2(n7206), .A(n7204), .ZN(n12758) );
  NAND2_X1 U9702 ( .A1(n13583), .A2(n13582), .ZN(n9771) );
  NAND2_X1 U9703 ( .A1(n13607), .A2(n9758), .ZN(n6663) );
  NAND3_X1 U9704 ( .A1(n7700), .A2(n9461), .A3(n9462), .ZN(n6672) );
  NAND2_X4 U9705 ( .A1(n13328), .A2(n9870), .ZN(n10089) );
  OAI211_X2 U9706 ( .C1(n13572), .C2(n6679), .A(n6677), .B(n7087), .ZN(n13451)
         );
  AOI21_X4 U9707 ( .B1(n13451), .B2(n13450), .A(n6456), .ZN(n13758) );
  OAI21_X1 U9708 ( .B1(n11294), .B2(n6685), .A(n6683), .ZN(n11689) );
  NAND2_X1 U9709 ( .A1(n11294), .A2(n6683), .ZN(n6682) );
  NAND2_X1 U9710 ( .A1(n9808), .A2(n9807), .ZN(n9809) );
  NAND2_X1 U9711 ( .A1(n9468), .A2(n6553), .ZN(n9606) );
  XNOR2_X2 U9712 ( .A(n13338), .B(n6693), .ZN(n13515) );
  INV_X2 U9713 ( .A(n13521), .ZN(n6693) );
  NAND2_X1 U9714 ( .A1(n6705), .A2(n6704), .ZN(n8062) );
  NAND3_X1 U9715 ( .A1(n7942), .A2(n10610), .A3(n7941), .ZN(n7980) );
  NAND2_X1 U9716 ( .A1(n8608), .A2(n6554), .ZN(n8901) );
  NAND2_X1 U9717 ( .A1(n8611), .A2(n6574), .ZN(n9027) );
  NAND3_X1 U9718 ( .A1(n7467), .A2(n7465), .A3(n6713), .ZN(n6712) );
  NAND2_X1 U9719 ( .A1(n6716), .A2(n6472), .ZN(n6852) );
  NAND3_X1 U9720 ( .A1(n13622), .A2(n13571), .A3(n6720), .ZN(n6719) );
  NAND4_X1 U9721 ( .A1(n13321), .A2(n13322), .A3(n13320), .A4(n13755), .ZN(
        n6726) );
  INV_X8 U9722 ( .A(n9464), .ZN(n7434) );
  NAND2_X1 U9723 ( .A1(n9464), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6729) );
  NAND3_X1 U9724 ( .A1(n6731), .A2(n6734), .A3(n6730), .ZN(n6736) );
  NAND2_X1 U9725 ( .A1(n12577), .A2(n6571), .ZN(n6730) );
  NAND2_X1 U9726 ( .A1(n12577), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n6733) );
  OR2_X1 U9727 ( .A1(n12599), .A2(n12591), .ZN(n6734) );
  NAND2_X1 U9728 ( .A1(n6735), .A2(n12607), .ZN(n7244) );
  XNOR2_X1 U9729 ( .A(n6736), .B(n12602), .ZN(n6735) );
  NAND2_X1 U9730 ( .A1(n12540), .A2(n12531), .ZN(n6743) );
  NAND2_X1 U9731 ( .A1(n12540), .A2(n6738), .ZN(n6737) );
  NAND3_X1 U9732 ( .A1(n6764), .A2(n6545), .A3(n6763), .ZN(n6762) );
  NAND2_X1 U9733 ( .A1(n6765), .A2(n13149), .ZN(n6764) );
  OAI21_X1 U9734 ( .B1(n13131), .B2(n6779), .A(n6777), .ZN(n6780) );
  AND2_X1 U9735 ( .A1(n6486), .A2(n6778), .ZN(n6777) );
  OR2_X1 U9736 ( .A1(n6781), .A2(n13132), .ZN(n6778) );
  AND2_X1 U9737 ( .A1(n6781), .A2(n13132), .ZN(n6779) );
  INV_X1 U9738 ( .A(n13130), .ZN(n6781) );
  XNOR2_X1 U9739 ( .A(n6782), .B(n10894), .ZN(n10666) );
  NAND2_X1 U9740 ( .A1(n14101), .A2(n6791), .ZN(n6789) );
  NAND2_X1 U9741 ( .A1(n6798), .A2(n6794), .ZN(n14195) );
  NAND2_X1 U9742 ( .A1(n6800), .A2(n13971), .ZN(n6797) );
  INV_X1 U9743 ( .A(n6800), .ZN(n6799) );
  INV_X1 U9744 ( .A(n6803), .ZN(n14167) );
  NOR2_X1 U9745 ( .A1(n9058), .A2(n6806), .ZN(n9223) );
  INV_X1 U9746 ( .A(n6815), .ZN(n6808) );
  NAND2_X1 U9747 ( .A1(n6809), .A2(n6812), .ZN(n11815) );
  NAND4_X1 U9748 ( .A1(n7546), .A2(n7547), .A3(n7949), .A4(n7972), .ZN(n6818)
         );
  NAND2_X1 U9749 ( .A1(n6818), .A2(n6556), .ZN(n7988) );
  NAND3_X1 U9750 ( .A1(n7546), .A2(n7547), .A3(n7949), .ZN(n6819) );
  NAND2_X1 U9751 ( .A1(n7557), .A2(n6828), .ZN(n6825) );
  NAND2_X1 U9752 ( .A1(n6825), .A2(n6826), .ZN(n8289) );
  NAND2_X1 U9753 ( .A1(n7560), .A2(n6834), .ZN(n6831) );
  NAND2_X1 U9754 ( .A1(n6831), .A2(n6832), .ZN(n8232) );
  INV_X1 U9755 ( .A(n8300), .ZN(n6837) );
  NAND2_X1 U9756 ( .A1(n8069), .A2(n6850), .ZN(n6849) );
  NAND2_X1 U9757 ( .A1(n6849), .A2(n7581), .ZN(n8108) );
  NAND2_X1 U9758 ( .A1(n8069), .A2(n8068), .ZN(n8071) );
  INV_X1 U9759 ( .A(n13526), .ZN(n6866) );
  OAI21_X1 U9760 ( .B1(n7429), .B2(n6874), .A(n6872), .ZN(n9119) );
  NAND2_X1 U9761 ( .A1(n7429), .A2(n6870), .ZN(n6869) );
  NAND2_X1 U9762 ( .A1(n7429), .A2(n7428), .ZN(n9103) );
  OAI21_X1 U9763 ( .B1(n9464), .B2(n10425), .A(n6875), .ZN(n8671) );
  NAND2_X1 U9764 ( .A1(n9464), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U9765 ( .A1(n9464), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U9766 ( .A1(n6878), .A2(n9987), .ZN(n9988) );
  NAND2_X1 U9767 ( .A1(n6880), .A2(n9943), .ZN(n6877) );
  NAND2_X1 U9768 ( .A1(n6880), .A2(n6527), .ZN(n6878) );
  NAND2_X1 U9769 ( .A1(n9942), .A2(n9943), .ZN(n9945) );
  NAND3_X1 U9770 ( .A1(n9942), .A2(n9943), .A3(n6881), .ZN(n6880) );
  NAND2_X1 U9771 ( .A1(n15155), .A2(n15154), .ZN(n6884) );
  NAND2_X1 U9772 ( .A1(n10503), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10506) );
  INV_X1 U9773 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U9774 ( .A1(n6892), .A2(n12096), .ZN(n12101) );
  NAND2_X1 U9775 ( .A1(n9827), .A2(n9826), .ZN(n11058) );
  NAND2_X1 U9776 ( .A1(n6900), .A2(n11058), .ZN(n6902) );
  NAND2_X1 U9777 ( .A1(n6902), .A2(n6901), .ZN(n11583) );
  OR2_X1 U9778 ( .A1(n7877), .A2(n7491), .ZN(n6901) );
  INV_X1 U9779 ( .A(n9830), .ZN(n13309) );
  NAND4_X4 U9780 ( .A1(n7162), .A2(n6904), .A3(n9498), .A4(n6905), .ZN(n10801)
         );
  NAND3_X2 U9781 ( .A1(n9522), .A2(n9523), .A3(n9521), .ZN(n10805) );
  INV_X1 U9782 ( .A(n7517), .ZN(n6914) );
  OAI21_X2 U9783 ( .B1(n13696), .B2(n6915), .A(n6913), .ZN(n13661) );
  NAND2_X1 U9784 ( .A1(n13681), .A2(n9844), .ZN(n13662) );
  NAND2_X1 U9785 ( .A1(n13696), .A2(n7517), .ZN(n13681) );
  OAI21_X2 U9786 ( .B1(n12041), .B2(n9841), .A(n9840), .ZN(n13696) );
  NAND2_X1 U9787 ( .A1(n12055), .A2(n12058), .ZN(n6917) );
  NAND2_X1 U9788 ( .A1(n6920), .A2(n12769), .ZN(n6919) );
  OAI21_X1 U9789 ( .B1(n13627), .B2(n6921), .A(n6924), .ZN(n13559) );
  INV_X1 U9790 ( .A(n6927), .ZN(n6921) );
  NAND2_X2 U9791 ( .A1(n6923), .A2(n6922), .ZN(n13551) );
  NAND4_X1 U9793 ( .A1(n7819), .A2(n8216), .A3(n7820), .A4(n6551), .ZN(n12927)
         );
  NOR2_X1 U9794 ( .A1(n12927), .A2(P3_IR_REG_30__SCAN_IN), .ZN(n7233) );
  NAND3_X1 U9795 ( .A1(n11175), .A2(n11181), .A3(n6931), .ZN(n11177) );
  XNOR2_X1 U9796 ( .A(n11164), .B(n11174), .ZN(n11181) );
  NAND2_X1 U9797 ( .A1(n6415), .A2(n12478), .ZN(n12463) );
  NAND2_X1 U9798 ( .A1(n11918), .A2(n6577), .ZN(n6936) );
  INV_X1 U9799 ( .A(n11536), .ZN(n6941) );
  NAND2_X1 U9800 ( .A1(n6949), .A2(n12463), .ZN(n6948) );
  INV_X1 U9801 ( .A(n6955), .ZN(n6954) );
  NAND3_X1 U9802 ( .A1(n6952), .A2(n6951), .A3(n6950), .ZN(n12553) );
  NAND2_X1 U9803 ( .A1(n10449), .A2(n10430), .ZN(n10392) );
  NAND2_X1 U9804 ( .A1(n10390), .A2(n10405), .ZN(n10430) );
  NAND2_X1 U9805 ( .A1(n11559), .A2(n6963), .ZN(n6959) );
  NAND2_X1 U9806 ( .A1(n6959), .A2(n6960), .ZN(n11841) );
  OAI21_X1 U9807 ( .B1(n15179), .B2(n15180), .A(n6480), .ZN(n6966) );
  INV_X1 U9808 ( .A(n6970), .ZN(n10479) );
  NAND2_X1 U9809 ( .A1(n6970), .A2(n6969), .ZN(n6968) );
  NAND2_X1 U9810 ( .A1(n10054), .A2(n10053), .ZN(n6970) );
  AOI21_X1 U9811 ( .B1(n10499), .B2(n6973), .A(n6972), .ZN(n11551) );
  NAND2_X1 U9812 ( .A1(n12082), .A2(n6414), .ZN(n6975) );
  NAND2_X1 U9813 ( .A1(n6975), .A2(n6976), .ZN(n7147) );
  NAND2_X1 U9814 ( .A1(n7600), .A2(n7598), .ZN(n13068) );
  AOI21_X1 U9815 ( .B1(n6989), .B2(n6988), .A(n6504), .ZN(n10868) );
  NAND2_X1 U9816 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  NAND2_X1 U9817 ( .A1(n10956), .A2(n10804), .ZN(n11012) );
  NOR2_X1 U9818 ( .A1(n11011), .A2(n11012), .ZN(n11010) );
  XNOR2_X1 U9819 ( .A(n10802), .B(n6990), .ZN(n11011) );
  NAND2_X1 U9820 ( .A1(n12982), .A2(n7005), .ZN(n7000) );
  NAND2_X1 U9821 ( .A1(n7009), .A2(n14961), .ZN(n14960) );
  OAI211_X1 U9822 ( .C1(n7009), .C2(n14961), .A(n14960), .B(n15308), .ZN(
        n15098) );
  NAND2_X1 U9823 ( .A1(n7012), .A2(n7010), .ZN(n8834) );
  NAND2_X1 U9824 ( .A1(n7013), .A2(n10304), .ZN(n10152) );
  NAND3_X1 U9825 ( .A1(n14321), .A2(n14326), .A3(n14527), .ZN(n7023) );
  NAND2_X1 U9826 ( .A1(n14766), .A2(n7030), .ZN(n7029) );
  NAND2_X1 U9827 ( .A1(n7025), .A2(n7024), .ZN(n7779) );
  NAND2_X1 U9828 ( .A1(n14766), .A2(n7026), .ZN(n7025) );
  NAND3_X1 U9829 ( .A1(n7362), .A2(n14769), .A3(n14768), .ZN(n7031) );
  INV_X1 U9830 ( .A(n9239), .ZN(n7038) );
  NAND3_X1 U9831 ( .A1(n7153), .A2(n9239), .A3(n11317), .ZN(n7036) );
  OAI21_X1 U9832 ( .B1(n11317), .B2(n7801), .A(n7153), .ZN(n11337) );
  NAND3_X1 U9833 ( .A1(n7036), .A2(n7034), .A3(n7032), .ZN(n9241) );
  NAND2_X1 U9834 ( .A1(n7153), .A2(n7033), .ZN(n7032) );
  INV_X1 U9835 ( .A(n7035), .ZN(n7034) );
  OAI21_X1 U9836 ( .B1(n7038), .B2(n14530), .A(n15227), .ZN(n7035) );
  NAND3_X2 U9837 ( .A1(n7040), .A2(n7039), .A3(n8622), .ZN(n8856) );
  OAI21_X1 U9838 ( .B1(n7043), .B2(n9243), .A(n9245), .ZN(n7042) );
  NAND2_X1 U9839 ( .A1(n14907), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U9840 ( .A1(n14901), .A2(n7049), .ZN(n7048) );
  NAND2_X1 U9841 ( .A1(n7048), .A2(n7052), .ZN(n14839) );
  NAND2_X1 U9842 ( .A1(n14901), .A2(n14902), .ZN(n7059) );
  OAI21_X1 U9843 ( .B1(n12148), .B2(n7064), .A(n7062), .ZN(n14731) );
  OAI22_X1 U9844 ( .A1(n12148), .A2(n7061), .B1(n7060), .B2(n7062), .ZN(n12137) );
  NAND2_X1 U9845 ( .A1(n12148), .A2(n7802), .ZN(n14758) );
  NAND2_X1 U9846 ( .A1(n9269), .A2(n7027), .ZN(n12148) );
  INV_X1 U9847 ( .A(n14578), .ZN(n15281) );
  NAND2_X1 U9848 ( .A1(n7359), .A2(n7360), .ZN(n9420) );
  AOI21_X1 U9849 ( .B1(n14839), .B2(n14399), .A(n9263), .ZN(n14824) );
  NAND2_X1 U9850 ( .A1(n8834), .A2(n7775), .ZN(n7774) );
  NAND2_X1 U9851 ( .A1(n7774), .A2(n7772), .ZN(n11377) );
  NAND2_X1 U9852 ( .A1(n14580), .A2(n10781), .ZN(n8758) );
  NAND2_X1 U9853 ( .A1(n14673), .A2(n14934), .ZN(n7140) );
  AOI21_X1 U9854 ( .B1(n14692), .B2(n15308), .A(n7113), .ZN(n7359) );
  OAI21_X1 U9855 ( .B1(n14670), .B2(n7141), .A(n7140), .ZN(n14676) );
  XNOR2_X2 U9856 ( .A(n8787), .B(n8809), .ZN(n15220) );
  OAI21_X1 U9857 ( .B1(n14648), .B2(n14647), .A(n6592), .ZN(n14660) );
  NOR2_X1 U9858 ( .A1(n10764), .A2(n10763), .ZN(n11108) );
  AOI21_X1 U9859 ( .B1(n10221), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10343), .ZN(
        n10216) );
  AOI21_X1 U9860 ( .B1(n10165), .B2(P1_REG1_REG_4__SCAN_IN), .A(n15204), .ZN(
        n10187) );
  NOR3_X1 U9861 ( .A1(n11971), .A2(n11797), .A3(n11796), .ZN(n14635) );
  NAND2_X1 U9862 ( .A1(n11249), .A2(n15440), .ZN(n11296) );
  NAND2_X1 U9863 ( .A1(n7152), .A2(n10986), .ZN(n10985) );
  NOR2_X2 U9864 ( .A1(n13652), .A2(n13814), .ZN(n7697) );
  NAND2_X2 U9865 ( .A1(n7701), .A2(n7702), .ZN(n13113) );
  NAND4_X1 U9866 ( .A1(n11695), .A2(n7689), .A3(n11698), .A4(n13734), .ZN(
        n13728) );
  NAND4_X1 U9867 ( .A1(n13459), .A2(n13460), .A3(n13458), .A4(n6465), .ZN(
        n13760) );
  NAND2_X1 U9868 ( .A1(n9823), .A2(n13300), .ZN(n10750) );
  CLKBUF_X1 U9869 ( .A(n7099), .Z(n7079) );
  NAND2_X1 U9870 ( .A1(n9524), .A2(n10805), .ZN(n10751) );
  NAND2_X1 U9871 ( .A1(n11629), .A2(n13310), .ZN(n11628) );
  NAND2_X1 U9872 ( .A1(n13864), .A2(n15448), .ZN(n7082) );
  INV_X1 U9873 ( .A(n9502), .ZN(n7702) );
  NAND2_X1 U9874 ( .A1(n11851), .A2(n9834), .ZN(n12041) );
  NAND2_X1 U9875 ( .A1(n12998), .A2(n12999), .ZN(n7600) );
  NAND2_X1 U9876 ( .A1(n11987), .A2(n11986), .ZN(n12081) );
  INV_X1 U9877 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7538) );
  OR2_X1 U9878 ( .A1(n7335), .A2(n6431), .ZN(n7332) );
  XNOR2_X1 U9879 ( .A(n9104), .B(SI_22_), .ZN(n9773) );
  XNOR2_X2 U9880 ( .A(n13792), .B(n13340), .ZN(n13571) );
  AOI21_X1 U9881 ( .B1(n13758), .B2(n13757), .A(n13756), .ZN(n13759) );
  NAND2_X1 U9882 ( .A1(n7082), .A2(n6585), .ZN(P2_U3496) );
  INV_X1 U9883 ( .A(n9461), .ZN(n9720) );
  NAND2_X1 U9884 ( .A1(n9461), .A2(n7090), .ZN(n9880) );
  NAND2_X1 U9885 ( .A1(n7716), .A2(n7717), .ZN(n13169) );
  AOI21_X1 U9886 ( .B1(n7107), .B2(n6550), .A(n7106), .ZN(n13282) );
  NAND2_X1 U9887 ( .A1(n12253), .A2(n12252), .ZN(n13031) );
  NAND2_X1 U9888 ( .A1(n8768), .A2(n8769), .ZN(n8782) );
  OAI21_X1 U9889 ( .B1(n8659), .B2(n7089), .A(n7088), .ZN(n8653) );
  NAND2_X2 U9890 ( .A1(n12204), .A2(n9480), .ZN(n9510) );
  INV_X1 U9891 ( .A(n8769), .ZN(n8766) );
  OR2_X1 U9892 ( .A1(n9751), .A2(n11048), .ZN(n7096) );
  MUX2_X1 U9893 ( .A(n13867), .B(n13866), .S(n15448), .Z(n13868) );
  NAND2_X1 U9894 ( .A1(n13104), .A2(n9859), .ZN(n15421) );
  NOR2_X1 U9895 ( .A1(n9509), .A2(n10076), .ZN(n7110) );
  NAND2_X1 U9896 ( .A1(n13485), .A2(n13687), .ZN(n7092) );
  NAND2_X1 U9897 ( .A1(n7147), .A2(n12225), .ZN(n13022) );
  NAND2_X1 U9898 ( .A1(n7092), .A2(n6532), .ZN(P2_U3237) );
  NAND2_X1 U9899 ( .A1(n11549), .A2(n11548), .ZN(n15161) );
  NAND4_X1 U9900 ( .A1(n9506), .A2(n9504), .A3(n7096), .A4(n9505), .ZN(n13355)
         );
  INV_X1 U9901 ( .A(n9480), .ZN(n9478) );
  INV_X1 U9902 ( .A(n10570), .ZN(n7135) );
  OR2_X1 U9903 ( .A1(n9811), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9527) );
  CLKBUF_X3 U9904 ( .A(n9751), .Z(n9811) );
  INV_X1 U9905 ( .A(n7100), .ZN(P2_U3528) );
  AOI21_X1 U9906 ( .B1(n13864), .B2(n15454), .A(n7101), .ZN(n7100) );
  NOR2_X1 U9907 ( .A1(n15454), .A2(n7102), .ZN(n7101) );
  NOR2_X1 U9908 ( .A1(n10089), .A2(n15336), .ZN(n7104) );
  NAND2_X1 U9909 ( .A1(n8645), .A2(n8752), .ZN(n8648) );
  NAND2_X1 U9910 ( .A1(n8910), .A2(n8889), .ZN(n8890) );
  NAND2_X1 U9911 ( .A1(n7353), .A2(n7519), .ZN(n8855) );
  NAND2_X1 U9912 ( .A1(n8644), .A2(SI_1_), .ZN(n8749) );
  OAI21_X1 U9913 ( .B1(n8659), .B2(n7139), .A(n7138), .ZN(n8644) );
  NAND2_X1 U9914 ( .A1(n8876), .A2(n8669), .ZN(n8928) );
  NAND2_X2 U9915 ( .A1(n10089), .A2(n7434), .ZN(n9536) );
  INV_X4 U9916 ( .A(n13277), .ZN(n13189) );
  NOR2_X1 U9917 ( .A1(n7881), .A2(n7110), .ZN(n9514) );
  NAND2_X1 U9918 ( .A1(n11690), .A2(n7127), .ZN(n11851) );
  AND2_X2 U9919 ( .A1(n7681), .A2(n9517), .ZN(n9585) );
  INV_X1 U9920 ( .A(n7079), .ZN(n7350) );
  NAND2_X1 U9921 ( .A1(n9278), .A2(n7126), .ZN(n14691) );
  NAND2_X1 U9922 ( .A1(n14691), .A2(n15321), .ZN(n7360) );
  AOI21_X1 U9923 ( .B1(n12137), .B2(n6436), .A(n9276), .ZN(n7126) );
  NAND2_X1 U9924 ( .A1(n14315), .A2(n14317), .ZN(n10668) );
  NOR2_X1 U9925 ( .A1(n6397), .A2(n14586), .ZN(n7433) );
  OAI21_X1 U9926 ( .B1(n8659), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n8642), .ZN(
        n8643) );
  XNOR2_X1 U9927 ( .A(n10486), .B(n15368), .ZN(n15155) );
  NAND2_X1 U9928 ( .A1(n8756), .A2(n8757), .ZN(n9230) );
  NAND2_X1 U9929 ( .A1(n14866), .A2(n14405), .ZN(n14840) );
  NAND2_X1 U9930 ( .A1(n8827), .A2(n6536), .ZN(n7353) );
  OAI21_X1 U9931 ( .B1(n8659), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n7115), .ZN(
        n8646) );
  OAI21_X1 U9932 ( .B1(n14991), .B2(n15289), .A(n14990), .ZN(n15116) );
  NAND2_X1 U9933 ( .A1(n8629), .A2(n7464), .ZN(n15134) );
  NAND4_X1 U9934 ( .A1(n8621), .A2(n8620), .A3(n9060), .A4(n9219), .ZN(n9296)
         );
  NOR2_X1 U9935 ( .A1(n6469), .A2(n7154), .ZN(n7153) );
  INV_X1 U9936 ( .A(n12137), .ZN(n7137) );
  INV_X1 U9937 ( .A(n11450), .ZN(n14180) );
  NAND2_X1 U9938 ( .A1(n9040), .A2(n9039), .ZN(n9058) );
  INV_X1 U9939 ( .A(n14090), .ZN(n10902) );
  NAND2_X1 U9940 ( .A1(n14279), .A2(n14280), .ZN(n14278) );
  INV_X1 U9941 ( .A(n8856), .ZN(n8857) );
  OAI211_X1 U9942 ( .C1(n7614), .C2(n7616), .A(n6506), .B(n7613), .ZN(n7619)
         );
  NAND3_X1 U9943 ( .A1(n14434), .A2(n14433), .A3(n6562), .ZN(n7117) );
  INV_X4 U9944 ( .A(n14448), .ZN(n14485) );
  NAND2_X1 U9945 ( .A1(n10784), .A2(n10783), .ZN(n10782) );
  NAND2_X1 U9946 ( .A1(n7164), .A2(n7163), .ZN(n13170) );
  NAND2_X2 U9947 ( .A1(n7405), .A2(n7407), .ZN(n10781) );
  NAND2_X4 U9948 ( .A1(n8755), .A2(n7434), .ZN(n14466) );
  INV_X2 U9949 ( .A(n10783), .ZN(n14527) );
  NAND2_X1 U9950 ( .A1(n7800), .A2(n9237), .ZN(n7154) );
  NAND2_X1 U9951 ( .A1(n10416), .A2(n10417), .ZN(n10633) );
  INV_X1 U9952 ( .A(n7492), .ZN(n7491) );
  INV_X1 U9953 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7682) );
  NAND2_X1 U9954 ( .A1(n7128), .A2(n13499), .ZN(n13769) );
  NAND2_X1 U9955 ( .A1(n7129), .A2(n13717), .ZN(n7128) );
  XNOR2_X1 U9956 ( .A(n13498), .B(n6723), .ZN(n7129) );
  NAND3_X1 U9957 ( .A1(n9514), .A2(n9513), .A3(n9512), .ZN(n10806) );
  NAND2_X1 U9958 ( .A1(n15121), .A2(n6403), .ZN(n7131) );
  NAND2_X1 U9959 ( .A1(n13117), .A2(n13118), .ZN(n7132) );
  NAND2_X1 U9960 ( .A1(n7631), .A2(n7633), .ZN(n12351) );
  NAND3_X1 U9961 ( .A1(n8589), .A2(n8591), .A3(n7133), .ZN(n8593) );
  NAND2_X1 U9962 ( .A1(n8916), .A2(n8915), .ZN(n15102) );
  AOI21_X2 U9963 ( .B1(n12311), .B2(n12310), .A(n7134), .ZN(n12402) );
  AOI21_X1 U9964 ( .B1(n7421), .B2(n7425), .A(n6438), .ZN(n7420) );
  AND2_X2 U9965 ( .A1(n9481), .A2(n9480), .ZN(n9503) );
  OAI21_X1 U9966 ( .B1(n7500), .B2(n7503), .A(n7507), .ZN(n13498) );
  NAND2_X1 U9967 ( .A1(n7149), .A2(n9259), .ZN(n14901) );
  NAND2_X1 U9968 ( .A1(n8659), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7138) );
  NAND3_X1 U9969 ( .A1(n7144), .A2(n7143), .A3(n14590), .ZN(n14588) );
  INV_X1 U9970 ( .A(n7494), .ZN(n7500) );
  AOI21_X1 U9971 ( .B1(n10204), .B2(n10200), .A(n10324), .ZN(n10201) );
  NOR2_X1 U9972 ( .A1(n7146), .A2(n12251), .ZN(n12252) );
  INV_X1 U9973 ( .A(n10803), .ZN(n7590) );
  NAND2_X1 U9974 ( .A1(n7608), .A2(n7606), .ZN(n11987) );
  INV_X1 U9975 ( .A(n7808), .ZN(n12138) );
  OR2_X1 U9976 ( .A1(n14713), .A2(n7155), .ZN(P1_U3265) );
  NOR2_X1 U9977 ( .A1(n7808), .A2(n14547), .ZN(n14711) );
  NAND2_X1 U9978 ( .A1(n9473), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9863) );
  NAND3_X1 U9979 ( .A1(n7161), .A2(n13767), .A3(n13766), .ZN(n13865) );
  NAND2_X1 U9980 ( .A1(n9497), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7162) );
  NAND2_X1 U9981 ( .A1(n7494), .A2(n7501), .ZN(n7499) );
  OAI21_X2 U9982 ( .B1(n11644), .B2(n7767), .A(n7764), .ZN(n12027) );
  NAND2_X1 U9983 ( .A1(n7779), .A2(n7778), .ZN(n14719) );
  AND2_X1 U9984 ( .A1(n7172), .A2(n10629), .ZN(n10520) );
  NAND2_X1 U9985 ( .A1(n12070), .A2(n7174), .ZN(n7173) );
  NAND2_X1 U9986 ( .A1(n8032), .A2(n7183), .ZN(n7180) );
  NAND2_X1 U9987 ( .A1(n7180), .A2(n7181), .ZN(n11596) );
  NAND2_X1 U9988 ( .A1(n12823), .A2(n7188), .ZN(n7187) );
  NAND2_X1 U9989 ( .A1(n7187), .A2(n6558), .ZN(n7731) );
  OAI22_X1 U9990 ( .A1(n12657), .A2(n7198), .B1(n7197), .B2(n7199), .ZN(n9390)
         );
  OAI21_X1 U9991 ( .B1(n12657), .B2(n12643), .A(n7199), .ZN(n7747) );
  NAND2_X1 U9992 ( .A1(n12657), .A2(n8520), .ZN(n12648) );
  INV_X1 U9993 ( .A(n7201), .ZN(n12703) );
  NAND2_X1 U9994 ( .A1(n7213), .A2(n7215), .ZN(n7208) );
  NOR2_X1 U9995 ( .A1(n11726), .A2(n11864), .ZN(n7217) );
  NAND3_X1 U9996 ( .A1(n11086), .A2(n10966), .A3(n10965), .ZN(n7219) );
  NAND3_X1 U9997 ( .A1(n7222), .A2(n7221), .A3(n9335), .ZN(n7220) );
  NAND2_X1 U9998 ( .A1(n10739), .A2(n9334), .ZN(n7222) );
  NAND2_X1 U9999 ( .A1(n12460), .A2(n10697), .ZN(n7223) );
  NAND3_X1 U10000 ( .A1(n7225), .A2(n7226), .A3(n7822), .ZN(n9354) );
  NAND2_X1 U10001 ( .A1(n12679), .A2(n7227), .ZN(n7225) );
  NOR2_X1 U10002 ( .A1(n7233), .A2(n7237), .ZN(n7236) );
  NAND2_X1 U10003 ( .A1(n12927), .A2(n7235), .ZN(n7234) );
  NOR2_X1 U10004 ( .A1(n12924), .A2(n7380), .ZN(n7235) );
  AND2_X1 U10005 ( .A1(n12924), .A2(n7380), .ZN(n7237) );
  NAND2_X1 U10006 ( .A1(n7251), .A2(n7247), .ZN(n12600) );
  NAND2_X1 U10007 ( .A1(n12532), .A2(n7249), .ZN(n7247) );
  NAND2_X1 U10008 ( .A1(n7254), .A2(n7255), .ZN(n12560) );
  INV_X1 U10009 ( .A(n12561), .ZN(n7253) );
  OAI21_X1 U10010 ( .B1(n10548), .B2(n7264), .A(n7261), .ZN(n11472) );
  OAI211_X1 U10011 ( .C1(n10548), .C2(n7260), .A(n7258), .B(n6538), .ZN(n7257)
         );
  NOR2_X2 U10012 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n7276) );
  NAND4_X1 U10013 ( .A1(n7284), .A2(n7281), .A3(n7279), .A4(n7278), .ZN(n8456)
         );
  NAND3_X1 U10014 ( .A1(n8440), .A2(n7287), .A3(n7282), .ZN(n7281) );
  NAND2_X1 U10015 ( .A1(n7288), .A2(n7289), .ZN(n8484) );
  NAND2_X1 U10016 ( .A1(n8469), .A2(n7291), .ZN(n7288) );
  INV_X1 U10018 ( .A(n7895), .ZN(n7298) );
  OAI21_X1 U10019 ( .B1(n8534), .B2(n7303), .A(n7299), .ZN(n7306) );
  NOR2_X1 U10020 ( .A1(n7304), .A2(n12352), .ZN(n7300) );
  NAND2_X1 U10021 ( .A1(n7306), .A2(n6524), .ZN(n8540) );
  NAND3_X1 U10022 ( .A1(n8517), .A2(n8515), .A3(n8516), .ZN(n7316) );
  NAND2_X1 U10023 ( .A1(n7318), .A2(n7885), .ZN(n7916) );
  NOR2_X1 U10024 ( .A1(n7931), .A2(n7317), .ZN(n10324) );
  INV_X1 U10025 ( .A(n7321), .ZN(n8599) );
  NAND2_X1 U10026 ( .A1(n7321), .A2(n8595), .ZN(n7320) );
  NAND2_X1 U10027 ( .A1(n12398), .A2(n7326), .ZN(n12336) );
  NAND2_X1 U10028 ( .A1(n12399), .A2(n7327), .ZN(n7323) );
  NAND3_X1 U10029 ( .A1(n7323), .A2(n7325), .A3(n7322), .ZN(n12408) );
  NAND3_X1 U10030 ( .A1(n12398), .A2(n7324), .A3(n7326), .ZN(n7325) );
  OAI21_X2 U10031 ( .B1(n10622), .B2(n7328), .A(n10516), .ZN(n10518) );
  AND2_X1 U10032 ( .A1(n7331), .A2(n7151), .ZN(n7700) );
  NAND2_X1 U10033 ( .A1(n9461), .A2(n7331), .ZN(n9463) );
  NOR2_X2 U10034 ( .A1(n9881), .A2(n9460), .ZN(n7331) );
  OAI21_X1 U10035 ( .B1(n13572), .B2(n7531), .A(n7529), .ZN(n13530) );
  NAND2_X1 U10036 ( .A1(n13865), .A2(n15454), .ZN(n7349) );
  NAND2_X1 U10037 ( .A1(n7349), .A2(n7348), .ZN(P2_U3527) );
  INV_X1 U10038 ( .A(n8825), .ZN(n7352) );
  NAND2_X1 U10039 ( .A1(n8908), .A2(n8909), .ZN(n11757) );
  MUX2_X1 U10040 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n9464), .Z(n7369) );
  INV_X2 U10041 ( .A(n7374), .ZN(n14359) );
  NAND2_X1 U10042 ( .A1(n7931), .A2(n7379), .ZN(n10321) );
  XNOR2_X2 U10043 ( .A(n7386), .B(n7385), .ZN(n12577) );
  NAND2_X1 U10044 ( .A1(n7626), .A2(n6557), .ZN(n7389) );
  INV_X1 U10045 ( .A(n14421), .ZN(n7391) );
  INV_X2 U10046 ( .A(n9298), .ZN(n8629) );
  OAI21_X2 U10047 ( .B1(n9299), .B2(n7393), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7392) );
  INV_X1 U10048 ( .A(n7616), .ZN(n7395) );
  NAND3_X1 U10049 ( .A1(n14445), .A2(n14447), .A3(n14444), .ZN(n7394) );
  NOR2_X1 U10050 ( .A1(n14358), .A2(n14357), .ZN(n14361) );
  INV_X1 U10051 ( .A(n14396), .ZN(n7403) );
  INV_X1 U10052 ( .A(n14397), .ZN(n7404) );
  OAI21_X1 U10053 ( .B1(n14336), .B2(n7409), .A(n7408), .ZN(n14342) );
  INV_X1 U10054 ( .A(n14342), .ZN(n14345) );
  NAND2_X1 U10055 ( .A1(n14462), .A2(n14485), .ZN(n7411) );
  NAND2_X1 U10056 ( .A1(n14482), .A2(n14507), .ZN(n7412) );
  NAND2_X1 U10057 ( .A1(n8876), .A2(n7421), .ZN(n7419) );
  NAND2_X1 U10058 ( .A1(n7419), .A2(n7420), .ZN(n8947) );
  NAND2_X1 U10059 ( .A1(n8927), .A2(n8931), .ZN(n7425) );
  OAI21_X2 U10060 ( .B1(n9146), .B2(n9145), .A(n9152), .ZN(n9164) );
  AND3_X2 U10061 ( .A1(n7431), .A2(n7430), .A3(n6397), .ZN(n7432) );
  NOR2_X4 U10062 ( .A1(n7433), .A2(n7432), .ZN(n11204) );
  NOR2_X2 U10063 ( .A1(n15108), .A2(n11760), .ZN(n12033) );
  INV_X1 U10064 ( .A(n7442), .ZN(n14808) );
  NAND2_X1 U10065 ( .A1(n14747), .A2(n6466), .ZN(n14735) );
  INV_X1 U10066 ( .A(n7453), .ZN(n14725) );
  NAND2_X1 U10067 ( .A1(n8629), .A2(n7811), .ZN(n7463) );
  NAND2_X1 U10068 ( .A1(n14158), .A2(n7472), .ZN(n7466) );
  NAND2_X1 U10069 ( .A1(n14158), .A2(n7470), .ZN(n7465) );
  NAND2_X1 U10070 ( .A1(n13355), .A2(n11051), .ZN(n10803) );
  OAI21_X1 U10071 ( .B1(n13305), .B2(n6448), .A(n9829), .ZN(n7492) );
  NAND2_X2 U10072 ( .A1(n7804), .A2(n8724), .ZN(n9228) );
  NOR2_X2 U10073 ( .A1(n10780), .A2(n10781), .ZN(n11506) );
  NAND2_X1 U10074 ( .A1(n8855), .A2(n8666), .ZN(n8874) );
  NAND2_X1 U10075 ( .A1(n7528), .A2(n11860), .ZN(n7527) );
  AOI21_X2 U10076 ( .B1(n7532), .B2(n7530), .A(n6467), .ZN(n7529) );
  INV_X1 U10077 ( .A(n7532), .ZN(n7531) );
  AND2_X4 U10078 ( .A1(n7536), .A2(n7535), .ZN(n8659) );
  NAND4_X1 U10079 ( .A1(n7538), .A2(n7539), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7535) );
  INV_X1 U10080 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U10081 ( .A1(n7544), .A2(n7924), .ZN(n7546) );
  INV_X1 U10082 ( .A(n7933), .ZN(n7544) );
  NAND2_X1 U10083 ( .A1(n7923), .A2(n7545), .ZN(n7547) );
  NAND2_X1 U10084 ( .A1(n7548), .A2(n7924), .ZN(n7950) );
  NAND2_X1 U10085 ( .A1(n8169), .A2(n7561), .ZN(n7560) );
  NAND2_X1 U10086 ( .A1(n7564), .A2(n8126), .ZN(n7565) );
  NAND2_X1 U10087 ( .A1(n8109), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U10088 ( .A1(n7565), .A2(n8129), .ZN(n8146) );
  NAND2_X1 U10089 ( .A1(n8366), .A2(n7571), .ZN(n7566) );
  NAND2_X1 U10090 ( .A1(n8366), .A2(n7575), .ZN(n8379) );
  OAI211_X1 U10091 ( .C1(n8366), .C2(n7573), .A(n7566), .B(n7567), .ZN(n12930)
         );
  NAND2_X1 U10092 ( .A1(n8366), .A2(n8365), .ZN(n8369) );
  NAND2_X1 U10093 ( .A1(n8290), .A2(n7578), .ZN(n7577) );
  NAND2_X1 U10094 ( .A1(n8300), .A2(n8290), .ZN(n8301) );
  NAND2_X1 U10095 ( .A1(n8071), .A2(n8070), .ZN(n8091) );
  OR2_X2 U10096 ( .A1(n13298), .A2(n15421), .ZN(n12272) );
  NAND2_X1 U10097 ( .A1(n11982), .A2(n11739), .ZN(n7607) );
  NAND2_X1 U10098 ( .A1(n11661), .A2(n6470), .ZN(n7608) );
  NAND2_X1 U10099 ( .A1(n11980), .A2(n11981), .ZN(n7609) );
  INV_X1 U10100 ( .A(n14398), .ZN(n7611) );
  NAND2_X1 U10101 ( .A1(n7618), .A2(n7612), .ZN(n7614) );
  NAND2_X1 U10102 ( .A1(n14447), .A2(n14446), .ZN(n7617) );
  NAND2_X1 U10103 ( .A1(n14440), .A2(n14441), .ZN(n14439) );
  NAND2_X1 U10104 ( .A1(n14429), .A2(n14430), .ZN(n14428) );
  NAND2_X1 U10105 ( .A1(n7622), .A2(n7624), .ZN(n14352) );
  NAND3_X1 U10106 ( .A1(n14347), .A2(n7623), .A3(n14346), .ZN(n7622) );
  NAND3_X1 U10107 ( .A1(n14418), .A2(n14417), .A3(n6539), .ZN(n7626) );
  NAND2_X1 U10108 ( .A1(n9223), .A2(n7628), .ZN(n9304) );
  NAND2_X1 U10109 ( .A1(n8756), .A2(n14580), .ZN(n7629) );
  NAND2_X1 U10110 ( .A1(n14472), .A2(n14308), .ZN(n14468) );
  INV_X2 U10111 ( .A(n14448), .ZN(n14483) );
  AND2_X1 U10112 ( .A1(n7629), .A2(n14448), .ZN(n14320) );
  OR2_X1 U10113 ( .A1(n12437), .A2(n12319), .ZN(n7631) );
  NAND2_X1 U10114 ( .A1(n7630), .A2(n7632), .ZN(n12354) );
  NAND2_X1 U10115 ( .A1(n12437), .A2(n7633), .ZN(n7630) );
  NAND2_X1 U10116 ( .A1(n12437), .A2(n12438), .ZN(n12436) );
  OAI21_X2 U10117 ( .B1(n7657), .B2(n7656), .A(n7653), .ZN(n12596) );
  NAND2_X1 U10118 ( .A1(n10636), .A2(n6548), .ZN(n7658) );
  NAND3_X1 U10119 ( .A1(n7658), .A2(n7659), .A3(n6561), .ZN(n7660) );
  INV_X1 U10120 ( .A(n7660), .ZN(n11480) );
  INV_X1 U10121 ( .A(n10541), .ZN(n7668) );
  INV_X1 U10122 ( .A(n10395), .ZN(n7667) );
  OAI211_X1 U10123 ( .C1(n10541), .C2(n7665), .A(n7664), .B(n6559), .ZN(n10882) );
  NAND2_X1 U10124 ( .A1(n12589), .A2(n7671), .ZN(n7670) );
  INV_X1 U10125 ( .A(n12601), .ZN(n7676) );
  OR2_X1 U10126 ( .A1(n12555), .A2(n12761), .ZN(n7680) );
  AND2_X2 U10127 ( .A1(n9499), .A2(n7685), .ZN(n9517) );
  INV_X1 U10128 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7685) );
  INV_X1 U10129 ( .A(n13517), .ZN(n7693) );
  OR2_X2 U10130 ( .A1(n13517), .A2(n13771), .ZN(n13506) );
  NOR2_X1 U10131 ( .A1(n13630), .A2(n7699), .ZN(n13601) );
  NOR2_X2 U10132 ( .A1(n13113), .A2(n11051), .ZN(n10986) );
  AOI21_X1 U10133 ( .B1(n13114), .B2(n13115), .A(n7704), .ZN(n7703) );
  OAI21_X1 U10134 ( .B1(n13114), .B2(n13115), .A(n13300), .ZN(n7706) );
  INV_X1 U10135 ( .A(n13128), .ZN(n7708) );
  OR2_X1 U10136 ( .A1(n7708), .A2(n13127), .ZN(n7709) );
  OR2_X1 U10137 ( .A1(n13135), .A2(n7712), .ZN(n7711) );
  INV_X1 U10138 ( .A(n13134), .ZN(n7712) );
  NAND3_X1 U10139 ( .A1(n13144), .A2(n6549), .A3(n13143), .ZN(n7713) );
  NAND3_X1 U10140 ( .A1(n13163), .A2(n6543), .A3(n13162), .ZN(n7716) );
  NAND2_X1 U10141 ( .A1(n8088), .A2(n7723), .ZN(n7722) );
  NAND2_X1 U10142 ( .A1(n12646), .A2(n7745), .ZN(n7741) );
  NAND2_X1 U10143 ( .A1(n7741), .A2(n7743), .ZN(n9429) );
  INV_X1 U10144 ( .A(n12192), .ZN(n7756) );
  INV_X1 U10145 ( .A(n8466), .ZN(n7760) );
  NAND2_X1 U10146 ( .A1(n12744), .A2(n7847), .ZN(n7762) );
  NAND2_X1 U10147 ( .A1(n9228), .A2(n11204), .ZN(n14315) );
  AND3_X2 U10148 ( .A1(n8617), .A2(n8618), .A3(n8809), .ZN(n7788) );
  AOI21_X1 U10149 ( .B1(n6446), .B2(n7794), .A(n7796), .ZN(P1_U3524) );
  AOI21_X1 U10150 ( .B1(n6446), .B2(n7795), .A(n7799), .ZN(P1_U3556) );
  NAND2_X1 U10151 ( .A1(n9235), .A2(n15281), .ZN(n7800) );
  INV_X1 U10152 ( .A(n7883), .ZN(n7801) );
  AND3_X2 U10153 ( .A1(n8721), .A2(n8722), .A3(n8723), .ZN(n7804) );
  OAI21_X2 U10154 ( .B1(n14732), .B2(n7060), .A(n7805), .ZN(n7808) );
  OAI21_X1 U10155 ( .B1(n10739), .B2(n6461), .A(n9334), .ZN(n11085) );
  NOR2_X2 U10156 ( .A1(n8056), .A2(n7890), .ZN(n7820) );
  NAND2_X1 U10157 ( .A1(n10951), .A2(n7828), .ZN(n7827) );
  NAND2_X1 U10158 ( .A1(n9355), .A2(n7873), .ZN(n7841) );
  NAND2_X1 U10159 ( .A1(n9355), .A2(n7832), .ZN(n7831) );
  NAND2_X1 U10160 ( .A1(n12714), .A2(n9347), .ZN(n7849) );
  NAND2_X1 U10161 ( .A1(n12828), .A2(n12759), .ZN(n7850) );
  NAND2_X1 U10162 ( .A1(n9342), .A2(n9341), .ZN(n11593) );
  NOR2_X1 U10163 ( .A1(n9344), .A2(n7858), .ZN(n7857) );
  INV_X1 U10164 ( .A(n9341), .ZN(n7858) );
  OAI21_X1 U10165 ( .B1(n13326), .B2(n7874), .A(n13288), .ZN(n13335) );
  NAND2_X1 U10166 ( .A1(n13326), .A2(n13287), .ZN(n13288) );
  INV_X1 U10167 ( .A(n14998), .ZN(n14755) );
  INV_X1 U10168 ( .A(n14689), .ZN(n14983) );
  NAND2_X1 U10169 ( .A1(n8108), .A2(n15539), .ZN(n8126) );
  NAND2_X1 U10170 ( .A1(n12765), .A2(n8491), .ZN(n12756) );
  NAND2_X1 U10171 ( .A1(n8364), .A2(n8363), .ZN(n8366) );
  OAI21_X1 U10172 ( .B1(n14332), .B2(n14331), .A(n14330), .ZN(n14334) );
  AND2_X1 U10173 ( .A1(n9870), .A2(n10088), .ZN(n13723) );
  OR2_X1 U10174 ( .A1(n9479), .A2(n10077), .ZN(n9528) );
  OR2_X1 U10175 ( .A1(n9136), .A2(n11327), .ZN(n8733) );
  OAI21_X1 U10176 ( .B1(n13471), .B2(n9861), .A(n13717), .ZN(n9874) );
  NAND2_X1 U10177 ( .A1(n9874), .A2(n9873), .ZN(n13487) );
  INV_X1 U10178 ( .A(n14691), .ZN(n14707) );
  NAND2_X1 U10179 ( .A1(n9209), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8743) );
  NOR2_X1 U10180 ( .A1(n12464), .A2(n12465), .ZN(n12492) );
  NAND2_X1 U10181 ( .A1(n15476), .A2(n12461), .ZN(n8421) );
  NAND2_X2 U10182 ( .A1(n12125), .A2(n8602), .ZN(n7918) );
  INV_X1 U10183 ( .A(n14841), .ZN(n14842) );
  INV_X1 U10184 ( .A(n12313), .ZN(n12863) );
  INV_X1 U10185 ( .A(n12340), .ZN(n12871) );
  AND2_X1 U10186 ( .A1(n11813), .A2(n11812), .ZN(n7860) );
  NAND2_X2 U10187 ( .A1(n11288), .A2(n15460), .ZN(n15472) );
  INV_X1 U10188 ( .A(n15514), .ZN(n9433) );
  INV_X2 U10189 ( .A(n15509), .ZN(n15510) );
  AND3_X1 U10190 ( .A1(n8571), .A2(n7301), .A3(n8570), .ZN(n7861) );
  INV_X1 U10191 ( .A(n13717), .ZN(n13701) );
  NAND2_X1 U10192 ( .A1(n15045), .A2(n15034), .ZN(n7862) );
  AND2_X1 U10193 ( .A1(n14131), .A2(n10286), .ZN(n7863) );
  OR2_X1 U10194 ( .A1(n14549), .A2(n9277), .ZN(n7864) );
  OR2_X1 U10195 ( .A1(n15327), .A2(n9324), .ZN(n7865) );
  OR2_X1 U10196 ( .A1(n14710), .A2(n14566), .ZN(n7867) );
  AND2_X1 U10197 ( .A1(n12300), .A2(n12452), .ZN(n7868) );
  AND2_X1 U10198 ( .A1(n12141), .A2(n6530), .ZN(n7869) );
  AND2_X1 U10199 ( .A1(n14850), .A2(n15043), .ZN(n7871) );
  AND2_X1 U10200 ( .A1(n14543), .A2(n14407), .ZN(n7872) );
  OR2_X1 U10201 ( .A1(n12449), .A2(n12645), .ZN(n7873) );
  AND2_X1 U10202 ( .A1(n13283), .A2(n13433), .ZN(n7874) );
  OR2_X1 U10203 ( .A1(n11233), .A2(n11232), .ZN(P1_U3291) );
  AND2_X1 U10204 ( .A1(n7434), .A2(P3_U3151), .ZN(n10509) );
  INV_X1 U10205 ( .A(n9870), .ZN(n10094) );
  OR2_X1 U10206 ( .A1(n11198), .A2(n9419), .ZN(n15323) );
  OR2_X1 U10207 ( .A1(n10275), .A2(n9419), .ZN(n15331) );
  INV_X1 U10208 ( .A(n15312), .ZN(n15107) );
  OR2_X1 U10209 ( .A1(n15269), .A2(n15289), .ZN(n14978) );
  NAND2_X1 U10210 ( .A1(n9281), .A2(n14111), .ZN(n15289) );
  AND2_X1 U10211 ( .A1(n13136), .A2(n11239), .ZN(n7877) );
  NOR2_X1 U10212 ( .A1(n13267), .A2(n13272), .ZN(n7878) );
  OR2_X1 U10213 ( .A1(n12406), .A2(n12668), .ZN(n7879) );
  AND2_X1 U10214 ( .A1(n12379), .A2(n12748), .ZN(n7880) );
  INV_X1 U10215 ( .A(n14547), .ZN(n12129) );
  NOR2_X1 U10216 ( .A1(n9751), .A2(n13370), .ZN(n7881) );
  NOR4_X1 U10217 ( .A1(n14542), .A2(n14827), .A3(n14541), .A4(n14865), .ZN(
        n7882) );
  AND2_X1 U10218 ( .A1(n15294), .A2(n15293), .ZN(n7884) );
  NAND2_X1 U10219 ( .A1(n14334), .A2(n14333), .ZN(n14336) );
  NAND2_X1 U10220 ( .A1(n14432), .A2(n14431), .ZN(n14433) );
  INV_X1 U10221 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8628) );
  INV_X1 U10222 ( .A(n12682), .ZN(n9350) );
  AND2_X1 U10223 ( .A1(n10966), .A2(n10965), .ZN(n9335) );
  INV_X1 U10224 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8581) );
  NOR2_X1 U10225 ( .A1(n12246), .A2(n12972), .ZN(n12251) );
  INV_X1 U10226 ( .A(n10806), .ZN(n9524) );
  OR2_X1 U10227 ( .A1(n9836), .A2(n9835), .ZN(n9841) );
  INV_X1 U10228 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8990) );
  INV_X1 U10229 ( .A(n11362), .ZN(n10513) );
  INV_X1 U10230 ( .A(n8256), .ZN(n8257) );
  INV_X1 U10231 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9724) );
  INV_X1 U10232 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n15549) );
  AOI21_X1 U10233 ( .B1(n9228), .B2(n14108), .A(n7863), .ZN(n10655) );
  OR2_X1 U10234 ( .A1(n14449), .A2(n14697), .ZN(n9201) );
  AOI21_X1 U10235 ( .B1(n7367), .B2(n9258), .A(n9257), .ZN(n9259) );
  INV_X1 U10236 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n15530) );
  INV_X1 U10237 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U10238 ( .A1(n7900), .A2(n8659), .ZN(n8642) );
  INV_X1 U10239 ( .A(n12781), .ZN(n11864) );
  INV_X1 U10240 ( .A(n11191), .ZN(n11188) );
  INV_X1 U10241 ( .A(n11719), .ZN(n11720) );
  INV_X1 U10242 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8157) );
  INV_X1 U10243 ( .A(n11564), .ZN(n11081) );
  INV_X1 U10244 ( .A(n12224), .ZN(n12225) );
  INV_X1 U10245 ( .A(n13762), .ZN(n13465) );
  INV_X1 U10246 ( .A(n13449), .ZN(n13476) );
  XNOR2_X1 U10247 ( .A(n13353), .B(n13119), .ZN(n13299) );
  INV_X1 U10248 ( .A(n9875), .ZN(n9877) );
  AND2_X1 U10249 ( .A1(n12175), .A2(n7866), .ZN(n12176) );
  NOR2_X1 U10250 ( .A1(n13993), .A2(n13992), .ZN(n13994) );
  OR2_X1 U10251 ( .A1(n10278), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9312) );
  INV_X1 U10252 ( .A(n14865), .ZN(n9050) );
  INV_X1 U10253 ( .A(n14304), .ZN(n9283) );
  AND2_X1 U10254 ( .A1(n8598), .A2(n8597), .ZN(n8600) );
  NAND2_X1 U10255 ( .A1(n10526), .A2(n10253), .ZN(n12429) );
  INV_X1 U10256 ( .A(n11927), .ZN(n12012) );
  INV_X1 U10257 ( .A(n15455), .ZN(n12581) );
  AND2_X1 U10258 ( .A1(n10137), .A2(n10128), .ZN(n10132) );
  NAND2_X1 U10259 ( .A1(n12620), .A2(n12704), .ZN(n12621) );
  INV_X1 U10260 ( .A(n12711), .ZN(n12739) );
  AND2_X1 U10261 ( .A1(n8458), .A2(n8459), .ZN(n11281) );
  INV_X1 U10262 ( .A(n12704), .ZN(n15467) );
  AND2_X1 U10263 ( .A1(n9408), .A2(n9357), .ZN(n15484) );
  INV_X1 U10264 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12924) );
  INV_X1 U10265 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13034) );
  OR2_X1 U10266 ( .A1(n10819), .A2(n13329), .ZN(n13074) );
  OR2_X1 U10267 ( .A1(n10819), .A2(n10818), .ZN(n10821) );
  INV_X1 U10268 ( .A(n9811), .ZN(n12282) );
  XNOR2_X1 U10269 ( .A(n13491), .B(n13476), .ZN(n13450) );
  OR2_X1 U10270 ( .A1(n10812), .A2(n9870), .ZN(n13676) );
  INV_X1 U10271 ( .A(n10815), .ZN(n9906) );
  INV_X1 U10272 ( .A(n13723), .ZN(n13678) );
  INV_X1 U10273 ( .A(n14567), .ZN(n14311) );
  INV_X1 U10274 ( .A(n14574), .ZN(n14360) );
  INV_X1 U10275 ( .A(n13994), .ZN(n13995) );
  OR2_X1 U10276 ( .A1(n14298), .A2(n15312), .ZN(n14227) );
  NAND2_X1 U10277 ( .A1(n14554), .A2(n9283), .ZN(n11201) );
  OR2_X1 U10278 ( .A1(n14753), .A2(n9136), .ZN(n8639) );
  AND2_X1 U10279 ( .A1(n10280), .A2(n10279), .ZN(n11199) );
  OR2_X1 U10280 ( .A1(n15269), .A2(n15310), .ZN(n14969) );
  INV_X1 U10281 ( .A(n14804), .ZN(n15017) );
  OR2_X1 U10282 ( .A1(n10001), .A2(n10282), .ZN(n10297) );
  INV_X1 U10283 ( .A(n8824), .ZN(n8826) );
  NAND2_X1 U10284 ( .A1(n8600), .A2(n9367), .ZN(n10233) );
  INV_X1 U10285 ( .A(n12443), .ZN(n12427) );
  AOI21_X1 U10286 ( .B1(n12613), .B2(n8355), .A(n8349), .ZN(n9426) );
  INV_X1 U10287 ( .A(n12597), .ZN(n12578) );
  AND2_X1 U10288 ( .A1(n10132), .A2(n12937), .ZN(n12607) );
  INV_X1 U10289 ( .A(n12726), .ZN(n12787) );
  INV_X1 U10290 ( .A(n12821), .ZN(n12840) );
  INV_X1 U10291 ( .A(n12843), .ZN(n12836) );
  AND2_X1 U10292 ( .A1(n9406), .A2(n9383), .ZN(n10625) );
  AND2_X1 U10293 ( .A1(n11357), .A2(n11347), .ZN(n12797) );
  INV_X1 U10294 ( .A(n12797), .ZN(n15501) );
  NAND2_X1 U10295 ( .A1(n9369), .A2(n9368), .ZN(n10621) );
  AND2_X1 U10296 ( .A1(n8198), .A2(n8182), .ZN(n8196) );
  OR2_X1 U10297 ( .A1(n13519), .A2(n9811), .ZN(n9817) );
  NAND2_X1 U10298 ( .A1(n10099), .A2(n10096), .ZN(n15395) );
  INV_X1 U10299 ( .A(n13430), .ZN(n15403) );
  INV_X1 U10300 ( .A(n13475), .ZN(n13470) );
  INV_X1 U10301 ( .A(n13676), .ZN(n13722) );
  OR2_X1 U10302 ( .A1(n13105), .A2(n9860), .ZN(n13717) );
  INV_X1 U10303 ( .A(n13549), .ZN(n13708) );
  NAND2_X1 U10304 ( .A1(n15416), .A2(n10820), .ZN(n13683) );
  INV_X1 U10305 ( .A(n13838), .ZN(n13789) );
  AND2_X1 U10306 ( .A1(n11267), .A2(n15422), .ZN(n13855) );
  INV_X1 U10307 ( .A(n13855), .ZN(n13835) );
  AND2_X1 U10308 ( .A1(n10972), .A2(n10814), .ZN(n10713) );
  AND2_X1 U10309 ( .A1(n9893), .A2(n9907), .ZN(n15412) );
  AND2_X1 U10310 ( .A1(n9463), .A2(n9887), .ZN(n9907) );
  AND2_X1 U10311 ( .A1(n9559), .A2(n9574), .ZN(n10268) );
  INV_X1 U10312 ( .A(n14295), .ZN(n14286) );
  OR2_X1 U10313 ( .A1(n14478), .A2(n10155), .ZN(n15310) );
  INV_X1 U10314 ( .A(n14298), .ZN(n14288) );
  OR2_X1 U10315 ( .A1(n14478), .A2(n9286), .ZN(n15312) );
  OR2_X1 U10316 ( .A1(n14059), .A2(n9136), .ZN(n9179) );
  INV_X1 U10317 ( .A(n14668), .ZN(n15210) );
  INV_X1 U10318 ( .A(n15277), .ZN(n15308) );
  AND2_X1 U10319 ( .A1(n14693), .A2(n15236), .ZN(n15260) );
  INV_X1 U10320 ( .A(n14906), .ZN(n14879) );
  OR2_X1 U10321 ( .A1(n14558), .A2(n9418), .ZN(n10275) );
  AND2_X1 U10322 ( .A1(n14305), .A2(n14308), .ZN(n15277) );
  INV_X1 U10323 ( .A(n15289), .ZN(n15321) );
  OR2_X1 U10324 ( .A1(n14558), .A2(n10293), .ZN(n11198) );
  NAND2_X1 U10325 ( .A1(n10041), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10001) );
  AND2_X1 U10326 ( .A1(n10137), .A2(n10136), .ZN(n15455) );
  INV_X1 U10327 ( .A(n12686), .ZN(n12873) );
  INV_X1 U10328 ( .A(n12414), .ZN(n12448) );
  NAND2_X1 U10329 ( .A1(n10245), .A2(n10252), .ZN(n12434) );
  INV_X1 U10330 ( .A(n12645), .ZN(n12620) );
  INV_X1 U10331 ( .A(n12749), .ZN(n12452) );
  INV_X1 U10332 ( .A(n12607), .ZN(n12024) );
  INV_X1 U10333 ( .A(n12590), .ZN(n12566) );
  OR2_X1 U10334 ( .A1(n11288), .A2(n10628), .ZN(n12726) );
  NAND2_X1 U10335 ( .A1(n15472), .A2(n15471), .ZN(n12790) );
  NAND2_X1 U10336 ( .A1(n15514), .A2(n15501), .ZN(n12843) );
  AND2_X2 U10337 ( .A1(n10625), .A2(n9388), .ZN(n15514) );
  NAND2_X1 U10338 ( .A1(n15510), .A2(n15501), .ZN(n12919) );
  NAND2_X1 U10339 ( .A1(n9413), .A2(n10252), .ZN(n15509) );
  INV_X1 U10340 ( .A(n12915), .ZN(n12894) );
  INV_X1 U10341 ( .A(SI_24_), .ZN(n11899) );
  INV_X1 U10342 ( .A(SI_19_), .ZN(n10874) );
  INV_X1 U10343 ( .A(SI_13_), .ZN(n10071) );
  INV_X1 U10344 ( .A(n11470), .ZN(n11479) );
  INV_X1 U10345 ( .A(n13804), .ZN(n13606) );
  NAND2_X1 U10346 ( .A1(n10858), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13085) );
  INV_X1 U10347 ( .A(n15405), .ZN(n11894) );
  INV_X1 U10348 ( .A(n13649), .ZN(n13735) );
  INV_X1 U10349 ( .A(n10996), .ZN(n11256) );
  NAND2_X1 U10350 ( .A1(n13687), .A2(n11046), .ZN(n13738) );
  NAND2_X1 U10351 ( .A1(n15454), .A2(n13851), .ZN(n13838) );
  INV_X1 U10352 ( .A(n15454), .ZN(n15452) );
  INV_X1 U10353 ( .A(n13587), .ZN(n13887) );
  NAND2_X1 U10354 ( .A1(n15448), .A2(n13851), .ZN(n13900) );
  INV_X1 U10355 ( .A(n15448), .ZN(n15446) );
  AND2_X2 U10356 ( .A1(n10974), .A2(n10713), .ZN(n15448) );
  NOR2_X1 U10357 ( .A1(n15419), .A2(n15412), .ZN(n15413) );
  INV_X1 U10358 ( .A(n15413), .ZN(n15515) );
  INV_X1 U10359 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13240) );
  INV_X1 U10360 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11671) );
  INV_X1 U10361 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10571) );
  INV_X1 U10362 ( .A(n14790), .ZN(n15021) );
  OR2_X1 U10363 ( .A1(n14298), .A2(n15310), .ZN(n14272) );
  INV_X1 U10364 ( .A(n15045), .ZN(n14855) );
  INV_X1 U10365 ( .A(n14042), .ZN(n14569) );
  INV_X1 U10366 ( .A(n15061), .ZN(n14858) );
  OR2_X1 U10367 ( .A1(n10156), .A2(n10064), .ZN(n14668) );
  OR2_X1 U10368 ( .A1(n10156), .A2(n10155), .ZN(n15221) );
  NAND2_X1 U10369 ( .A1(n10063), .A2(n10061), .ZN(n15226) );
  AND2_X1 U10370 ( .A1(n12148), .A2(n12147), .ZN(n15008) );
  INV_X1 U10371 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11496) );
  INV_X1 U10372 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10686) );
  AND2_X2 U10373 ( .A1(n9915), .A2(n12922), .ZN(P3_U3897) );
  NOR3_X1 U10374 ( .A1(n10093), .A2(n10092), .A3(P2_U3088), .ZN(P2_U3947) );
  INV_X1 U10375 ( .A(n14600), .ZN(P1_U4016) );
  NOR2_X1 U10376 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n7889) );
  NOR2_X1 U10377 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n7888) );
  NOR2_X1 U10378 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n7887) );
  NAND4_X1 U10379 ( .A1(n7889), .A2(n7888), .A3(n7887), .A4(n8581), .ZN(n7890)
         );
  NAND2_X1 U10380 ( .A1(n8590), .A2(n8580), .ZN(n7891) );
  INV_X1 U10382 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10536) );
  OR2_X1 U10383 ( .A1(n8390), .A2(n7317), .ZN(n7898) );
  INV_X1 U10384 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10632) );
  OR2_X1 U10385 ( .A1(n7982), .A2(n10632), .ZN(n7897) );
  OAI21_X1 U10386 ( .B1(P2_DATAO_REG_0__SCAN_IN), .B2(n7900), .A(n7919), .ZN(
        n7902) );
  MUX2_X1 U10387 ( .A(n7902), .B(SI_0_), .S(n7434), .Z(n12951) );
  MUX2_X1 U10388 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12951), .S(n7918), .Z(n10629)
         );
  NAND2_X2 U10389 ( .A1(n7918), .A2(n9464), .ZN(n8171) );
  XNOR2_X1 U10390 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7921) );
  XNOR2_X1 U10391 ( .A(n7919), .B(n7921), .ZN(n9930) );
  OR2_X1 U10392 ( .A1(n8171), .A2(n9930), .ZN(n7906) );
  INV_X1 U10393 ( .A(SI_1_), .ZN(n9931) );
  OR2_X1 U10394 ( .A1(n7918), .A2(n10321), .ZN(n7904) );
  NAND2_X1 U10395 ( .A1(n8386), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7911) );
  INV_X1 U10396 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n7907) );
  INV_X1 U10397 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10527) );
  OR2_X1 U10398 ( .A1(n7982), .A2(n10527), .ZN(n7909) );
  INV_X1 U10399 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15491) );
  OR2_X1 U10400 ( .A1(n8390), .A2(n15491), .ZN(n7908) );
  NAND2_X1 U10402 ( .A1(n8386), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7915) );
  OR2_X1 U10403 ( .A1(n7982), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n7914) );
  OR2_X1 U10404 ( .A1(n8372), .A2(n10743), .ZN(n7913) );
  INV_X1 U10405 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10391) );
  OR2_X1 U10406 ( .A1(n8390), .A2(n10391), .ZN(n7912) );
  NAND2_X1 U10407 ( .A1(n7916), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7917) );
  XNOR2_X1 U10408 ( .A(n7917), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10455) );
  INV_X1 U10409 ( .A(n7919), .ZN(n7920) );
  NAND2_X1 U10410 ( .A1(n7921), .A2(n7920), .ZN(n7923) );
  INV_X1 U10411 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U10412 ( .A1(n9926), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7922) );
  XNOR2_X1 U10413 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7933) );
  NAND2_X1 U10414 ( .A1(n9927), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7924) );
  XNOR2_X1 U10415 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7949) );
  XNOR2_X1 U10416 ( .A(n7950), .B(n7949), .ZN(n9923) );
  OR2_X1 U10417 ( .A1(n8171), .A2(n9923), .ZN(n7926) );
  OR2_X1 U10418 ( .A1(n8382), .A2(SI_3_), .ZN(n7925) );
  OAI211_X1 U10419 ( .C1(n10455), .C2(n7918), .A(n7926), .B(n7925), .ZN(n11412) );
  NAND2_X1 U10420 ( .A1(n8386), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7930) );
  INV_X1 U10421 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15459) );
  OR2_X1 U10422 ( .A1(n7982), .A2(n15459), .ZN(n7929) );
  INV_X1 U10423 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10329) );
  OR2_X1 U10424 ( .A1(n8372), .A2(n10329), .ZN(n7928) );
  INV_X1 U10425 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15474) );
  OR2_X1 U10426 ( .A1(n8390), .A2(n15474), .ZN(n7927) );
  NAND4_X2 U10427 ( .A1(n7930), .A2(n7929), .A3(n7928), .A4(n7927), .ZN(n15480) );
  XNOR2_X1 U10428 ( .A(n7932), .B(n7933), .ZN(n9919) );
  OR2_X1 U10429 ( .A1(n8171), .A2(n9919), .ZN(n7935) );
  OR2_X1 U10430 ( .A1(n8382), .A2(SI_2_), .ZN(n7934) );
  OAI211_X1 U10431 ( .C1(n6399), .C2(n7918), .A(n7935), .B(n7934), .ZN(n15458)
         );
  NAND2_X1 U10432 ( .A1(n15480), .A2(n15458), .ZN(n8430) );
  AND2_X1 U10433 ( .A1(n8555), .A2(n8430), .ZN(n8432) );
  NAND2_X1 U10434 ( .A1(n15457), .A2(n8432), .ZN(n7939) );
  INV_X1 U10435 ( .A(n8555), .ZN(n7936) );
  OR2_X1 U10436 ( .A1(n15480), .A2(n15458), .ZN(n10736) );
  OR2_X1 U10437 ( .A1(n10836), .A2(n11412), .ZN(n8556) );
  INV_X1 U10438 ( .A(n7937), .ZN(n7938) );
  NAND2_X1 U10439 ( .A1(n7939), .A2(n7938), .ZN(n10829) );
  NAND2_X1 U10440 ( .A1(n7997), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7948) );
  INV_X1 U10441 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n7940) );
  OR2_X1 U10442 ( .A1(n7960), .A2(n7940), .ZN(n7947) );
  NAND2_X1 U10443 ( .A1(n7963), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n7943) );
  AND2_X1 U10444 ( .A1(n7980), .A2(n7943), .ZN(n11091) );
  OR2_X1 U10445 ( .A1(n8080), .A2(n11091), .ZN(n7946) );
  INV_X1 U10446 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n7944) );
  OR2_X1 U10447 ( .A1(n8372), .A2(n7944), .ZN(n7945) );
  NAND4_X1 U10448 ( .A1(n7948), .A2(n7947), .A3(n7946), .A4(n7945), .ZN(n12459) );
  INV_X1 U10449 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U10450 ( .A1(n9925), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10451 ( .A1(n9977), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7952) );
  XNOR2_X1 U10452 ( .A(n7988), .B(n7987), .ZN(n9921) );
  OR2_X1 U10453 ( .A1(n8171), .A2(n9921), .ZN(n7958) );
  OR2_X1 U10454 ( .A1(n8382), .A2(SI_5_), .ZN(n7957) );
  INV_X1 U10455 ( .A(n7968), .ZN(n7954) );
  NAND2_X1 U10456 ( .A1(n7954), .A2(n7953), .ZN(n8057) );
  NAND2_X1 U10457 ( .A1(n8057), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7955) );
  XNOR2_X1 U10458 ( .A(n7955), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10412) );
  OR2_X1 U10459 ( .A1(n7918), .A2(n10412), .ZN(n7956) );
  INV_X1 U10460 ( .A(n11093), .ZN(n11129) );
  NAND2_X1 U10461 ( .A1(n12459), .A2(n11129), .ZN(n8441) );
  INV_X1 U10462 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n7959) );
  INV_X1 U10463 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n7961) );
  OR2_X1 U10464 ( .A1(n7960), .A2(n7961), .ZN(n7966) );
  NAND2_X1 U10465 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7962) );
  AND2_X1 U10466 ( .A1(n7963), .A2(n7962), .ZN(n11405) );
  INV_X1 U10467 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10409) );
  OR2_X1 U10468 ( .A1(n8372), .A2(n10409), .ZN(n7964) );
  NAND2_X1 U10469 ( .A1(n7968), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7969) );
  MUX2_X1 U10470 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7969), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7970) );
  NAND2_X1 U10471 ( .A1(n7970), .A2(n8057), .ZN(n10410) );
  INV_X1 U10472 ( .A(n10410), .ZN(n10443) );
  OR2_X1 U10473 ( .A1(n8382), .A2(SI_4_), .ZN(n7974) );
  XNOR2_X1 U10474 ( .A(n7971), .B(n7972), .ZN(n9917) );
  OR2_X1 U10475 ( .A1(n8171), .A2(n9917), .ZN(n7973) );
  OAI211_X1 U10476 ( .C1(n10443), .C2(n7918), .A(n7974), .B(n7973), .ZN(n11406) );
  NAND2_X1 U10477 ( .A1(n12460), .A2(n11406), .ZN(n8442) );
  NAND2_X1 U10478 ( .A1(n10829), .A2(n7975), .ZN(n7979) );
  INV_X1 U10479 ( .A(n8441), .ZN(n7976) );
  OR2_X1 U10480 ( .A1(n12459), .A2(n11129), .ZN(n8448) );
  OAI21_X1 U10481 ( .B1(n7976), .B2(n11082), .A(n8448), .ZN(n7977) );
  INV_X1 U10482 ( .A(n7977), .ZN(n7978) );
  NAND2_X1 U10483 ( .A1(n7979), .A2(n7978), .ZN(n10963) );
  NAND2_X1 U10484 ( .A1(n7997), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7986) );
  INV_X1 U10485 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15518) );
  OR2_X1 U10486 ( .A1(n7960), .A2(n15518), .ZN(n7985) );
  NAND2_X1 U10487 ( .A1(n7980), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7981) );
  AND2_X1 U10488 ( .A1(n8000), .A2(n7981), .ZN(n11098) );
  OR2_X1 U10489 ( .A1(n8080), .A2(n11098), .ZN(n7984) );
  INV_X1 U10490 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10401) );
  OR2_X1 U10491 ( .A1(n8372), .A2(n10401), .ZN(n7983) );
  NAND2_X1 U10492 ( .A1(n7988), .A2(n7987), .ZN(n7991) );
  INV_X1 U10493 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10494 ( .A1(n7989), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7990) );
  XNOR2_X1 U10495 ( .A(n9975), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7992) );
  XNOR2_X1 U10496 ( .A(n8007), .B(n7992), .ZN(n9928) );
  OR2_X1 U10497 ( .A1(n9928), .A2(n8171), .ZN(n7996) );
  INV_X1 U10498 ( .A(SI_6_), .ZN(n9929) );
  OR2_X1 U10499 ( .A1(n6612), .A2(n9929), .ZN(n7995) );
  NAND2_X1 U10500 ( .A1(n8010), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10501 ( .A1(n8217), .A2(n10640), .ZN(n7994) );
  OR2_X1 U10502 ( .A1(n12458), .A2(n11121), .ZN(n8450) );
  NAND2_X1 U10503 ( .A1(n12458), .A2(n11121), .ZN(n8449) );
  INV_X1 U10504 ( .A(n10966), .ZN(n10962) );
  NAND2_X1 U10505 ( .A1(n10963), .A2(n10962), .ZN(n10961) );
  NAND2_X1 U10506 ( .A1(n10961), .A2(n8450), .ZN(n10949) );
  NAND2_X1 U10507 ( .A1(n7997), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U10508 ( .A1(n8000), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8001) );
  AND2_X1 U10509 ( .A1(n8018), .A2(n8001), .ZN(n11418) );
  OR2_X1 U10510 ( .A1(n8080), .A2(n11418), .ZN(n8004) );
  INV_X1 U10511 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8002) );
  OR2_X1 U10512 ( .A1(n8372), .A2(n8002), .ZN(n8003) );
  NAND4_X1 U10513 ( .A1(n8006), .A2(n8005), .A3(n8004), .A4(n8003), .ZN(n12457) );
  NAND2_X1 U10514 ( .A1(n9979), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8008) );
  XNOR2_X1 U10515 ( .A(n8026), .B(n8025), .ZN(n9935) );
  NAND2_X1 U10516 ( .A1(n9935), .A2(n8381), .ZN(n8016) );
  INV_X1 U10517 ( .A(SI_7_), .ZN(n9934) );
  INV_X1 U10518 ( .A(n8010), .ZN(n8012) );
  NAND2_X1 U10519 ( .A1(n8012), .A2(n8011), .ZN(n8028) );
  NAND2_X1 U10520 ( .A1(n8028), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8014) );
  XNOR2_X1 U10521 ( .A(n8014), .B(n8013), .ZN(n10878) );
  AOI22_X1 U10522 ( .A1(n8218), .A2(n9934), .B1(n8217), .B2(n10878), .ZN(n8015) );
  NAND2_X1 U10523 ( .A1(n8016), .A2(n8015), .ZN(n11419) );
  NAND2_X1 U10524 ( .A1(n12457), .A2(n11419), .ZN(n8454) );
  INV_X1 U10525 ( .A(n11164), .ZN(n10948) );
  NAND2_X1 U10526 ( .A1(n10949), .A2(n10948), .ZN(n10947) );
  NAND2_X1 U10527 ( .A1(n10947), .A2(n8453), .ZN(n11278) );
  NAND2_X1 U10528 ( .A1(n7997), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8024) );
  INV_X1 U10529 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8017) );
  OR2_X1 U10530 ( .A1(n7960), .A2(n8017), .ZN(n8023) );
  NAND2_X1 U10531 ( .A1(n8018), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8019) );
  AND2_X1 U10532 ( .A1(n8044), .A2(n8019), .ZN(n11432) );
  OR2_X1 U10533 ( .A1(n8080), .A2(n11432), .ZN(n8022) );
  INV_X1 U10534 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n8020) );
  OR2_X1 U10535 ( .A1(n8372), .A2(n8020), .ZN(n8021) );
  NAND4_X1 U10536 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8021), .ZN(n12456) );
  NAND2_X1 U10537 ( .A1(n9994), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8027) );
  XNOR2_X1 U10538 ( .A(n7094), .B(P1_DATAO_REG_8__SCAN_IN), .ZN(n8033) );
  XNOR2_X1 U10539 ( .A(n8035), .B(n8033), .ZN(n9965) );
  NAND2_X1 U10540 ( .A1(n9965), .A2(n8381), .ZN(n8031) );
  NAND2_X1 U10541 ( .A1(n8038), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8029) );
  AOI22_X1 U10542 ( .A1(n8218), .A2(SI_8_), .B1(n11470), .B2(n8217), .ZN(n8030) );
  NAND2_X1 U10543 ( .A1(n8031), .A2(n8030), .ZN(n11436) );
  OR2_X1 U10544 ( .A1(n11353), .A2(n11436), .ZN(n8458) );
  NAND2_X1 U10545 ( .A1(n11353), .A2(n11436), .ZN(n8459) );
  NAND2_X1 U10546 ( .A1(n11278), .A2(n11281), .ZN(n8032) );
  INV_X1 U10547 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U10548 ( .A1(n7094), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10549 ( .A1(n8037), .A2(n8036), .ZN(n8053) );
  XNOR2_X1 U10550 ( .A(n8053), .B(n8052), .ZN(n9964) );
  NAND2_X1 U10551 ( .A1(n9964), .A2(n8381), .ZN(n8042) );
  OAI21_X1 U10552 ( .B1(n8038), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8040) );
  XNOR2_X1 U10553 ( .A(n8040), .B(n8039), .ZN(n11486) );
  INV_X1 U10554 ( .A(SI_9_), .ZN(n9963) );
  AOI22_X1 U10555 ( .A1(n11486), .A2(n8217), .B1(n8218), .B2(n9963), .ZN(n8041) );
  NAND2_X1 U10556 ( .A1(n8042), .A2(n8041), .ZN(n11570) );
  NAND2_X1 U10557 ( .A1(n7997), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8049) );
  INV_X1 U10558 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15628) );
  OR2_X1 U10559 ( .A1(n7960), .A2(n15628), .ZN(n8048) );
  NAND2_X1 U10560 ( .A1(n8044), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8045) );
  AND2_X1 U10561 ( .A1(n8062), .A2(n8045), .ZN(n11192) );
  OR2_X1 U10562 ( .A1(n8080), .A2(n11192), .ZN(n8047) );
  INV_X1 U10563 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11568) );
  OR2_X1 U10564 ( .A1(n8372), .A2(n11568), .ZN(n8046) );
  NAND2_X1 U10565 ( .A1(n11570), .A2(n11365), .ZN(n8050) );
  OR2_X1 U10566 ( .A1(n11570), .A2(n11365), .ZN(n8051) );
  NAND2_X1 U10567 ( .A1(n8053), .A2(n8052), .ZN(n8055) );
  NAND2_X1 U10568 ( .A1(n10043), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U10569 ( .A1(n8055), .A2(n8054), .ZN(n8069) );
  XNOR2_X1 U10570 ( .A(n8069), .B(n8068), .ZN(n9974) );
  NAND2_X1 U10571 ( .A1(n9974), .A2(n8381), .ZN(n8061) );
  OAI21_X1 U10572 ( .B1(n8057), .B2(n8056), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8059) );
  XNOR2_X1 U10573 ( .A(n8059), .B(n8058), .ZN(n11917) );
  AOI22_X1 U10574 ( .A1(n8218), .A2(n9973), .B1(n8217), .B2(n11917), .ZN(n8060) );
  NAND2_X1 U10575 ( .A1(n8061), .A2(n8060), .ZN(n11677) );
  NAND2_X1 U10576 ( .A1(n7997), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8067) );
  INV_X1 U10577 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11369) );
  OR2_X1 U10578 ( .A1(n7960), .A2(n11369), .ZN(n8066) );
  NAND2_X1 U10579 ( .A1(n8062), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8063) );
  AND2_X1 U10580 ( .A1(n8081), .A2(n8063), .ZN(n11617) );
  OR2_X1 U10581 ( .A1(n8080), .A2(n11617), .ZN(n8065) );
  INV_X1 U10582 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11673) );
  OR2_X1 U10583 ( .A1(n8372), .A2(n11673), .ZN(n8064) );
  NAND4_X1 U10584 ( .A1(n8067), .A2(n8066), .A3(n8065), .A4(n8064), .ZN(n12455) );
  OR2_X1 U10585 ( .A1(n11677), .A2(n12455), .ZN(n8466) );
  NAND2_X1 U10586 ( .A1(n11677), .A2(n12455), .ZN(n8467) );
  INV_X1 U10587 ( .A(n11596), .ZN(n8088) );
  NAND2_X1 U10588 ( .A1(n7098), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8070) );
  XNOR2_X1 U10589 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .ZN(n8072) );
  XNOR2_X1 U10590 ( .A(n8091), .B(n8072), .ZN(n9992) );
  NAND2_X1 U10591 ( .A1(n9992), .A2(n8381), .ZN(n8079) );
  INV_X1 U10592 ( .A(n8591), .ZN(n8074) );
  NAND2_X1 U10593 ( .A1(n8074), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8075) );
  MUX2_X1 U10594 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8075), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n8077) );
  NAND2_X1 U10595 ( .A1(n8591), .A2(n8076), .ZN(n8113) );
  NAND2_X1 U10596 ( .A1(n8077), .A2(n8113), .ZN(n11927) );
  AOI22_X1 U10597 ( .A1(n8218), .A2(n9991), .B1(n8217), .B2(n11927), .ZN(n8078) );
  NAND2_X1 U10598 ( .A1(n8081), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10599 ( .A1(n8100), .A2(n8082), .ZN(n11788) );
  NAND2_X1 U10600 ( .A1(n8355), .A2(n11788), .ZN(n8086) );
  INV_X1 U10601 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11786) );
  OR2_X1 U10602 ( .A1(n8390), .A2(n11786), .ZN(n8085) );
  INV_X1 U10603 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n11599) );
  OR2_X1 U10604 ( .A1(n7960), .A2(n11599), .ZN(n8084) );
  INV_X1 U10605 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n12001) );
  OR2_X1 U10606 ( .A1(n8372), .A2(n12001), .ZN(n8083) );
  NAND2_X1 U10607 ( .A1(n11787), .A2(n11955), .ZN(n8473) );
  NAND2_X1 U10608 ( .A1(n8470), .A2(n8473), .ZN(n11595) );
  NAND2_X1 U10609 ( .A1(n10425), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10610 ( .A1(n10151), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10611 ( .A1(n15618), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10612 ( .A1(n8106), .A2(n8092), .ZN(n8093) );
  NAND2_X1 U10613 ( .A1(n8094), .A2(n8093), .ZN(n8095) );
  NAND2_X1 U10614 ( .A1(n8107), .A2(n8095), .ZN(n9998) );
  OR2_X1 U10615 ( .A1(n9998), .A2(n8171), .ZN(n8098) );
  NAND2_X1 U10616 ( .A1(n8113), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8096) );
  XNOR2_X1 U10617 ( .A(n8096), .B(P3_IR_REG_12__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U10618 ( .A1(n8218), .A2(SI_12_), .B1(n8217), .B2(n12021), .ZN(
        n8097) );
  NAND2_X1 U10619 ( .A1(n8100), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U10620 ( .A1(n8118), .A2(n8101), .ZN(n11961) );
  NAND2_X1 U10621 ( .A1(n8355), .A2(n11961), .ZN(n8105) );
  INV_X1 U10622 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n11964) );
  OR2_X1 U10623 ( .A1(n7960), .A2(n11964), .ZN(n8104) );
  INV_X1 U10624 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12004) );
  OR2_X1 U10625 ( .A1(n8390), .A2(n12004), .ZN(n8103) );
  INV_X1 U10626 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11958) );
  OR2_X1 U10627 ( .A1(n8372), .A2(n11958), .ZN(n8102) );
  NAND2_X1 U10628 ( .A1(n11909), .A2(n12454), .ZN(n8474) );
  INV_X1 U10629 ( .A(n8110), .ZN(n8111) );
  NAND2_X1 U10630 ( .A1(n8111), .A2(n10274), .ZN(n8112) );
  NAND2_X1 U10631 ( .A1(n8127), .A2(n8112), .ZN(n10070) );
  OR2_X1 U10632 ( .A1(n10070), .A2(n8171), .ZN(n8116) );
  NAND2_X1 U10633 ( .A1(n8586), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8114) );
  XNOR2_X1 U10634 ( .A(n8114), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U10635 ( .A1(n8218), .A2(SI_13_), .B1(n8217), .B2(n12498), .ZN(
        n8115) );
  INV_X1 U10636 ( .A(n12110), .ZN(n11726) );
  NAND2_X1 U10637 ( .A1(n8118), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10638 ( .A1(n8140), .A2(n8119), .ZN(n12109) );
  NAND2_X1 U10639 ( .A1(n8355), .A2(n12109), .ZN(n8123) );
  NAND2_X1 U10640 ( .A1(n7997), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8122) );
  INV_X1 U10641 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12074) );
  OR2_X1 U10642 ( .A1(n7960), .A2(n12074), .ZN(n8121) );
  INV_X1 U10643 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15554) );
  OR2_X1 U10644 ( .A1(n8372), .A2(n15554), .ZN(n8120) );
  NAND4_X1 U10645 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), .ZN(n12781) );
  NAND2_X1 U10646 ( .A1(n11726), .A2(n12781), .ZN(n8124) );
  NAND2_X1 U10647 ( .A1(n12110), .A2(n11864), .ZN(n8125) );
  NAND2_X1 U10648 ( .A1(n10539), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10649 ( .A1(n10571), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8128) );
  OR2_X1 U10650 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  NAND2_X1 U10651 ( .A1(n8146), .A2(n8131), .ZN(n10272) );
  NAND2_X1 U10652 ( .A1(n10272), .A2(n8381), .ZN(n8137) );
  INV_X1 U10653 ( .A(n8586), .ZN(n8133) );
  NAND2_X1 U10654 ( .A1(n8133), .A2(n8132), .ZN(n8148) );
  NAND2_X1 U10655 ( .A1(n8148), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8135) );
  INV_X1 U10656 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8134) );
  XNOR2_X1 U10657 ( .A(n8135), .B(n8134), .ZN(n12505) );
  AOI22_X1 U10658 ( .A1(n8217), .A2(n12505), .B1(n8218), .B2(n10271), .ZN(
        n8136) );
  NAND2_X1 U10659 ( .A1(n8386), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U10660 ( .A1(n8385), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8138) );
  AND2_X1 U10661 ( .A1(n8139), .A2(n8138), .ZN(n8144) );
  NAND2_X1 U10662 ( .A1(n8140), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10663 ( .A1(n8158), .A2(n8141), .ZN(n12786) );
  NAND2_X1 U10664 ( .A1(n12786), .A2(n8355), .ZN(n8143) );
  NAND2_X1 U10665 ( .A1(n7997), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10666 ( .A1(n12916), .A2(n12058), .ZN(n8480) );
  INV_X1 U10667 ( .A(n12916), .ZN(n11871) );
  NAND2_X1 U10668 ( .A1(n11871), .A2(n12769), .ZN(n8479) );
  NAND2_X1 U10669 ( .A1(n8480), .A2(n8479), .ZN(n12778) );
  INV_X1 U10670 ( .A(n12778), .ZN(n12779) );
  NAND2_X1 U10671 ( .A1(n8146), .A2(n8145), .ZN(n8164) );
  NAND2_X1 U10672 ( .A1(n10826), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10673 ( .A1(n10827), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10674 ( .A1(n8165), .A2(n8147), .ZN(n8162) );
  XNOR2_X1 U10675 ( .A(n8164), .B(n8162), .ZN(n10475) );
  NAND2_X1 U10676 ( .A1(n10475), .A2(n8381), .ZN(n8156) );
  NAND2_X1 U10677 ( .A1(n8150), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8149) );
  MUX2_X1 U10678 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8149), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n8153) );
  INV_X1 U10679 ( .A(n8150), .ZN(n8152) );
  INV_X1 U10680 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10681 ( .A1(n8152), .A2(n8151), .ZN(n8183) );
  NAND2_X1 U10682 ( .A1(n8153), .A2(n8183), .ZN(n12531) );
  OAI22_X1 U10683 ( .A1(n12531), .A2(n7918), .B1(n6612), .B2(n10477), .ZN(
        n8154) );
  INV_X1 U10684 ( .A(n8154), .ZN(n8155) );
  INV_X1 U10685 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12835) );
  NAND2_X1 U10686 ( .A1(n8158), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10687 ( .A1(n8175), .A2(n8159), .ZN(n12773) );
  NAND2_X1 U10688 ( .A1(n12773), .A2(n8355), .ZN(n8161) );
  AOI22_X1 U10689 ( .A1(n7997), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n8386), .B2(
        P3_REG0_REG_15__SCAN_IN), .ZN(n8160) );
  OAI211_X1 U10690 ( .C1(n8372), .C2(n12835), .A(n8161), .B(n8160), .ZN(n12782) );
  OR2_X1 U10691 ( .A1(n12908), .A2(n12383), .ZN(n8486) );
  NAND2_X1 U10692 ( .A1(n12908), .A2(n12383), .ZN(n8491) );
  NAND2_X1 U10693 ( .A1(n12766), .A2(n12767), .ZN(n12765) );
  INV_X1 U10694 ( .A(n8162), .ZN(n8163) );
  NAND2_X1 U10695 ( .A1(n8164), .A2(n8163), .ZN(n8166) );
  NAND2_X1 U10696 ( .A1(n8166), .A2(n8165), .ZN(n8169) );
  NAND2_X1 U10697 ( .A1(n10569), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10698 ( .A1(n10618), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8167) );
  OR2_X1 U10699 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  NAND2_X1 U10700 ( .A1(n8181), .A2(n8170), .ZN(n10511) );
  OR2_X1 U10701 ( .A1(n10511), .A2(n8171), .ZN(n8174) );
  NAND2_X1 U10702 ( .A1(n8183), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8172) );
  XNOR2_X1 U10703 ( .A(n8172), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U10704 ( .A1(n12555), .A2(n8217), .B1(n8218), .B2(SI_16_), .ZN(
        n8173) );
  INV_X1 U10705 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U10706 ( .A1(n8175), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8176) );
  NAND2_X1 U10707 ( .A1(n8189), .A2(n8176), .ZN(n12762) );
  NAND2_X1 U10708 ( .A1(n12762), .A2(n8355), .ZN(n8178) );
  AOI22_X1 U10709 ( .A1(n7997), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n8386), .B2(
        P3_REG0_REG_16__SCAN_IN), .ZN(n8177) );
  XNOR2_X1 U10710 ( .A(n12902), .B(n12770), .ZN(n12757) );
  NAND2_X1 U10711 ( .A1(n12756), .A2(n12757), .ZN(n8179) );
  NAND2_X1 U10712 ( .A1(n12902), .A2(n12748), .ZN(n8492) );
  NAND2_X1 U10713 ( .A1(n8179), .A2(n8492), .ZN(n12744) );
  NAND2_X1 U10714 ( .A1(n10686), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U10715 ( .A1(n10760), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8182) );
  XNOR2_X1 U10716 ( .A(n8197), .B(n8196), .ZN(n10684) );
  NAND2_X1 U10717 ( .A1(n10684), .A2(n8381), .ZN(n8188) );
  NAND2_X1 U10718 ( .A1(n8200), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8185) );
  NOR2_X1 U10719 ( .A1(n6612), .A2(SI_17_), .ZN(n8186) );
  AOI21_X1 U10720 ( .B1(n12576), .B2(n8217), .A(n8186), .ZN(n8187) );
  NAND2_X1 U10721 ( .A1(n8189), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10722 ( .A1(n8205), .A2(n8190), .ZN(n12750) );
  NAND2_X1 U10723 ( .A1(n12750), .A2(n8355), .ZN(n8195) );
  INV_X1 U10724 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12752) );
  NAND2_X1 U10725 ( .A1(n8385), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U10726 ( .A1(n8386), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8191) );
  OAI211_X1 U10727 ( .C1(n8390), .C2(n12752), .A(n8192), .B(n8191), .ZN(n8193)
         );
  INV_X1 U10728 ( .A(n8193), .ZN(n8194) );
  XNOR2_X1 U10729 ( .A(n12392), .B(n12759), .ZN(n12745) );
  OR2_X1 U10730 ( .A1(n12392), .A2(n12759), .ZN(n8420) );
  NAND2_X1 U10731 ( .A1(n15608), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8213) );
  INV_X1 U10732 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11172) );
  NAND2_X1 U10733 ( .A1(n11172), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8199) );
  XNOR2_X1 U10734 ( .A(n8212), .B(n6566), .ZN(n10841) );
  NAND2_X1 U10735 ( .A1(n10841), .A2(n8381), .ZN(n8204) );
  OAI21_X1 U10736 ( .B1(n8200), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8201) );
  XNOR2_X1 U10737 ( .A(n8201), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12599) );
  NOR2_X1 U10738 ( .A1(n6612), .A2(n10844), .ZN(n8202) );
  AOI21_X1 U10739 ( .B1(n12599), .B2(n8217), .A(n8202), .ZN(n8203) );
  INV_X1 U10740 ( .A(n8222), .ZN(n8223) );
  NAND2_X1 U10741 ( .A1(n8205), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U10742 ( .A1(n8223), .A2(n8206), .ZN(n12734) );
  NAND2_X1 U10743 ( .A1(n12734), .A2(n8355), .ZN(n8211) );
  INV_X1 U10744 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12735) );
  NAND2_X1 U10745 ( .A1(n8385), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U10746 ( .A1(n8386), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8207) );
  OAI211_X1 U10747 ( .C1(n8390), .C2(n12735), .A(n8208), .B(n8207), .ZN(n8209)
         );
  INV_X1 U10748 ( .A(n8209), .ZN(n8210) );
  NAND2_X1 U10749 ( .A1(n12738), .A2(n12749), .ZN(n8498) );
  INV_X1 U10750 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U10751 ( .A1(n11235), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8231) );
  INV_X1 U10752 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11234) );
  NAND2_X1 U10753 ( .A1(n11234), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8214) );
  XNOR2_X1 U10754 ( .A(n8230), .B(n8229), .ZN(n10873) );
  NAND2_X1 U10755 ( .A1(n10873), .A2(n8381), .ZN(n8220) );
  AOI22_X1 U10756 ( .A1(n8218), .A2(n10874), .B1(n12596), .B2(n8217), .ZN(
        n8219) );
  NAND2_X1 U10757 ( .A1(n8223), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U10758 ( .A1(n8235), .A2(n8224), .ZN(n12724) );
  INV_X1 U10759 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12721) );
  NAND2_X1 U10760 ( .A1(n8385), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10761 ( .A1(n8386), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8225) );
  OAI211_X1 U10762 ( .C1(n8390), .C2(n12721), .A(n8226), .B(n8225), .ZN(n8227)
         );
  AOI21_X1 U10763 ( .B1(n12724), .B2(n8355), .A(n8227), .ZN(n12430) );
  NAND2_X1 U10764 ( .A1(n12893), .A2(n12732), .ZN(n8552) );
  INV_X1 U10765 ( .A(n8552), .ZN(n8228) );
  NAND2_X1 U10766 ( .A1(n8232), .A2(n8231), .ZN(n8258) );
  XNOR2_X1 U10767 ( .A(n8258), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8242) );
  XNOR2_X1 U10768 ( .A(n8242), .B(n11374), .ZN(n11360) );
  NAND2_X1 U10769 ( .A1(n11360), .A2(n8381), .ZN(n8234) );
  OR2_X1 U10770 ( .A1(n6612), .A2(n11363), .ZN(n8233) );
  NAND2_X1 U10771 ( .A1(n8235), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U10772 ( .A1(n8251), .A2(n8236), .ZN(n12708) );
  NAND2_X1 U10773 ( .A1(n12708), .A2(n8355), .ZN(n8241) );
  INV_X1 U10774 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12707) );
  INV_X1 U10775 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n15579) );
  OR2_X1 U10776 ( .A1(n8372), .A2(n15579), .ZN(n8238) );
  INV_X1 U10777 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n15630) );
  OR2_X1 U10778 ( .A1(n7960), .A2(n15630), .ZN(n8237) );
  OAI211_X1 U10779 ( .C1(n8390), .C2(n12707), .A(n8238), .B(n8237), .ZN(n8239)
         );
  INV_X1 U10780 ( .A(n8239), .ZN(n8240) );
  INV_X1 U10781 ( .A(n8242), .ZN(n8243) );
  NAND2_X1 U10782 ( .A1(n8243), .A2(n11374), .ZN(n8245) );
  NAND2_X1 U10783 ( .A1(n8258), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10784 ( .A1(n8245), .A2(n8244), .ZN(n8247) );
  INV_X1 U10785 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11499) );
  NAND2_X1 U10786 ( .A1(n11499), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8259) );
  INV_X1 U10787 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11498) );
  NAND2_X1 U10788 ( .A1(n11498), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10789 ( .A1(n8259), .A2(n8260), .ZN(n8246) );
  XNOR2_X1 U10790 ( .A(n8247), .B(n8246), .ZN(n11563) );
  NAND2_X1 U10791 ( .A1(n11563), .A2(n8381), .ZN(n8249) );
  INV_X1 U10792 ( .A(SI_21_), .ZN(n11566) );
  OR2_X1 U10793 ( .A1(n6612), .A2(n11566), .ZN(n8248) );
  NAND2_X1 U10794 ( .A1(n8251), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U10795 ( .A1(n8265), .A2(n8252), .ZN(n12698) );
  INV_X1 U10796 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U10797 ( .A1(n8385), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10798 ( .A1(n8386), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8253) );
  OAI211_X1 U10799 ( .C1(n8390), .C2(n12697), .A(n8254), .B(n8253), .ZN(n8255)
         );
  NAND2_X1 U10800 ( .A1(n12879), .A2(n12681), .ZN(n8510) );
  OR2_X1 U10801 ( .A1(n12879), .A2(n12681), .ZN(n8509) );
  NAND3_X1 U10802 ( .A1(n8259), .A2(P1_DATAO_REG_20__SCAN_IN), .A3(n11374), 
        .ZN(n8261) );
  AND2_X1 U10803 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  XNOR2_X1 U10804 ( .A(n11671), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8273) );
  XNOR2_X1 U10805 ( .A(n8272), .B(n8273), .ZN(n11263) );
  NAND2_X1 U10806 ( .A1(n11263), .A2(n8381), .ZN(n8264) );
  INV_X1 U10807 ( .A(SI_22_), .ZN(n8703) );
  OR2_X1 U10808 ( .A1(n6612), .A2(n8703), .ZN(n8263) );
  NAND2_X1 U10809 ( .A1(n8265), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10810 ( .A1(n8277), .A2(n8266), .ZN(n12685) );
  NAND2_X1 U10811 ( .A1(n12685), .A2(n8355), .ZN(n8271) );
  INV_X1 U10812 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12684) );
  NAND2_X1 U10813 ( .A1(n8385), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U10814 ( .A1(n8386), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8267) );
  OAI211_X1 U10815 ( .C1(n8390), .C2(n12684), .A(n8268), .B(n8267), .ZN(n8269)
         );
  INV_X1 U10816 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U10817 ( .A1(n11671), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8274) );
  XNOR2_X1 U10818 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8286) );
  XNOR2_X1 U10819 ( .A(n8287), .B(n8286), .ZN(n11516) );
  NAND2_X1 U10820 ( .A1(n11516), .A2(n8381), .ZN(n8276) );
  INV_X1 U10821 ( .A(SI_23_), .ZN(n11519) );
  OR2_X1 U10822 ( .A1(n6612), .A2(n11519), .ZN(n8275) );
  NAND2_X1 U10823 ( .A1(n8277), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U10824 ( .A1(n6499), .A2(n8278), .ZN(n12671) );
  NAND2_X1 U10825 ( .A1(n12671), .A2(n8355), .ZN(n8284) );
  INV_X1 U10826 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10827 ( .A1(n8385), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U10828 ( .A1(n8386), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8279) );
  OAI211_X1 U10829 ( .C1(n8390), .C2(n8281), .A(n8280), .B(n8279), .ZN(n8282)
         );
  INV_X1 U10830 ( .A(n8282), .ZN(n8283) );
  NAND2_X1 U10831 ( .A1(n12340), .A2(n12682), .ZN(n8518) );
  NAND2_X1 U10832 ( .A1(n8285), .A2(n8518), .ZN(n12666) );
  INV_X1 U10833 ( .A(n12666), .ZN(n8516) );
  INV_X1 U10834 ( .A(n8285), .ZN(n8519) );
  INV_X1 U10835 ( .A(n8289), .ZN(n8288) );
  INV_X1 U10836 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U10837 ( .A1(n8289), .A2(n11996), .ZN(n8290) );
  INV_X1 U10838 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15647) );
  XNOR2_X1 U10839 ( .A(n8301), .B(n15647), .ZN(n11896) );
  NAND2_X1 U10840 ( .A1(n11896), .A2(n8381), .ZN(n8292) );
  OR2_X1 U10841 ( .A1(n6612), .A2(n11899), .ZN(n8291) );
  NAND2_X1 U10842 ( .A1(n6499), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10843 ( .A1(n8307), .A2(n8293), .ZN(n12659) );
  NAND2_X1 U10844 ( .A1(n12659), .A2(n8355), .ZN(n8299) );
  INV_X1 U10845 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10846 ( .A1(n8385), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10847 ( .A1(n8386), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8294) );
  OAI211_X1 U10848 ( .C1(n8390), .C2(n8296), .A(n8295), .B(n8294), .ZN(n8297)
         );
  INV_X1 U10849 ( .A(n8297), .ZN(n8298) );
  NAND2_X1 U10850 ( .A1(n8299), .A2(n8298), .ZN(n12668) );
  OR2_X1 U10851 ( .A1(n12406), .A2(n12644), .ZN(n8521) );
  NAND2_X1 U10852 ( .A1(n12406), .A2(n12644), .ZN(n8520) );
  INV_X1 U10853 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13917) );
  XNOR2_X1 U10854 ( .A(n13917), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8302) );
  XNOR2_X1 U10855 ( .A(n8315), .B(n8302), .ZN(n12945) );
  NAND2_X1 U10856 ( .A1(n12945), .A2(n8381), .ZN(n8304) );
  INV_X1 U10857 ( .A(SI_25_), .ZN(n12946) );
  OR2_X1 U10858 ( .A1(n6612), .A2(n12946), .ZN(n8303) );
  INV_X1 U10859 ( .A(n8307), .ZN(n8306) );
  INV_X1 U10860 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U10861 ( .A1(n8307), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U10862 ( .A1(n8320), .A2(n8308), .ZN(n12649) );
  NAND2_X1 U10863 ( .A1(n12649), .A2(n8355), .ZN(n8313) );
  INV_X1 U10864 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n15575) );
  NAND2_X1 U10865 ( .A1(n7997), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U10866 ( .A1(n8386), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8309) );
  OAI211_X1 U10867 ( .C1(n15575), .C2(n8372), .A(n8310), .B(n8309), .ZN(n8311)
         );
  INV_X1 U10868 ( .A(n8311), .ZN(n8312) );
  OR2_X1 U10869 ( .A1(n12313), .A2(n12656), .ZN(n8526) );
  NAND2_X1 U10870 ( .A1(n12313), .A2(n12656), .ZN(n8527) );
  NAND2_X1 U10871 ( .A1(n8526), .A2(n8527), .ZN(n12643) );
  INV_X1 U10872 ( .A(n12643), .ZN(n12647) );
  NAND2_X1 U10873 ( .A1(n13917), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8314) );
  INV_X1 U10874 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15145) );
  NAND2_X1 U10875 ( .A1(n15145), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8316) );
  XNOR2_X1 U10876 ( .A(n11945), .B(P1_DATAO_REG_26__SCAN_IN), .ZN(n8317) );
  XNOR2_X1 U10877 ( .A(n8329), .B(n8317), .ZN(n12940) );
  NAND2_X1 U10878 ( .A1(n12940), .A2(n8381), .ZN(n8319) );
  OR2_X1 U10879 ( .A1(n6612), .A2(n12942), .ZN(n8318) );
  NAND2_X1 U10880 ( .A1(n8320), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10881 ( .A1(n8334), .A2(n8321), .ZN(n12640) );
  NAND2_X1 U10882 ( .A1(n12640), .A2(n8355), .ZN(n8326) );
  INV_X1 U10883 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n15617) );
  NAND2_X1 U10884 ( .A1(n7997), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10885 ( .A1(n8386), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8322) );
  OAI211_X1 U10886 ( .C1(n15617), .C2(n8372), .A(n8323), .B(n8322), .ZN(n8324)
         );
  INV_X1 U10887 ( .A(n8324), .ZN(n8325) );
  AND2_X1 U10888 ( .A1(n11945), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8328) );
  INV_X1 U10889 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U10890 ( .A1(n11948), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8327) );
  XNOR2_X1 U10891 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8330) );
  XNOR2_X1 U10892 ( .A(n8341), .B(n8330), .ZN(n12936) );
  NAND2_X1 U10893 ( .A1(n12936), .A2(n8381), .ZN(n8332) );
  INV_X1 U10894 ( .A(SI_27_), .ZN(n12939) );
  OR2_X1 U10895 ( .A1(n6612), .A2(n12939), .ZN(n8331) );
  INV_X1 U10896 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U10897 ( .A1(n8345), .A2(n8335), .ZN(n12627) );
  INV_X1 U10898 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n15563) );
  NAND2_X1 U10899 ( .A1(n7997), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10900 ( .A1(n8385), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8336) );
  OAI211_X1 U10901 ( .C1(n7960), .C2(n15563), .A(n8337), .B(n8336), .ZN(n8338)
         );
  NAND2_X1 U10902 ( .A1(n12793), .A2(n12357), .ZN(n9391) );
  AND2_X1 U10903 ( .A1(n15530), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8340) );
  INV_X1 U10904 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15143) );
  INV_X1 U10905 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12205) );
  XNOR2_X1 U10906 ( .A(n12205), .B(P1_DATAO_REG_28__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U10907 ( .A1(n12123), .A2(n8381), .ZN(n8344) );
  INV_X1 U10908 ( .A(SI_28_), .ZN(n12126) );
  OR2_X1 U10909 ( .A1(n6612), .A2(n12126), .ZN(n8343) );
  NAND2_X1 U10910 ( .A1(n8345), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U10911 ( .A1(n12143), .A2(n8346), .ZN(n12613) );
  INV_X1 U10912 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U10913 ( .A1(n8386), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10914 ( .A1(n8385), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8347) );
  OAI211_X1 U10915 ( .C1(n12612), .C2(n8390), .A(n8348), .B(n8347), .ZN(n8349)
         );
  INV_X1 U10916 ( .A(n9429), .ZN(n8361) );
  AND2_X1 U10917 ( .A1(n12205), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8351) );
  INV_X1 U10918 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U10919 ( .A1(n9186), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8350) );
  XNOR2_X1 U10920 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8363) );
  XNOR2_X1 U10921 ( .A(n8362), .B(n8363), .ZN(n12932) );
  NAND2_X1 U10922 ( .A1(n12932), .A2(n8381), .ZN(n8354) );
  INV_X1 U10923 ( .A(SI_29_), .ZN(n12935) );
  OR2_X1 U10924 ( .A1(n6612), .A2(n12935), .ZN(n8353) );
  INV_X1 U10925 ( .A(n12143), .ZN(n8356) );
  NAND2_X1 U10926 ( .A1(n8356), .A2(n8355), .ZN(n8393) );
  INV_X1 U10927 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U10928 ( .A1(n8386), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10929 ( .A1(n7997), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8357) );
  OAI211_X1 U10930 ( .C1(n9430), .C2(n8372), .A(n8358), .B(n8357), .ZN(n8359)
         );
  INV_X1 U10931 ( .A(n8359), .ZN(n8360) );
  NAND2_X1 U10932 ( .A1(n8361), .A2(n8544), .ZN(n8410) );
  INV_X1 U10933 ( .A(n8362), .ZN(n8364) );
  INV_X1 U10934 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12289) );
  NAND2_X1 U10935 ( .A1(n12289), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8365) );
  INV_X1 U10936 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n15631) );
  NAND2_X1 U10937 ( .A1(n15631), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8378) );
  INV_X1 U10938 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U10939 ( .A1(n14465), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10940 ( .A1(n8378), .A2(n8367), .ZN(n8368) );
  NAND2_X1 U10941 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  NAND2_X1 U10942 ( .A1(n8379), .A2(n8370), .ZN(n12206) );
  INV_X1 U10943 ( .A(SI_30_), .ZN(n12208) );
  INV_X1 U10944 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10945 ( .A1(n8386), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8374) );
  INV_X1 U10946 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n8371) );
  OR2_X1 U10947 ( .A1(n8372), .A2(n8371), .ZN(n8373) );
  OAI211_X1 U10948 ( .C1(n8390), .C2(n8375), .A(n8374), .B(n8373), .ZN(n8376)
         );
  INV_X1 U10949 ( .A(n8376), .ZN(n8377) );
  NAND2_X1 U10950 ( .A1(n8393), .A2(n8377), .ZN(n12450) );
  INV_X1 U10951 ( .A(n12450), .ZN(n8541) );
  XNOR2_X1 U10952 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8380) );
  NAND2_X1 U10953 ( .A1(n12930), .A2(n8381), .ZN(n8384) );
  INV_X1 U10954 ( .A(SI_31_), .ZN(n12925) );
  OR2_X1 U10955 ( .A1(n6612), .A2(n12925), .ZN(n8383) );
  AOI21_X1 U10956 ( .B1(n12848), .B2(n8541), .A(n8542), .ZN(n8395) );
  NAND2_X1 U10957 ( .A1(n12850), .A2(n12355), .ZN(n8543) );
  INV_X1 U10958 ( .A(n8543), .ZN(n8394) );
  INV_X1 U10959 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10960 ( .A1(n8385), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10961 ( .A1(n8386), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8387) );
  OAI211_X1 U10962 ( .C1(n8390), .C2(n8389), .A(n8388), .B(n8387), .ZN(n8391)
         );
  INV_X1 U10963 ( .A(n8391), .ZN(n8392) );
  NAND2_X1 U10964 ( .A1(n8393), .A2(n8392), .ZN(n12451) );
  INV_X1 U10965 ( .A(n8414), .ZN(n8545) );
  NOR4_X1 U10966 ( .A1(n8395), .A2(n12593), .A3(n8394), .A4(n8545), .ZN(n8409)
         );
  NAND2_X1 U10967 ( .A1(n12848), .A2(n8543), .ZN(n8403) );
  NOR2_X1 U10968 ( .A1(n8542), .A2(n12596), .ZN(n8412) );
  OAI21_X1 U10969 ( .B1(n12450), .B2(n8403), .A(n8412), .ZN(n8407) );
  NAND2_X1 U10970 ( .A1(n8416), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10971 ( .A1(n8397), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8398) );
  MUX2_X1 U10972 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8398), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8399) );
  NAND2_X1 U10973 ( .A1(n11081), .A2(n10513), .ZN(n9357) );
  INV_X1 U10974 ( .A(n9357), .ZN(n8406) );
  NAND2_X1 U10975 ( .A1(n12848), .A2(n12451), .ZN(n8546) );
  NAND2_X1 U10976 ( .A1(n8546), .A2(n12450), .ZN(n8400) );
  NAND3_X1 U10977 ( .A1(n8400), .A2(n8542), .A3(n12596), .ZN(n8405) );
  AND2_X1 U10978 ( .A1(n12450), .A2(n12593), .ZN(n8401) );
  AND2_X1 U10979 ( .A1(n8546), .A2(n8401), .ZN(n8413) );
  NAND2_X1 U10980 ( .A1(n8543), .A2(n12451), .ZN(n8402) );
  NAND3_X1 U10981 ( .A1(n8413), .A2(n8403), .A3(n8402), .ZN(n8404) );
  NAND4_X1 U10982 ( .A1(n8407), .A2(n8406), .A3(n8405), .A4(n8404), .ZN(n8408)
         );
  AOI21_X1 U10983 ( .B1(n8410), .B2(n8409), .A(n8408), .ZN(n8579) );
  INV_X1 U10984 ( .A(n8410), .ZN(n8411) );
  OAI21_X1 U10985 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8578) );
  AND2_X1 U10986 ( .A1(n8546), .A2(n8414), .ZN(n8571) );
  INV_X1 U10987 ( .A(n8532), .ZN(n8415) );
  INV_X1 U10988 ( .A(n12633), .ZN(n12636) );
  AND2_X1 U10989 ( .A1(n8418), .A2(n9385), .ZN(n8419) );
  NAND2_X1 U10990 ( .A1(n8552), .A2(n8419), .ZN(n8501) );
  INV_X1 U10991 ( .A(n8420), .ZN(n8497) );
  OR2_X1 U10992 ( .A1(n11570), .A2(n11431), .ZN(n9339) );
  INV_X1 U10993 ( .A(n9339), .ZN(n8464) );
  MUX2_X1 U10994 ( .A(n11431), .B(n11570), .S(n9385), .Z(n8463) );
  INV_X1 U10995 ( .A(n8421), .ZN(n8424) );
  NAND2_X1 U10996 ( .A1(n15481), .A2(n10946), .ZN(n8554) );
  INV_X1 U10997 ( .A(n8554), .ZN(n8422) );
  OAI21_X1 U10998 ( .B1(n9326), .B2(n8422), .A(n8428), .ZN(n8423) );
  MUX2_X1 U10999 ( .A(n8424), .B(n8423), .S(n9385), .Z(n8438) );
  NAND2_X1 U11000 ( .A1(n8425), .A2(n11564), .ZN(n8427) );
  INV_X1 U11001 ( .A(n11264), .ZN(n9401) );
  NAND3_X1 U11002 ( .A1(n15481), .A2(n10946), .A3(n9401), .ZN(n8426) );
  NAND2_X1 U11003 ( .A1(n8427), .A2(n8426), .ZN(n8429) );
  NAND2_X1 U11004 ( .A1(n8429), .A2(n8428), .ZN(n8431) );
  NAND2_X1 U11005 ( .A1(n10736), .A2(n8430), .ZN(n9329) );
  INV_X1 U11006 ( .A(n9329), .ZN(n15464) );
  NAND2_X1 U11007 ( .A1(n8431), .A2(n15464), .ZN(n8437) );
  NAND2_X1 U11008 ( .A1(n8556), .A2(n10736), .ZN(n8434) );
  INV_X1 U11009 ( .A(n8432), .ZN(n8433) );
  MUX2_X1 U11010 ( .A(n8434), .B(n8433), .S(n9385), .Z(n8435) );
  INV_X1 U11011 ( .A(n8435), .ZN(n8436) );
  OAI21_X1 U11012 ( .B1(n8438), .B2(n8437), .A(n8436), .ZN(n8440) );
  INV_X1 U11013 ( .A(n9333), .ZN(n10833) );
  MUX2_X1 U11014 ( .A(n8555), .B(n8556), .S(n9385), .Z(n8439) );
  NAND2_X1 U11015 ( .A1(n8441), .A2(n8449), .ZN(n8443) );
  NAND2_X1 U11016 ( .A1(n8443), .A2(n10126), .ZN(n8447) );
  INV_X1 U11017 ( .A(n8442), .ZN(n8445) );
  NOR2_X1 U11018 ( .A1(n8443), .A2(n11082), .ZN(n8444) );
  MUX2_X1 U11019 ( .A(n8445), .B(n8444), .S(n10126), .Z(n8446) );
  AOI21_X1 U11020 ( .B1(n8450), .B2(n8448), .A(n10126), .ZN(n8452) );
  MUX2_X1 U11021 ( .A(n8450), .B(n8449), .S(n9385), .Z(n8451) );
  MUX2_X1 U11022 ( .A(n8454), .B(n8453), .S(n9385), .Z(n8455) );
  NAND3_X1 U11023 ( .A1(n8456), .A2(n11281), .A3(n8455), .ZN(n8461) );
  NAND2_X1 U11024 ( .A1(n11570), .A2(n11431), .ZN(n8457) );
  INV_X1 U11025 ( .A(n11349), .ZN(n11351) );
  MUX2_X1 U11026 ( .A(n8459), .B(n8458), .S(n9385), .Z(n8460) );
  NAND3_X1 U11027 ( .A1(n8461), .A2(n11351), .A3(n8460), .ZN(n8462) );
  OAI21_X1 U11028 ( .B1(n8464), .B2(n8463), .A(n8462), .ZN(n8465) );
  NAND2_X1 U11029 ( .A1(n8466), .A2(n8467), .ZN(n9340) );
  INV_X1 U11030 ( .A(n9340), .ZN(n11367) );
  NAND2_X1 U11031 ( .A1(n8465), .A2(n11367), .ZN(n8469) );
  MUX2_X1 U11032 ( .A(n8467), .B(n8466), .S(n9385), .Z(n8468) );
  NAND2_X1 U11033 ( .A1(n8475), .A2(n8470), .ZN(n8471) );
  NAND2_X1 U11034 ( .A1(n8471), .A2(n10126), .ZN(n8472) );
  AOI21_X1 U11035 ( .B1(n8474), .B2(n8473), .A(n10126), .ZN(n8476) );
  XNOR2_X1 U11036 ( .A(n12110), .B(n11864), .ZN(n12067) );
  INV_X1 U11037 ( .A(n12067), .ZN(n12071) );
  MUX2_X1 U11038 ( .A(n11726), .B(n9385), .S(n11864), .Z(n8477) );
  OAI21_X1 U11039 ( .B1(n10126), .B2(n12110), .A(n8477), .ZN(n8478) );
  NAND2_X1 U11040 ( .A1(n12779), .A2(n8478), .ZN(n8482) );
  MUX2_X1 U11041 ( .A(n8480), .B(n8479), .S(n9385), .Z(n8481) );
  NAND2_X1 U11042 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NAND2_X1 U11043 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U11044 ( .A1(n8485), .A2(n12767), .ZN(n8490) );
  OAI21_X1 U11045 ( .B1(n12902), .B2(n12748), .A(n8486), .ZN(n8487) );
  NAND2_X1 U11046 ( .A1(n8487), .A2(n10126), .ZN(n8489) );
  INV_X1 U11047 ( .A(n8492), .ZN(n8488) );
  AOI21_X1 U11048 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8495) );
  AOI21_X1 U11049 ( .B1(n8492), .B2(n8491), .A(n10126), .ZN(n8494) );
  INV_X1 U11050 ( .A(n12902), .ZN(n12384) );
  NAND3_X1 U11051 ( .A1(n12384), .A2(n9385), .A3(n12770), .ZN(n8493) );
  OAI21_X1 U11052 ( .B1(n8495), .B2(n8494), .A(n8493), .ZN(n8496) );
  AOI22_X1 U11053 ( .A1(n8501), .A2(n8497), .B1(n8496), .B2(n7847), .ZN(n8503)
         );
  AND3_X1 U11054 ( .A1(n8498), .A2(n12759), .A3(n12392), .ZN(n8500) );
  NAND3_X1 U11055 ( .A1(n8553), .A2(n8498), .A3(n10126), .ZN(n8499) );
  OAI21_X1 U11056 ( .B1(n8501), .B2(n8500), .A(n8499), .ZN(n8502) );
  MUX2_X1 U11057 ( .A(n8552), .B(n8553), .S(n9385), .Z(n8504) );
  NOR2_X1 U11058 ( .A1(n12884), .A2(n10126), .ZN(n8506) );
  AND2_X1 U11059 ( .A1(n12884), .A2(n10126), .ZN(n8505) );
  MUX2_X1 U11060 ( .A(n8506), .B(n8505), .S(n12718), .Z(n8507) );
  NAND2_X1 U11061 ( .A1(n8509), .A2(n8510), .ZN(n12692) );
  INV_X1 U11062 ( .A(n8514), .ZN(n8508) );
  INV_X1 U11063 ( .A(n12676), .ZN(n12678) );
  MUX2_X1 U11064 ( .A(n8510), .B(n8509), .S(n10126), .Z(n8511) );
  NAND3_X1 U11065 ( .A1(n8512), .A2(n12678), .A3(n8511), .ZN(n8517) );
  MUX2_X1 U11066 ( .A(n8514), .B(n7733), .S(n10126), .Z(n8515) );
  INV_X1 U11067 ( .A(n8520), .ZN(n8524) );
  NAND2_X1 U11068 ( .A1(n8520), .A2(n8519), .ZN(n8522) );
  NAND2_X1 U11069 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  MUX2_X1 U11070 ( .A(n8524), .B(n8523), .S(n10126), .Z(n8525) );
  MUX2_X1 U11071 ( .A(n8527), .B(n8526), .S(n9385), .Z(n8528) );
  NAND3_X1 U11072 ( .A1(n12636), .A2(n8529), .A3(n8528), .ZN(n8534) );
  INV_X1 U11073 ( .A(n8530), .ZN(n8531) );
  MUX2_X1 U11074 ( .A(n8532), .B(n8531), .S(n9385), .Z(n8533) );
  INV_X1 U11075 ( .A(n12625), .ZN(n8536) );
  INV_X1 U11076 ( .A(n12793), .ZN(n12629) );
  NOR2_X1 U11077 ( .A1(n12357), .A2(n9385), .ZN(n8535) );
  NAND2_X1 U11078 ( .A1(n8539), .A2(n8537), .ZN(n12352) );
  NAND2_X1 U11079 ( .A1(n8571), .A2(n8540), .ZN(n8551) );
  NAND3_X1 U11080 ( .A1(n7543), .A2(n9385), .A3(n8543), .ZN(n8550) );
  INV_X1 U11081 ( .A(n8544), .ZN(n8547) );
  OAI211_X1 U11082 ( .C1(n8551), .C2(n8550), .A(n8549), .B(n6484), .ZN(n8576)
         );
  INV_X1 U11083 ( .A(n12692), .ZN(n12689) );
  NAND2_X1 U11084 ( .A1(n8553), .A2(n8552), .ZN(n12722) );
  NOR2_X1 U11085 ( .A1(n9333), .A2(n9329), .ZN(n8558) );
  NAND2_X1 U11086 ( .A1(n8425), .A2(n8554), .ZN(n10533) );
  NOR2_X1 U11087 ( .A1(n9326), .A2(n10533), .ZN(n8557) );
  NAND2_X1 U11088 ( .A1(n8556), .A2(n8555), .ZN(n9332) );
  INV_X1 U11089 ( .A(n9332), .ZN(n10738) );
  NAND4_X1 U11090 ( .A1(n8558), .A2(n8557), .A3(n10738), .A4(n11086), .ZN(
        n8559) );
  NOR2_X1 U11091 ( .A1(n8559), .A2(n10966), .ZN(n8560) );
  NAND4_X1 U11092 ( .A1(n8560), .A2(n11351), .A3(n10948), .A4(n11281), .ZN(
        n8561) );
  NOR2_X1 U11093 ( .A1(n8561), .A2(n9340), .ZN(n8562) );
  NAND3_X1 U11094 ( .A1(n11951), .A2(n8087), .A3(n8562), .ZN(n8563) );
  NOR3_X1 U11095 ( .A1(n12778), .A2(n12067), .A3(n8563), .ZN(n8564) );
  NAND4_X1 U11096 ( .A1(n12711), .A2(n12767), .A3(n8564), .A4(n12757), .ZN(
        n8565) );
  OR4_X1 U11097 ( .A1(n12676), .A2(n12745), .A3(n12722), .A4(n8565), .ZN(n8566) );
  NOR2_X1 U11098 ( .A1(n8566), .A2(n12666), .ZN(n8568) );
  INV_X1 U11099 ( .A(n12702), .ZN(n8567) );
  NAND4_X1 U11100 ( .A1(n12658), .A2(n12689), .A3(n8568), .A4(n8567), .ZN(
        n8569) );
  NOR4_X1 U11101 ( .A1(n12625), .A2(n12633), .A3(n12643), .A4(n8569), .ZN(
        n8570) );
  XNOR2_X1 U11102 ( .A(n8572), .B(n12596), .ZN(n8573) );
  NAND2_X1 U11103 ( .A1(n8573), .A2(n10512), .ZN(n8575) );
  NAND2_X1 U11104 ( .A1(n8576), .A2(n15462), .ZN(n8574) );
  OAI211_X1 U11105 ( .C1(n10515), .C2(n8576), .A(n8575), .B(n8574), .ZN(n8577)
         );
  AOI21_X1 U11106 ( .B1(n8579), .B2(n8578), .A(n8577), .ZN(n8606) );
  INV_X1 U11107 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8583) );
  NAND4_X1 U11108 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n8584)
         );
  NOR2_X1 U11109 ( .A1(n8215), .A2(n8584), .ZN(n8589) );
  INV_X1 U11110 ( .A(n8589), .ZN(n8585) );
  OR2_X1 U11111 ( .A1(n10124), .A2(P3_U3151), .ZN(n11517) );
  OR2_X1 U11112 ( .A1(n10515), .A2(n10126), .ZN(n10532) );
  INV_X1 U11113 ( .A(n10532), .ZN(n8601) );
  NAND2_X1 U11114 ( .A1(n8593), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8592) );
  MUX2_X1 U11115 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8592), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8594) );
  NAND2_X2 U11116 ( .A1(n8594), .A2(n8599), .ZN(n11897) );
  INV_X1 U11117 ( .A(n11897), .ZN(n8598) );
  XNOR2_X2 U11118 ( .A(n8596), .B(n8595), .ZN(n12949) );
  INV_X1 U11119 ( .A(n12949), .ZN(n8597) );
  NAND2_X1 U11120 ( .A1(n8601), .A2(n10252), .ZN(n10237) );
  NOR3_X1 U11121 ( .A1(n10237), .A2(n11473), .A3(n12125), .ZN(n8604) );
  OAI21_X1 U11122 ( .B1(n11517), .B2(n11264), .A(P3_B_REG_SCAN_IN), .ZN(n8603)
         );
  OR2_X1 U11123 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  OAI21_X1 U11124 ( .B1(n8606), .B2(n11517), .A(n8605), .ZN(P3_U3296) );
  INV_X1 U11125 ( .A(n8817), .ZN(n8607) );
  NAND2_X1 U11126 ( .A1(n8607), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8844) );
  INV_X1 U11127 ( .A(n8844), .ZN(n8608) );
  INV_X1 U11128 ( .A(n8938), .ZN(n8610) );
  INV_X1 U11129 ( .A(n9089), .ZN(n8614) );
  AND2_X1 U11130 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n8613) );
  INV_X1 U11131 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14254) );
  INV_X1 U11132 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9122) );
  INV_X1 U11133 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U11134 ( .A1(n9135), .A2(n14162), .ZN(n8616) );
  NAND2_X1 U11135 ( .A1(n9156), .A2(n8616), .ZN(n14753) );
  NOR2_X1 U11136 ( .A1(n9037), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n8619) );
  NOR2_X1 U11137 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n8621) );
  NOR2_X2 U11138 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8620) );
  INV_X2 U11139 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9060) );
  INV_X1 U11140 ( .A(n9038), .ZN(n8625) );
  NAND3_X1 U11141 ( .A1(n8627), .A2(n8626), .A3(n8625), .ZN(n9298) );
  XNOR2_X2 U11142 ( .A(n8630), .B(n15135), .ZN(n12203) );
  XNOR2_X2 U11143 ( .A(n8632), .B(n8631), .ZN(n12290) );
  INV_X1 U11144 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8636) );
  NAND2_X2 U11145 ( .A1(n12290), .A2(n8633), .ZN(n8759) );
  NAND2_X1 U11146 ( .A1(n9210), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U11147 ( .A1(n9209), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8634) );
  OAI211_X1 U11148 ( .C1(n9213), .C2(n8636), .A(n8635), .B(n8634), .ZN(n8637)
         );
  INV_X1 U11149 ( .A(n8637), .ZN(n8638) );
  INV_X1 U11150 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9969) );
  INV_X1 U11151 ( .A(SI_2_), .ZN(n8640) );
  NAND2_X1 U11152 ( .A1(n8646), .A2(n8640), .ZN(n8752) );
  INV_X1 U11153 ( .A(n8644), .ZN(n8641) );
  NAND2_X1 U11154 ( .A1(n8641), .A2(n9931), .ZN(n8725) );
  INV_X1 U11155 ( .A(SI_0_), .ZN(n8736) );
  NOR2_X2 U11156 ( .A1(n8643), .A2(n8736), .ZN(n8727) );
  NAND3_X1 U11157 ( .A1(n8752), .A2(n8725), .A3(n8727), .ZN(n8649) );
  INV_X1 U11158 ( .A(n8749), .ZN(n8645) );
  INV_X1 U11159 ( .A(n8646), .ZN(n8647) );
  NAND2_X1 U11160 ( .A1(n8647), .A2(SI_2_), .ZN(n8751) );
  INV_X1 U11161 ( .A(n8653), .ZN(n8651) );
  INV_X1 U11162 ( .A(SI_3_), .ZN(n8650) );
  NAND2_X1 U11163 ( .A1(n8651), .A2(n8650), .ZN(n8765) );
  INV_X1 U11164 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U11165 ( .A(n9972), .B(n9977), .S(n8659), .Z(n8654) );
  INV_X1 U11166 ( .A(SI_4_), .ZN(n8652) );
  NAND2_X1 U11167 ( .A1(n8654), .A2(n8652), .ZN(n8784) );
  NAND2_X1 U11168 ( .A1(n8653), .A2(SI_3_), .ZN(n8781) );
  INV_X1 U11169 ( .A(n8781), .ZN(n8657) );
  INV_X1 U11170 ( .A(n8654), .ZN(n8655) );
  NAND2_X1 U11171 ( .A1(n8655), .A2(SI_4_), .ZN(n8783) );
  INV_X1 U11172 ( .A(n8783), .ZN(n8656) );
  MUX2_X1 U11173 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8659), .Z(n8660) );
  NAND2_X1 U11174 ( .A1(n8660), .A2(SI_5_), .ZN(n8662) );
  OAI21_X1 U11175 ( .B1(SI_5_), .B2(n8660), .A(n8662), .ZN(n8804) );
  INV_X1 U11176 ( .A(n8804), .ZN(n8661) );
  NAND2_X1 U11177 ( .A1(n8803), .A2(n8661), .ZN(n8806) );
  NAND2_X1 U11178 ( .A1(n8665), .A2(SI_8_), .ZN(n8666) );
  MUX2_X1 U11179 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n7434), .Z(n8667) );
  NAND2_X1 U11180 ( .A1(n8667), .A2(SI_9_), .ZN(n8669) );
  OAI21_X1 U11181 ( .B1(SI_9_), .B2(n8667), .A(n8669), .ZN(n8668) );
  INV_X1 U11182 ( .A(n8668), .ZN(n8873) );
  INV_X1 U11183 ( .A(n8671), .ZN(n8670) );
  NAND2_X1 U11184 ( .A1(n8670), .A2(n9991), .ZN(n8931) );
  NAND2_X1 U11185 ( .A1(n8672), .A2(n9973), .ZN(n8927) );
  INV_X1 U11186 ( .A(n8929), .ZN(n8674) );
  XNOR2_X1 U11187 ( .A(n8676), .B(n9999), .ZN(n8933) );
  INV_X1 U11188 ( .A(n8933), .ZN(n8673) );
  INV_X1 U11189 ( .A(n8676), .ZN(n8677) );
  MUX2_X1 U11190 ( .A(n15539), .B(n10274), .S(n7434), .Z(n8678) );
  XNOR2_X1 U11191 ( .A(n8678), .B(SI_13_), .ZN(n8946) );
  NAND2_X1 U11192 ( .A1(n8947), .A2(n8946), .ZN(n8680) );
  NAND2_X1 U11193 ( .A1(n8678), .A2(n10071), .ZN(n8679) );
  MUX2_X1 U11194 ( .A(n10539), .B(n10571), .S(n7434), .Z(n8966) );
  NOR2_X1 U11195 ( .A1(n8681), .A2(SI_14_), .ZN(n8683) );
  XNOR2_X1 U11196 ( .A(n8684), .B(SI_15_), .ZN(n8980) );
  NAND2_X1 U11197 ( .A1(n8681), .A2(SI_14_), .ZN(n8682) );
  MUX2_X1 U11198 ( .A(n10569), .B(n10618), .S(n7434), .Z(n8686) );
  XNOR2_X1 U11199 ( .A(n8686), .B(SI_16_), .ZN(n9012) );
  NAND2_X1 U11200 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  MUX2_X1 U11201 ( .A(n10686), .B(n10760), .S(n7434), .Z(n8999) );
  NOR2_X1 U11202 ( .A1(n8688), .A2(SI_17_), .ZN(n8689) );
  MUX2_X1 U11203 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7434), .Z(n9051) );
  INV_X1 U11204 ( .A(n9051), .ZN(n8690) );
  MUX2_X1 U11205 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n7434), .Z(n8692) );
  NAND2_X1 U11206 ( .A1(n8692), .A2(SI_19_), .ZN(n9056) );
  OAI21_X1 U11207 ( .B1(n10844), .B2(n8690), .A(n9056), .ZN(n8691) );
  NOR2_X1 U11208 ( .A1(n9051), .A2(SI_18_), .ZN(n8695) );
  INV_X1 U11209 ( .A(n8692), .ZN(n8693) );
  NAND2_X1 U11210 ( .A1(n8693), .A2(n10874), .ZN(n9055) );
  INV_X1 U11211 ( .A(n9055), .ZN(n8694) );
  MUX2_X1 U11212 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7434), .Z(n9075) );
  MUX2_X1 U11213 ( .A(n11374), .B(n15584), .S(n7434), .Z(n9098) );
  INV_X1 U11214 ( .A(n9098), .ZN(n9071) );
  NOR2_X1 U11215 ( .A1(n9071), .A2(SI_20_), .ZN(n8697) );
  NOR2_X1 U11216 ( .A1(n9098), .A2(n11363), .ZN(n8700) );
  INV_X1 U11217 ( .A(n8698), .ZN(n8699) );
  AOI22_X1 U11218 ( .A1(n8700), .A2(n8699), .B1(SI_21_), .B2(n9075), .ZN(n9102) );
  MUX2_X1 U11219 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n7434), .Z(n9772) );
  NAND2_X1 U11220 ( .A1(n9772), .A2(SI_22_), .ZN(n8701) );
  INV_X1 U11221 ( .A(n9772), .ZN(n8704) );
  MUX2_X1 U11222 ( .A(n11496), .B(n8705), .S(n7434), .Z(n9117) );
  NOR2_X1 U11223 ( .A1(n8707), .A2(SI_23_), .ZN(n8706) );
  XNOR2_X1 U11224 ( .A(n9146), .B(SI_24_), .ZN(n9130) );
  INV_X1 U11225 ( .A(n9130), .ZN(n8708) );
  MUX2_X1 U11226 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n7434), .Z(n9147) );
  NAND2_X1 U11227 ( .A1(n8708), .A2(n9147), .ZN(n8710) );
  NAND2_X1 U11228 ( .A1(n9146), .A2(SI_24_), .ZN(n8709) );
  NAND2_X1 U11229 ( .A1(n8710), .A2(n8709), .ZN(n8714) );
  MUX2_X1 U11230 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n7434), .Z(n8711) );
  NAND2_X1 U11231 ( .A1(n8711), .A2(SI_25_), .ZN(n9150) );
  INV_X1 U11232 ( .A(n8711), .ZN(n8712) );
  NAND2_X1 U11233 ( .A1(n8712), .A2(n12946), .ZN(n9148) );
  NAND2_X1 U11234 ( .A1(n9150), .A2(n9148), .ZN(n8713) );
  XNOR2_X2 U11235 ( .A(n8714), .B(n8713), .ZN(n13915) );
  NAND2_X1 U11236 ( .A1(n13915), .A2(n6409), .ZN(n8720) );
  OR2_X1 U11237 ( .A1(n14466), .A2(n15145), .ZN(n8719) );
  NAND2_X1 U11238 ( .A1(n9209), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8724) );
  INV_X1 U11239 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11207) );
  NAND2_X1 U11240 ( .A1(n8794), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8722) );
  INV_X1 U11241 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14582) );
  NAND2_X1 U11242 ( .A1(n8749), .A2(n8725), .ZN(n8729) );
  INV_X1 U11243 ( .A(n8729), .ZN(n8726) );
  NAND2_X1 U11244 ( .A1(n8726), .A2(n8727), .ZN(n8750) );
  INV_X1 U11245 ( .A(n8727), .ZN(n8728) );
  NAND2_X1 U11246 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U11247 ( .A1(n8750), .A2(n8730), .ZN(n9968) );
  MUX2_X1 U11248 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8731), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8732) );
  INV_X1 U11249 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n11328) );
  INV_X1 U11250 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11327) );
  NOR2_X1 U11251 ( .A1(n7434), .A2(n8736), .ZN(n8737) );
  XNOR2_X1 U11252 ( .A(n8737), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15151) );
  MUX2_X1 U11253 ( .A(n7040), .B(n15151), .S(n8755), .Z(n11333) );
  INV_X1 U11254 ( .A(n14315), .ZN(n8738) );
  AOI21_X2 U11255 ( .B1(n14317), .B2(n10152), .A(n8738), .ZN(n14321) );
  INV_X1 U11256 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8739) );
  OR2_X1 U11257 ( .A1(n9136), .A2(n8739), .ZN(n8741) );
  INV_X1 U11258 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10173) );
  OR2_X1 U11259 ( .A1(n8759), .A2(n10173), .ZN(n8740) );
  AND2_X1 U11260 ( .A1(n8741), .A2(n8740), .ZN(n8745) );
  INV_X1 U11261 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8742) );
  OR2_X1 U11262 ( .A1(n9213), .A2(n8742), .ZN(n8744) );
  INV_X1 U11263 ( .A(n14580), .ZN(n8757) );
  NAND2_X1 U11264 ( .A1(n8746), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8747) );
  MUX2_X1 U11265 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8747), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n8748) );
  NAND2_X1 U11266 ( .A1(n8750), .A2(n8749), .ZN(n8754) );
  NAND2_X1 U11267 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  XNOR2_X1 U11268 ( .A(n8754), .B(n8753), .ZN(n9519) );
  INV_X1 U11269 ( .A(n9519), .ZN(n9970) );
  OR2_X1 U11270 ( .A1(n14580), .A2(n8756), .ZN(n14318) );
  NAND2_X1 U11271 ( .A1(n9209), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8764) );
  INV_X1 U11272 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11510) );
  OR2_X1 U11273 ( .A1(n8759), .A2(n11510), .ZN(n8763) );
  INV_X1 U11274 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8760) );
  OR2_X1 U11275 ( .A1(n9213), .A2(n8760), .ZN(n8762) );
  OR2_X1 U11276 ( .A1(n14466), .A2(n7089), .ZN(n8775) );
  NAND2_X1 U11277 ( .A1(n8781), .A2(n8765), .ZN(n8767) );
  NAND2_X1 U11278 ( .A1(n8766), .A2(n8767), .ZN(n8770) );
  INV_X1 U11279 ( .A(n8767), .ZN(n8768) );
  NAND2_X1 U11280 ( .A1(n8770), .A2(n8782), .ZN(n9967) );
  OR2_X1 U11281 ( .A1(n14463), .A2(n9967), .ZN(n8774) );
  NAND2_X1 U11282 ( .A1(n8856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8771) );
  MUX2_X1 U11283 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8771), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8772) );
  NAND2_X1 U11284 ( .A1(n8772), .A2(n8808), .ZN(n14621) );
  OR2_X1 U11285 ( .A1(n6397), .A2(n14621), .ZN(n8773) );
  NAND2_X1 U11286 ( .A1(n14579), .A2(n15275), .ZN(n14326) );
  NAND2_X1 U11287 ( .A1(n9209), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8780) );
  INV_X1 U11288 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11320) );
  OR2_X1 U11289 ( .A1(n8759), .A2(n11320), .ZN(n8779) );
  XNOR2_X1 U11290 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11322) );
  OR2_X1 U11291 ( .A1(n9136), .A2(n11322), .ZN(n8778) );
  INV_X1 U11292 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8776) );
  OR2_X1 U11293 ( .A1(n9213), .A2(n8776), .ZN(n8777) );
  NAND2_X1 U11294 ( .A1(n8782), .A2(n8781), .ZN(n8786) );
  NAND2_X1 U11295 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  XNOR2_X1 U11296 ( .A(n8786), .B(n8785), .ZN(n9971) );
  NAND2_X1 U11297 ( .A1(n14450), .A2(n9971), .ZN(n8790) );
  NAND2_X1 U11298 ( .A1(n8808), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8787) );
  OR2_X1 U11299 ( .A1(n6397), .A2(n15220), .ZN(n8789) );
  OR2_X1 U11300 ( .A1(n14466), .A2(n9972), .ZN(n8788) );
  AND3_X2 U11301 ( .A1(n8790), .A2(n8789), .A3(n8788), .ZN(n15246) );
  NAND2_X1 U11302 ( .A1(n15250), .A2(n15246), .ZN(n8791) );
  INV_X1 U11303 ( .A(n15250), .ZN(n15247) );
  NAND2_X1 U11304 ( .A1(n15247), .A2(n15285), .ZN(n8792) );
  NAND2_X1 U11305 ( .A1(n8793), .A2(n8792), .ZN(n15245) );
  NAND2_X1 U11306 ( .A1(n14453), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8802) );
  INV_X1 U11307 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10177) );
  OR2_X1 U11308 ( .A1(n8759), .A2(n10177), .ZN(n8801) );
  INV_X1 U11309 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11310 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n8795) );
  NAND2_X1 U11311 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  NAND2_X1 U11312 ( .A1(n8817), .A2(n8797), .ZN(n14186) );
  OR2_X1 U11313 ( .A1(n9136), .A2(n14186), .ZN(n8800) );
  INV_X1 U11314 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8798) );
  OR2_X1 U11315 ( .A1(n14455), .A2(n8798), .ZN(n8799) );
  NAND4_X1 U11316 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(n14578) );
  INV_X1 U11317 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U11318 ( .A1(n8805), .A2(n8804), .ZN(n8807) );
  AND2_X1 U11319 ( .A1(n8806), .A2(n8807), .ZN(n9932) );
  NAND2_X1 U11320 ( .A1(n9932), .A2(n14450), .ZN(n8814) );
  INV_X1 U11321 ( .A(n8808), .ZN(n8810) );
  NAND2_X1 U11322 ( .A1(n8810), .A2(n8809), .ZN(n8829) );
  NAND2_X1 U11323 ( .A1(n8829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8812) );
  INV_X1 U11324 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8811) );
  XNOR2_X1 U11325 ( .A(n8812), .B(n8811), .ZN(n10176) );
  OR2_X1 U11326 ( .A1(n8755), .A2(n10176), .ZN(n8813) );
  NAND2_X1 U11327 ( .A1(n15281), .A2(n6407), .ZN(n8815) );
  NAND2_X1 U11328 ( .A1(n9209), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8823) );
  INV_X1 U11329 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8816) );
  OR2_X1 U11330 ( .A1(n8759), .A2(n8816), .ZN(n8822) );
  INV_X1 U11331 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n15520) );
  NAND2_X1 U11332 ( .A1(n8817), .A2(n15520), .ZN(n8818) );
  NAND2_X1 U11333 ( .A1(n8844), .A2(n8818), .ZN(n11454) );
  OR2_X1 U11334 ( .A1(n9136), .A2(n11454), .ZN(n8821) );
  INV_X1 U11335 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8819) );
  OR2_X1 U11336 ( .A1(n9213), .A2(n8819), .ZN(n8820) );
  NAND4_X1 U11337 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n14577) );
  NAND2_X1 U11338 ( .A1(n8826), .A2(n8825), .ZN(n8828) );
  NAND2_X1 U11339 ( .A1(n8828), .A2(n8827), .ZN(n9980) );
  OR2_X1 U11340 ( .A1(n9980), .A2(n14463), .ZN(n8832) );
  NAND2_X1 U11341 ( .A1(n8839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8830) );
  XNOR2_X1 U11342 ( .A(n8830), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U11343 ( .A1(n9063), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9062), .B2(
        n10220), .ZN(n8831) );
  NAND2_X1 U11344 ( .A1(n14577), .A2(n15298), .ZN(n8833) );
  OR2_X1 U11345 ( .A1(n8836), .A2(n8835), .ZN(n8837) );
  AND2_X1 U11346 ( .A1(n8838), .A2(n8837), .ZN(n9993) );
  NAND2_X1 U11347 ( .A1(n9993), .A2(n14450), .ZN(n8842) );
  OAI21_X1 U11348 ( .B1(n8839), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8840) );
  XNOR2_X1 U11349 ( .A(n8840), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U11350 ( .A1(n9063), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9062), .B2(
        n10221), .ZN(n8841) );
  NAND2_X1 U11351 ( .A1(n8842), .A2(n8841), .ZN(n14348) );
  NAND2_X1 U11352 ( .A1(n14453), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8850) );
  INV_X1 U11353 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10222) );
  OR2_X1 U11354 ( .A1(n8759), .A2(n10222), .ZN(n8849) );
  INV_X1 U11355 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11356 ( .A1(n8844), .A2(n8843), .ZN(n8845) );
  NAND2_X1 U11357 ( .A1(n8864), .A2(n8845), .ZN(n15235) );
  OR2_X1 U11358 ( .A1(n9136), .A2(n15235), .ZN(n8848) );
  INV_X1 U11359 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n8846) );
  OR2_X1 U11360 ( .A1(n14455), .A2(n8846), .ZN(n8847) );
  NOR2_X1 U11361 ( .A1(n14348), .A2(n15313), .ZN(n8851) );
  OR2_X1 U11362 ( .A1(n8853), .A2(n8852), .ZN(n8854) );
  NAND2_X1 U11363 ( .A1(n8855), .A2(n8854), .ZN(n10007) );
  OR2_X1 U11364 ( .A1(n10007), .A2(n14463), .ZN(n8862) );
  INV_X1 U11365 ( .A(n9040), .ZN(n8859) );
  NAND2_X1 U11366 ( .A1(n8859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8858) );
  MUX2_X1 U11367 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8858), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n8860) );
  AOI22_X1 U11368 ( .A1(n9063), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9062), .B2(
        n10312), .ZN(n8861) );
  NAND2_X1 U11369 ( .A1(n9209), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8870) );
  INV_X1 U11370 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10223) );
  OR2_X1 U11371 ( .A1(n8759), .A2(n10223), .ZN(n8869) );
  INV_X1 U11372 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U11373 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  NAND2_X1 U11374 ( .A1(n8881), .A2(n8865), .ZN(n11379) );
  OR2_X1 U11375 ( .A1(n9136), .A2(n11379), .ZN(n8868) );
  INV_X1 U11376 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8866) );
  OR2_X1 U11377 ( .A1(n9213), .A2(n8866), .ZN(n8867) );
  XNOR2_X1 U11378 ( .A(n15316), .B(n11933), .ZN(n14524) );
  INV_X1 U11379 ( .A(n14524), .ZN(n8871) );
  INV_X1 U11380 ( .A(n15316), .ZN(n9242) );
  NAND2_X1 U11381 ( .A1(n9242), .A2(n14575), .ZN(n8872) );
  OR2_X1 U11382 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  NAND2_X1 U11383 ( .A1(n8876), .A2(n8875), .ZN(n10044) );
  OR2_X1 U11384 ( .A1(n10044), .A2(n14463), .ZN(n8879) );
  NAND2_X1 U11385 ( .A1(n9002), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8877) );
  XNOR2_X1 U11386 ( .A(n8877), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U11387 ( .A1(n9063), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9062), .B2(
        n10317), .ZN(n8878) );
  NAND2_X1 U11388 ( .A1(n14453), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8886) );
  INV_X1 U11389 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10463) );
  OR2_X1 U11390 ( .A1(n8759), .A2(n10463), .ZN(n8885) );
  NAND2_X1 U11391 ( .A1(n8881), .A2(n8880), .ZN(n8882) );
  NAND2_X1 U11392 ( .A1(n8901), .A2(n8882), .ZN(n11648) );
  OR2_X1 U11393 ( .A1(n9136), .A2(n11648), .ZN(n8884) );
  INV_X1 U11394 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10458) );
  OR2_X1 U11395 ( .A1(n14455), .A2(n10458), .ZN(n8883) );
  XNOR2_X1 U11396 ( .A(n14355), .B(n15311), .ZN(n14535) );
  NAND2_X1 U11397 ( .A1(n14355), .A2(n15311), .ZN(n8887) );
  NAND2_X1 U11398 ( .A1(n8928), .A2(n8888), .ZN(n8910) );
  NAND2_X1 U11399 ( .A1(n8890), .A2(n9973), .ZN(n8891) );
  INV_X1 U11400 ( .A(n9002), .ZN(n8893) );
  INV_X1 U11401 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11402 ( .A1(n8893), .A2(n8892), .ZN(n8895) );
  NAND2_X1 U11403 ( .A1(n8895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8894) );
  MUX2_X1 U11404 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8894), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n8898) );
  INV_X1 U11405 ( .A(n8895), .ZN(n8897) );
  INV_X1 U11406 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8896) );
  AOI22_X1 U11407 ( .A1(n9063), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9062), 
        .B2(n10559), .ZN(n8899) );
  NAND2_X1 U11408 ( .A1(n9209), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8907) );
  INV_X1 U11409 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11763) );
  OR2_X1 U11410 ( .A1(n8759), .A2(n11763), .ZN(n8906) );
  NAND2_X1 U11411 ( .A1(n8901), .A2(n8900), .ZN(n8902) );
  NAND2_X1 U11412 ( .A1(n8919), .A2(n8902), .ZN(n12181) );
  OR2_X1 U11413 ( .A1(n9136), .A2(n12181), .ZN(n8905) );
  INV_X1 U11414 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8903) );
  OR2_X1 U11415 ( .A1(n9213), .A2(n8903), .ZN(n8904) );
  NAND4_X1 U11416 ( .A1(n8907), .A2(n8906), .A3(n8905), .A4(n8904), .ZN(n14574) );
  NAND2_X1 U11417 ( .A1(n15108), .A2(n14360), .ZN(n8908) );
  NAND2_X1 U11418 ( .A1(n10422), .A2(n14450), .ZN(n8916) );
  NAND2_X1 U11419 ( .A1(n8987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8914) );
  XNOR2_X1 U11420 ( .A(n8914), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U11421 ( .A1(n9063), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9062), 
        .B2(n10768), .ZN(n8915) );
  NAND2_X1 U11422 ( .A1(n9209), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8925) );
  INV_X1 U11423 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8917) );
  OR2_X1 U11424 ( .A1(n8759), .A2(n8917), .ZN(n8924) );
  INV_X1 U11425 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11426 ( .A1(n8919), .A2(n8918), .ZN(n8920) );
  NAND2_X1 U11427 ( .A1(n8938), .A2(n8920), .ZN(n14263) );
  OR2_X1 U11428 ( .A1(n9136), .A2(n14263), .ZN(n8923) );
  INV_X1 U11429 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8921) );
  OR2_X1 U11430 ( .A1(n9213), .A2(n8921), .ZN(n8922) );
  NAND4_X1 U11431 ( .A1(n8925), .A2(n8924), .A3(n8923), .A4(n8922), .ZN(n15092) );
  INV_X1 U11432 ( .A(n15092), .ZN(n14364) );
  OR2_X1 U11433 ( .A1(n7165), .A2(n14364), .ZN(n8926) );
  NAND2_X1 U11434 ( .A1(n8928), .A2(n8927), .ZN(n8930) );
  NAND2_X1 U11435 ( .A1(n8930), .A2(n8929), .ZN(n8932) );
  NAND2_X1 U11436 ( .A1(n8932), .A2(n8931), .ZN(n8934) );
  XNOR2_X1 U11437 ( .A(n8934), .B(n8933), .ZN(n10150) );
  NAND2_X1 U11438 ( .A1(n10150), .A2(n14450), .ZN(n8937) );
  NAND2_X1 U11439 ( .A1(n8935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8948) );
  XNOR2_X1 U11440 ( .A(n8948), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U11441 ( .A1(n9063), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9062), 
        .B2(n10769), .ZN(n8936) );
  NAND2_X1 U11442 ( .A1(n9210), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8944) );
  INV_X1 U11443 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11110) );
  OR2_X1 U11444 ( .A1(n14455), .A2(n11110), .ZN(n8943) );
  INV_X1 U11445 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n14149) );
  NAND2_X1 U11446 ( .A1(n8938), .A2(n14149), .ZN(n8939) );
  NAND2_X1 U11447 ( .A1(n8956), .A2(n8939), .ZN(n14965) );
  OR2_X1 U11448 ( .A1(n9136), .A2(n14965), .ZN(n8942) );
  INV_X1 U11449 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8940) );
  OR2_X1 U11450 ( .A1(n9213), .A2(n8940), .ZN(n8941) );
  NAND4_X1 U11451 ( .A1(n8944), .A2(n8943), .A3(n8942), .A4(n8941), .ZN(n14946) );
  XNOR2_X1 U11452 ( .A(n14972), .B(n14946), .ZN(n14961) );
  INV_X1 U11453 ( .A(n14946), .ZN(n15083) );
  OR2_X1 U11454 ( .A1(n14972), .A2(n15083), .ZN(n8945) );
  NAND2_X1 U11455 ( .A1(n14960), .A2(n8945), .ZN(n14945) );
  XNOR2_X1 U11456 ( .A(n8947), .B(n8946), .ZN(n10184) );
  NAND2_X1 U11457 ( .A1(n10184), .A2(n14450), .ZN(n8954) );
  NAND2_X1 U11458 ( .A1(n8948), .A2(n8984), .ZN(n8949) );
  NAND2_X1 U11459 ( .A1(n8949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8951) );
  INV_X1 U11460 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U11461 ( .A1(n8951), .A2(n8950), .ZN(n8969) );
  OR2_X1 U11462 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  AOI22_X1 U11463 ( .A1(n9063), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9062), 
        .B2(n11112), .ZN(n8953) );
  NAND2_X1 U11464 ( .A1(n9209), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8962) );
  INV_X1 U11465 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11104) );
  OR2_X1 U11466 ( .A1(n8759), .A2(n11104), .ZN(n8961) );
  NAND2_X1 U11467 ( .A1(n8956), .A2(n8955), .ZN(n8957) );
  NAND2_X1 U11468 ( .A1(n8973), .A2(n8957), .ZN(n14947) );
  OR2_X1 U11469 ( .A1(n9136), .A2(n14947), .ZN(n8960) );
  INV_X1 U11470 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8958) );
  OR2_X1 U11471 ( .A1(n9213), .A2(n8958), .ZN(n8959) );
  NAND4_X1 U11472 ( .A1(n8962), .A2(n8961), .A3(n8960), .A4(n8959), .ZN(n15091) );
  XNOR2_X1 U11473 ( .A(n15086), .B(n15091), .ZN(n14944) );
  NAND2_X1 U11474 ( .A1(n14945), .A2(n14944), .ZN(n14943) );
  INV_X1 U11475 ( .A(n15091), .ZN(n15075) );
  OR2_X1 U11476 ( .A1(n15086), .A2(n15075), .ZN(n8963) );
  NAND2_X1 U11477 ( .A1(n8964), .A2(n10271), .ZN(n8965) );
  NAND2_X1 U11478 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U11479 ( .A1(n8969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8970) );
  AOI22_X1 U11480 ( .A1(n11801), .A2(n9062), .B1(n9063), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11481 ( .A1(n14453), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8978) );
  INV_X1 U11482 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8972) );
  OR2_X1 U11483 ( .A1(n8759), .A2(n8972), .ZN(n8977) );
  INV_X1 U11484 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11111) );
  OR2_X1 U11485 ( .A1(n14455), .A2(n11111), .ZN(n8976) );
  NAND2_X1 U11486 ( .A1(n8973), .A2(n6711), .ZN(n8974) );
  NAND2_X1 U11487 ( .A1(n8991), .A2(n8974), .ZN(n14936) );
  OR2_X1 U11488 ( .A1(n9136), .A2(n14936), .ZN(n8975) );
  NAND2_X1 U11489 ( .A1(n15078), .A2(n15082), .ZN(n14389) );
  AND2_X2 U11490 ( .A1(n14390), .A2(n14389), .ZN(n14930) );
  INV_X1 U11491 ( .A(n8980), .ZN(n8981) );
  INV_X1 U11492 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8983) );
  NAND3_X1 U11493 ( .A1(n8985), .A2(n8984), .A3(n8983), .ZN(n8986) );
  OAI21_X1 U11494 ( .B1(n8987), .B2(n8986), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8988) );
  XNOR2_X1 U11495 ( .A(n8988), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U11496 ( .A1(n9063), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9062), 
        .B2(n11976), .ZN(n8989) );
  NAND2_X1 U11497 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  AND2_X1 U11498 ( .A1(n9025), .A2(n8992), .ZN(n14919) );
  NAND2_X1 U11499 ( .A1(n9216), .A2(n14919), .ZN(n8998) );
  INV_X1 U11500 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8993) );
  OR2_X1 U11501 ( .A1(n14455), .A2(n8993), .ZN(n8997) );
  INV_X1 U11502 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11803) );
  OR2_X1 U11503 ( .A1(n8759), .A2(n11803), .ZN(n8996) );
  INV_X1 U11504 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8994) );
  OR2_X1 U11505 ( .A1(n9213), .A2(n8994), .ZN(n8995) );
  XNOR2_X1 U11506 ( .A(n8999), .B(SI_17_), .ZN(n9000) );
  XNOR2_X1 U11507 ( .A(n9001), .B(n9000), .ZN(n10685) );
  NAND2_X1 U11508 ( .A1(n10685), .A2(n6409), .ZN(n9006) );
  NOR2_X1 U11509 ( .A1(n9002), .A2(n9038), .ZN(n9014) );
  NAND2_X1 U11510 ( .A1(n9014), .A2(n9003), .ZN(n9017) );
  NAND2_X1 U11511 ( .A1(n9017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9004) );
  XNOR2_X1 U11512 ( .A(n9004), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14644) );
  AOI22_X1 U11513 ( .A1(n9063), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9062), 
        .B2(n14644), .ZN(n9005) );
  NAND2_X1 U11514 ( .A1(n9027), .A2(n9007), .ZN(n9008) );
  AND2_X1 U11515 ( .A1(n9045), .A2(n9008), .ZN(n14881) );
  NAND2_X1 U11516 ( .A1(n14881), .A2(n9216), .ZN(n9011) );
  AOI22_X1 U11517 ( .A1(n14453), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n9210), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U11518 ( .A1(n9209), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9009) );
  XNOR2_X1 U11519 ( .A(n9013), .B(n9012), .ZN(n10568) );
  NAND2_X1 U11520 ( .A1(n10568), .A2(n6409), .ZN(n9020) );
  INV_X1 U11521 ( .A(n9014), .ZN(n9015) );
  NAND2_X1 U11522 ( .A1(n9015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9016) );
  MUX2_X1 U11523 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9016), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9018) );
  AOI22_X1 U11524 ( .A1(n9063), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9062), 
        .B2(n14636), .ZN(n9019) );
  INV_X1 U11525 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9021) );
  OR2_X1 U11526 ( .A1(n14455), .A2(n9021), .ZN(n9023) );
  INV_X1 U11527 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14895) );
  OR2_X1 U11528 ( .A1(n8759), .A2(n14895), .ZN(n9022) );
  AND2_X1 U11529 ( .A1(n9023), .A2(n9022), .ZN(n9030) );
  INV_X1 U11530 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U11531 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  NAND2_X1 U11532 ( .A1(n9027), .A2(n9026), .ZN(n14894) );
  OR2_X1 U11533 ( .A1(n14894), .A2(n9136), .ZN(n9029) );
  NAND2_X1 U11534 ( .A1(n14453), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9028) );
  OR2_X1 U11535 ( .A1(n15064), .A2(n15053), .ZN(n9031) );
  OAI211_X1 U11536 ( .C1(n15057), .C2(n15061), .A(n14872), .B(n9031), .ZN(
        n9032) );
  INV_X1 U11537 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U11538 ( .A1(n15064), .A2(n15053), .ZN(n14873) );
  NAND2_X1 U11539 ( .A1(n14873), .A2(n14858), .ZN(n9035) );
  NOR2_X1 U11540 ( .A1(n14858), .A2(n14884), .ZN(n9034) );
  AOI22_X1 U11541 ( .A1(n15057), .A2(n9035), .B1(n9034), .B2(n15064), .ZN(
        n9036) );
  XNOR2_X1 U11542 ( .A(n9052), .B(n9051), .ZN(n11171) );
  NAND2_X1 U11543 ( .A1(n11171), .A2(n6409), .ZN(n9043) );
  NAND2_X1 U11544 ( .A1(n9058), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9041) );
  XNOR2_X1 U11545 ( .A(n9041), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14664) );
  AOI22_X1 U11546 ( .A1(n9063), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9062), 
        .B2(n14664), .ZN(n9042) );
  INV_X1 U11547 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U11548 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U11549 ( .A1(n9089), .A2(n9046), .ZN(n14859) );
  OR2_X1 U11550 ( .A1(n14859), .A2(n9136), .ZN(n9049) );
  AOI22_X1 U11551 ( .A1(n9209), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9210), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11552 ( .A1(n14453), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11553 ( .A1(n15045), .A2(n15054), .ZN(n14404) );
  NAND2_X1 U11554 ( .A1(n14405), .A2(n14404), .ZN(n14865) );
  NAND2_X1 U11555 ( .A1(n9053), .A2(SI_18_), .ZN(n9054) );
  NAND2_X1 U11556 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U11557 ( .A1(n9734), .A2(n6409), .ZN(n9065) );
  NAND2_X1 U11558 ( .A1(n9218), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9061) );
  XNOR2_X2 U11559 ( .A(n9061), .B(n9060), .ZN(n14934) );
  AOI22_X1 U11560 ( .A1(n9063), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14672), 
        .B2(n9062), .ZN(n9064) );
  XNOR2_X1 U11561 ( .A(n9089), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n14845) );
  NAND2_X1 U11562 ( .A1(n14845), .A2(n9216), .ZN(n9070) );
  INV_X1 U11563 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15646) );
  NAND2_X1 U11564 ( .A1(n9210), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11565 ( .A1(n14453), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9066) );
  OAI211_X1 U11566 ( .C1(n15646), .C2(n14455), .A(n9067), .B(n9066), .ZN(n9068) );
  INV_X1 U11567 ( .A(n9068), .ZN(n9069) );
  NAND2_X1 U11568 ( .A1(n9099), .A2(n9071), .ZN(n9074) );
  OR2_X1 U11569 ( .A1(n9072), .A2(n11363), .ZN(n9073) );
  NAND2_X1 U11570 ( .A1(n9074), .A2(n9073), .ZN(n9077) );
  XNOR2_X1 U11571 ( .A(n9075), .B(SI_21_), .ZN(n9076) );
  NAND2_X1 U11572 ( .A1(n11497), .A2(n6409), .ZN(n9079) );
  OR2_X1 U11573 ( .A1(n14466), .A2(n11498), .ZN(n9078) );
  NAND2_X2 U11574 ( .A1(n9079), .A2(n9078), .ZN(n14790) );
  INV_X1 U11575 ( .A(n9080), .ZN(n9090) );
  INV_X1 U11576 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15581) );
  NAND2_X1 U11577 ( .A1(n9090), .A2(n15581), .ZN(n9081) );
  NAND2_X1 U11578 ( .A1(n9106), .A2(n9081), .ZN(n14818) );
  INV_X1 U11579 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11580 ( .A1(n9209), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11581 ( .A1(n9210), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9082) );
  OAI211_X1 U11582 ( .C1(n9084), .C2(n9213), .A(n9083), .B(n9082), .ZN(n9085)
         );
  INV_X1 U11583 ( .A(n9085), .ZN(n9086) );
  INV_X1 U11584 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n14103) );
  INV_X1 U11585 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9088) );
  OAI21_X1 U11586 ( .B1(n9089), .B2(n14103), .A(n9088), .ZN(n9091) );
  NAND2_X1 U11587 ( .A1(n9091), .A2(n9090), .ZN(n14228) );
  OR2_X1 U11588 ( .A1(n14228), .A2(n9136), .ZN(n9097) );
  INV_X1 U11589 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11590 ( .A1(n9210), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11591 ( .A1(n9209), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9092) );
  OAI211_X1 U11592 ( .C1(n9213), .C2(n9094), .A(n9093), .B(n9092), .ZN(n9095)
         );
  INV_X1 U11593 ( .A(n9095), .ZN(n9096) );
  XNOR2_X1 U11594 ( .A(n9099), .B(n9098), .ZN(n11372) );
  NAND2_X1 U11595 ( .A1(n11372), .A2(n6409), .ZN(n9101) );
  OR2_X1 U11596 ( .A1(n14466), .A2(n11374), .ZN(n9100) );
  AOI22_X1 U11597 ( .A1(n14790), .A2(n15027), .B1(n14848), .B2(n15030), .ZN(
        n14768) );
  NAND2_X1 U11598 ( .A1(n9103), .A2(n9102), .ZN(n9104) );
  XNOR2_X1 U11599 ( .A(n9105), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15150) );
  NAND2_X1 U11600 ( .A1(n9106), .A2(n14254), .ZN(n9107) );
  NAND2_X1 U11601 ( .A1(n9123), .A2(n9107), .ZN(n14801) );
  OR2_X1 U11602 ( .A1(n14801), .A2(n9136), .ZN(n9112) );
  INV_X1 U11603 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15578) );
  NAND2_X1 U11604 ( .A1(n14453), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11605 ( .A1(n9210), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9108) );
  OAI211_X1 U11606 ( .C1(n14455), .C2(n15578), .A(n9109), .B(n9108), .ZN(n9110) );
  INV_X1 U11607 ( .A(n9110), .ZN(n9111) );
  OR2_X1 U11608 ( .A1(n14804), .A2(n14572), .ZN(n14769) );
  XNOR2_X1 U11609 ( .A(n14804), .B(n14010), .ZN(n14791) );
  OR2_X1 U11610 ( .A1(n15030), .A2(n14848), .ZN(n14789) );
  NAND2_X1 U11611 ( .A1(n14789), .A2(n15027), .ZN(n9115) );
  NAND2_X1 U11612 ( .A1(n14573), .A2(n15035), .ZN(n9113) );
  NOR2_X1 U11613 ( .A1(n15030), .A2(n9113), .ZN(n9114) );
  AOI21_X1 U11614 ( .B1(n15021), .B2(n9115), .A(n9114), .ZN(n9116) );
  NAND2_X1 U11615 ( .A1(n14791), .A2(n9116), .ZN(n14767) );
  XNOR2_X1 U11616 ( .A(n9117), .B(SI_23_), .ZN(n9118) );
  XNOR2_X1 U11617 ( .A(n9119), .B(n9118), .ZN(n11494) );
  NAND2_X1 U11618 ( .A1(n11494), .A2(n6409), .ZN(n9121) );
  OR2_X1 U11619 ( .A1(n14466), .A2(n11496), .ZN(n9120) );
  NAND2_X1 U11620 ( .A1(n9123), .A2(n9122), .ZN(n9124) );
  AND2_X1 U11621 ( .A1(n9133), .A2(n9124), .ZN(n14778) );
  INV_X1 U11622 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U11623 ( .A1(n9209), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11624 ( .A1(n9210), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9125) );
  OAI211_X1 U11625 ( .C1(n9127), .C2(n9213), .A(n9126), .B(n9125), .ZN(n9128)
         );
  XNOR2_X1 U11626 ( .A(n15009), .B(n14251), .ZN(n14542) );
  AOI21_X1 U11627 ( .B1(n14767), .B2(n14769), .A(n14542), .ZN(n9129) );
  XNOR2_X1 U11628 ( .A(n9130), .B(n9147), .ZN(n11995) );
  NAND2_X1 U11629 ( .A1(n11995), .A2(n6409), .ZN(n9132) );
  OR2_X1 U11630 ( .A1(n14466), .A2(n15647), .ZN(n9131) );
  INV_X1 U11631 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14208) );
  NAND2_X1 U11632 ( .A1(n9133), .A2(n14208), .ZN(n9134) );
  NAND2_X1 U11633 ( .A1(n9135), .A2(n9134), .ZN(n14209) );
  OR2_X1 U11634 ( .A1(n14209), .A2(n9136), .ZN(n9142) );
  INV_X1 U11635 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U11636 ( .A1(n9209), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U11637 ( .A1(n9210), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9137) );
  OAI211_X1 U11638 ( .C1(n9139), .C2(n9213), .A(n9138), .B(n9137), .ZN(n9140)
         );
  INV_X1 U11639 ( .A(n9140), .ZN(n9141) );
  INV_X1 U11640 ( .A(n14570), .ZN(n14160) );
  XNOR2_X1 U11641 ( .A(n14998), .B(n14042), .ZN(n14746) );
  INV_X1 U11642 ( .A(n9147), .ZN(n9144) );
  OAI21_X1 U11643 ( .B1(n9144), .B2(n11899), .A(n9150), .ZN(n9145) );
  NOR2_X1 U11644 ( .A1(n9147), .A2(SI_24_), .ZN(n9151) );
  INV_X1 U11645 ( .A(n9148), .ZN(n9149) );
  AOI21_X1 U11646 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(n9152) );
  MUX2_X1 U11647 ( .A(n11945), .B(n11948), .S(n7434), .Z(n9163) );
  XNOR2_X1 U11648 ( .A(n9163), .B(SI_26_), .ZN(n9153) );
  XNOR2_X1 U11649 ( .A(n9164), .B(n9153), .ZN(n11944) );
  NAND2_X1 U11650 ( .A1(n11944), .A2(n6409), .ZN(n9155) );
  OR2_X1 U11651 ( .A1(n14466), .A2(n11945), .ZN(n9154) );
  INV_X1 U11652 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U11653 ( .A1(n9156), .A2(n14285), .ZN(n9157) );
  INV_X1 U11654 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U11655 ( .A1(n9210), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11656 ( .A1(n9209), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9158) );
  OAI211_X1 U11657 ( .C1(n9213), .C2(n9160), .A(n9159), .B(n9158), .ZN(n9161)
         );
  INV_X1 U11658 ( .A(n9161), .ZN(n9162) );
  NAND2_X1 U11659 ( .A1(n9164), .A2(n12942), .ZN(n9165) );
  MUX2_X1 U11660 ( .A(n15143), .B(n15530), .S(n7434), .Z(n9181) );
  XNOR2_X1 U11661 ( .A(n9181), .B(SI_27_), .ZN(n9167) );
  NAND2_X1 U11662 ( .A1(n12064), .A2(n6409), .ZN(n9169) );
  OR2_X1 U11663 ( .A1(n14466), .A2(n15143), .ZN(n9168) );
  INV_X1 U11664 ( .A(n9172), .ZN(n9170) );
  NAND2_X1 U11665 ( .A1(n9170), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9193) );
  INV_X1 U11666 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U11667 ( .A1(n9172), .A2(n9171), .ZN(n9173) );
  NAND2_X1 U11668 ( .A1(n9193), .A2(n9173), .ZN(n14059) );
  INV_X1 U11669 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U11670 ( .A1(n9209), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U11671 ( .A1(n9210), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9174) );
  OAI211_X1 U11672 ( .C1(n9176), .C2(n9213), .A(n9175), .B(n9174), .ZN(n9177)
         );
  INV_X1 U11673 ( .A(n9177), .ZN(n9178) );
  NAND2_X1 U11674 ( .A1(n9184), .A2(n12939), .ZN(n9183) );
  INV_X1 U11675 ( .A(n9181), .ZN(n9182) );
  NAND2_X1 U11676 ( .A1(n9183), .A2(n9182), .ZN(n9185) );
  MUX2_X1 U11677 ( .A(n12205), .B(n9186), .S(n7434), .Z(n9187) );
  NAND2_X1 U11678 ( .A1(n9187), .A2(n12126), .ZN(n9205) );
  INV_X1 U11679 ( .A(n9187), .ZN(n9188) );
  NAND2_X1 U11680 ( .A1(n9188), .A2(SI_28_), .ZN(n9189) );
  NAND2_X1 U11681 ( .A1(n9205), .A2(n9189), .ZN(n9203) );
  NAND2_X1 U11682 ( .A1(n12269), .A2(n6409), .ZN(n9191) );
  OR2_X1 U11683 ( .A1(n14466), .A2(n12205), .ZN(n9190) );
  INV_X1 U11684 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9192) );
  NAND2_X1 U11685 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  NAND2_X1 U11686 ( .A1(n14708), .A2(n9216), .ZN(n9200) );
  INV_X1 U11687 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U11688 ( .A1(n9209), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U11689 ( .A1(n9210), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9195) );
  OAI211_X1 U11690 ( .C1(n9197), .C2(n9213), .A(n9196), .B(n9195), .ZN(n9198)
         );
  INV_X1 U11691 ( .A(n9198), .ZN(n9199) );
  NAND2_X1 U11692 ( .A1(n12130), .A2(n7867), .ZN(n9202) );
  INV_X1 U11693 ( .A(n14566), .ZN(n14697) );
  NAND2_X1 U11694 ( .A1(n9202), .A2(n9201), .ZN(n9217) );
  MUX2_X1 U11695 ( .A(n12289), .B(n13240), .S(n7434), .Z(n12193) );
  XNOR2_X1 U11696 ( .A(n12193), .B(SI_29_), .ZN(n12196) );
  NAND2_X1 U11697 ( .A1(n13239), .A2(n6409), .ZN(n9207) );
  OR2_X1 U11698 ( .A1(n14466), .A2(n12289), .ZN(n9206) );
  INV_X1 U11699 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U11700 ( .A1(n9209), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U11701 ( .A1(n9210), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9211) );
  OAI211_X1 U11702 ( .C1(n9214), .C2(n9213), .A(n9212), .B(n9211), .ZN(n9215)
         );
  XNOR2_X1 U11703 ( .A(n14486), .B(n14484), .ZN(n14549) );
  XNOR2_X1 U11704 ( .A(n9217), .B(n14549), .ZN(n14692) );
  NAND2_X1 U11705 ( .A1(n14304), .A2(n14672), .ZN(n14305) );
  NAND2_X1 U11706 ( .A1(n9227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9222) );
  INV_X1 U11707 ( .A(n9223), .ZN(n9224) );
  NAND2_X1 U11708 ( .A1(n9224), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9225) );
  INV_X1 U11709 ( .A(n11375), .ZN(n14476) );
  NAND2_X1 U11710 ( .A1(n9285), .A2(n14476), .ZN(n14308) );
  INV_X1 U11711 ( .A(n11333), .ZN(n10304) );
  NAND2_X1 U11712 ( .A1(n14581), .A2(n10304), .ZN(n10670) );
  NAND2_X1 U11713 ( .A1(n10668), .A2(n10670), .ZN(n10669) );
  OR2_X1 U11714 ( .A1(n9228), .A2(n14131), .ZN(n9229) );
  NAND2_X1 U11715 ( .A1(n10669), .A2(n9229), .ZN(n10784) );
  NAND2_X1 U11716 ( .A1(n10782), .A2(n9230), .ZN(n11502) );
  NAND2_X1 U11717 ( .A1(n14327), .A2(n14326), .ZN(n14526) );
  NAND2_X1 U11718 ( .A1(n11502), .A2(n14526), .ZN(n11317) );
  NAND2_X1 U11719 ( .A1(n15250), .A2(n15285), .ZN(n9232) );
  NAND2_X1 U11720 ( .A1(n14578), .A2(n6407), .ZN(n9231) );
  OR2_X1 U11721 ( .A1(n15250), .A2(n15285), .ZN(n9233) );
  INV_X1 U11722 ( .A(n9233), .ZN(n9235) );
  NAND2_X1 U11723 ( .A1(n9233), .A2(n14578), .ZN(n9234) );
  INV_X1 U11724 ( .A(n15275), .ZN(n14094) );
  OR2_X1 U11725 ( .A1(n14579), .A2(n14094), .ZN(n11316) );
  XNOR2_X1 U11726 ( .A(n14577), .B(n15298), .ZN(n14530) );
  INV_X1 U11727 ( .A(n14577), .ZN(n9238) );
  NAND2_X1 U11728 ( .A1(n9238), .A2(n15298), .ZN(n9239) );
  XNOR2_X1 U11729 ( .A(n14348), .B(n15313), .ZN(n15227) );
  NAND2_X1 U11730 ( .A1(n15303), .A2(n15313), .ZN(n9240) );
  NAND2_X1 U11731 ( .A1(n9241), .A2(n9240), .ZN(n11376) );
  NAND2_X1 U11732 ( .A1(n11376), .A2(n14524), .ZN(n9244) );
  NAND2_X1 U11733 ( .A1(n9242), .A2(n11933), .ZN(n9243) );
  NAND2_X1 U11734 ( .A1(n7437), .A2(n15311), .ZN(n9245) );
  NAND2_X1 U11735 ( .A1(n14359), .A2(n14360), .ZN(n9246) );
  INV_X1 U11736 ( .A(n14539), .ZN(n9248) );
  NAND2_X1 U11737 ( .A1(n12026), .A2(n9248), .ZN(n9250) );
  OR2_X1 U11738 ( .A1(n7165), .A2(n15092), .ZN(n9249) );
  INV_X1 U11739 ( .A(n14961), .ZN(n9251) );
  OR2_X1 U11740 ( .A1(n14972), .A2(n14946), .ZN(n9252) );
  INV_X1 U11741 ( .A(n14944), .ZN(n9253) );
  INV_X1 U11742 ( .A(n15082), .ZN(n9254) );
  NAND2_X1 U11743 ( .A1(n15078), .A2(n9254), .ZN(n9255) );
  INV_X1 U11744 ( .A(n14930), .ZN(n14927) );
  INV_X1 U11745 ( .A(n9255), .ZN(n14908) );
  NOR2_X1 U11746 ( .A1(n14927), .A2(n14908), .ZN(n9258) );
  INV_X1 U11747 ( .A(n15074), .ZN(n14897) );
  NOR2_X1 U11748 ( .A1(n15071), .A2(n14897), .ZN(n9257) );
  XNOR2_X1 U11749 ( .A(n15064), .B(n15053), .ZN(n14902) );
  OR2_X1 U11750 ( .A1(n15064), .A2(n14884), .ZN(n9260) );
  NAND2_X1 U11751 ( .A1(n15057), .A2(n14858), .ZN(n9261) );
  OR2_X1 U11752 ( .A1(n15045), .A2(n15034), .ZN(n9262) );
  INV_X1 U11753 ( .A(n15043), .ZN(n14833) );
  NOR2_X1 U11754 ( .A1(n14850), .A2(n14833), .ZN(n9263) );
  XNOR2_X1 U11755 ( .A(n15030), .B(n14848), .ZN(n14827) );
  NAND2_X1 U11756 ( .A1(n15030), .A2(n15035), .ZN(n9264) );
  OR2_X1 U11757 ( .A1(n14804), .A2(n14010), .ZN(n9266) );
  OAI21_X1 U11758 ( .B1(n15021), .B2(n15027), .A(n9266), .ZN(n9265) );
  NOR2_X1 U11759 ( .A1(n14790), .A2(n14573), .ZN(n14786) );
  AOI22_X1 U11760 ( .A1(n14786), .A2(n9266), .B1(n14010), .B2(n14804), .ZN(
        n9267) );
  INV_X1 U11761 ( .A(n14251), .ZN(n14571) );
  NAND2_X1 U11762 ( .A1(n15009), .A2(n14571), .ZN(n9268) );
  INV_X1 U11763 ( .A(n12146), .ZN(n9269) );
  OR2_X1 U11764 ( .A1(n15006), .A2(n14570), .ZN(n9270) );
  INV_X1 U11765 ( .A(n14746), .ZN(n14759) );
  NAND2_X1 U11766 ( .A1(n14998), .A2(n14569), .ZN(n9271) );
  NAND2_X1 U11767 ( .A1(n14994), .A2(n14568), .ZN(n9272) );
  INV_X1 U11768 ( .A(n14549), .ZN(n9275) );
  NAND2_X1 U11769 ( .A1(n14449), .A2(n14566), .ZN(n12127) );
  INV_X1 U11770 ( .A(n12127), .ZN(n9273) );
  OR2_X1 U11771 ( .A1(n14449), .A2(n14566), .ZN(n12128) );
  OR2_X1 U11772 ( .A1(n14985), .A2(n14567), .ZN(n12135) );
  NAND2_X1 U11773 ( .A1(n12128), .A2(n12135), .ZN(n9277) );
  AOI21_X1 U11774 ( .B1(n12127), .B2(n9277), .A(n9275), .ZN(n9274) );
  AOI21_X1 U11775 ( .B1(n9275), .B2(n12127), .A(n9274), .ZN(n9276) );
  NAND2_X1 U11776 ( .A1(n14304), .A2(n14479), .ZN(n9281) );
  NAND2_X1 U11777 ( .A1(n14304), .A2(n14934), .ZN(n9280) );
  INV_X1 U11778 ( .A(n9293), .ZN(n9282) );
  OR2_X1 U11779 ( .A1(n9282), .A2(n14934), .ZN(n9284) );
  NAND2_X1 U11780 ( .A1(n14304), .A2(n9285), .ZN(n14478) );
  INV_X1 U11781 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9289) );
  INV_X1 U11782 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14686) );
  OR2_X1 U11783 ( .A1(n8759), .A2(n14686), .ZN(n9288) );
  NAND2_X1 U11784 ( .A1(n14453), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9287) );
  OAI211_X1 U11785 ( .C1(n14455), .C2(n9289), .A(n9288), .B(n9287), .ZN(n14564) );
  INV_X1 U11786 ( .A(n9286), .ZN(n10155) );
  INV_X1 U11787 ( .A(P1_B_REG_SCAN_IN), .ZN(n9291) );
  NOR2_X1 U11788 ( .A1(n6410), .A2(n9291), .ZN(n9292) );
  NOR2_X1 U11789 ( .A1(n15310), .A2(n9292), .ZN(n14678) );
  NAND2_X1 U11790 ( .A1(n14564), .A2(n14678), .ZN(n14694) );
  OAI21_X1 U11791 ( .B1(n14697), .B2(n15312), .A(n14694), .ZN(n9294) );
  OR2_X2 U11792 ( .A1(n14131), .A2(n10304), .ZN(n10780) );
  INV_X1 U11793 ( .A(n15102), .ZN(n14363) );
  NAND2_X1 U11794 ( .A1(n12033), .A2(n14363), .ZN(n12032) );
  OR2_X2 U11795 ( .A1(n12032), .A2(n14972), .ZN(n14962) );
  INV_X1 U11796 ( .A(n15078), .ZN(n14932) );
  INV_X1 U11797 ( .A(n15071), .ZN(n14921) );
  INV_X1 U11798 ( .A(n15009), .ZN(n14780) );
  AND2_X2 U11799 ( .A1(n14799), .A2(n14780), .ZN(n14777) );
  INV_X1 U11800 ( .A(n15006), .ZN(n14214) );
  NAND2_X2 U11801 ( .A1(n9293), .A2(n11375), .ZN(n10283) );
  NOR2_X2 U11802 ( .A1(n12140), .A2(n14486), .ZN(n14685) );
  AOI211_X1 U11803 ( .C1(n14486), .C2(n12140), .A(n10283), .B(n14685), .ZN(
        n14704) );
  AOI211_X2 U11804 ( .C1(n14486), .C2(n15315), .A(n9294), .B(n14704), .ZN(
        n9295) );
  AND2_X1 U11805 ( .A1(n11375), .A2(n14934), .ZN(n9307) );
  OAI21_X1 U11806 ( .B1(n9058), .B2(n9296), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9297) );
  MUX2_X1 U11807 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9297), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9300) );
  NAND2_X1 U11808 ( .A1(n9301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U11809 ( .A1(n9299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9303) );
  OAI211_X1 U11810 ( .C1(n14478), .C2(n9307), .A(n10288), .B(n10041), .ZN(
        n10301) );
  NAND3_X1 U11811 ( .A1(n11998), .A2(P1_B_REG_SCAN_IN), .A3(n15149), .ZN(n9310) );
  INV_X1 U11812 ( .A(n9311), .ZN(n11946) );
  NAND2_X1 U11813 ( .A1(n11946), .A2(n11998), .ZN(n10003) );
  NAND2_X1 U11814 ( .A1(n9312), .A2(n10003), .ZN(n9418) );
  NOR4_X1 U11815 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9316) );
  NOR4_X1 U11816 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9315) );
  NOR4_X1 U11817 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9314) );
  NOR4_X1 U11818 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9313) );
  NAND4_X1 U11819 ( .A1(n9316), .A2(n9315), .A3(n9314), .A4(n9313), .ZN(n9322)
         );
  NOR2_X1 U11820 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n9320) );
  NOR4_X1 U11821 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9319) );
  NOR4_X1 U11822 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9318) );
  NOR4_X1 U11823 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9317) );
  NAND4_X1 U11824 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(n9321)
         );
  NOR2_X1 U11825 ( .A1(n9322), .A2(n9321), .ZN(n10276) );
  NAND2_X1 U11826 ( .A1(n11946), .A2(n15149), .ZN(n10279) );
  OAI21_X1 U11827 ( .B1(n10278), .B2(P1_D_REG_1__SCAN_IN), .A(n10279), .ZN(
        n9323) );
  OAI211_X1 U11828 ( .C1(n10276), .C2(n10278), .A(n10300), .B(n9323), .ZN(
        n9419) );
  NAND2_X1 U11829 ( .A1(n9420), .A2(n15327), .ZN(n9325) );
  INV_X1 U11830 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11831 ( .A1(n9325), .A2(n7865), .ZN(P1_U3557) );
  NAND2_X1 U11832 ( .A1(n15481), .A2(n10629), .ZN(n10575) );
  NAND2_X1 U11833 ( .A1(n9326), .A2(n10575), .ZN(n9328) );
  INV_X1 U11834 ( .A(n15476), .ZN(n10579) );
  OR2_X1 U11835 ( .A1(n12461), .A2(n10579), .ZN(n9327) );
  NAND2_X1 U11836 ( .A1(n15463), .A2(n9329), .ZN(n9331) );
  OR2_X1 U11837 ( .A1(n15480), .A2(n10587), .ZN(n9330) );
  NAND2_X1 U11838 ( .A1(n9331), .A2(n9330), .ZN(n10739) );
  INV_X1 U11839 ( .A(n11412), .ZN(n10613) );
  AND2_X1 U11840 ( .A1(n10836), .A2(n10613), .ZN(n10830) );
  INV_X1 U11841 ( .A(n11406), .ZN(n10697) );
  OR2_X1 U11842 ( .A1(n12459), .A2(n11093), .ZN(n10965) );
  INV_X1 U11843 ( .A(n11121), .ZN(n11100) );
  NAND2_X1 U11844 ( .A1(n12458), .A2(n11100), .ZN(n9336) );
  NAND2_X1 U11845 ( .A1(n12457), .A2(n6932), .ZN(n9337) );
  OR2_X1 U11846 ( .A1(n11436), .A2(n12456), .ZN(n9338) );
  INV_X1 U11847 ( .A(n12455), .ZN(n11352) );
  OR2_X1 U11848 ( .A1(n11677), .A2(n11352), .ZN(n9341) );
  NOR2_X1 U11849 ( .A1(n11787), .A2(n11908), .ZN(n9344) );
  NAND2_X1 U11850 ( .A1(n11787), .A2(n11908), .ZN(n9343) );
  NOR2_X1 U11851 ( .A1(n12908), .A2(n12782), .ZN(n9345) );
  INV_X1 U11852 ( .A(n12908), .ZN(n12059) );
  INV_X1 U11853 ( .A(n12392), .ZN(n12828) );
  NOR2_X1 U11854 ( .A1(n12893), .A2(n12430), .ZN(n9346) );
  NOR2_X1 U11855 ( .A1(n9346), .A2(n12711), .ZN(n9348) );
  INV_X1 U11856 ( .A(n9346), .ZN(n9347) );
  OR2_X1 U11857 ( .A1(n12738), .A2(n12452), .ZN(n12713) );
  NAND2_X1 U11858 ( .A1(n12722), .A2(n12713), .ZN(n12714) );
  NAND2_X1 U11859 ( .A1(n12686), .A2(n12695), .ZN(n9349) );
  NAND2_X1 U11860 ( .A1(n12340), .A2(n9350), .ZN(n9351) );
  NAND2_X1 U11861 ( .A1(n12313), .A2(n9352), .ZN(n9353) );
  NAND2_X1 U11862 ( .A1(n9354), .A2(n9353), .ZN(n12635) );
  INV_X1 U11863 ( .A(n12635), .ZN(n9355) );
  NAND2_X1 U11864 ( .A1(n12449), .A2(n12645), .ZN(n9356) );
  NAND2_X1 U11865 ( .A1(n12593), .A2(n11264), .ZN(n9408) );
  NAND3_X1 U11866 ( .A1(n9424), .A2(n12784), .A3(n9359), .ZN(n9363) );
  INV_X1 U11867 ( .A(n12125), .ZN(n9427) );
  NAND2_X1 U11868 ( .A1(n9427), .A2(n11473), .ZN(n10130) );
  AND2_X1 U11869 ( .A1(n7918), .A2(n10130), .ZN(n9360) );
  NAND2_X1 U11870 ( .A1(n9363), .A2(n9362), .ZN(n12610) );
  XNOR2_X1 U11871 ( .A(n11897), .B(P3_B_REG_SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11872 ( .A1(n9364), .A2(n12949), .ZN(n9365) );
  INV_X1 U11873 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9366) );
  NAND2_X1 U11874 ( .A1(n10010), .A2(n9366), .ZN(n9369) );
  INV_X1 U11875 ( .A(n9367), .ZN(n12944) );
  NAND2_X1 U11876 ( .A1(n12944), .A2(n12949), .ZN(n9368) );
  INV_X1 U11877 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U11878 ( .A1(n6449), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U11879 ( .A1(n12944), .A2(n11897), .ZN(n9371) );
  NAND2_X1 U11880 ( .A1(n10621), .A2(n10622), .ZN(n9406) );
  NOR2_X1 U11881 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .ZN(
        n9376) );
  NOR4_X1 U11882 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9375) );
  NOR4_X1 U11883 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9374) );
  NOR4_X1 U11884 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9373) );
  NAND4_X1 U11885 ( .A1(n9376), .A2(n9375), .A3(n9374), .A4(n9373), .ZN(n9382)
         );
  NOR4_X1 U11886 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9380) );
  NOR4_X1 U11887 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9379) );
  NOR4_X1 U11888 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9378) );
  NOR4_X1 U11889 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9377) );
  NAND4_X1 U11890 ( .A1(n9380), .A2(n9379), .A3(n9378), .A4(n9377), .ZN(n9381)
         );
  OAI21_X1 U11891 ( .B1(n9382), .B2(n9381), .A(n10010), .ZN(n9407) );
  AND2_X1 U11892 ( .A1(n9407), .A2(n10252), .ZN(n9383) );
  AND2_X1 U11893 ( .A1(n11564), .A2(n11362), .ZN(n9394) );
  OAI211_X1 U11894 ( .C1(n11264), .C2(n9394), .A(n9408), .B(n10515), .ZN(n9384) );
  NAND3_X1 U11895 ( .A1(n10621), .A2(n10126), .A3(n9384), .ZN(n9387) );
  NAND2_X1 U11896 ( .A1(n9385), .A2(n10515), .ZN(n10235) );
  NAND3_X1 U11897 ( .A1(n12596), .A2(n11264), .A3(n10513), .ZN(n9399) );
  NAND2_X1 U11898 ( .A1(n9399), .A2(n10126), .ZN(n10619) );
  NAND2_X1 U11899 ( .A1(n10622), .A2(n10623), .ZN(n9386) );
  NAND2_X1 U11900 ( .A1(n9387), .A2(n9386), .ZN(n9388) );
  MUX2_X1 U11901 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n12610), .S(n15514), .Z(
        n9389) );
  INV_X1 U11902 ( .A(n9389), .ZN(n9404) );
  INV_X1 U11903 ( .A(n9391), .ZN(n9392) );
  NOR2_X1 U11904 ( .A1(n9390), .A2(n9392), .ZN(n9393) );
  INV_X1 U11905 ( .A(n9394), .ZN(n9395) );
  XNOR2_X1 U11906 ( .A(n11264), .B(n9395), .ZN(n9397) );
  NAND2_X1 U11907 ( .A1(n12596), .A2(n11564), .ZN(n9396) );
  NAND2_X1 U11908 ( .A1(n9397), .A2(n9396), .ZN(n10241) );
  NOR2_X1 U11909 ( .A1(n12829), .A2(n10515), .ZN(n9398) );
  NAND2_X1 U11910 ( .A1(n10241), .A2(n9398), .ZN(n9400) );
  AND2_X1 U11911 ( .A1(n9400), .A2(n9399), .ZN(n11357) );
  NAND2_X1 U11912 ( .A1(n15462), .A2(n9401), .ZN(n11347) );
  INV_X1 U11913 ( .A(n12614), .ZN(n9423) );
  OAI22_X1 U11914 ( .A1(n12617), .A2(n12843), .B1(n9423), .B2(n12821), .ZN(
        n9402) );
  INV_X1 U11915 ( .A(n9402), .ZN(n9403) );
  NAND2_X1 U11916 ( .A1(n9404), .A2(n9403), .ZN(P3_U3487) );
  INV_X1 U11917 ( .A(n10241), .ZN(n9412) );
  INV_X1 U11918 ( .A(n9407), .ZN(n9405) );
  INV_X1 U11919 ( .A(n10622), .ZN(n12923) );
  INV_X1 U11920 ( .A(n10621), .ZN(n12921) );
  NAND3_X1 U11921 ( .A1(n12923), .A2(n12921), .A3(n9407), .ZN(n10247) );
  INV_X1 U11922 ( .A(n9408), .ZN(n9409) );
  NAND2_X1 U11923 ( .A1(n9409), .A2(n10512), .ZN(n10244) );
  AND2_X1 U11924 ( .A1(n10244), .A2(n10532), .ZN(n9410) );
  MUX2_X1 U11925 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n12610), .S(n15510), .Z(
        n9414) );
  INV_X1 U11926 ( .A(n9414), .ZN(n9417) );
  OAI22_X1 U11927 ( .A1(n12617), .A2(n12919), .B1(n9423), .B2(n12894), .ZN(
        n9415) );
  INV_X1 U11928 ( .A(n9415), .ZN(n9416) );
  NAND2_X1 U11929 ( .A1(n9417), .A2(n9416), .ZN(P3_U3455) );
  INV_X1 U11930 ( .A(n9418), .ZN(n10293) );
  NAND2_X1 U11931 ( .A1(n9420), .A2(n6403), .ZN(n9422) );
  NAND2_X1 U11932 ( .A1(n15323), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U11933 ( .A1(n9422), .A2(n9421), .ZN(P1_U3525) );
  NAND2_X1 U11934 ( .A1(n9424), .A2(n7876), .ZN(n9425) );
  INV_X1 U11935 ( .A(n9426), .ZN(n12619) );
  AOI21_X1 U11936 ( .B1(n9427), .B2(P3_B_REG_SCAN_IN), .A(n15469), .ZN(n12142)
         );
  AOI22_X1 U11937 ( .A1(n12704), .A2(n12619), .B1(n12451), .B2(n12142), .ZN(
        n9428) );
  XNOR2_X1 U11938 ( .A(n9429), .B(n6524), .ZN(n12192) );
  INV_X1 U11939 ( .A(n12850), .ZN(n12187) );
  INV_X1 U11940 ( .A(n9431), .ZN(n9432) );
  OAI21_X1 U11941 ( .B1(n12849), .B2(n9433), .A(n9432), .ZN(P3_U3488) );
  INV_X1 U11942 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n15532) );
  NOR2_X1 U11943 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .ZN(n9436) );
  NAND4_X1 U11944 ( .A1(n9436), .A2(n9435), .A3(n9434), .A4(n9685), .ZN(n9711)
         );
  NAND3_X1 U11945 ( .A1(n9586), .A2(n9438), .A3(n9437), .ZN(n9439) );
  NAND2_X1 U11946 ( .A1(n9880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9442) );
  XNOR2_X2 U11947 ( .A(n9442), .B(n9441), .ZN(n13666) );
  NAND2_X1 U11948 ( .A1(n13111), .A2(n6398), .ZN(n11267) );
  INV_X1 U11949 ( .A(n9457), .ZN(n9445) );
  NAND2_X1 U11950 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n9447) );
  NAND3_X1 U11951 ( .A1(n9445), .A2(P2_IR_REG_31__SCAN_IN), .A3(n9447), .ZN(
        n9454) );
  NAND2_X1 U11952 ( .A1(n9818), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9444) );
  OAI211_X1 U11953 ( .C1(n9445), .C2(n9818), .A(n9447), .B(n9444), .ZN(n9452)
         );
  OAI211_X1 U11954 ( .C1(n9446), .C2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_19__SCAN_IN), .B(n9876), .ZN(n9450) );
  INV_X1 U11955 ( .A(n9447), .ZN(n9448) );
  NAND3_X1 U11956 ( .A1(n9448), .A2(P2_IR_REG_19__SCAN_IN), .A3(n9818), .ZN(
        n9449) );
  NAND2_X1 U11957 ( .A1(n9450), .A2(n9449), .ZN(n9451) );
  AOI21_X1 U11958 ( .B1(n9452), .B2(n13905), .A(n9451), .ZN(n9453) );
  OAI21_X1 U11959 ( .B1(n9880), .B2(n9454), .A(n9453), .ZN(n9455) );
  NAND3_X1 U11960 ( .A1(n7090), .A2(n9884), .A3(n9459), .ZN(n9460) );
  NAND2_X1 U11961 ( .A1(n12064), .A2(n13262), .ZN(n9466) );
  NAND2_X1 U11962 ( .A1(n6400), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9465) );
  INV_X1 U11963 ( .A(n9550), .ZN(n9467) );
  NAND2_X1 U11964 ( .A1(n9467), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9567) );
  INV_X1 U11965 ( .A(n9567), .ZN(n9468) );
  INV_X1 U11966 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15516) );
  INV_X1 U11967 ( .A(n9490), .ZN(n9473) );
  INV_X1 U11968 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U11969 ( .A1(n9490), .A2(n9474), .ZN(n9475) );
  NAND2_X1 U11970 ( .A1(n9863), .A2(n9475), .ZN(n13489) );
  NAND2_X1 U11971 ( .A1(n13099), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U11972 ( .A1(n12277), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9482) );
  OAI211_X1 U11973 ( .C1(n15532), .C2(n9479), .A(n9483), .B(n9482), .ZN(n9484)
         );
  INV_X1 U11974 ( .A(n9484), .ZN(n9485) );
  NAND2_X1 U11975 ( .A1(n11944), .A2(n13262), .ZN(n9488) );
  NAND2_X1 U11976 ( .A1(n6400), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9487) );
  INV_X1 U11977 ( .A(n13771), .ZN(n13231) );
  NAND2_X1 U11978 ( .A1(n9810), .A2(n15516), .ZN(n9489) );
  NAND2_X1 U11979 ( .A1(n13502), .A2(n12282), .ZN(n9495) );
  INV_X1 U11980 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13504) );
  NAND2_X1 U11981 ( .A1(n12277), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9492) );
  NAND2_X1 U11982 ( .A1(n12278), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9491) );
  OAI211_X1 U11983 ( .C1(n9814), .C2(n13504), .A(n9492), .B(n9491), .ZN(n9493)
         );
  INV_X1 U11984 ( .A(n9493), .ZN(n9494) );
  INV_X1 U11985 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9496) );
  INV_X1 U11986 ( .A(n9751), .ZN(n9497) );
  INV_X1 U11987 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10072) );
  OR2_X1 U11988 ( .A1(n9509), .A2(n10072), .ZN(n9498) );
  INV_X1 U11989 ( .A(n13328), .ZN(n13438) );
  NOR2_X1 U11990 ( .A1(n7434), .A2(n9926), .ZN(n9500) );
  OAI21_X1 U11991 ( .B1(n10089), .B2(n13362), .A(n9501), .ZN(n9502) );
  INV_X1 U11992 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10142) );
  INV_X1 U11993 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11048) );
  NAND2_X1 U11994 ( .A1(n7434), .A2(SI_0_), .ZN(n9507) );
  XNOR2_X1 U11995 ( .A(n9507), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13919) );
  OR2_X1 U11996 ( .A1(n10801), .A2(n13113), .ZN(n9508) );
  INV_X1 U11997 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13370) );
  INV_X1 U11998 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10076) );
  INV_X1 U11999 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9511) );
  OR2_X1 U12000 ( .A1(n9510), .A2(n9511), .ZN(n9513) );
  NAND2_X1 U12001 ( .A1(n13099), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U12002 ( .A1(n9515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9516) );
  MUX2_X1 U12003 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9516), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n9518) );
  INV_X1 U12004 ( .A(n9517), .ZN(n9532) );
  INV_X1 U12005 ( .A(n13372), .ZN(n10104) );
  INV_X1 U12006 ( .A(n9536), .ZN(n9520) );
  NAND2_X1 U12007 ( .A1(n9520), .A2(n9519), .ZN(n9522) );
  OR2_X1 U12008 ( .A1(n13354), .A2(n10805), .ZN(n9525) );
  NAND2_X1 U12009 ( .A1(n13099), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9530) );
  INV_X1 U12010 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9526) );
  OR2_X1 U12011 ( .A1(n13100), .A2(n9526), .ZN(n9529) );
  INV_X1 U12012 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U12013 ( .A1(n9556), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U12014 ( .A1(n9532), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9531) );
  MUX2_X1 U12015 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9531), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9533) );
  NAND2_X1 U12016 ( .A1(n9735), .A2(n13389), .ZN(n9534) );
  INV_X1 U12017 ( .A(n13299), .ZN(n10752) );
  OR2_X1 U12018 ( .A1(n13353), .A2(n13119), .ZN(n9537) );
  NAND2_X1 U12019 ( .A1(n12277), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9541) );
  INV_X1 U12020 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11004) );
  OAI21_X1 U12021 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n9550), .ZN(n11005) );
  OR2_X1 U12022 ( .A1(n9811), .A2(n11005), .ZN(n9539) );
  INV_X1 U12023 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10081) );
  OR2_X1 U12024 ( .A1(n9479), .A2(n10081), .ZN(n9538) );
  NAND2_X1 U12025 ( .A1(n9543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9542) );
  MUX2_X1 U12026 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9542), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9546) );
  INV_X1 U12027 ( .A(n9543), .ZN(n9545) );
  INV_X1 U12028 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U12029 ( .A1(n9545), .A2(n9544), .ZN(n9558) );
  NAND2_X1 U12030 ( .A1(n9546), .A2(n9558), .ZN(n15336) );
  NAND2_X1 U12031 ( .A1(n6400), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9547) );
  XNOR2_X1 U12032 ( .A(n13352), .B(n6405), .ZN(n13304) );
  INV_X1 U12033 ( .A(n13304), .ZN(n11000) );
  NAND2_X1 U12034 ( .A1(n10993), .A2(n11000), .ZN(n10995) );
  OR2_X1 U12035 ( .A1(n13352), .A2(n6405), .ZN(n9548) );
  NAND2_X1 U12036 ( .A1(n10995), .A2(n9548), .ZN(n11055) );
  NAND2_X1 U12037 ( .A1(n12277), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9555) );
  INV_X1 U12038 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11063) );
  OR2_X1 U12039 ( .A1(n9814), .A2(n11063), .ZN(n9554) );
  INV_X1 U12040 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U12041 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  NAND2_X1 U12042 ( .A1(n9567), .A2(n9551), .ZN(n11067) );
  OR2_X1 U12043 ( .A1(n9811), .A2(n11067), .ZN(n9553) );
  INV_X1 U12044 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10083) );
  OR2_X1 U12045 ( .A1(n9479), .A2(n10083), .ZN(n9552) );
  NAND4_X1 U12046 ( .A1(n9555), .A2(n9554), .A3(n9553), .A4(n9552), .ZN(n13351) );
  NAND2_X1 U12047 ( .A1(n9558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9557) );
  MUX2_X1 U12048 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9557), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9559) );
  AOI22_X1 U12049 ( .A1(n9556), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9735), .B2(
        n10268), .ZN(n9561) );
  NAND2_X1 U12050 ( .A1(n9932), .A2(n13262), .ZN(n9560) );
  INV_X1 U12051 ( .A(n13129), .ZN(n11274) );
  XNOR2_X1 U12052 ( .A(n13351), .B(n11274), .ZN(n13302) );
  NAND2_X1 U12053 ( .A1(n11055), .A2(n13302), .ZN(n11054) );
  OR2_X1 U12054 ( .A1(n13351), .A2(n13129), .ZN(n9562) );
  NAND2_X1 U12055 ( .A1(n11054), .A2(n9562), .ZN(n11238) );
  OR2_X1 U12056 ( .A1(n9980), .A2(n13091), .ZN(n9565) );
  NAND2_X1 U12057 ( .A1(n9574), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9563) );
  XNOR2_X1 U12058 ( .A(n9563), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U12059 ( .A1(n6400), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9735), .B2(
        n10111), .ZN(n9564) );
  NAND2_X1 U12060 ( .A1(n9565), .A2(n9564), .ZN(n13133) );
  NAND2_X1 U12061 ( .A1(n12277), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9572) );
  INV_X1 U12062 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11248) );
  OR2_X1 U12063 ( .A1(n9814), .A2(n11248), .ZN(n9571) );
  INV_X1 U12064 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U12065 ( .A1(n9567), .A2(n9566), .ZN(n9568) );
  NAND2_X1 U12066 ( .A1(n9579), .A2(n9568), .ZN(n11250) );
  OR2_X1 U12067 ( .A1(n9811), .A2(n11250), .ZN(n9570) );
  INV_X1 U12068 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10085) );
  OR2_X1 U12069 ( .A1(n9479), .A2(n10085), .ZN(n9569) );
  XNOR2_X1 U12070 ( .A(n13133), .B(n13350), .ZN(n13305) );
  INV_X1 U12071 ( .A(n13305), .ZN(n11242) );
  INV_X1 U12072 ( .A(n13133), .ZN(n15440) );
  INV_X1 U12073 ( .A(n13350), .ZN(n11056) );
  NAND2_X1 U12074 ( .A1(n15440), .A2(n11056), .ZN(n9573) );
  NAND2_X1 U12075 ( .A1(n11237), .A2(n9573), .ZN(n11294) );
  NAND2_X1 U12076 ( .A1(n9993), .A2(n13262), .ZN(n9577) );
  OAI21_X1 U12077 ( .B1(n9574), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9575) );
  XNOR2_X1 U12078 ( .A(n9575), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U12079 ( .A1(n6400), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9735), .B2(
        n10114), .ZN(n9576) );
  NAND2_X1 U12080 ( .A1(n12277), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9584) );
  INV_X1 U12081 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10113) );
  OR2_X1 U12082 ( .A1(n9814), .A2(n10113), .ZN(n9583) );
  INV_X1 U12083 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U12084 ( .A1(n9579), .A2(n9578), .ZN(n9580) );
  NAND2_X1 U12085 ( .A1(n9604), .A2(n9580), .ZN(n11222) );
  OR2_X1 U12086 ( .A1(n9811), .A2(n11222), .ZN(n9582) );
  INV_X1 U12087 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15552) );
  OR2_X1 U12088 ( .A1(n9479), .A2(n15552), .ZN(n9581) );
  XNOR2_X1 U12089 ( .A(n13136), .B(n13349), .ZN(n13306) );
  OR2_X1 U12090 ( .A1(n10044), .A2(n13091), .ZN(n9589) );
  NAND2_X1 U12091 ( .A1(n9585), .A2(n9586), .ZN(n9617) );
  NAND2_X1 U12092 ( .A1(n9617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9587) );
  XNOR2_X1 U12093 ( .A(n9587), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U12094 ( .A1(n6400), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9735), .B2(
        n10370), .ZN(n9588) );
  NAND2_X1 U12095 ( .A1(n13099), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9596) );
  INV_X1 U12096 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9590) );
  OR2_X1 U12097 ( .A1(n13100), .A2(n9590), .ZN(n9595) );
  INV_X1 U12098 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U12099 ( .A1(n9606), .A2(n9591), .ZN(n9592) );
  NAND2_X1 U12100 ( .A1(n9621), .A2(n9592), .ZN(n11668) );
  OR2_X1 U12101 ( .A1(n9811), .A2(n11668), .ZN(n9594) );
  INV_X1 U12102 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10363) );
  OR2_X1 U12103 ( .A1(n9479), .A2(n10363), .ZN(n9593) );
  NAND4_X1 U12104 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n13347) );
  OR2_X1 U12105 ( .A1(n10007), .A2(n13091), .ZN(n9601) );
  INV_X1 U12106 ( .A(n9585), .ZN(n9597) );
  NAND2_X1 U12107 ( .A1(n9597), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9598) );
  MUX2_X1 U12108 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9598), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9599) );
  NAND2_X1 U12109 ( .A1(n9599), .A2(n9617), .ZN(n10359) );
  INV_X1 U12110 ( .A(n10359), .ZN(n10367) );
  AOI22_X1 U12111 ( .A1(n9556), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9735), .B2(
        n10367), .ZN(n9600) );
  NAND2_X1 U12112 ( .A1(n13099), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9610) );
  INV_X1 U12113 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9602) );
  OR2_X1 U12114 ( .A1(n13100), .A2(n9602), .ZN(n9609) );
  NAND2_X1 U12115 ( .A1(n9604), .A2(n9603), .ZN(n9605) );
  NAND2_X1 U12116 ( .A1(n9606), .A2(n9605), .ZN(n11580) );
  OR2_X1 U12117 ( .A1(n9811), .A2(n11580), .ZN(n9608) );
  INV_X1 U12118 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10358) );
  OR2_X1 U12119 ( .A1(n9479), .A2(n10358), .ZN(n9607) );
  NAND4_X1 U12120 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n13348) );
  OAI22_X1 U12121 ( .A1(n13148), .A2(n13347), .B1(n13145), .B2(n13348), .ZN(
        n9611) );
  NOR2_X1 U12122 ( .A1(n13136), .A2(n13349), .ZN(n11571) );
  NOR2_X1 U12123 ( .A1(n9611), .A2(n11571), .ZN(n9612) );
  NAND2_X1 U12124 ( .A1(n13145), .A2(n13348), .ZN(n11621) );
  INV_X1 U12125 ( .A(n13347), .ZN(n11692) );
  NAND2_X1 U12126 ( .A1(n11621), .A2(n11692), .ZN(n9613) );
  NAND2_X1 U12127 ( .A1(n13148), .A2(n9613), .ZN(n9615) );
  NAND3_X1 U12128 ( .A1(n13145), .A2(n13347), .A3(n13348), .ZN(n9614) );
  AND2_X1 U12129 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  NAND2_X1 U12130 ( .A1(n9712), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9618) );
  XNOR2_X1 U12131 ( .A(n9618), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U12132 ( .A1(n6400), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9735), 
        .B2(n10591), .ZN(n9619) );
  NAND2_X1 U12133 ( .A1(n12277), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9627) );
  INV_X1 U12134 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11699) );
  OR2_X1 U12135 ( .A1(n9814), .A2(n11699), .ZN(n9626) );
  NAND2_X1 U12136 ( .A1(n9621), .A2(n9620), .ZN(n9622) );
  NAND2_X1 U12137 ( .A1(n9637), .A2(n9622), .ZN(n11744) );
  OR2_X1 U12138 ( .A1(n9811), .A2(n11744), .ZN(n9625) );
  INV_X1 U12139 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9623) );
  OR2_X1 U12140 ( .A1(n9479), .A2(n9623), .ZN(n9624) );
  NAND4_X1 U12141 ( .A1(n9627), .A2(n9626), .A3(n9625), .A4(n9624), .ZN(n13346) );
  INV_X1 U12142 ( .A(n13311), .ZN(n9628) );
  NAND2_X1 U12143 ( .A1(n13152), .A2(n13346), .ZN(n9629) );
  INV_X1 U12144 ( .A(n9712), .ZN(n9632) );
  INV_X1 U12145 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U12146 ( .A1(n9632), .A2(n9631), .ZN(n9645) );
  NAND2_X1 U12147 ( .A1(n9645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9633) );
  XNOR2_X1 U12148 ( .A(n9633), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U12149 ( .A1(n9556), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9735), 
        .B2(n10724), .ZN(n9634) );
  NAND2_X1 U12150 ( .A1(n13099), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9642) );
  INV_X1 U12151 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15641) );
  OR2_X1 U12152 ( .A1(n13100), .A2(n15641), .ZN(n9641) );
  INV_X1 U12153 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12154 ( .A1(n9637), .A2(n9636), .ZN(n9638) );
  NAND2_X1 U12155 ( .A1(n9665), .A2(n9638), .ZN(n11989) );
  OR2_X1 U12156 ( .A1(n9811), .A2(n11989), .ZN(n9640) );
  INV_X1 U12157 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10717) );
  OR2_X1 U12158 ( .A1(n9479), .A2(n10717), .ZN(n9639) );
  NAND4_X1 U12159 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(n13345) );
  AND2_X1 U12160 ( .A1(n7105), .A2(n13345), .ZN(n9644) );
  OR2_X1 U12161 ( .A1(n7105), .A2(n13345), .ZN(n9643) );
  NAND2_X1 U12162 ( .A1(n10150), .A2(n13262), .ZN(n9652) );
  NAND2_X1 U12163 ( .A1(n9647), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9646) );
  MUX2_X1 U12164 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9646), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9650) );
  INV_X1 U12165 ( .A(n9647), .ZN(n9649) );
  INV_X1 U12166 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U12167 ( .A1(n9649), .A2(n9648), .ZN(n9659) );
  NAND2_X1 U12168 ( .A1(n9650), .A2(n9659), .ZN(n11138) );
  INV_X1 U12169 ( .A(n11138), .ZN(n11133) );
  AOI22_X1 U12170 ( .A1(n6400), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11133), 
        .B2(n9735), .ZN(n9651) );
  NAND2_X1 U12171 ( .A1(n12277), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9657) );
  INV_X1 U12172 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9653) );
  OR2_X1 U12173 ( .A1(n9814), .A2(n9653), .ZN(n9656) );
  XNOR2_X1 U12174 ( .A(n9665), .B(n10722), .ZN(n12085) );
  OR2_X1 U12175 ( .A1(n9811), .A2(n12085), .ZN(n9655) );
  INV_X1 U12176 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10716) );
  OR2_X1 U12177 ( .A1(n9479), .A2(n10716), .ZN(n9654) );
  NAND4_X1 U12178 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n13721) );
  XNOR2_X1 U12179 ( .A(n13846), .B(n13721), .ZN(n13313) );
  INV_X1 U12180 ( .A(n13313), .ZN(n12043) );
  NAND2_X1 U12181 ( .A1(n10184), .A2(n13262), .ZN(n9662) );
  NAND2_X1 U12182 ( .A1(n9659), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9658) );
  MUX2_X1 U12183 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9658), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9660) );
  AOI22_X1 U12184 ( .A1(n11608), .A2(n9735), .B1(n6400), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U12185 ( .A1(n13099), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9671) );
  INV_X1 U12186 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9663) );
  OR2_X1 U12187 ( .A1(n13100), .A2(n9663), .ZN(n9670) );
  OAI21_X1 U12188 ( .B1(n9665), .B2(n10722), .A(n9664), .ZN(n9666) );
  NAND2_X1 U12189 ( .A1(n9666), .A2(n9677), .ZN(n13730) );
  OR2_X1 U12190 ( .A1(n9751), .A2(n13730), .ZN(n9669) );
  INV_X1 U12191 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9667) );
  OR2_X1 U12192 ( .A1(n9479), .A2(n9667), .ZN(n9668) );
  NAND4_X1 U12193 ( .A1(n9671), .A2(n9670), .A3(n9669), .A4(n9668), .ZN(n13344) );
  OR2_X1 U12194 ( .A1(n13839), .A2(n13344), .ZN(n9672) );
  NAND2_X1 U12195 ( .A1(n13839), .A2(n13344), .ZN(n9673) );
  NAND2_X1 U12196 ( .A1(n9684), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9674) );
  XNOR2_X1 U12197 ( .A(n9674), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U12198 ( .A1(n11687), .A2(n9735), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n6400), .ZN(n9675) );
  NAND2_X1 U12199 ( .A1(n13099), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9682) );
  INV_X1 U12200 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n13898) );
  OR2_X1 U12201 ( .A1(n13100), .A2(n13898), .ZN(n9681) );
  INV_X1 U12202 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n15606) );
  NAND2_X1 U12203 ( .A1(n9677), .A2(n15606), .ZN(n9678) );
  NAND2_X1 U12204 ( .A1(n9690), .A2(n9678), .ZN(n13709) );
  OR2_X1 U12205 ( .A1(n9811), .A2(n13709), .ZN(n9680) );
  INV_X1 U12206 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n13836) );
  OR2_X1 U12207 ( .A1(n9479), .A2(n13836), .ZN(n9679) );
  NAND4_X1 U12208 ( .A1(n9682), .A2(n9681), .A3(n9680), .A4(n9679), .ZN(n13724) );
  OR2_X1 U12209 ( .A1(n13707), .A2(n13724), .ZN(n9683) );
  NAND2_X1 U12210 ( .A1(n10825), .A2(n13262), .ZN(n9689) );
  OAI21_X1 U12211 ( .B1(n9684), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U12212 ( .A1(n9686), .A2(n9685), .ZN(n9699) );
  OR2_X1 U12213 ( .A1(n9686), .A2(n9685), .ZN(n9687) );
  AOI22_X1 U12214 ( .A1(n11887), .A2(n9735), .B1(P1_DATAO_REG_15__SCAN_IN), 
        .B2(n6400), .ZN(n9688) );
  NAND2_X1 U12215 ( .A1(n9690), .A2(n6689), .ZN(n9691) );
  NAND2_X1 U12216 ( .A1(n9704), .A2(n9691), .ZN(n13684) );
  OR2_X1 U12217 ( .A1(n13684), .A2(n9811), .ZN(n9697) );
  NAND2_X1 U12218 ( .A1(n13099), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9696) );
  INV_X1 U12219 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9692) );
  OR2_X1 U12220 ( .A1(n13100), .A2(n9692), .ZN(n9695) );
  INV_X1 U12221 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9693) );
  OR2_X1 U12222 ( .A1(n9479), .A2(n9693), .ZN(n9694) );
  NAND4_X1 U12223 ( .A1(n9697), .A2(n9696), .A3(n9695), .A4(n9694), .ZN(n13343) );
  INV_X1 U12224 ( .A(n13343), .ZN(n9843) );
  OR2_X1 U12225 ( .A1(n13828), .A2(n13343), .ZN(n9698) );
  NAND2_X1 U12226 ( .A1(n10568), .A2(n13262), .ZN(n9702) );
  NAND2_X1 U12227 ( .A1(n9699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9700) );
  XNOR2_X1 U12228 ( .A(n9700), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U12229 ( .A1(n13407), .A2(n9735), .B1(P1_DATAO_REG_16__SCAN_IN), 
        .B2(n6400), .ZN(n9701) );
  NAND2_X1 U12230 ( .A1(n9704), .A2(n9703), .ZN(n9705) );
  NAND2_X1 U12231 ( .A1(n6493), .A2(n9705), .ZN(n13660) );
  NAND2_X1 U12232 ( .A1(n13099), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U12233 ( .A1(n12277), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9706) );
  AND2_X1 U12234 ( .A1(n9707), .A2(n9706), .ZN(n9709) );
  INV_X1 U12235 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n15531) );
  OR2_X1 U12236 ( .A1(n9479), .A2(n15531), .ZN(n9708) );
  OAI211_X1 U12237 ( .C1(n13660), .C2(n9811), .A(n9709), .B(n9708), .ZN(n13641) );
  XNOR2_X1 U12238 ( .A(n13180), .B(n13641), .ZN(n13667) );
  NAND2_X1 U12239 ( .A1(n13180), .A2(n13641), .ZN(n9710) );
  NAND2_X1 U12240 ( .A1(n10685), .A2(n13262), .ZN(n9715) );
  OAI21_X1 U12241 ( .B1(n9712), .B2(n9711), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9713) );
  XNOR2_X1 U12242 ( .A(n9713), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13410) );
  AOI22_X1 U12243 ( .A1(n6400), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9735), 
        .B2(n13410), .ZN(n9714) );
  INV_X1 U12244 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13647) );
  INV_X1 U12245 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U12246 ( .A1(n6493), .A2(n9716), .ZN(n9717) );
  NAND2_X1 U12247 ( .A1(n9725), .A2(n9717), .ZN(n13646) );
  OR2_X1 U12248 ( .A1(n13646), .A2(n9811), .ZN(n9719) );
  AOI22_X1 U12249 ( .A1(n12277), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n12278), 
        .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n9718) );
  OAI211_X1 U12250 ( .C1(n9814), .C2(n13647), .A(n9719), .B(n9718), .ZN(n13342) );
  NAND2_X1 U12251 ( .A1(n11171), .A2(n13262), .ZN(n9723) );
  NAND2_X1 U12252 ( .A1(n9720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9721) );
  XNOR2_X1 U12253 ( .A(n9721), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13422) );
  AOI22_X1 U12254 ( .A1(n6400), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9735), 
        .B2(n13422), .ZN(n9722) );
  NAND2_X2 U12255 ( .A1(n9723), .A2(n9722), .ZN(n13814) );
  NAND2_X1 U12256 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  AND2_X1 U12257 ( .A1(n9738), .A2(n9726), .ZN(n13631) );
  NAND2_X1 U12258 ( .A1(n13631), .A2(n12282), .ZN(n9731) );
  INV_X1 U12259 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13415) );
  NAND2_X1 U12260 ( .A1(n12277), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U12261 ( .A1(n12278), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9727) );
  OAI211_X1 U12262 ( .C1(n13415), .C2(n9814), .A(n9728), .B(n9727), .ZN(n9729)
         );
  INV_X1 U12263 ( .A(n9729), .ZN(n9730) );
  NAND2_X1 U12264 ( .A1(n9731), .A2(n9730), .ZN(n13642) );
  NOR2_X1 U12265 ( .A1(n13814), .A2(n13642), .ZN(n13620) );
  NAND2_X1 U12266 ( .A1(n13819), .A2(n13342), .ZN(n13619) );
  NAND2_X1 U12267 ( .A1(n13619), .A2(n13294), .ZN(n9733) );
  NOR2_X1 U12268 ( .A1(n13619), .A2(n13294), .ZN(n9732) );
  AOI21_X1 U12269 ( .B1(n13814), .B2(n9733), .A(n9732), .ZN(n9745) );
  AOI22_X1 U12270 ( .A1(n6400), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13433), 
        .B2(n9735), .ZN(n9736) );
  NAND2_X1 U12271 ( .A1(n9738), .A2(n6692), .ZN(n9739) );
  NAND2_X1 U12272 ( .A1(n9749), .A2(n9739), .ZN(n13616) );
  OR2_X1 U12273 ( .A1(n13616), .A2(n9811), .ZN(n9744) );
  INV_X1 U12274 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13427) );
  NAND2_X1 U12275 ( .A1(n12278), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U12276 ( .A1(n12277), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9740) );
  OAI211_X1 U12277 ( .C1(n9814), .C2(n13427), .A(n9741), .B(n9740), .ZN(n9742)
         );
  INV_X1 U12278 ( .A(n9742), .ZN(n9743) );
  NAND2_X1 U12279 ( .A1(n9744), .A2(n9743), .ZN(n13598) );
  NAND2_X1 U12280 ( .A1(n13809), .A2(n13598), .ZN(n13296) );
  OAI211_X1 U12281 ( .C1(n13644), .C2(n13620), .A(n9745), .B(n13296), .ZN(
        n9746) );
  OR2_X1 U12282 ( .A1(n13809), .A2(n13598), .ZN(n13297) );
  NAND2_X1 U12283 ( .A1(n11372), .A2(n13262), .ZN(n9748) );
  NAND2_X1 U12284 ( .A1(n6400), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U12285 ( .A1(n9749), .A2(n13044), .ZN(n9750) );
  NAND2_X1 U12286 ( .A1(n9762), .A2(n9750), .ZN(n13603) );
  OR2_X1 U12287 ( .A1(n13603), .A2(n9751), .ZN(n9757) );
  INV_X1 U12288 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U12289 ( .A1(n12278), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9753) );
  NAND2_X1 U12290 ( .A1(n12277), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9752) );
  OAI211_X1 U12291 ( .C1(n9814), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9755)
         );
  INV_X1 U12292 ( .A(n9755), .ZN(n9756) );
  NAND2_X1 U12293 ( .A1(n9757), .A2(n9756), .ZN(n13341) );
  NAND2_X1 U12294 ( .A1(n13804), .A2(n13341), .ZN(n9758) );
  OR2_X1 U12295 ( .A1(n13804), .A2(n13341), .ZN(n9759) );
  NAND2_X1 U12296 ( .A1(n11497), .A2(n13262), .ZN(n9761) );
  NAND2_X1 U12297 ( .A1(n9556), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U12298 ( .A1(n9762), .A2(n15549), .ZN(n9763) );
  AND2_X1 U12299 ( .A1(n9777), .A2(n9763), .ZN(n13588) );
  NAND2_X1 U12300 ( .A1(n13588), .A2(n12282), .ZN(n9769) );
  INV_X1 U12301 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9766) );
  NAND2_X1 U12302 ( .A1(n12278), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U12303 ( .A1(n12277), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9764) );
  OAI211_X1 U12304 ( .C1(n9814), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9767)
         );
  INV_X1 U12305 ( .A(n9767), .ZN(n9768) );
  XNOR2_X1 U12306 ( .A(n13587), .B(n13599), .ZN(n13576) );
  OR2_X1 U12307 ( .A1(n13587), .A2(n13599), .ZN(n9770) );
  XNOR2_X1 U12308 ( .A(n9773), .B(n9772), .ZN(n11669) );
  NAND2_X1 U12309 ( .A1(n6400), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9774) );
  NAND2_X2 U12310 ( .A1(n9775), .A2(n9774), .ZN(n13792) );
  INV_X1 U12311 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U12312 ( .A1(n9777), .A2(n9776), .ZN(n9778) );
  NAND2_X1 U12313 ( .A1(n9788), .A2(n9778), .ZN(n13567) );
  OR2_X1 U12314 ( .A1(n13567), .A2(n9811), .ZN(n9783) );
  INV_X1 U12315 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13568) );
  NAND2_X1 U12316 ( .A1(n12278), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9780) );
  NAND2_X1 U12317 ( .A1(n12277), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9779) );
  OAI211_X1 U12318 ( .C1(n9814), .C2(n13568), .A(n9780), .B(n9779), .ZN(n9781)
         );
  INV_X1 U12319 ( .A(n9781), .ZN(n9782) );
  NAND2_X1 U12320 ( .A1(n13792), .A2(n13340), .ZN(n9784) );
  NAND2_X1 U12321 ( .A1(n11494), .A2(n13262), .ZN(n9786) );
  NAND2_X1 U12322 ( .A1(n6400), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9785) );
  INV_X1 U12323 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U12324 ( .A1(n9788), .A2(n9787), .ZN(n9789) );
  NAND2_X1 U12325 ( .A1(n9797), .A2(n9789), .ZN(n13545) );
  OR2_X1 U12326 ( .A1(n13545), .A2(n9811), .ZN(n9794) );
  INV_X1 U12327 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13546) );
  NAND2_X1 U12328 ( .A1(n12278), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U12329 ( .A1(n12277), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9790) );
  OAI211_X1 U12330 ( .C1(n9814), .C2(n13546), .A(n9791), .B(n9790), .ZN(n9792)
         );
  INV_X1 U12331 ( .A(n9792), .ZN(n9793) );
  NAND2_X1 U12332 ( .A1(n11995), .A2(n13262), .ZN(n9796) );
  NAND2_X1 U12333 ( .A1(n6400), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9795) );
  NAND2_X1 U12334 ( .A1(n9797), .A2(n13034), .ZN(n9798) );
  AND2_X1 U12335 ( .A1(n9808), .A2(n9798), .ZN(n13534) );
  NAND2_X1 U12336 ( .A1(n13534), .A2(n12282), .ZN(n9804) );
  INV_X1 U12337 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9801) );
  NAND2_X1 U12338 ( .A1(n12278), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U12339 ( .A1(n12277), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9799) );
  OAI211_X1 U12340 ( .C1(n9814), .C2(n9801), .A(n9800), .B(n9799), .ZN(n9802)
         );
  INV_X1 U12341 ( .A(n9802), .ZN(n9803) );
  XNOR2_X1 U12342 ( .A(n13535), .B(n13339), .ZN(n13526) );
  NAND2_X1 U12343 ( .A1(n13915), .A2(n13262), .ZN(n9806) );
  NAND2_X1 U12344 ( .A1(n6400), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9805) );
  NAND2_X2 U12345 ( .A1(n9806), .A2(n9805), .ZN(n13521) );
  INV_X1 U12346 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U12347 ( .A1(n9810), .A2(n9809), .ZN(n13519) );
  INV_X1 U12348 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13518) );
  NAND2_X1 U12349 ( .A1(n12277), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U12350 ( .A1(n12278), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9812) );
  OAI211_X1 U12351 ( .C1(n9814), .C2(n13518), .A(n9813), .B(n9812), .ZN(n9815)
         );
  INV_X1 U12352 ( .A(n9815), .ZN(n9816) );
  XOR2_X1 U12353 ( .A(n13450), .B(n13451), .Z(n13492) );
  INV_X1 U12354 ( .A(n13148), .ZN(n11626) );
  AND2_X2 U12355 ( .A1(n11624), .A2(n11626), .ZN(n11695) );
  INV_X1 U12356 ( .A(n13152), .ZN(n11698) );
  INV_X1 U12357 ( .A(n13839), .ZN(n13734) );
  INV_X1 U12358 ( .A(n13819), .ZN(n13650) );
  NAND2_X1 U12359 ( .A1(n13658), .A2(n13650), .ZN(n13652) );
  OR2_X2 U12360 ( .A1(n13564), .A2(n13880), .ZN(n13543) );
  NOR2_X2 U12361 ( .A1(n13543), .A2(n13535), .ZN(n13532) );
  NAND2_X1 U12362 ( .A1(n13506), .A2(n13491), .ZN(n9820) );
  NAND2_X1 U12363 ( .A1(n9820), .A2(n13840), .ZN(n9821) );
  INV_X1 U12364 ( .A(n11051), .ZN(n15420) );
  INV_X1 U12365 ( .A(n13113), .ZN(n11257) );
  OR2_X1 U12366 ( .A1(n10801), .A2(n11257), .ZN(n10975) );
  NAND2_X1 U12367 ( .A1(n10976), .A2(n10975), .ZN(n9823) );
  NAND2_X1 U12368 ( .A1(n10750), .A2(n10751), .ZN(n9824) );
  NAND2_X1 U12369 ( .A1(n9824), .A2(n13299), .ZN(n10749) );
  INV_X1 U12370 ( .A(n13119), .ZN(n11029) );
  OR2_X1 U12371 ( .A1(n13353), .A2(n11029), .ZN(n10999) );
  NAND2_X1 U12372 ( .A1(n10749), .A2(n10999), .ZN(n9825) );
  NAND2_X1 U12373 ( .A1(n9825), .A2(n13304), .ZN(n10998) );
  OR2_X1 U12374 ( .A1(n13352), .A2(n7686), .ZN(n11059) );
  NAND2_X1 U12375 ( .A1(n10998), .A2(n11059), .ZN(n9827) );
  INV_X1 U12376 ( .A(n13302), .ZN(n9826) );
  OR2_X1 U12377 ( .A1(n13351), .A2(n11274), .ZN(n11241) );
  INV_X1 U12378 ( .A(n13136), .ZN(n11462) );
  NAND2_X1 U12379 ( .A1(n11462), .A2(n13349), .ZN(n9829) );
  INV_X1 U12380 ( .A(n13349), .ZN(n11239) );
  INV_X1 U12381 ( .A(n13145), .ZN(n11581) );
  NAND2_X1 U12382 ( .A1(n11581), .A2(n13348), .ZN(n9831) );
  XNOR2_X1 U12383 ( .A(n13148), .B(n13347), .ZN(n13310) );
  NAND2_X1 U12384 ( .A1(n11626), .A2(n13347), .ZN(n9832) );
  NAND2_X1 U12385 ( .A1(n11698), .A2(n13346), .ZN(n9833) );
  INV_X1 U12386 ( .A(n13315), .ZN(n11859) );
  INV_X1 U12387 ( .A(n13345), .ZN(n12045) );
  NAND2_X1 U12388 ( .A1(n7105), .A2(n12045), .ZN(n9834) );
  AND2_X1 U12389 ( .A1(n13839), .A2(n13695), .ZN(n9836) );
  INV_X1 U12390 ( .A(n13721), .ZN(n11852) );
  AND2_X1 U12391 ( .A1(n13846), .A2(n11852), .ZN(n9835) );
  XNOR2_X1 U12392 ( .A(n13707), .B(n13724), .ZN(n13703) );
  OR2_X1 U12393 ( .A1(n13846), .A2(n11852), .ZN(n13693) );
  NAND2_X1 U12394 ( .A1(n13693), .A2(n13695), .ZN(n9838) );
  INV_X1 U12395 ( .A(n13846), .ZN(n12091) );
  AND2_X1 U12396 ( .A1(n13344), .A2(n13721), .ZN(n9837) );
  AOI22_X1 U12397 ( .A1(n9838), .A2(n13734), .B1(n12091), .B2(n9837), .ZN(
        n9839) );
  INV_X1 U12398 ( .A(n13724), .ZN(n13677) );
  NAND2_X1 U12399 ( .A1(n13707), .A2(n13677), .ZN(n9842) );
  OR2_X1 U12400 ( .A1(n13828), .A2(n9843), .ZN(n9844) );
  INV_X1 U12401 ( .A(n13641), .ZN(n13679) );
  OR2_X1 U12402 ( .A1(n13180), .A2(n13679), .ZN(n9845) );
  INV_X1 U12403 ( .A(n13342), .ZN(n13060) );
  NAND2_X1 U12404 ( .A1(n13819), .A2(n13060), .ZN(n9846) );
  NAND2_X1 U12405 ( .A1(n13640), .A2(n9846), .ZN(n9848) );
  OR2_X1 U12406 ( .A1(n13819), .A2(n13060), .ZN(n9847) );
  NAND2_X1 U12407 ( .A1(n13814), .A2(n13294), .ZN(n9849) );
  INV_X1 U12408 ( .A(n13598), .ZN(n13192) );
  AND2_X1 U12409 ( .A1(n13809), .A2(n13192), .ZN(n9850) );
  INV_X1 U12410 ( .A(n13599), .ZN(n13558) );
  OR2_X1 U12411 ( .A1(n13804), .A2(n13581), .ZN(n13295) );
  OAI21_X1 U12412 ( .B1(n13587), .B2(n13558), .A(n13295), .ZN(n9854) );
  NAND2_X1 U12413 ( .A1(n13804), .A2(n13581), .ZN(n13557) );
  INV_X1 U12414 ( .A(n13557), .ZN(n13575) );
  NAND2_X1 U12415 ( .A1(n13557), .A2(n13599), .ZN(n9851) );
  AOI22_X1 U12416 ( .A1(n13575), .A2(n13558), .B1(n9851), .B2(n13587), .ZN(
        n9852) );
  AND2_X1 U12417 ( .A1(n9852), .A2(n13571), .ZN(n9853) );
  INV_X1 U12418 ( .A(n13340), .ZN(n13580) );
  INV_X1 U12419 ( .A(n13561), .ZN(n13293) );
  NOR2_X1 U12420 ( .A1(n13880), .A2(n13293), .ZN(n9856) );
  NAND2_X1 U12421 ( .A1(n13880), .A2(n13293), .ZN(n9855) );
  INV_X1 U12422 ( .A(n13339), .ZN(n13196) );
  AND2_X1 U12423 ( .A1(n13535), .A2(n13196), .ZN(n9857) );
  OR2_X1 U12424 ( .A1(n13771), .A2(n13232), .ZN(n13292) );
  NAND2_X1 U12425 ( .A1(n13771), .A2(n13232), .ZN(n13291) );
  NOR2_X1 U12426 ( .A1(n9859), .A2(n13666), .ZN(n13105) );
  AND2_X1 U12427 ( .A1(n13323), .A2(n13298), .ZN(n9860) );
  INV_X1 U12428 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U12429 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  NAND2_X1 U12430 ( .A1(n12276), .A2(n12282), .ZN(n9869) );
  INV_X1 U12431 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15576) );
  NAND2_X1 U12432 ( .A1(n9503), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12433 ( .A1(n12277), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9865) );
  OAI211_X1 U12434 ( .C1(n15576), .C2(n9479), .A(n9866), .B(n9865), .ZN(n9867)
         );
  INV_X1 U12435 ( .A(n9867), .ZN(n9868) );
  INV_X1 U12436 ( .A(n10812), .ZN(n10088) );
  AOI211_X1 U12437 ( .C1(n13835), .C2(n13492), .A(n13493), .B(n13487), .ZN(
        n13866) );
  INV_X1 U12438 ( .A(n11997), .ZN(n9895) );
  INV_X1 U12439 ( .A(n9880), .ZN(n9883) );
  NAND2_X1 U12440 ( .A1(n9883), .A2(n9882), .ZN(n9888) );
  INV_X1 U12441 ( .A(n9888), .ZN(n9885) );
  NAND2_X1 U12442 ( .A1(n9885), .A2(n9884), .ZN(n9890) );
  NAND2_X1 U12443 ( .A1(n9890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9886) );
  MUX2_X1 U12444 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9886), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9887) );
  XNOR2_X1 U12445 ( .A(n11997), .B(P2_B_REG_SCAN_IN), .ZN(n9892) );
  NAND2_X1 U12446 ( .A1(n9888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9889) );
  MUX2_X1 U12447 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9889), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9891) );
  NAND2_X1 U12448 ( .A1(n9892), .A2(n13918), .ZN(n9893) );
  INV_X1 U12449 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15414) );
  NAND2_X1 U12450 ( .A1(n15412), .A2(n15414), .ZN(n9894) );
  NOR2_X1 U12451 ( .A1(n15415), .A2(n10820), .ZN(n9912) );
  NOR4_X1 U12452 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9899) );
  NOR4_X1 U12453 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9898) );
  NOR4_X1 U12454 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n9897) );
  NOR4_X1 U12455 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n9896) );
  AND4_X1 U12456 ( .A1(n9899), .A2(n9898), .A3(n9897), .A4(n9896), .ZN(n9904)
         );
  NOR2_X1 U12457 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n15545) );
  NOR4_X1 U12458 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9902) );
  NOR4_X1 U12459 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9901) );
  NOR4_X1 U12460 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9900) );
  AND4_X1 U12461 ( .A1(n15545), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9903)
         );
  NAND2_X1 U12462 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  OR2_X1 U12463 ( .A1(n10812), .A2(n13286), .ZN(n10815) );
  INV_X1 U12464 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15418) );
  NAND2_X1 U12465 ( .A1(n15412), .A2(n15418), .ZN(n9909) );
  NAND2_X1 U12466 ( .A1(n11949), .A2(n13918), .ZN(n9908) );
  NAND2_X1 U12467 ( .A1(n9910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9911) );
  AND2_X1 U12468 ( .A1(n10972), .A2(n15416), .ZN(n15417) );
  MUX2_X1 U12469 ( .A(n15532), .B(n13866), .S(n15454), .Z(n9914) );
  INV_X1 U12470 ( .A(n13491), .ZN(n13869) );
  NAND2_X1 U12471 ( .A1(n13491), .A2(n13789), .ZN(n9913) );
  NAND2_X1 U12472 ( .A1(n9914), .A2(n9913), .ZN(P2_U3526) );
  INV_X4 U12473 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U12474 ( .A(n10233), .ZN(n9915) );
  AOI222_X1 U12475 ( .A1(n9917), .A2(n12929), .B1(n10443), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n10509), .ZN(n9918) );
  INV_X1 U12476 ( .A(n9918), .ZN(P3_U3291) );
  AOI222_X1 U12477 ( .A1(n9919), .A2(n12929), .B1(n6399), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_2_), .C2(n10509), .ZN(n9920) );
  INV_X1 U12478 ( .A(n9920), .ZN(P3_U3293) );
  AOI222_X1 U12479 ( .A1(n9921), .A2(n12929), .B1(n10412), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_5_), .C2(n10509), .ZN(n9922) );
  INV_X1 U12480 ( .A(n9922), .ZN(P3_U3290) );
  AOI222_X1 U12481 ( .A1(n9923), .A2(n12929), .B1(n10455), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n10509), .ZN(n9924) );
  INV_X1 U12482 ( .A(n9924), .ZN(P3_U3292) );
  INV_X2 U12483 ( .A(n13910), .ZN(n13916) );
  INV_X1 U12484 ( .A(n13389), .ZN(n13382) );
  OAI222_X1 U12485 ( .A1(n13916), .A2(n9925), .B1(n13913), .B2(n9967), .C1(
        n13382), .C2(P2_U3088), .ZN(P2_U3324) );
  OAI222_X1 U12486 ( .A1(n13916), .A2(n9926), .B1(n13913), .B2(n9968), .C1(
        n13362), .C2(P2_U3088), .ZN(P2_U3326) );
  OAI222_X1 U12487 ( .A1(n13916), .A2(n9927), .B1(n13913), .B2(n9970), .C1(
        P2_U3088), .C2(n13372), .ZN(P2_U3325) );
  INV_X2 U12488 ( .A(n10509), .ZN(n12941) );
  INV_X1 U12489 ( .A(n12929), .ZN(n12948) );
  INV_X1 U12490 ( .A(n10640), .ZN(n10634) );
  OAI222_X1 U12491 ( .A1(n12941), .A2(n9929), .B1(n12948), .B2(n9928), .C1(
        P3_U3151), .C2(n10634), .ZN(P3_U3289) );
  OAI222_X1 U12492 ( .A1(n12941), .A2(n9931), .B1(n12948), .B2(n9930), .C1(
        n10321), .C2(P3_U3151), .ZN(P3_U3294) );
  INV_X1 U12493 ( .A(n9932), .ZN(n9982) );
  AOI22_X1 U12494 ( .A1(n10268), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n13910), .ZN(n9933) );
  OAI21_X1 U12495 ( .B1(n9982), .B2(n13913), .A(n9933), .ZN(P2_U3322) );
  OAI222_X1 U12496 ( .A1(n10878), .A2(P3_U3151), .B1(n12948), .B2(n9935), .C1(
        n9934), .C2(n12941), .ZN(P3_U3288) );
  NAND2_X1 U12497 ( .A1(n9948), .A2(n9949), .ZN(n9937) );
  INV_X1 U12498 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14583) );
  NAND2_X1 U12499 ( .A1(n14583), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U12500 ( .A1(n9937), .A2(n9936), .ZN(n9947) );
  NAND2_X1 U12501 ( .A1(n14602), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U12502 ( .A1(n10336), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U12503 ( .A1(n9947), .A2(n9946), .ZN(n9940) );
  NAND2_X1 U12504 ( .A1(n9940), .A2(n9939), .ZN(n9941) );
  NAND2_X1 U12505 ( .A1(n9941), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n9943) );
  INV_X1 U12506 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9944) );
  XNOR2_X1 U12507 ( .A(n9988), .B(n9944), .ZN(n9983) );
  XNOR2_X1 U12508 ( .A(n9983), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n9961) );
  XNOR2_X1 U12509 ( .A(n9945), .B(n6881), .ZN(n9955) );
  XNOR2_X1 U12510 ( .A(n9947), .B(n9946), .ZN(n15202) );
  NAND2_X1 U12511 ( .A1(n15202), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n9952) );
  XNOR2_X1 U12512 ( .A(n9948), .B(n9949), .ZN(n9951) );
  INV_X1 U12513 ( .A(n9949), .ZN(n9950) );
  OAI21_X1 U12514 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n10069), .A(n9950), .ZN(
        n15153) );
  NAND2_X1 U12515 ( .A1(n15153), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n15669) );
  XNOR2_X1 U12516 ( .A(n9951), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15668) );
  NOR2_X1 U12517 ( .A1(n15669), .A2(n15668), .ZN(n15667) );
  AOI21_X1 U12518 ( .B1(n9951), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n15667), .ZN(
        n15201) );
  NAND2_X1 U12519 ( .A1(n9952), .A2(n15201), .ZN(n9954) );
  OR2_X1 U12520 ( .A1(n15202), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U12521 ( .A1(n9954), .A2(n9953), .ZN(n9956) );
  NAND2_X1 U12522 ( .A1(n9955), .A2(n9956), .ZN(n15664) );
  NAND2_X1 U12523 ( .A1(n15664), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n9959) );
  INV_X1 U12524 ( .A(n9955), .ZN(n9958) );
  INV_X1 U12525 ( .A(n9956), .ZN(n9957) );
  NAND2_X1 U12526 ( .A1(n9958), .A2(n9957), .ZN(n15665) );
  NAND2_X1 U12527 ( .A1(n9959), .A2(n15665), .ZN(n9960) );
  NAND2_X1 U12528 ( .A1(n9961), .A2(n9960), .ZN(n9986) );
  OAI21_X1 U12529 ( .B1(n9961), .B2(n9960), .A(n9986), .ZN(n9962) );
  INV_X1 U12530 ( .A(n9962), .ZN(SUB_1596_U59) );
  OAI222_X1 U12531 ( .A1(n11486), .A2(P3_U3151), .B1(n12948), .B2(n9964), .C1(
        n9963), .C2(n12941), .ZN(P3_U3286) );
  INV_X1 U12532 ( .A(n9965), .ZN(n9966) );
  OAI222_X1 U12533 ( .A1(n12941), .A2(n6615), .B1(n12948), .B2(n9966), .C1(
        n11479), .C2(P3_U3151), .ZN(P3_U3287) );
  AND2_X1 U12534 ( .A1(n7434), .A2(P1_U3086), .ZN(n10140) );
  INV_X2 U12535 ( .A(n10140), .ZN(n15144) );
  NOR2_X1 U12536 ( .A1(n7434), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15139) );
  INV_X2 U12537 ( .A(n15139), .ZN(n15147) );
  OAI222_X1 U12538 ( .A1(P1_U3086), .A2(n14621), .B1(n15144), .B2(n7089), .C1(
        n15147), .C2(n9967), .ZN(P1_U3352) );
  OAI222_X1 U12539 ( .A1(P1_U3086), .A2(n14586), .B1(n15144), .B2(n7139), .C1(
        n15147), .C2(n9968), .ZN(P1_U3354) );
  OAI222_X1 U12540 ( .A1(n14605), .A2(P1_U3086), .B1(n15147), .B2(n9970), .C1(
        n9969), .C2(n15144), .ZN(P1_U3353) );
  INV_X1 U12541 ( .A(n9971), .ZN(n9976) );
  OAI222_X1 U12542 ( .A1(n15220), .A2(P1_U3086), .B1(n15147), .B2(n9976), .C1(
        n9972), .C2(n15144), .ZN(P1_U3351) );
  OAI222_X1 U12543 ( .A1(n11917), .A2(P3_U3151), .B1(n12948), .B2(n9974), .C1(
        n9973), .C2(n12941), .ZN(P3_U3285) );
  INV_X1 U12544 ( .A(n10111), .ZN(n15351) );
  OAI222_X1 U12545 ( .A1(P2_U3088), .A2(n15351), .B1(n13916), .B2(n9975), .C1(
        n13913), .C2(n9980), .ZN(P2_U3321) );
  OAI222_X1 U12546 ( .A1(n13916), .A2(n9977), .B1(n13913), .B2(n9976), .C1(
        P2_U3088), .C2(n15336), .ZN(P2_U3323) );
  INV_X1 U12547 ( .A(n10220), .ZN(n9978) );
  OAI222_X1 U12548 ( .A1(n15147), .A2(n9980), .B1(n15144), .B2(n9979), .C1(
        n9978), .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U12549 ( .A1(n15147), .A2(n9982), .B1(n15144), .B2(n9981), .C1(
        n10176), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U12550 ( .A(n9983), .ZN(n9984) );
  NAND2_X1 U12551 ( .A1(n9984), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U12552 ( .A1(n9986), .A2(n9985), .ZN(n10049) );
  OAI21_X1 U12553 ( .B1(n9988), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9987), .ZN(
        n9989) );
  NAND2_X1 U12554 ( .A1(n9989), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U12555 ( .A1(n10053), .A2(n9990), .ZN(n10052) );
  INV_X1 U12556 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10190) );
  XNOR2_X1 U12557 ( .A(n10052), .B(n10190), .ZN(n10047) );
  XNOR2_X1 U12558 ( .A(n10049), .B(n10047), .ZN(n10046) );
  INV_X1 U12559 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10270) );
  XNOR2_X1 U12560 ( .A(n10046), .B(n10270), .ZN(SUB_1596_U58) );
  OAI222_X1 U12561 ( .A1(P3_U3151), .A2(n11927), .B1(n12948), .B2(n9992), .C1(
        n9991), .C2(n12941), .ZN(P3_U3284) );
  INV_X1 U12562 ( .A(n9993), .ZN(n9995) );
  INV_X1 U12563 ( .A(n10221), .ZN(n10357) );
  OAI222_X1 U12564 ( .A1(n15147), .A2(n9995), .B1(n10357), .B2(P1_U3086), .C1(
        n9994), .C2(n15144), .ZN(P1_U3348) );
  INV_X1 U12565 ( .A(n10114), .ZN(n15365) );
  INV_X1 U12566 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9996) );
  OAI222_X1 U12567 ( .A1(P2_U3088), .A2(n15365), .B1(n13916), .B2(n9996), .C1(
        n13913), .C2(n9995), .ZN(P2_U3320) );
  INV_X1 U12568 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15593) );
  NAND2_X1 U12569 ( .A1(n10836), .A2(P3_U3897), .ZN(n9997) );
  OAI21_X1 U12570 ( .B1(P3_U3897), .B2(n15593), .A(n9997), .ZN(P3_U3494) );
  INV_X1 U12571 ( .A(n10312), .ZN(n10218) );
  OAI222_X1 U12572 ( .A1(n15147), .A2(n10007), .B1(n10218), .B2(P1_U3086), 
        .C1(n7094), .C2(n15144), .ZN(P1_U3347) );
  INV_X1 U12573 ( .A(n12021), .ZN(n12476) );
  OAI222_X1 U12574 ( .A1(n12941), .A2(n9999), .B1(n12948), .B2(n9998), .C1(
        n12476), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12575 ( .A(n10288), .ZN(n10282) );
  INV_X1 U12576 ( .A(n10297), .ZN(n10000) );
  INV_X1 U12577 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n15640) );
  INV_X1 U12578 ( .A(n10279), .ZN(n10002) );
  INV_X1 U12579 ( .A(n10001), .ZN(n10004) );
  AOI22_X1 U12580 ( .A1(n15270), .A2(n15640), .B1(n10002), .B2(n10004), .ZN(
        P1_U3446) );
  INV_X1 U12581 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10006) );
  INV_X1 U12582 ( .A(n10003), .ZN(n10005) );
  AOI22_X1 U12583 ( .A1(n15270), .A2(n10006), .B1(n10005), .B2(n10004), .ZN(
        P1_U3445) );
  INV_X1 U12584 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10008) );
  OAI222_X1 U12585 ( .A1(P2_U3088), .A2(n10359), .B1(n13916), .B2(n10008), 
        .C1(n13913), .C2(n10007), .ZN(P2_U3319) );
  INV_X1 U12586 ( .A(n12922), .ZN(n10009) );
  NOR2_X1 U12587 ( .A1(n10010), .A2(n10009), .ZN(n10019) );
  CLKBUF_X1 U12588 ( .A(n10019), .Z(n10040) );
  INV_X1 U12589 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10011) );
  NOR2_X1 U12590 ( .A1(n10040), .A2(n10011), .ZN(P3_U3256) );
  INV_X1 U12591 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10012) );
  NOR2_X1 U12592 ( .A1(n10040), .A2(n10012), .ZN(P3_U3257) );
  INV_X1 U12593 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U12594 ( .A1(n10040), .A2(n10013), .ZN(P3_U3250) );
  INV_X1 U12595 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U12596 ( .A1(n10040), .A2(n10014), .ZN(P3_U3249) );
  INV_X1 U12597 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10015) );
  NOR2_X1 U12598 ( .A1(n10040), .A2(n10015), .ZN(P3_U3248) );
  INV_X1 U12599 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U12600 ( .A1(n10040), .A2(n10016), .ZN(P3_U3247) );
  INV_X1 U12601 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U12602 ( .A1(n10040), .A2(n10017), .ZN(P3_U3246) );
  INV_X1 U12603 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U12604 ( .A1(n10040), .A2(n10018), .ZN(P3_U3252) );
  INV_X1 U12605 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10020) );
  NOR2_X1 U12606 ( .A1(n10040), .A2(n10020), .ZN(P3_U3258) );
  INV_X1 U12607 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10021) );
  NOR2_X1 U12608 ( .A1(n10019), .A2(n10021), .ZN(P3_U3243) );
  INV_X1 U12609 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n15644) );
  NOR2_X1 U12610 ( .A1(n10019), .A2(n15644), .ZN(P3_U3242) );
  INV_X1 U12611 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U12612 ( .A1(n10019), .A2(n10022), .ZN(P3_U3241) );
  INV_X1 U12613 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10023) );
  NOR2_X1 U12614 ( .A1(n10019), .A2(n10023), .ZN(P3_U3240) );
  INV_X1 U12615 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U12616 ( .A1(n10019), .A2(n10024), .ZN(P3_U3239) );
  INV_X1 U12617 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10025) );
  NOR2_X1 U12618 ( .A1(n10019), .A2(n10025), .ZN(P3_U3238) );
  INV_X1 U12619 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U12620 ( .A1(n10019), .A2(n10026), .ZN(P3_U3237) );
  INV_X1 U12621 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10027) );
  NOR2_X1 U12622 ( .A1(n10019), .A2(n10027), .ZN(P3_U3236) );
  INV_X1 U12623 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U12624 ( .A1(n10040), .A2(n10028), .ZN(P3_U3251) );
  INV_X1 U12625 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15548) );
  NOR2_X1 U12626 ( .A1(n10019), .A2(n15548), .ZN(P3_U3234) );
  INV_X1 U12627 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U12628 ( .A1(n10040), .A2(n10029), .ZN(P3_U3254) );
  INV_X1 U12629 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U12630 ( .A1(n10040), .A2(n10030), .ZN(P3_U3253) );
  INV_X1 U12631 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U12632 ( .A1(n10040), .A2(n10031), .ZN(P3_U3261) );
  INV_X1 U12633 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U12634 ( .A1(n10019), .A2(n10032), .ZN(P3_U3235) );
  INV_X1 U12635 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10033) );
  NOR2_X1 U12636 ( .A1(n10019), .A2(n10033), .ZN(P3_U3245) );
  INV_X1 U12637 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U12638 ( .A1(n10040), .A2(n10034), .ZN(P3_U3263) );
  INV_X1 U12639 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U12640 ( .A1(n10040), .A2(n10035), .ZN(P3_U3262) );
  INV_X1 U12641 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10036) );
  NOR2_X1 U12642 ( .A1(n10040), .A2(n10036), .ZN(P3_U3260) );
  INV_X1 U12643 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10037) );
  NOR2_X1 U12644 ( .A1(n10040), .A2(n10037), .ZN(P3_U3255) );
  INV_X1 U12645 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U12646 ( .A1(n10040), .A2(n10038), .ZN(P3_U3244) );
  INV_X1 U12647 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U12648 ( .A1(n10040), .A2(n10039), .ZN(P3_U3259) );
  OR2_X1 U12649 ( .A1(n10041), .A2(P1_U3086), .ZN(n14561) );
  NAND2_X1 U12650 ( .A1(n10297), .A2(n14561), .ZN(n10063) );
  INV_X1 U12651 ( .A(n14478), .ZN(n10294) );
  NAND2_X1 U12652 ( .A1(n10294), .A2(n10041), .ZN(n10042) );
  NAND2_X1 U12653 ( .A1(n10042), .A2(n6397), .ZN(n10061) );
  INV_X1 U12654 ( .A(n15226), .ZN(n14653) );
  NOR2_X1 U12655 ( .A1(n14653), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12656 ( .A(n10317), .ZN(n10464) );
  OAI222_X1 U12657 ( .A1(n15147), .A2(n10044), .B1(n10464), .B2(P1_U3086), 
        .C1(n10043), .C2(n15144), .ZN(P1_U3346) );
  INV_X1 U12658 ( .A(n10370), .ZN(n15390) );
  INV_X1 U12659 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10045) );
  OAI222_X1 U12660 ( .A1(P2_U3088), .A2(n15390), .B1(n13916), .B2(n10045), 
        .C1(n13913), .C2(n10044), .ZN(P2_U3318) );
  NAND2_X1 U12661 ( .A1(n10046), .A2(n10270), .ZN(n10051) );
  INV_X1 U12662 ( .A(n10047), .ZN(n10048) );
  OR2_X1 U12663 ( .A1(n10049), .A2(n10048), .ZN(n10050) );
  NAND2_X1 U12664 ( .A1(n10051), .A2(n10050), .ZN(n10482) );
  XNOR2_X1 U12665 ( .A(n10482), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n10056) );
  INV_X1 U12666 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10480) );
  XNOR2_X1 U12667 ( .A(n10480), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n10478) );
  XNOR2_X1 U12668 ( .A(n10479), .B(n10478), .ZN(n10055) );
  NAND2_X1 U12669 ( .A1(n10056), .A2(n10055), .ZN(n10485) );
  OAI21_X1 U12670 ( .B1(n10056), .B2(n10055), .A(n10485), .ZN(n10057) );
  INV_X1 U12671 ( .A(n10057), .ZN(SUB_1596_U57) );
  INV_X1 U12672 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n15567) );
  NAND2_X1 U12673 ( .A1(n11365), .A2(P3_U3897), .ZN(n10058) );
  OAI21_X1 U12674 ( .B1(P3_U3897), .B2(n15567), .A(n10058), .ZN(P3_U3500) );
  INV_X1 U12675 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15565) );
  NAND2_X1 U12676 ( .A1(n11955), .A2(P3_U3897), .ZN(n10059) );
  OAI21_X1 U12677 ( .B1(P3_U3897), .B2(n15565), .A(n10059), .ZN(P3_U3502) );
  MUX2_X1 U12678 ( .A(n10571), .B(n15082), .S(P1_U4016), .Z(n10060) );
  INV_X1 U12679 ( .A(n10060), .ZN(P1_U3574) );
  INV_X1 U12680 ( .A(n10061), .ZN(n10062) );
  NAND2_X1 U12681 ( .A1(n10063), .A2(n10062), .ZN(n10156) );
  INV_X1 U12682 ( .A(n6410), .ZN(n10064) );
  INV_X1 U12683 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10287) );
  NAND3_X1 U12684 ( .A1(n15210), .A2(n7069), .A3(n10287), .ZN(n10068) );
  INV_X1 U12685 ( .A(n10156), .ZN(n10170) );
  OAI21_X1 U12686 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n6410), .A(n10155), .ZN(
        n14601) );
  AOI21_X1 U12687 ( .B1(n6410), .B2(n10287), .A(n14601), .ZN(n10065) );
  MUX2_X1 U12688 ( .A(n14601), .B(n10065), .S(n7040), .Z(n10066) );
  AOI22_X1 U12689 ( .A1(n10170), .A2(n10066), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10067) );
  OAI211_X1 U12690 ( .C1(n15226), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        P1_U3243) );
  INV_X1 U12691 ( .A(n12498), .ZN(n12478) );
  OAI222_X1 U12692 ( .A1(n12941), .A2(n10071), .B1(n12948), .B2(n10070), .C1(
        n12478), .C2(P3_U3151), .ZN(P3_U3282) );
  AND2_X1 U12693 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10073) );
  NAND2_X1 U12694 ( .A1(n10074), .A2(n10073), .ZN(n13366) );
  INV_X1 U12695 ( .A(n13362), .ZN(n10101) );
  NAND2_X1 U12696 ( .A1(n10101), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10075) );
  NAND2_X1 U12697 ( .A1(n13366), .A2(n10075), .ZN(n13376) );
  MUX2_X1 U12698 ( .A(n10076), .B(P2_REG1_REG_2__SCAN_IN), .S(n13372), .Z(
        n13377) );
  NAND2_X1 U12699 ( .A1(n13376), .A2(n13377), .ZN(n13391) );
  NAND2_X1 U12700 ( .A1(n10104), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13390) );
  NAND2_X1 U12701 ( .A1(n13391), .A2(n13390), .ZN(n10079) );
  MUX2_X1 U12702 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10077), .S(n13389), .Z(
        n10078) );
  NAND2_X1 U12703 ( .A1(n10079), .A2(n10078), .ZN(n13394) );
  NAND2_X1 U12704 ( .A1(n13389), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U12705 ( .A1(n13394), .A2(n10080), .ZN(n15342) );
  MUX2_X1 U12706 ( .A(n10081), .B(P2_REG1_REG_4__SCAN_IN), .S(n15336), .Z(
        n15343) );
  NAND2_X1 U12707 ( .A1(n15342), .A2(n15343), .ZN(n15341) );
  INV_X1 U12708 ( .A(n15336), .ZN(n10108) );
  NAND2_X1 U12709 ( .A1(n10108), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U12710 ( .A1(n15341), .A2(n10082), .ZN(n10263) );
  MUX2_X1 U12711 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10083), .S(n10268), .Z(
        n10264) );
  NAND2_X1 U12712 ( .A1(n10263), .A2(n10264), .ZN(n10262) );
  NAND2_X1 U12713 ( .A1(n10268), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U12714 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10085), .S(n10111), .Z(
        n15361) );
  XNOR2_X1 U12715 ( .A(n10114), .B(n15552), .ZN(n15374) );
  NAND2_X1 U12716 ( .A1(n10114), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U12717 ( .A1(n10087), .A2(n10086), .ZN(n10362) );
  XNOR2_X1 U12718 ( .A(n10359), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n10361) );
  XNOR2_X1 U12719 ( .A(n10362), .B(n10361), .ZN(n10122) );
  NAND2_X1 U12720 ( .A1(n10088), .A2(n11491), .ZN(n10090) );
  NAND2_X1 U12721 ( .A1(n10090), .A2(n10089), .ZN(n10091) );
  OAI21_X1 U12722 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10099) );
  NAND2_X1 U12723 ( .A1(n10094), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13911) );
  NOR2_X1 U12724 ( .A1(n13911), .A2(n13438), .ZN(n10095) );
  NAND2_X1 U12725 ( .A1(n10099), .A2(n10095), .ZN(n13430) );
  OR2_X1 U12726 ( .A1(n10099), .A2(P2_U3088), .ZN(n15399) );
  INV_X1 U12727 ( .A(n15399), .ZN(n15334) );
  NOR2_X1 U12728 ( .A1(n10094), .A2(P2_U3088), .ZN(n10096) );
  NAND2_X1 U12729 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11401) );
  OAI21_X1 U12730 ( .B1(n15395), .B2(n10359), .A(n11401), .ZN(n10097) );
  AOI21_X1 U12731 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(n15334), .A(n10097), .ZN(
        n10121) );
  NOR2_X1 U12732 ( .A1(n13328), .A2(P2_U3088), .ZN(n12065) );
  AND2_X1 U12733 ( .A1(n12065), .A2(n10094), .ZN(n10098) );
  INV_X1 U12734 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10100) );
  AND2_X1 U12735 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n13361) );
  NAND2_X1 U12736 ( .A1(n10101), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U12737 ( .A1(n13359), .A2(n10102), .ZN(n13374) );
  INV_X1 U12738 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n15528) );
  MUX2_X1 U12739 ( .A(n15528), .B(P2_REG2_REG_2__SCAN_IN), .S(n13372), .Z(
        n10103) );
  NAND2_X1 U12740 ( .A1(n10104), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13384) );
  INV_X1 U12741 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11077) );
  MUX2_X1 U12742 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11077), .S(n13389), .Z(
        n10105) );
  NAND2_X1 U12743 ( .A1(n10106), .A2(n10105), .ZN(n13388) );
  NAND2_X1 U12744 ( .A1(n13389), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U12745 ( .A1(n13388), .A2(n10107), .ZN(n15345) );
  MUX2_X1 U12746 ( .A(n11004), .B(P2_REG2_REG_4__SCAN_IN), .S(n15336), .Z(
        n15346) );
  NAND2_X1 U12747 ( .A1(n10108), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U12748 ( .A1(n15344), .A2(n10109), .ZN(n10260) );
  MUX2_X1 U12749 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11063), .S(n10268), .Z(
        n10261) );
  NAND2_X1 U12750 ( .A1(n10260), .A2(n10261), .ZN(n10259) );
  NAND2_X1 U12751 ( .A1(n10268), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U12752 ( .A1(n10259), .A2(n10110), .ZN(n15357) );
  MUX2_X1 U12753 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11248), .S(n10111), .Z(
        n15358) );
  NAND2_X1 U12754 ( .A1(n15357), .A2(n15358), .ZN(n15356) );
  NAND2_X1 U12755 ( .A1(n10111), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10112) );
  NAND2_X1 U12756 ( .A1(n15356), .A2(n10112), .ZN(n15371) );
  MUX2_X1 U12757 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10113), .S(n10114), .Z(
        n15372) );
  NAND2_X1 U12758 ( .A1(n10114), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U12759 ( .A1(n15370), .A2(n10118), .ZN(n10116) );
  INV_X1 U12760 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11589) );
  MUX2_X1 U12761 ( .A(n11589), .B(P2_REG2_REG_8__SCAN_IN), .S(n10359), .Z(
        n10115) );
  NAND2_X1 U12762 ( .A1(n10116), .A2(n10115), .ZN(n10369) );
  MUX2_X1 U12763 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11589), .S(n10359), .Z(
        n10117) );
  NAND3_X1 U12764 ( .A1(n15370), .A2(n10118), .A3(n10117), .ZN(n10119) );
  NAND3_X1 U12765 ( .A1(n15405), .A2(n10369), .A3(n10119), .ZN(n10120) );
  OAI211_X1 U12766 ( .C1(n10122), .C2(n13430), .A(n10121), .B(n10120), .ZN(
        P2_U3222) );
  INV_X1 U12767 ( .A(P3_U3897), .ZN(n12453) );
  INV_X1 U12768 ( .A(n10252), .ZN(n10123) );
  NAND2_X1 U12769 ( .A1(n10123), .A2(n11517), .ZN(n10137) );
  INV_X1 U12770 ( .A(n10124), .ZN(n10125) );
  OR2_X1 U12771 ( .A1(n10126), .A2(n10125), .ZN(n10127) );
  NAND2_X1 U12772 ( .A1(n10127), .A2(n7918), .ZN(n10136) );
  INV_X1 U12773 ( .A(n10136), .ZN(n10128) );
  INV_X1 U12774 ( .A(n10132), .ZN(n10129) );
  MUX2_X1 U12775 ( .A(n12453), .B(n10129), .S(n12125), .Z(n12597) );
  INV_X1 U12776 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10202) );
  INV_X1 U12777 ( .A(n10130), .ZN(n10131) );
  NAND2_X1 U12778 ( .A1(P3_U3897), .A2(n12125), .ZN(n12605) );
  NAND3_X1 U12779 ( .A1(n12566), .A2(n12024), .A3(n12605), .ZN(n10135) );
  MUX2_X1 U12780 ( .A(n7317), .B(n10536), .S(n12937), .Z(n10133) );
  NAND2_X1 U12781 ( .A1(n10133), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10322) );
  OAI21_X1 U12782 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n10133), .A(n10322), .ZN(
        n10134) );
  NAND2_X1 U12783 ( .A1(n10135), .A2(n10134), .ZN(n10139) );
  AOI22_X1 U12784 ( .A1(n15455), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10138) );
  OAI211_X1 U12785 ( .C1(n12597), .C2(n10202), .A(n10139), .B(n10138), .ZN(
        P3_U3182) );
  AOI22_X1 U12786 ( .A1(n10559), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10140), .ZN(n10141) );
  OAI21_X1 U12787 ( .B1(n10256), .B2(n15147), .A(n10141), .ZN(P1_U3345) );
  INV_X1 U12788 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10143) );
  OAI22_X1 U12789 ( .A1(n11894), .A2(n10143), .B1(n10142), .B2(n13430), .ZN(
        n10146) );
  NAND2_X1 U12790 ( .A1(n15405), .A2(n10143), .ZN(n10144) );
  OAI211_X1 U12791 ( .C1(n13430), .C2(P2_REG1_REG_0__SCAN_IN), .A(n10144), .B(
        n15395), .ZN(n10145) );
  MUX2_X1 U12792 ( .A(n10146), .B(n10145), .S(P2_IR_REG_0__SCAN_IN), .Z(n10149) );
  INV_X1 U12793 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10147) );
  OAI22_X1 U12794 ( .A1(n15399), .A2(n10147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11048), .ZN(n10148) );
  OR2_X1 U12795 ( .A1(n10149), .A2(n10148), .ZN(P2_U3214) );
  INV_X1 U12796 ( .A(n10150), .ZN(n10214) );
  INV_X1 U12797 ( .A(n10769), .ZN(n11109) );
  OAI222_X1 U12798 ( .A1(n15147), .A2(n10214), .B1(n15144), .B2(n10151), .C1(
        n11109), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U12799 ( .A1(n15289), .A2(n15277), .ZN(n10153) );
  NAND2_X1 U12800 ( .A1(n14581), .A2(n11333), .ZN(n14313) );
  NAND2_X1 U12801 ( .A1(n10152), .A2(n14313), .ZN(n14525) );
  AOI222_X1 U12802 ( .A1(n10153), .A2(n14525), .B1(n10304), .B2(n9293), .C1(
        n9228), .C2(n15090), .ZN(n15272) );
  NAND2_X1 U12803 ( .A1(n15331), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10154) );
  OAI21_X1 U12804 ( .B1(n15272), .B2(n15331), .A(n10154), .ZN(P1_U3528) );
  INV_X1 U12805 ( .A(n15221), .ZN(n14654) );
  NAND2_X1 U12806 ( .A1(n14654), .A2(n10220), .ZN(n10157) );
  NAND2_X1 U12807 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11453) );
  OAI211_X1 U12808 ( .C1(n15226), .C2(n10480), .A(n10157), .B(n11453), .ZN(
        n10183) );
  INV_X1 U12809 ( .A(n10176), .ZN(n10188) );
  INV_X1 U12810 ( .A(n15220), .ZN(n10165) );
  INV_X1 U12811 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10158) );
  AND2_X1 U12812 ( .A1(n7069), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14590) );
  INV_X1 U12813 ( .A(n14586), .ZN(n14585) );
  NAND2_X1 U12814 ( .A1(n14585), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U12815 ( .A1(n14588), .A2(n10159), .ZN(n14607) );
  INV_X1 U12816 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10160) );
  MUX2_X1 U12817 ( .A(n10160), .B(P1_REG1_REG_2__SCAN_IN), .S(n14605), .Z(
        n10161) );
  INV_X1 U12818 ( .A(n14605), .ZN(n14604) );
  NAND2_X1 U12819 ( .A1(n14604), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14618) );
  NAND2_X1 U12820 ( .A1(n14619), .A2(n14618), .ZN(n10164) );
  INV_X1 U12821 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10162) );
  MUX2_X1 U12822 ( .A(n10162), .B(P1_REG1_REG_3__SCAN_IN), .S(n14621), .Z(
        n10163) );
  NAND2_X1 U12823 ( .A1(n10164), .A2(n10163), .ZN(n15207) );
  OR2_X1 U12824 ( .A1(n14621), .A2(n10162), .ZN(n15206) );
  INV_X1 U12825 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15325) );
  MUX2_X1 U12826 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n15325), .S(n15220), .Z(
        n15205) );
  AOI21_X1 U12827 ( .B1(n15207), .B2(n15206), .A(n15205), .ZN(n15204) );
  MUX2_X1 U12828 ( .A(n8798), .B(P1_REG1_REG_5__SCAN_IN), .S(n10176), .Z(
        n10186) );
  NAND2_X1 U12829 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  OAI21_X1 U12830 ( .B1(n10188), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10185), .ZN(
        n10168) );
  INV_X1 U12831 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15328) );
  MUX2_X1 U12832 ( .A(n15328), .B(P1_REG1_REG_6__SCAN_IN), .S(n10220), .Z(
        n10167) );
  INV_X1 U12833 ( .A(n10346), .ZN(n10166) );
  AOI211_X1 U12834 ( .C1(n10168), .C2(n10167), .A(n10166), .B(n14668), .ZN(
        n10182) );
  NOR2_X1 U12835 ( .A1(n9286), .A2(n6410), .ZN(n10169) );
  INV_X1 U12836 ( .A(n15217), .ZN(n14657) );
  MUX2_X1 U12837 ( .A(n11207), .B(P1_REG2_REG_1__SCAN_IN), .S(n14586), .Z(
        n14592) );
  AND2_X1 U12838 ( .A1(n7069), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U12839 ( .A1(n14592), .A2(n10171), .ZN(n14591) );
  NAND2_X1 U12840 ( .A1(n14585), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U12841 ( .A1(n14591), .A2(n10172), .ZN(n14609) );
  MUX2_X1 U12842 ( .A(n10173), .B(P1_REG2_REG_2__SCAN_IN), .S(n14605), .Z(
        n14610) );
  NAND2_X1 U12843 ( .A1(n14609), .A2(n14610), .ZN(n14624) );
  NAND2_X1 U12844 ( .A1(n14604), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14623) );
  NAND2_X1 U12845 ( .A1(n14624), .A2(n14623), .ZN(n10175) );
  MUX2_X1 U12846 ( .A(n11510), .B(P1_REG2_REG_3__SCAN_IN), .S(n14621), .Z(
        n10174) );
  NAND2_X1 U12847 ( .A1(n10175), .A2(n10174), .ZN(n15214) );
  OR2_X1 U12848 ( .A1(n14621), .A2(n11510), .ZN(n15213) );
  MUX2_X1 U12849 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11320), .S(n15220), .Z(
        n15212) );
  AOI21_X1 U12850 ( .B1(n15214), .B2(n15213), .A(n15212), .ZN(n15211) );
  NOR2_X1 U12851 ( .A1(n15220), .A2(n11320), .ZN(n10193) );
  MUX2_X1 U12852 ( .A(n10177), .B(P1_REG2_REG_5__SCAN_IN), .S(n10176), .Z(
        n10192) );
  NAND2_X1 U12853 ( .A1(n10188), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10179) );
  MUX2_X1 U12854 ( .A(n8816), .B(P1_REG2_REG_6__SCAN_IN), .S(n10220), .Z(
        n10178) );
  AOI21_X1 U12855 ( .B1(n10191), .B2(n10179), .A(n10178), .ZN(n10219) );
  AND3_X1 U12856 ( .A1(n10191), .A2(n10179), .A3(n10178), .ZN(n10180) );
  NOR3_X1 U12857 ( .A1(n14657), .A2(n10219), .A3(n10180), .ZN(n10181) );
  OR3_X1 U12858 ( .A1(n10183), .A2(n10182), .A3(n10181), .ZN(P1_U3249) );
  INV_X1 U12859 ( .A(n10184), .ZN(n10273) );
  INV_X1 U12860 ( .A(n11112), .ZN(n11162) );
  OAI222_X1 U12861 ( .A1(n15147), .A2(n10273), .B1(n15144), .B2(n15539), .C1(
        n11162), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI21_X1 U12862 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(n10198) );
  NAND2_X1 U12863 ( .A1(n14654), .A2(n10188), .ZN(n10189) );
  NAND2_X1 U12864 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14182) );
  OAI211_X1 U12865 ( .C1(n15226), .C2(n10190), .A(n10189), .B(n14182), .ZN(
        n10197) );
  INV_X1 U12866 ( .A(n10191), .ZN(n10195) );
  NOR3_X1 U12867 ( .A1(n15211), .A2(n10193), .A3(n10192), .ZN(n10194) );
  NOR3_X1 U12868 ( .A1(n14657), .A2(n10195), .A3(n10194), .ZN(n10196) );
  AOI211_X1 U12869 ( .C1(n15210), .C2(n10198), .A(n10197), .B(n10196), .ZN(
        n10199) );
  INV_X1 U12870 ( .A(n10199), .ZN(P1_U3248) );
  NAND2_X1 U12871 ( .A1(n10202), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U12872 ( .A1(n10201), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10326) );
  OAI21_X1 U12873 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(n10201), .A(n10326), .ZN(
        n10210) );
  NAND2_X1 U12874 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10202), .ZN(n10203) );
  NOR3_X1 U12875 ( .A1(n10536), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n10330) );
  AOI21_X1 U12876 ( .B1(n10204), .B2(n10203), .A(n10330), .ZN(n10205) );
  NAND2_X1 U12877 ( .A1(n10205), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10332) );
  OAI21_X1 U12878 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10205), .A(n10332), .ZN(
        n10206) );
  AND2_X1 U12879 ( .A1(n12607), .A2(n10206), .ZN(n10209) );
  INV_X1 U12880 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10207) );
  OAI22_X1 U12881 ( .A1(n12581), .A2(n10207), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10527), .ZN(n10208) );
  AOI211_X1 U12882 ( .C1(n12590), .C2(n10210), .A(n10209), .B(n10208), .ZN(
        n10213) );
  INV_X1 U12883 ( .A(n12605), .ZN(n12491) );
  XNOR2_X1 U12884 ( .A(n10323), .B(n10322), .ZN(n10211) );
  NAND2_X1 U12885 ( .A1(n12491), .A2(n10211), .ZN(n10212) );
  OAI211_X1 U12886 ( .C1(n12597), .C2(n10321), .A(n10213), .B(n10212), .ZN(
        P3_U3183) );
  OAI222_X1 U12887 ( .A1(P2_U3088), .A2(n11138), .B1(n13916), .B2(n15618), 
        .C1(n13913), .C2(n10214), .ZN(P2_U3315) );
  NAND2_X1 U12888 ( .A1(n10220), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10345) );
  MUX2_X1 U12889 ( .A(n8846), .B(P1_REG1_REG_7__SCAN_IN), .S(n10221), .Z(
        n10344) );
  AOI21_X1 U12890 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(n10343) );
  INV_X1 U12891 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15332) );
  MUX2_X1 U12892 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n15332), .S(n10312), .Z(
        n10215) );
  NAND2_X1 U12893 ( .A1(n10216), .A2(n10215), .ZN(n10311) );
  OAI21_X1 U12894 ( .B1(n10216), .B2(n10215), .A(n10311), .ZN(n10230) );
  AND2_X1 U12895 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11828) );
  AOI21_X1 U12896 ( .B1(n14653), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11828), .ZN(
        n10217) );
  OAI21_X1 U12897 ( .B1(n10218), .B2(n15221), .A(n10217), .ZN(n10229) );
  AOI21_X1 U12898 ( .B1(n10220), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10219), .ZN(
        n10350) );
  MUX2_X1 U12899 ( .A(n10222), .B(P1_REG2_REG_7__SCAN_IN), .S(n10221), .Z(
        n10351) );
  NOR2_X1 U12900 ( .A1(n10357), .A2(n10222), .ZN(n10225) );
  MUX2_X1 U12901 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10223), .S(n10312), .Z(
        n10224) );
  INV_X1 U12902 ( .A(n10309), .ZN(n10227) );
  NOR3_X1 U12903 ( .A1(n10349), .A2(n10225), .A3(n10224), .ZN(n10226) );
  NOR3_X1 U12904 ( .A1(n10227), .A2(n10226), .A3(n14657), .ZN(n10228) );
  AOI211_X1 U12905 ( .C1(n15210), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10231) );
  INV_X1 U12906 ( .A(n10231), .ZN(P1_U3251) );
  NAND2_X1 U12907 ( .A1(n10247), .A2(n10241), .ZN(n10236) );
  INV_X1 U12908 ( .A(n10244), .ZN(n10232) );
  NAND2_X1 U12909 ( .A1(n10250), .A2(n10232), .ZN(n10234) );
  NAND4_X1 U12910 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10240) );
  INV_X1 U12911 ( .A(n10237), .ZN(n10238) );
  AND2_X1 U12912 ( .A1(n10250), .A2(n10238), .ZN(n10239) );
  AOI21_X1 U12913 ( .B1(n10240), .B2(P3_STATE_REG_SCAN_IN), .A(n10239), .ZN(
        n10609) );
  AND2_X1 U12914 ( .A1(n10609), .A2(n12922), .ZN(n10590) );
  INV_X1 U12915 ( .A(n12829), .ZN(n15475) );
  NAND2_X1 U12916 ( .A1(n10241), .A2(n15475), .ZN(n10242) );
  OR2_X1 U12917 ( .A1(n10247), .A2(n10242), .ZN(n10243) );
  OAI21_X1 U12918 ( .B1(n10250), .B2(n10244), .A(n10243), .ZN(n10245) );
  INV_X1 U12919 ( .A(n10248), .ZN(n10246) );
  OR2_X1 U12920 ( .A1(n10247), .A2(n10246), .ZN(n10249) );
  INV_X1 U12921 ( .A(n12461), .ZN(n15466) );
  INV_X1 U12922 ( .A(n10250), .ZN(n10526) );
  INV_X1 U12923 ( .A(n10515), .ZN(n10251) );
  NAND2_X1 U12924 ( .A1(n10252), .A2(n10251), .ZN(n10524) );
  NOR2_X1 U12925 ( .A1(n10524), .A2(n15469), .ZN(n10253) );
  OAI22_X1 U12926 ( .A1(n12448), .A2(n10946), .B1(n15466), .B2(n12429), .ZN(
        n10254) );
  AOI21_X1 U12927 ( .B1(n12439), .B2(n10533), .A(n10254), .ZN(n10255) );
  OAI21_X1 U12928 ( .B1(n10590), .B2(n10632), .A(n10255), .ZN(P3_U3172) );
  INV_X1 U12929 ( .A(n10591), .ZN(n10258) );
  INV_X1 U12930 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10257) );
  OAI222_X1 U12931 ( .A1(P2_U3088), .A2(n10258), .B1(n13916), .B2(n10257), 
        .C1(n13913), .C2(n10256), .ZN(P2_U3317) );
  OAI211_X1 U12932 ( .C1(n10261), .C2(n10260), .A(n15405), .B(n10259), .ZN(
        n10266) );
  OAI211_X1 U12933 ( .C1(n10264), .C2(n10263), .A(n15403), .B(n10262), .ZN(
        n10265) );
  NAND2_X1 U12934 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  AND2_X1 U12935 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10927) );
  AOI211_X1 U12936 ( .C1(n6638), .C2(n10268), .A(n10267), .B(n10927), .ZN(
        n10269) );
  OAI21_X1 U12937 ( .B1(n10270), .B2(n15399), .A(n10269), .ZN(P2_U3219) );
  OAI222_X1 U12938 ( .A1(n12505), .A2(P3_U3151), .B1(n12948), .B2(n10272), 
        .C1(n10271), .C2(n12941), .ZN(P3_U3281) );
  INV_X1 U12939 ( .A(n11608), .ZN(n11146) );
  OAI222_X1 U12940 ( .A1(P2_U3088), .A2(n11146), .B1(n13916), .B2(n10274), 
        .C1(n13913), .C2(n10273), .ZN(P2_U3314) );
  INV_X1 U12941 ( .A(n10275), .ZN(n10281) );
  AND2_X1 U12942 ( .A1(n10276), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10277) );
  OR2_X1 U12943 ( .A1(n10278), .A2(n10277), .ZN(n10280) );
  NAND2_X1 U12944 ( .A1(n10281), .A2(n11199), .ZN(n14298) );
  AND2_X2 U12945 ( .A1(n14479), .A2(n10288), .ZN(n10286) );
  OAI22_X1 U12946 ( .A1(n11333), .A2(n14020), .B1(n10288), .B2(n7040), .ZN(
        n10285) );
  AOI21_X1 U12947 ( .B1(n14581), .B2(n14108), .A(n10285), .ZN(n10292) );
  NAND2_X1 U12948 ( .A1(n14581), .A2(n10286), .ZN(n10291) );
  OAI22_X1 U12949 ( .A1(n11333), .A2(n14011), .B1(n10288), .B2(n10287), .ZN(
        n10289) );
  INV_X1 U12950 ( .A(n10289), .ZN(n10290) );
  NAND2_X1 U12951 ( .A1(n10291), .A2(n10290), .ZN(n10650) );
  NAND2_X1 U12952 ( .A1(n10292), .A2(n10650), .ZN(n10653) );
  OAI21_X1 U12953 ( .B1(n10292), .B2(n10650), .A(n10653), .ZN(n14596) );
  NAND2_X1 U12954 ( .A1(n10293), .A2(n11199), .ZN(n10299) );
  NOR2_X1 U12955 ( .A1(n10297), .A2(n10299), .ZN(n10296) );
  NOR2_X1 U12956 ( .A1(n15315), .A2(n10294), .ZN(n10295) );
  NAND2_X1 U12957 ( .A1(n14596), .A2(n14281), .ZN(n10306) );
  INV_X1 U12958 ( .A(n10296), .ZN(n10298) );
  NAND2_X1 U12959 ( .A1(n10300), .A2(n10299), .ZN(n10303) );
  INV_X1 U12960 ( .A(n10301), .ZN(n10302) );
  NAND2_X1 U12961 ( .A1(n10303), .A2(n10302), .ZN(n10912) );
  OR2_X1 U12962 ( .A1(n10912), .A2(P1_U3086), .ZN(n14132) );
  AOI22_X1 U12963 ( .A1(n10304), .A2(n14300), .B1(n14132), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10305) );
  OAI211_X1 U12964 ( .C1(n7111), .C2(n14272), .A(n10306), .B(n10305), .ZN(
        P1_U3232) );
  NAND2_X1 U12965 ( .A1(n10312), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10308) );
  MUX2_X1 U12966 ( .A(n10463), .B(P1_REG2_REG_9__SCAN_IN), .S(n10317), .Z(
        n10307) );
  NAND3_X1 U12967 ( .A1(n10309), .A2(n10308), .A3(n10307), .ZN(n10310) );
  NAND2_X1 U12968 ( .A1(n10310), .A2(n15217), .ZN(n10320) );
  XNOR2_X1 U12969 ( .A(n10317), .B(n10458), .ZN(n10314) );
  OAI21_X1 U12970 ( .B1(n10312), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10311), .ZN(
        n10313) );
  OAI21_X1 U12971 ( .B1(n10314), .B2(n10313), .A(n10462), .ZN(n10315) );
  NAND2_X1 U12972 ( .A1(n10315), .A2(n15210), .ZN(n10319) );
  AND2_X1 U12973 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14218) );
  INV_X1 U12974 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10932) );
  NOR2_X1 U12975 ( .A1(n15226), .A2(n10932), .ZN(n10316) );
  AOI211_X1 U12976 ( .C1(n14654), .C2(n10317), .A(n14218), .B(n10316), .ZN(
        n10318) );
  OAI211_X1 U12977 ( .C1(n10467), .C2(n10320), .A(n10319), .B(n10318), .ZN(
        P1_U3252) );
  MUX2_X1 U12978 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12937), .Z(n10380) );
  XNOR2_X1 U12979 ( .A(n10380), .B(n6399), .ZN(n10382) );
  XOR2_X1 U12980 ( .A(n10382), .B(n10383), .Z(n10342) );
  XNOR2_X1 U12981 ( .A(n6399), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10328) );
  INV_X1 U12982 ( .A(n10324), .ZN(n10325) );
  NAND2_X1 U12983 ( .A1(n10326), .A2(n10325), .ZN(n10327) );
  NAND2_X1 U12984 ( .A1(n10327), .A2(n10328), .ZN(n10389) );
  OAI21_X1 U12985 ( .B1(n10328), .B2(n10327), .A(n10389), .ZN(n10339) );
  MUX2_X1 U12986 ( .A(n10329), .B(P3_REG1_REG_2__SCAN_IN), .S(n10402), .Z(
        n10334) );
  INV_X1 U12987 ( .A(n10330), .ZN(n10331) );
  NAND2_X1 U12988 ( .A1(n10332), .A2(n10331), .ZN(n10333) );
  NAND2_X1 U12989 ( .A1(n10333), .A2(n10334), .ZN(n10404) );
  OAI21_X1 U12990 ( .B1(n10334), .B2(n10333), .A(n10404), .ZN(n10335) );
  AND2_X1 U12991 ( .A1(n12607), .A2(n10335), .ZN(n10338) );
  OAI22_X1 U12992 ( .A1(n12581), .A2(n10336), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15459), .ZN(n10337) );
  AOI211_X1 U12993 ( .C1(n12590), .C2(n10339), .A(n10338), .B(n10337), .ZN(
        n10341) );
  NAND2_X1 U12994 ( .A1(n12578), .A2(n6399), .ZN(n10340) );
  OAI211_X1 U12995 ( .C1(n10342), .C2(n12605), .A(n10341), .B(n10340), .ZN(
        P3_U3184) );
  INV_X1 U12996 ( .A(n10343), .ZN(n10348) );
  NAND3_X1 U12997 ( .A1(n10346), .A2(n10345), .A3(n10344), .ZN(n10347) );
  NAND3_X1 U12998 ( .A1(n10348), .A2(n15210), .A3(n10347), .ZN(n10356) );
  NAND2_X1 U12999 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11936) );
  AOI211_X1 U13000 ( .C1(n10351), .C2(n10350), .A(n10349), .B(n14657), .ZN(
        n10352) );
  INV_X1 U13001 ( .A(n10352), .ZN(n10353) );
  NAND2_X1 U13002 ( .A1(n11936), .A2(n10353), .ZN(n10354) );
  AOI21_X1 U13003 ( .B1(n14653), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10354), .ZN(
        n10355) );
  OAI211_X1 U13004 ( .C1(n15221), .C2(n10357), .A(n10356), .B(n10355), .ZN(
        P1_U3250) );
  INV_X1 U13005 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10379) );
  NOR2_X1 U13006 ( .A1(n10359), .A2(n10358), .ZN(n10360) );
  XNOR2_X1 U13007 ( .A(n10370), .B(n10363), .ZN(n15379) );
  NOR2_X1 U13008 ( .A1(n10370), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10365) );
  XNOR2_X1 U13009 ( .A(n10591), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n10364) );
  OAI21_X1 U13010 ( .B1(n15381), .B2(n10365), .A(n10364), .ZN(n10366) );
  NAND3_X1 U13011 ( .A1(n6641), .A2(n15403), .A3(n10366), .ZN(n10378) );
  NAND2_X1 U13012 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11743)
         );
  MUX2_X1 U13013 ( .A(n11699), .B(P2_REG2_REG_10__SCAN_IN), .S(n10591), .Z(
        n10372) );
  NAND2_X1 U13014 ( .A1(n10367), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U13015 ( .A1(n10369), .A2(n10368), .ZN(n15384) );
  INV_X1 U13016 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11632) );
  MUX2_X1 U13017 ( .A(n11632), .B(P2_REG2_REG_9__SCAN_IN), .S(n10370), .Z(
        n15383) );
  OR2_X1 U13018 ( .A1(n10370), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10371) );
  AOI21_X1 U13019 ( .B1(n10372), .B2(n10373), .A(n11894), .ZN(n10374) );
  NAND2_X1 U13020 ( .A1(n10374), .A2(n10593), .ZN(n10375) );
  NAND2_X1 U13021 ( .A1(n11743), .A2(n10375), .ZN(n10376) );
  AOI21_X1 U13022 ( .B1(n6638), .B2(n10591), .A(n10376), .ZN(n10377) );
  OAI211_X1 U13023 ( .C1(n15399), .C2(n10379), .A(n10378), .B(n10377), .ZN(
        P2_U3224) );
  MUX2_X1 U13024 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12937), .Z(n10638) );
  XNOR2_X1 U13025 ( .A(n10638), .B(n10640), .ZN(n10641) );
  INV_X1 U13026 ( .A(n10380), .ZN(n10381) );
  AOI22_X1 U13027 ( .A1(n10383), .A2(n10382), .B1(n6399), .B2(n10381), .ZN(
        n10446) );
  MUX2_X1 U13028 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12937), .Z(n10384) );
  XOR2_X1 U13029 ( .A(n10455), .B(n10384), .Z(n10447) );
  INV_X1 U13030 ( .A(n10455), .ZN(n10405) );
  OAI22_X1 U13031 ( .A1(n10446), .A2(n10447), .B1(n10384), .B2(n10405), .ZN(
        n10427) );
  MUX2_X1 U13032 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12937), .Z(n10385) );
  XNOR2_X1 U13033 ( .A(n10385), .B(n10443), .ZN(n10428) );
  INV_X1 U13034 ( .A(n10385), .ZN(n10386) );
  AOI22_X1 U13035 ( .A1(n10427), .A2(n10428), .B1(n10443), .B2(n10386), .ZN(
        n10548) );
  MUX2_X1 U13036 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12937), .Z(n10387) );
  XOR2_X1 U13037 ( .A(n10412), .B(n10387), .Z(n10549) );
  INV_X1 U13038 ( .A(n10412), .ZN(n10547) );
  XOR2_X1 U13039 ( .A(n10641), .B(n10642), .Z(n10421) );
  OR2_X1 U13040 ( .A1(n6399), .A2(n15474), .ZN(n10388) );
  NAND2_X1 U13041 ( .A1(n10389), .A2(n10388), .ZN(n10390) );
  XNOR2_X1 U13042 ( .A(n10410), .B(n7959), .ZN(n10429) );
  NAND2_X1 U13043 ( .A1(n10392), .A2(n10429), .ZN(n10433) );
  NAND2_X1 U13044 ( .A1(n10410), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U13045 ( .A1(n10433), .A2(n10393), .ZN(n10394) );
  OAI21_X1 U13046 ( .B1(n10394), .B2(n10547), .A(n10395), .ZN(n10541) );
  INV_X1 U13047 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11090) );
  INV_X1 U13048 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11096) );
  XNOR2_X1 U13049 ( .A(n10640), .B(n11096), .ZN(n10396) );
  NAND3_X1 U13050 ( .A1(n10543), .A2(n10396), .A3(n10395), .ZN(n10397) );
  NAND2_X1 U13051 ( .A1(n6587), .A2(n10397), .ZN(n10400) );
  AND2_X1 U13052 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11023) );
  AOI21_X1 U13053 ( .B1(n15455), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11023), .ZN(
        n10398) );
  OAI21_X1 U13054 ( .B1(n12597), .B2(n10634), .A(n10398), .ZN(n10399) );
  AOI21_X1 U13055 ( .B1(n10400), .B2(n12590), .A(n10399), .ZN(n10420) );
  MUX2_X1 U13056 ( .A(n10401), .B(P3_REG1_REG_6__SCAN_IN), .S(n10640), .Z(
        n10417) );
  OR2_X1 U13057 ( .A1(n6399), .A2(n10329), .ZN(n10403) );
  NAND2_X1 U13058 ( .A1(n10404), .A2(n10403), .ZN(n10406) );
  NAND2_X1 U13059 ( .A1(n10448), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U13060 ( .A1(n10406), .A2(n10405), .ZN(n10407) );
  NAND2_X1 U13061 ( .A1(n10408), .A2(n10407), .ZN(n10436) );
  MUX2_X1 U13062 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10409), .S(n10410), .Z(
        n10437) );
  NAND2_X1 U13063 ( .A1(n10436), .A2(n10437), .ZN(n10435) );
  NAND2_X1 U13064 ( .A1(n10410), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U13065 ( .A1(n10435), .A2(n10411), .ZN(n10413) );
  XNOR2_X1 U13066 ( .A(n10413), .B(n10412), .ZN(n10540) );
  NAND2_X1 U13067 ( .A1(n10540), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U13068 ( .A1(n10413), .A2(n10547), .ZN(n10414) );
  NAND2_X1 U13069 ( .A1(n10415), .A2(n10414), .ZN(n10416) );
  OAI21_X1 U13070 ( .B1(n10417), .B2(n10416), .A(n10633), .ZN(n10418) );
  NAND2_X1 U13071 ( .A1(n10418), .A2(n12607), .ZN(n10419) );
  OAI211_X1 U13072 ( .C1(n10421), .C2(n12605), .A(n10420), .B(n10419), .ZN(
        P3_U3188) );
  INV_X1 U13073 ( .A(n10768), .ZN(n10424) );
  INV_X1 U13074 ( .A(n10422), .ZN(n10426) );
  OAI222_X1 U13075 ( .A1(n10424), .A2(P1_U3086), .B1(n15147), .B2(n10426), 
        .C1(n10423), .C2(n15144), .ZN(P1_U3344) );
  INV_X1 U13076 ( .A(n10724), .ZN(n10718) );
  OAI222_X1 U13077 ( .A1(n10718), .A2(P2_U3088), .B1(n13913), .B2(n10426), 
        .C1(n10425), .C2(n13916), .ZN(P2_U3316) );
  XOR2_X1 U13078 ( .A(n10428), .B(n10427), .Z(n10445) );
  INV_X1 U13079 ( .A(n10429), .ZN(n10431) );
  NAND3_X1 U13080 ( .A1(n10449), .A2(n10431), .A3(n10430), .ZN(n10432) );
  AND2_X1 U13081 ( .A1(n10433), .A2(n10432), .ZN(n10441) );
  NAND2_X1 U13082 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10698) );
  INV_X1 U13083 ( .A(n10698), .ZN(n10434) );
  AOI21_X1 U13084 ( .B1(n15455), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10434), .ZN(
        n10440) );
  OAI21_X1 U13085 ( .B1(n10437), .B2(n10436), .A(n10435), .ZN(n10438) );
  NAND2_X1 U13086 ( .A1(n12607), .A2(n10438), .ZN(n10439) );
  OAI211_X1 U13087 ( .C1(n12566), .C2(n10441), .A(n10440), .B(n10439), .ZN(
        n10442) );
  AOI21_X1 U13088 ( .B1(n10443), .B2(n12578), .A(n10442), .ZN(n10444) );
  OAI21_X1 U13089 ( .B1(n10445), .B2(n12605), .A(n10444), .ZN(P3_U3186) );
  XOR2_X1 U13090 ( .A(n10447), .B(n10446), .Z(n10457) );
  XOR2_X1 U13091 ( .A(P3_REG1_REG_3__SCAN_IN), .B(n10448), .Z(n10453) );
  AOI22_X1 U13092 ( .A1(n15455), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10452) );
  OAI21_X1 U13093 ( .B1(n6594), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10449), .ZN(
        n10450) );
  NAND2_X1 U13094 ( .A1(n12590), .A2(n10450), .ZN(n10451) );
  OAI211_X1 U13095 ( .C1(n12024), .C2(n10453), .A(n10452), .B(n10451), .ZN(
        n10454) );
  AOI21_X1 U13096 ( .B1(n10455), .B2(n12578), .A(n10454), .ZN(n10456) );
  OAI21_X1 U13097 ( .B1(n10457), .B2(n12605), .A(n10456), .ZN(P3_U3185) );
  NAND2_X1 U13098 ( .A1(n10464), .A2(n10458), .ZN(n10460) );
  INV_X1 U13099 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10459) );
  XNOR2_X1 U13100 ( .A(n10559), .B(n10459), .ZN(n10461) );
  AOI21_X1 U13101 ( .B1(n10462), .B2(n10460), .A(n10461), .ZN(n10474) );
  NAND2_X1 U13102 ( .A1(n10562), .A2(n15210), .ZN(n10473) );
  INV_X1 U13103 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U13104 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12180)
         );
  OAI21_X1 U13105 ( .B1(n15226), .B2(n10933), .A(n12180), .ZN(n10471) );
  NOR2_X1 U13106 ( .A1(n10464), .A2(n10463), .ZN(n10466) );
  MUX2_X1 U13107 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11763), .S(n10559), .Z(
        n10465) );
  INV_X1 U13108 ( .A(n10557), .ZN(n10469) );
  NOR3_X1 U13109 ( .A1(n10467), .A2(n10466), .A3(n10465), .ZN(n10468) );
  NOR3_X1 U13110 ( .A1(n10469), .A2(n10468), .A3(n14657), .ZN(n10470) );
  AOI211_X1 U13111 ( .C1(n14654), .C2(n10559), .A(n10471), .B(n10470), .ZN(
        n10472) );
  OAI21_X1 U13112 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(P1_U3253) );
  INV_X1 U13113 ( .A(n10475), .ZN(n10476) );
  OAI222_X1 U13114 ( .A1(n12941), .A2(n10477), .B1(n12948), .B2(n10476), .C1(
        P3_U3151), .C2(n12531), .ZN(P3_U3280) );
  INV_X1 U13115 ( .A(n10489), .ZN(n10481) );
  XNOR2_X1 U13116 ( .A(n10481), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15154) );
  INV_X1 U13117 ( .A(n10482), .ZN(n10483) );
  NAND2_X1 U13118 ( .A1(n10483), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U13119 ( .A1(n10485), .A2(n10484), .ZN(n10486) );
  INV_X1 U13120 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15368) );
  NAND2_X1 U13121 ( .A1(n10486), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10487) );
  INV_X1 U13122 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U13123 ( .A1(n10489), .A2(n10488), .ZN(n10493) );
  INV_X1 U13124 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10490) );
  NAND2_X1 U13125 ( .A1(n10493), .A2(n10492), .ZN(n10499) );
  INV_X1 U13126 ( .A(n10499), .ZN(n10497) );
  INV_X1 U13127 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U13128 ( .A1(n10494), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10930) );
  INV_X1 U13129 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10495) );
  NAND2_X1 U13130 ( .A1(n10495), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10496) );
  AND2_X1 U13131 ( .A1(n10930), .A2(n10496), .ZN(n10498) );
  NAND2_X1 U13132 ( .A1(n10497), .A2(n6974), .ZN(n10500) );
  NAND2_X1 U13133 ( .A1(n10500), .A2(n10931), .ZN(n10501) );
  NAND2_X1 U13134 ( .A1(n10502), .A2(n10501), .ZN(n10504) );
  INV_X1 U13135 ( .A(n10503), .ZN(n10508) );
  INV_X1 U13136 ( .A(n10504), .ZN(n10505) );
  OAI21_X1 U13137 ( .B1(n10506), .B2(n10505), .A(P2_ADDR_REG_8__SCAN_IN), .ZN(
        n10507) );
  OAI21_X1 U13138 ( .B1(n15158), .B2(n10508), .A(n10507), .ZN(SUB_1596_U55) );
  AOI22_X1 U13139 ( .A1(n12555), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_16_), .B2(
        n10509), .ZN(n10510) );
  OAI21_X1 U13140 ( .B1(n10511), .B2(n12948), .A(n10510), .ZN(P3_U3279) );
  OR2_X1 U13141 ( .A1(n11564), .A2(n10513), .ZN(n10514) );
  XNOR2_X1 U13142 ( .A(n6610), .B(n10579), .ZN(n10517) );
  NAND2_X1 U13143 ( .A1(n10517), .A2(n15466), .ZN(n10572) );
  NAND3_X1 U13144 ( .A1(n11174), .A2(n12461), .A3(n10579), .ZN(n10519) );
  NAND2_X1 U13145 ( .A1(n10572), .A2(n10519), .ZN(n10523) );
  INV_X1 U13146 ( .A(n9326), .ZN(n10521) );
  NOR3_X1 U13147 ( .A1(n10521), .A2(n11174), .A3(n10520), .ZN(n10522) );
  AOI211_X1 U13148 ( .C1(n10581), .C2(n6610), .A(n15477), .B(n10523), .ZN(
        n10574) );
  AOI211_X1 U13149 ( .C1(n15477), .C2(n10523), .A(n10522), .B(n10574), .ZN(
        n10531) );
  NOR2_X1 U13150 ( .A1(n15467), .A2(n10524), .ZN(n10525) );
  NAND2_X1 U13151 ( .A1(n10526), .A2(n10525), .ZN(n12443) );
  INV_X1 U13152 ( .A(n15480), .ZN(n10608) );
  OAI22_X1 U13153 ( .A1(n7172), .A2(n12443), .B1(n12429), .B2(n10608), .ZN(
        n10529) );
  NOR2_X1 U13154 ( .A1(n10590), .A2(n10527), .ZN(n10528) );
  AOI211_X1 U13155 ( .C1(n10579), .C2(n12414), .A(n10529), .B(n10528), .ZN(
        n10530) );
  OAI21_X1 U13156 ( .B1(n10531), .B2(n12434), .A(n10530), .ZN(P3_U3162) );
  NAND3_X1 U13157 ( .A1(n10533), .A2(n15475), .A3(n10532), .ZN(n10535) );
  NAND2_X1 U13158 ( .A1(n12461), .A2(n15479), .ZN(n10534) );
  NAND2_X1 U13159 ( .A1(n10535), .A2(n10534), .ZN(n10944) );
  INV_X1 U13160 ( .A(n10944), .ZN(n10627) );
  MUX2_X1 U13161 ( .A(n10627), .B(n10536), .S(n9433), .Z(n10537) );
  OAI21_X1 U13162 ( .B1(n10946), .B2(n12821), .A(n10537), .ZN(P3_U3459) );
  INV_X1 U13163 ( .A(n11801), .ZN(n10538) );
  OAI222_X1 U13164 ( .A1(n15147), .A2(n10570), .B1(n15144), .B2(n10539), .C1(
        n10538), .C2(P1_U3086), .ZN(P1_U3341) );
  XNOR2_X1 U13165 ( .A(n10540), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n10553) );
  AND2_X1 U13166 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10852) );
  AOI21_X1 U13167 ( .B1(n15455), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10852), .ZN(
        n10546) );
  NAND2_X1 U13168 ( .A1(n10541), .A2(n11090), .ZN(n10542) );
  NAND2_X1 U13169 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  NAND2_X1 U13170 ( .A1(n12590), .A2(n10544), .ZN(n10545) );
  OAI211_X1 U13171 ( .C1(n12597), .C2(n10547), .A(n10546), .B(n10545), .ZN(
        n10552) );
  XOR2_X1 U13172 ( .A(n10549), .B(n10548), .Z(n10550) );
  NOR2_X1 U13173 ( .A1(n10550), .A2(n12605), .ZN(n10551) );
  AOI211_X1 U13174 ( .C1(n12607), .C2(n10553), .A(n10552), .B(n10551), .ZN(
        n10554) );
  INV_X1 U13175 ( .A(n10554), .ZN(P3_U3187) );
  NAND2_X1 U13176 ( .A1(n10559), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10556) );
  MUX2_X1 U13177 ( .A(n8917), .B(P1_REG2_REG_11__SCAN_IN), .S(n10768), .Z(
        n10555) );
  NAND3_X1 U13178 ( .A1(n10557), .A2(n10556), .A3(n10555), .ZN(n10558) );
  NAND2_X1 U13179 ( .A1(n10558), .A2(n15217), .ZN(n10567) );
  NOR2_X1 U13180 ( .A1(n10768), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10761) );
  AOI21_X1 U13181 ( .B1(n10768), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10761), 
        .ZN(n10560) );
  NAND2_X1 U13182 ( .A1(n10559), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10561) );
  AOI21_X1 U13183 ( .B1(n10562), .B2(n10561), .A(n10560), .ZN(n10563) );
  OAI21_X1 U13184 ( .B1(n10762), .B2(n10563), .A(n15210), .ZN(n10566) );
  INV_X1 U13185 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U13186 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n14262)
         );
  OAI21_X1 U13187 ( .B1(n15226), .B2(n11554), .A(n14262), .ZN(n10564) );
  AOI21_X1 U13188 ( .B1(n14654), .B2(n10768), .A(n10564), .ZN(n10565) );
  OAI211_X1 U13189 ( .C1(n10767), .C2(n10567), .A(n10566), .B(n10565), .ZN(
        P1_U3254) );
  INV_X1 U13190 ( .A(n10568), .ZN(n10617) );
  INV_X1 U13191 ( .A(n14636), .ZN(n11810) );
  OAI222_X1 U13192 ( .A1(n15147), .A2(n10617), .B1(n15144), .B2(n10569), .C1(
        n11810), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13193 ( .A(n11687), .ZN(n11609) );
  OAI222_X1 U13194 ( .A1(P2_U3088), .A2(n11609), .B1(n13916), .B2(n10571), 
        .C1(n13913), .C2(n10570), .ZN(P2_U3313) );
  XNOR2_X1 U13195 ( .A(n10518), .B(n10587), .ZN(n10603) );
  XNOR2_X1 U13196 ( .A(n10603), .B(n15480), .ZN(n10583) );
  INV_X1 U13197 ( .A(n10572), .ZN(n10573) );
  NOR3_X1 U13198 ( .A1(n10574), .A2(n10583), .A3(n10573), .ZN(n10585) );
  NAND3_X1 U13199 ( .A1(n11174), .A2(n15477), .A3(n10579), .ZN(n10578) );
  NAND2_X1 U13200 ( .A1(n10575), .A2(n15476), .ZN(n10576) );
  NAND2_X1 U13201 ( .A1(n10576), .A2(n12461), .ZN(n10577) );
  OAI211_X1 U13202 ( .C1(n11174), .C2(n10579), .A(n10578), .B(n10577), .ZN(
        n10580) );
  OAI21_X1 U13203 ( .B1(n11174), .B2(n10581), .A(n10580), .ZN(n10582) );
  INV_X1 U13204 ( .A(n10606), .ZN(n10584) );
  OAI21_X1 U13205 ( .B1(n10585), .B2(n10584), .A(n12439), .ZN(n10589) );
  INV_X1 U13206 ( .A(n10836), .ZN(n15468) );
  OAI22_X1 U13207 ( .A1(n15466), .A2(n12443), .B1(n12429), .B2(n15468), .ZN(
        n10586) );
  AOI21_X1 U13208 ( .B1(n10587), .B2(n12414), .A(n10586), .ZN(n10588) );
  OAI211_X1 U13209 ( .C1(n10590), .C2(n15459), .A(n10589), .B(n10588), .ZN(
        P3_U3177) );
  XNOR2_X1 U13210 ( .A(n10724), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n10719) );
  XNOR2_X1 U13211 ( .A(n6463), .B(n10719), .ZN(n10602) );
  NAND2_X1 U13212 ( .A1(n10591), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10592) );
  INV_X1 U13213 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10594) );
  MUX2_X1 U13214 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10594), .S(n10724), .Z(
        n10595) );
  OAI21_X1 U13215 ( .B1(n10596), .B2(n10595), .A(n10728), .ZN(n10600) );
  NOR2_X1 U13216 ( .A1(n15399), .A2(n6889), .ZN(n10599) );
  AND2_X1 U13217 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11991) );
  INV_X1 U13218 ( .A(n11991), .ZN(n10597) );
  OAI21_X1 U13219 ( .B1(n15395), .B2(n10718), .A(n10597), .ZN(n10598) );
  AOI211_X1 U13220 ( .C1(n10600), .C2(n15405), .A(n10599), .B(n10598), .ZN(
        n10601) );
  OAI21_X1 U13221 ( .B1(n10602), .B2(n13430), .A(n10601), .ZN(P2_U3225) );
  NAND2_X1 U13222 ( .A1(n10603), .A2(n10608), .ZN(n10604) );
  AOI21_X1 U13223 ( .B1(n10606), .B2(n10604), .A(n10605), .ZN(n10616) );
  NAND2_X1 U13224 ( .A1(n10690), .A2(n12439), .ZN(n10615) );
  INV_X1 U13225 ( .A(n12460), .ZN(n10850) );
  OAI22_X1 U13226 ( .A1(n10850), .A2(n12429), .B1(n12443), .B2(n10608), .ZN(
        n10612) );
  MUX2_X1 U13227 ( .A(P3_U3151), .B(n12441), .S(n10610), .Z(n10611) );
  AOI211_X1 U13228 ( .C1(n10613), .C2(n12414), .A(n10612), .B(n10611), .ZN(
        n10614) );
  OAI21_X1 U13229 ( .B1(n10616), .B2(n10615), .A(n10614), .ZN(P3_U3158) );
  INV_X1 U13230 ( .A(n13407), .ZN(n13398) );
  OAI222_X1 U13231 ( .A1(P2_U3088), .A2(n13398), .B1(n13916), .B2(n10618), 
        .C1(n13913), .C2(n10617), .ZN(P2_U3311) );
  INV_X1 U13232 ( .A(n10619), .ZN(n10620) );
  OAI22_X1 U13233 ( .A1(n10623), .A2(n10622), .B1(n10621), .B2(n10620), .ZN(
        n10624) );
  INV_X1 U13234 ( .A(n10624), .ZN(n10626) );
  MUX2_X1 U13235 ( .A(n7317), .B(n10627), .S(n15472), .Z(n10631) );
  INV_X1 U13236 ( .A(n15462), .ZN(n15486) );
  NAND2_X1 U13237 ( .A1(n15486), .A2(n12829), .ZN(n10628) );
  NAND2_X1 U13238 ( .A1(n12787), .A2(n10629), .ZN(n10630) );
  OAI211_X1 U13239 ( .C1(n15460), .C2(n10632), .A(n10631), .B(n10630), .ZN(
        P3_U3233) );
  INV_X1 U13240 ( .A(n10878), .ZN(n10635) );
  XOR2_X1 U13241 ( .A(P3_REG1_REG_7__SCAN_IN), .B(n10875), .Z(n10648) );
  OAI21_X1 U13242 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n10636), .A(n10886), .ZN(
        n10646) );
  NAND2_X1 U13243 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U13244 ( .A1(n15455), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n10637) );
  OAI211_X1 U13245 ( .C1(n12597), .C2(n10878), .A(n11165), .B(n10637), .ZN(
        n10645) );
  MUX2_X1 U13246 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12937), .Z(n10879) );
  XNOR2_X1 U13247 ( .A(n10879), .B(n10878), .ZN(n10880) );
  INV_X1 U13248 ( .A(n10638), .ZN(n10639) );
  XOR2_X1 U13249 ( .A(n10880), .B(n10881), .Z(n10643) );
  NOR2_X1 U13250 ( .A1(n10643), .A2(n12605), .ZN(n10644) );
  AOI211_X1 U13251 ( .C1(n12590), .C2(n10646), .A(n10645), .B(n10644), .ZN(
        n10647) );
  OAI21_X1 U13252 ( .B1(n10648), .B2(n12024), .A(n10647), .ZN(P3_U3189) );
  OR2_X1 U13253 ( .A1(n11204), .A2(n14011), .ZN(n10649) );
  XNOR2_X1 U13254 ( .A(n10654), .B(n10655), .ZN(n14128) );
  INV_X1 U13255 ( .A(n10650), .ZN(n10651) );
  NAND2_X1 U13256 ( .A1(n10651), .A2(n14111), .ZN(n10652) );
  NAND2_X1 U13257 ( .A1(n10653), .A2(n10652), .ZN(n14129) );
  NAND2_X1 U13258 ( .A1(n14128), .A2(n14129), .ZN(n10658) );
  INV_X1 U13259 ( .A(n10654), .ZN(n10656) );
  NAND2_X1 U13260 ( .A1(n10656), .A2(n10655), .ZN(n10657) );
  NAND2_X1 U13261 ( .A1(n14580), .A2(n10286), .ZN(n10660) );
  NAND2_X1 U13262 ( .A1(n10781), .A2(n10284), .ZN(n10659) );
  NAND2_X1 U13263 ( .A1(n10660), .A2(n10659), .ZN(n10661) );
  AND2_X1 U13264 ( .A1(n10781), .A2(n10286), .ZN(n10662) );
  AOI21_X1 U13265 ( .B1(n14580), .B2(n14108), .A(n10662), .ZN(n10896) );
  XNOR2_X1 U13266 ( .A(n10895), .B(n10896), .ZN(n10894) );
  INV_X1 U13267 ( .A(n14579), .ZN(n15282) );
  INV_X1 U13268 ( .A(n14227), .ZN(n14275) );
  NAND2_X1 U13269 ( .A1(n14275), .A2(n9228), .ZN(n10664) );
  AOI22_X1 U13270 ( .A1(n10781), .A2(n14300), .B1(n14132), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10663) );
  OAI211_X1 U13271 ( .C1(n15282), .C2(n14272), .A(n10664), .B(n10663), .ZN(
        n10665) );
  AOI21_X1 U13272 ( .B1(n10666), .B2(n14281), .A(n10665), .ZN(n10667) );
  INV_X1 U13273 ( .A(n10667), .ZN(P1_U3237) );
  INV_X1 U13274 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10680) );
  OAI21_X1 U13275 ( .B1(n10668), .B2(n10670), .A(n10669), .ZN(n10671) );
  INV_X1 U13276 ( .A(n10671), .ZN(n11210) );
  INV_X1 U13277 ( .A(n10668), .ZN(n14528) );
  AOI21_X1 U13278 ( .B1(n14528), .B2(n14581), .A(n15277), .ZN(n10675) );
  OR2_X1 U13279 ( .A1(n11204), .A2(n11333), .ZN(n10672) );
  NAND2_X1 U13280 ( .A1(n10672), .A2(n10780), .ZN(n10676) );
  XOR2_X1 U13281 ( .A(n9228), .B(n10676), .Z(n10673) );
  NOR2_X1 U13282 ( .A1(n10673), .A2(n15277), .ZN(n10674) );
  OAI22_X1 U13283 ( .A1(n15107), .A2(n10675), .B1(n10674), .B2(n14581), .ZN(
        n11206) );
  NOR2_X1 U13284 ( .A1(n11204), .A2(n15302), .ZN(n10677) );
  NOR2_X1 U13285 ( .A1(n10676), .A2(n10283), .ZN(n11202) );
  AOI211_X1 U13286 ( .C1(n15090), .C2(n14580), .A(n10677), .B(n11202), .ZN(
        n10678) );
  OAI211_X1 U13287 ( .C1(n15289), .C2(n11210), .A(n11206), .B(n10678), .ZN(
        n10681) );
  NAND2_X1 U13288 ( .A1(n10681), .A2(n6403), .ZN(n10679) );
  OAI21_X1 U13289 ( .B1(n6403), .B2(n10680), .A(n10679), .ZN(P1_U3462) );
  INV_X2 U13290 ( .A(n15331), .ZN(n15327) );
  NAND2_X1 U13291 ( .A1(n10681), .A2(n15327), .ZN(n10682) );
  OAI21_X1 U13292 ( .B1(n15327), .B2(n10158), .A(n10682), .ZN(P1_U3529) );
  INV_X1 U13293 ( .A(SI_17_), .ZN(n10683) );
  OAI222_X1 U13294 ( .A1(P3_U3151), .A2(n12576), .B1(n12948), .B2(n10684), 
        .C1(n10683), .C2(n12941), .ZN(P3_U3278) );
  INV_X1 U13295 ( .A(n10685), .ZN(n10759) );
  INV_X1 U13296 ( .A(n14644), .ZN(n14645) );
  OAI222_X1 U13297 ( .A1(n15147), .A2(n10759), .B1(n15144), .B2(n10686), .C1(
        n14645), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13298 ( .A(n10687), .ZN(n10688) );
  NAND2_X1 U13299 ( .A1(n10688), .A2(n10836), .ZN(n10689) );
  XNOR2_X1 U13300 ( .A(n12293), .B(n10697), .ZN(n10691) );
  NAND2_X1 U13301 ( .A1(n10691), .A2(n10850), .ZN(n10845) );
  INV_X1 U13302 ( .A(n10691), .ZN(n10692) );
  NAND2_X1 U13303 ( .A1(n10692), .A2(n12460), .ZN(n10693) );
  NAND2_X1 U13304 ( .A1(n10845), .A2(n10693), .ZN(n10695) );
  INV_X1 U13305 ( .A(n10846), .ZN(n10694) );
  AOI21_X1 U13306 ( .B1(n10696), .B2(n10695), .A(n10694), .ZN(n10703) );
  INV_X1 U13307 ( .A(n11405), .ZN(n10701) );
  INV_X1 U13308 ( .A(n12459), .ZN(n11018) );
  AOI22_X1 U13309 ( .A1(n12427), .A2(n10836), .B1(n12414), .B2(n10697), .ZN(
        n10699) );
  OAI211_X1 U13310 ( .C1(n11018), .C2(n12429), .A(n10699), .B(n10698), .ZN(
        n10700) );
  AOI21_X1 U13311 ( .B1(n10701), .B2(n12441), .A(n10700), .ZN(n10702) );
  OAI21_X1 U13312 ( .B1(n10703), .B2(n12434), .A(n10702), .ZN(P3_U3170) );
  NAND2_X1 U13313 ( .A1(n7079), .A2(n7590), .ZN(n10704) );
  AND2_X1 U13314 ( .A1(n10705), .A2(n10704), .ZN(n11255) );
  OAI22_X1 U13315 ( .A1(n6906), .A2(n13676), .B1(n9524), .B2(n13678), .ZN(
        n10707) );
  NOR2_X1 U13316 ( .A1(n11255), .A2(n15422), .ZN(n10706) );
  AOI211_X1 U13317 ( .C1(n13717), .C2(n10708), .A(n10707), .B(n10706), .ZN(
        n11258) );
  NAND2_X1 U13318 ( .A1(n11051), .A2(n13113), .ZN(n10709) );
  NAND2_X1 U13319 ( .A1(n13840), .A2(n10709), .ZN(n10710) );
  OR2_X1 U13320 ( .A1(n10710), .A2(n10986), .ZN(n11259) );
  OAI211_X1 U13321 ( .C1(n11255), .C2(n11267), .A(n11258), .B(n11259), .ZN(
        n10778) );
  AND2_X1 U13322 ( .A1(n15415), .A2(n15416), .ZN(n10711) );
  OAI22_X1 U13323 ( .A1(n13900), .A2(n11257), .B1(n15448), .B2(n9496), .ZN(
        n10714) );
  AOI21_X1 U13324 ( .B1(n10778), .B2(n15448), .A(n10714), .ZN(n10715) );
  INV_X1 U13325 ( .A(n10715), .ZN(P2_U3433) );
  XNOR2_X1 U13326 ( .A(n11138), .B(n10716), .ZN(n10721) );
  OAI22_X1 U13327 ( .A1(n6463), .A2(n10719), .B1(n10718), .B2(n10717), .ZN(
        n10720) );
  NOR2_X1 U13328 ( .A1(n10720), .A2(n10721), .ZN(n11135) );
  AOI21_X1 U13329 ( .B1(n10721), .B2(n10720), .A(n11135), .ZN(n10735) );
  NOR2_X1 U13330 ( .A1(n10722), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12087) );
  NOR2_X1 U13331 ( .A1(n15395), .A2(n11138), .ZN(n10723) );
  AOI211_X1 U13332 ( .C1(n15334), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n12087), 
        .B(n10723), .ZN(n10734) );
  INV_X1 U13333 ( .A(n10728), .ZN(n10726) );
  MUX2_X1 U13334 ( .A(n9653), .B(P2_REG2_REG_12__SCAN_IN), .S(n11138), .Z(
        n10729) );
  OR2_X1 U13335 ( .A1(n10724), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10727) );
  INV_X1 U13336 ( .A(n10727), .ZN(n10725) );
  NOR3_X1 U13337 ( .A1(n10726), .A2(n10729), .A3(n10725), .ZN(n10732) );
  NAND2_X1 U13338 ( .A1(n10728), .A2(n10727), .ZN(n10730) );
  NAND2_X1 U13339 ( .A1(n10730), .A2(n10729), .ZN(n11140) );
  INV_X1 U13340 ( .A(n11140), .ZN(n10731) );
  OAI21_X1 U13341 ( .B1(n10732), .B2(n10731), .A(n15405), .ZN(n10733) );
  OAI211_X1 U13342 ( .C1(n10735), .C2(n13430), .A(n10734), .B(n10733), .ZN(
        P2_U3226) );
  NAND2_X1 U13343 ( .A1(n15457), .A2(n15464), .ZN(n15456) );
  NAND2_X1 U13344 ( .A1(n15456), .A2(n10736), .ZN(n10737) );
  XNOR2_X1 U13345 ( .A(n10737), .B(n10738), .ZN(n11416) );
  OR2_X1 U13346 ( .A1(n10739), .A2(n10738), .ZN(n10832) );
  NAND2_X1 U13347 ( .A1(n10739), .A2(n10738), .ZN(n10740) );
  NAND3_X1 U13348 ( .A1(n10832), .A2(n12784), .A3(n10740), .ZN(n10742) );
  AOI22_X1 U13349 ( .A1(n15479), .A2(n12460), .B1(n15480), .B2(n12704), .ZN(
        n10741) );
  NAND2_X1 U13350 ( .A1(n10742), .A2(n10741), .ZN(n11413) );
  AOI21_X1 U13351 ( .B1(n11416), .B2(n15501), .A(n11413), .ZN(n11044) );
  INV_X1 U13352 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10743) );
  OAI22_X1 U13353 ( .A1(n12821), .A2(n11412), .B1(n15514), .B2(n10743), .ZN(
        n10744) );
  INV_X1 U13354 ( .A(n10744), .ZN(n10745) );
  OAI21_X1 U13355 ( .B1(n11044), .B2(n9433), .A(n10745), .ZN(P3_U3462) );
  OAI21_X1 U13356 ( .B1(n10747), .B2(n10752), .A(n10746), .ZN(n11073) );
  AOI211_X1 U13357 ( .C1(n13119), .C2(n10985), .A(n13542), .B(n10748), .ZN(
        n11074) );
  NAND3_X1 U13358 ( .A1(n10750), .A2(n10752), .A3(n10751), .ZN(n10753) );
  NAND2_X1 U13359 ( .A1(n10749), .A2(n10753), .ZN(n10754) );
  NAND2_X1 U13360 ( .A1(n10754), .A2(n13717), .ZN(n10756) );
  AOI22_X1 U13361 ( .A1(n13722), .A2(n13354), .B1(n13352), .B2(n13723), .ZN(
        n10755) );
  NAND2_X1 U13362 ( .A1(n10756), .A2(n10755), .ZN(n11075) );
  AOI211_X1 U13363 ( .C1(n13835), .C2(n11073), .A(n11074), .B(n11075), .ZN(
        n10797) );
  OAI22_X1 U13364 ( .A1(n13900), .A2(n11029), .B1(n15448), .B2(n9526), .ZN(
        n10757) );
  INV_X1 U13365 ( .A(n10757), .ZN(n10758) );
  OAI21_X1 U13366 ( .B1(n10797), .B2(n15446), .A(n10758), .ZN(P2_U3439) );
  INV_X1 U13367 ( .A(n13410), .ZN(n15394) );
  OAI222_X1 U13368 ( .A1(P2_U3088), .A2(n15394), .B1(n13916), .B2(n10760), 
        .C1(n13913), .C2(n10759), .ZN(P2_U3310) );
  NOR2_X1 U13369 ( .A1(n10762), .A2(n10761), .ZN(n10764) );
  XNOR2_X1 U13370 ( .A(n10769), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n10763) );
  AOI21_X1 U13371 ( .B1(n10764), .B2(n10763), .A(n11108), .ZN(n10776) );
  NOR2_X1 U13372 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14149), .ZN(n10766) );
  NOR2_X1 U13373 ( .A1(n15221), .A2(n11109), .ZN(n10765) );
  AOI211_X1 U13374 ( .C1(n14653), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10766), 
        .B(n10765), .ZN(n10775) );
  INV_X1 U13375 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10770) );
  MUX2_X1 U13376 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10770), .S(n10769), .Z(
        n10771) );
  NAND2_X1 U13377 ( .A1(n10772), .A2(n10771), .ZN(n11151) );
  OAI21_X1 U13378 ( .B1(n10772), .B2(n10771), .A(n11151), .ZN(n10773) );
  NAND2_X1 U13379 ( .A1(n10773), .A2(n15217), .ZN(n10774) );
  OAI211_X1 U13380 ( .C1(n10776), .C2(n14668), .A(n10775), .B(n10774), .ZN(
        P1_U3255) );
  OAI22_X1 U13381 ( .A1(n13838), .A2(n11257), .B1(n15454), .B2(n10072), .ZN(
        n10777) );
  AOI21_X1 U13382 ( .B1(n10778), .B2(n15454), .A(n10777), .ZN(n10779) );
  INV_X1 U13383 ( .A(n10779), .ZN(P2_U3500) );
  AOI211_X1 U13384 ( .C1(n10781), .C2(n10780), .A(n10283), .B(n11506), .ZN(
        n11229) );
  AOI21_X1 U13385 ( .B1(n10781), .B2(n15315), .A(n11229), .ZN(n10794) );
  OAI21_X1 U13386 ( .B1(n10784), .B2(n10783), .A(n10782), .ZN(n10785) );
  NAND2_X1 U13387 ( .A1(n10785), .A2(n15321), .ZN(n10792) );
  OAI21_X1 U13388 ( .B1(n14321), .B2(n14527), .A(n10786), .ZN(n10790) );
  NAND2_X1 U13389 ( .A1(n9228), .A2(n15107), .ZN(n10788) );
  NAND2_X1 U13390 ( .A1(n14579), .A2(n15090), .ZN(n10787) );
  NAND2_X1 U13391 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  AOI21_X1 U13392 ( .B1(n10790), .B2(n15308), .A(n10789), .ZN(n10791) );
  NAND2_X1 U13393 ( .A1(n10792), .A2(n10791), .ZN(n11231) );
  INV_X1 U13394 ( .A(n11231), .ZN(n10793) );
  NAND2_X1 U13395 ( .A1(n10794), .A2(n10793), .ZN(n10798) );
  NAND2_X1 U13396 ( .A1(n10798), .A2(n15327), .ZN(n10795) );
  OAI21_X1 U13397 ( .B1(n15327), .B2(n10160), .A(n10795), .ZN(P1_U3530) );
  AOI22_X1 U13398 ( .A1(n13789), .A2(n13119), .B1(n15452), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10796) );
  OAI21_X1 U13399 ( .B1(n10797), .B2(n15452), .A(n10796), .ZN(P2_U3502) );
  NAND2_X1 U13400 ( .A1(n10798), .A2(n6403), .ZN(n10799) );
  OAI21_X1 U13401 ( .B1(n6403), .B2(n8742), .A(n10799), .ZN(P1_U3465) );
  NAND2_X1 U13402 ( .A1(n13354), .A2(n12272), .ZN(n10807) );
  NAND2_X1 U13403 ( .A1(n10808), .A2(n10807), .ZN(n10859) );
  OAI21_X1 U13404 ( .B1(n10808), .B2(n10807), .A(n10859), .ZN(n10809) );
  AOI21_X1 U13405 ( .B1(n10810), .B2(n10809), .A(n10861), .ZN(n10824) );
  NAND3_X1 U13406 ( .A1(n15416), .A2(n10812), .A3(n15439), .ZN(n10813) );
  NAND2_X1 U13407 ( .A1(n15416), .A2(n13286), .ZN(n13329) );
  NAND2_X1 U13408 ( .A1(n10819), .A2(n10814), .ZN(n10816) );
  NAND2_X1 U13409 ( .A1(n10816), .A2(n10815), .ZN(n10857) );
  INV_X1 U13410 ( .A(n15416), .ZN(n15419) );
  OR2_X1 U13411 ( .A1(n10857), .A2(n15419), .ZN(n11016) );
  AOI22_X1 U13412 ( .A1(n13083), .A2(n10801), .B1(n11016), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13413 ( .A1(n13061), .A2(n13723), .ZN(n13081) );
  INV_X1 U13414 ( .A(n13081), .ZN(n13052) );
  INV_X1 U13415 ( .A(n15421), .ZN(n10817) );
  AND2_X1 U13416 ( .A1(n10817), .A2(n13298), .ZN(n10990) );
  NAND2_X1 U13417 ( .A1(n15416), .A2(n10990), .ZN(n10818) );
  AOI22_X1 U13418 ( .A1(n13052), .A2(n13353), .B1(n10805), .B2(n13087), .ZN(
        n10822) );
  OAI211_X1 U13419 ( .C1(n10824), .C2(n13089), .A(n10823), .B(n10822), .ZN(
        P2_U3209) );
  INV_X1 U13420 ( .A(n10825), .ZN(n10828) );
  OAI222_X1 U13421 ( .A1(n7072), .A2(P1_U3086), .B1(n15147), .B2(n10828), .C1(
        n10826), .C2(n15144), .ZN(P1_U3340) );
  INV_X1 U13422 ( .A(n11887), .ZN(n11611) );
  OAI222_X1 U13423 ( .A1(n11611), .A2(P2_U3088), .B1(n13913), .B2(n10828), 
        .C1(n10827), .C2(n13916), .ZN(P2_U3312) );
  NAND2_X1 U13424 ( .A1(n10829), .A2(n10833), .ZN(n11083) );
  OAI21_X1 U13425 ( .B1(n10829), .B2(n10833), .A(n11083), .ZN(n11410) );
  INV_X1 U13426 ( .A(n10830), .ZN(n10831) );
  NAND2_X1 U13427 ( .A1(n10832), .A2(n10831), .ZN(n10834) );
  XNOR2_X1 U13428 ( .A(n10834), .B(n10833), .ZN(n10835) );
  NAND2_X1 U13429 ( .A1(n10835), .A2(n12784), .ZN(n10838) );
  AOI22_X1 U13430 ( .A1(n15479), .A2(n12459), .B1(n10836), .B2(n12704), .ZN(
        n10837) );
  NAND2_X1 U13431 ( .A1(n10838), .A2(n10837), .ZN(n11407) );
  AOI21_X1 U13432 ( .B1(n15501), .B2(n11410), .A(n11407), .ZN(n11040) );
  OAI22_X1 U13433 ( .A1(n12821), .A2(n11406), .B1(n15514), .B2(n10409), .ZN(
        n10839) );
  INV_X1 U13434 ( .A(n10839), .ZN(n10840) );
  OAI21_X1 U13435 ( .B1(n11040), .B2(n9433), .A(n10840), .ZN(P3_U3463) );
  INV_X1 U13436 ( .A(n10841), .ZN(n10843) );
  INV_X1 U13437 ( .A(n12599), .ZN(n10842) );
  OAI222_X1 U13438 ( .A1(n12941), .A2(n10844), .B1(n12948), .B2(n10843), .C1(
        P3_U3151), .C2(n10842), .ZN(P3_U3277) );
  INV_X1 U13439 ( .A(n12441), .ZN(n11433) );
  XNOR2_X1 U13440 ( .A(n12293), .B(n11093), .ZN(n11019) );
  XNOR2_X1 U13441 ( .A(n11019), .B(n12459), .ZN(n10848) );
  NAND2_X1 U13442 ( .A1(n10847), .A2(n10848), .ZN(n11179) );
  OAI21_X1 U13443 ( .B1(n10848), .B2(n10847), .A(n11179), .ZN(n10849) );
  NAND2_X1 U13444 ( .A1(n10849), .A2(n12439), .ZN(n10854) );
  INV_X1 U13445 ( .A(n12429), .ZN(n12445) );
  OAI22_X1 U13446 ( .A1(n12448), .A2(n11129), .B1(n10850), .B2(n12443), .ZN(
        n10851) );
  AOI211_X1 U13447 ( .C1(n12445), .C2(n12458), .A(n10852), .B(n10851), .ZN(
        n10853) );
  OAI211_X1 U13448 ( .C1(n11091), .C2(n11433), .A(n10854), .B(n10853), .ZN(
        P3_U3167) );
  INV_X1 U13449 ( .A(n10855), .ZN(n10856) );
  OR2_X1 U13450 ( .A1(n10857), .A2(n10856), .ZN(n10858) );
  INV_X1 U13451 ( .A(n10859), .ZN(n10860) );
  NAND2_X1 U13452 ( .A1(n13353), .A2(n12272), .ZN(n10862) );
  XNOR2_X1 U13453 ( .A(n13119), .B(n7171), .ZN(n10863) );
  XNOR2_X1 U13454 ( .A(n10862), .B(n10863), .ZN(n11026) );
  INV_X1 U13455 ( .A(n10862), .ZN(n10864) );
  INV_X2 U13456 ( .A(n10917), .ZN(n13542) );
  AND2_X1 U13457 ( .A1(n13352), .A2(n13542), .ZN(n10866) );
  XNOR2_X1 U13458 ( .A(n6405), .B(n7171), .ZN(n10865) );
  NOR2_X1 U13459 ( .A1(n10865), .A2(n10866), .ZN(n10920) );
  AOI21_X1 U13460 ( .B1(n10866), .B2(n10865), .A(n10920), .ZN(n10867) );
  OAI21_X1 U13461 ( .B1(n10868), .B2(n10867), .A(n10922), .ZN(n10869) );
  NAND2_X1 U13462 ( .A1(n10869), .A2(n13042), .ZN(n10872) );
  AND2_X1 U13463 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n15335) );
  INV_X1 U13464 ( .A(n13083), .ZN(n12994) );
  INV_X1 U13465 ( .A(n13353), .ZN(n10997) );
  INV_X1 U13466 ( .A(n13351), .ZN(n11240) );
  OAI22_X1 U13467 ( .A1(n12994), .A2(n10997), .B1(n11240), .B2(n13081), .ZN(
        n10870) );
  AOI211_X1 U13468 ( .C1(n6405), .C2(n13087), .A(n15335), .B(n10870), .ZN(
        n10871) );
  OAI211_X1 U13469 ( .C1(n13085), .C2(n11005), .A(n10872), .B(n10871), .ZN(
        P2_U3202) );
  OAI222_X1 U13470 ( .A1(n12941), .A2(n10874), .B1(n12948), .B2(n10873), .C1(
        n12596), .C2(P3_U3151), .ZN(P3_U3276) );
  MUX2_X1 U13471 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n8020), .S(n11470), .Z(
        n10877) );
  AOI21_X1 U13472 ( .B1(n10877), .B2(n10876), .A(n6593), .ZN(n10893) );
  MUX2_X1 U13473 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12937), .Z(n11468) );
  XNOR2_X1 U13474 ( .A(n11470), .B(n11468), .ZN(n11471) );
  XNOR2_X1 U13475 ( .A(n11472), .B(n11471), .ZN(n10891) );
  INV_X1 U13476 ( .A(n10882), .ZN(n10884) );
  INV_X1 U13477 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10883) );
  XNOR2_X1 U13478 ( .A(n11470), .B(n10883), .ZN(n10885) );
  AND3_X1 U13479 ( .A1(n10886), .A2(n10885), .A3(n10884), .ZN(n10887) );
  OAI21_X1 U13480 ( .B1(n11478), .B2(n10887), .A(n12590), .ZN(n10889) );
  AND2_X1 U13481 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11429) );
  AOI21_X1 U13482 ( .B1(n15455), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11429), .ZN(
        n10888) );
  OAI211_X1 U13483 ( .C1(n12597), .C2(n11479), .A(n10889), .B(n10888), .ZN(
        n10890) );
  AOI21_X1 U13484 ( .B1(n12491), .B2(n10891), .A(n10890), .ZN(n10892) );
  OAI21_X1 U13485 ( .B1(n10893), .B2(n12024), .A(n10892), .ZN(P3_U3190) );
  INV_X1 U13486 ( .A(n10895), .ZN(n10897) );
  NAND2_X1 U13487 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  NAND2_X1 U13488 ( .A1(n14579), .A2(n10286), .ZN(n10900) );
  NAND2_X1 U13489 ( .A1(n14094), .A2(n10284), .ZN(n10899) );
  NAND2_X1 U13490 ( .A1(n10900), .A2(n10899), .ZN(n10901) );
  XNOR2_X1 U13491 ( .A(n10901), .B(n14051), .ZN(n10904) );
  AOI22_X1 U13492 ( .A1(n14579), .A2(n14108), .B1(n14094), .B2(n10286), .ZN(
        n10903) );
  XNOR2_X1 U13493 ( .A(n10904), .B(n10903), .ZN(n14090) );
  OR2_X1 U13494 ( .A1(n10904), .A2(n10903), .ZN(n10905) );
  NAND2_X1 U13495 ( .A1(n14092), .A2(n10905), .ZN(n11445) );
  NAND2_X1 U13496 ( .A1(n15250), .A2(n10286), .ZN(n10907) );
  OR2_X1 U13497 ( .A1(n15246), .A2(n14011), .ZN(n10906) );
  NAND2_X1 U13498 ( .A1(n10907), .A2(n10906), .ZN(n10908) );
  XNOR2_X1 U13499 ( .A(n10908), .B(n14111), .ZN(n11440) );
  NAND2_X1 U13500 ( .A1(n15250), .A2(n14108), .ZN(n10910) );
  OR2_X1 U13501 ( .A1(n15246), .A2(n14020), .ZN(n10909) );
  NAND2_X1 U13502 ( .A1(n10910), .A2(n10909), .ZN(n11439) );
  INV_X1 U13503 ( .A(n11439), .ZN(n11441) );
  XNOR2_X1 U13504 ( .A(n11440), .B(n11441), .ZN(n10911) );
  XNOR2_X1 U13505 ( .A(n11445), .B(n10911), .ZN(n10916) );
  NAND2_X1 U13506 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15224) );
  OAI21_X1 U13507 ( .B1(n14286), .B2(n11322), .A(n15224), .ZN(n10913) );
  AOI21_X1 U13508 ( .B1(n15285), .B2(n14300), .A(n10913), .ZN(n10915) );
  INV_X1 U13509 ( .A(n14272), .ZN(n14133) );
  AOI22_X1 U13510 ( .A1(n14133), .A2(n14578), .B1(n14275), .B2(n14579), .ZN(
        n10914) );
  OAI211_X1 U13511 ( .C1(n10916), .C2(n14302), .A(n10915), .B(n10914), .ZN(
        P1_U3230) );
  AND2_X1 U13512 ( .A1(n13351), .A2(n13542), .ZN(n10919) );
  XNOR2_X1 U13513 ( .A(n13129), .B(n7171), .ZN(n10918) );
  NOR2_X1 U13514 ( .A1(n10918), .A2(n10919), .ZN(n11211) );
  AOI21_X1 U13515 ( .B1(n10919), .B2(n10918), .A(n11211), .ZN(n10924) );
  INV_X1 U13516 ( .A(n10920), .ZN(n10921) );
  OAI21_X1 U13517 ( .B1(n10924), .B2(n10923), .A(n11213), .ZN(n10925) );
  NAND2_X1 U13518 ( .A1(n10925), .A2(n13042), .ZN(n10929) );
  INV_X1 U13519 ( .A(n13352), .ZN(n11057) );
  OAI22_X1 U13520 ( .A1(n12994), .A2(n11057), .B1(n11056), .B2(n13081), .ZN(
        n10926) );
  AOI211_X1 U13521 ( .C1(n13129), .C2(n13087), .A(n10927), .B(n10926), .ZN(
        n10928) );
  OAI211_X1 U13522 ( .C1(n13085), .C2(n11067), .A(n10929), .B(n10928), .ZN(
        P2_U3199) );
  XNOR2_X1 U13523 ( .A(n10932), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n10935) );
  XNOR2_X1 U13524 ( .A(n11551), .B(n10933), .ZN(n11550) );
  INV_X1 U13525 ( .A(n11550), .ZN(n10934) );
  XNOR2_X1 U13526 ( .A(n10934), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n10941) );
  INV_X1 U13527 ( .A(n10941), .ZN(n10939) );
  INV_X1 U13528 ( .A(n10935), .ZN(n10936) );
  XNOR2_X1 U13529 ( .A(n10937), .B(n10936), .ZN(n15156) );
  NAND2_X1 U13530 ( .A1(n10939), .A2(n10938), .ZN(n11548) );
  NAND2_X1 U13531 ( .A1(n11548), .A2(n11547), .ZN(n10942) );
  XNOR2_X1 U13532 ( .A(n10942), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  NOR2_X1 U13533 ( .A1(n15510), .A2(n6622), .ZN(n10943) );
  AOI21_X1 U13534 ( .B1(n15510), .B2(n10944), .A(n10943), .ZN(n10945) );
  OAI21_X1 U13535 ( .B1(n10946), .B2(n12894), .A(n10945), .ZN(P3_U3390) );
  OAI21_X1 U13536 ( .B1(n10949), .B2(n10948), .A(n10947), .ZN(n11423) );
  OAI211_X1 U13537 ( .C1(n10951), .C2(n11164), .A(n10950), .B(n12784), .ZN(
        n10953) );
  AOI22_X1 U13538 ( .A1(n12704), .A2(n12458), .B1(n12456), .B2(n15479), .ZN(
        n10952) );
  NAND2_X1 U13539 ( .A1(n10953), .A2(n10952), .ZN(n11420) );
  AOI21_X1 U13540 ( .B1(n15501), .B2(n11423), .A(n11420), .ZN(n11037) );
  OAI22_X1 U13541 ( .A1(n12821), .A2(n11419), .B1(n15514), .B2(n8002), .ZN(
        n10954) );
  INV_X1 U13542 ( .A(n10954), .ZN(n10955) );
  OAI21_X1 U13543 ( .B1(n11037), .B2(n9433), .A(n10955), .ZN(P3_U3466) );
  INV_X1 U13544 ( .A(n10956), .ZN(n10957) );
  INV_X1 U13545 ( .A(n13087), .ZN(n13049) );
  OAI21_X1 U13546 ( .B1(n10957), .B2(n13089), .A(n13049), .ZN(n10958) );
  AOI22_X1 U13547 ( .A1(n10958), .A2(n11051), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n11016), .ZN(n10960) );
  NAND4_X1 U13548 ( .A1(n13042), .A2(n13542), .A3(n7148), .A4(n10803), .ZN(
        n10959) );
  OAI211_X1 U13549 ( .C1(n6602), .C2(n13081), .A(n10960), .B(n10959), .ZN(
        P2_U3204) );
  OAI21_X1 U13550 ( .B1(n10963), .B2(n10962), .A(n10961), .ZN(n10964) );
  INV_X1 U13551 ( .A(n10964), .ZN(n11103) );
  OR2_X1 U13552 ( .A1(n11085), .A2(n11086), .ZN(n11087) );
  NAND2_X1 U13553 ( .A1(n11087), .A2(n10965), .ZN(n10967) );
  XNOR2_X1 U13554 ( .A(n10967), .B(n10966), .ZN(n10969) );
  OAI22_X1 U13555 ( .A1(n11018), .A2(n15467), .B1(n6933), .B2(n15469), .ZN(
        n10968) );
  AOI21_X1 U13556 ( .B1(n10969), .B2(n12784), .A(n10968), .ZN(n11097) );
  OAI21_X1 U13557 ( .B1(n12797), .B2(n11103), .A(n11097), .ZN(n11123) );
  OAI22_X1 U13558 ( .A1(n12821), .A2(n11121), .B1(n15514), .B2(n10401), .ZN(
        n10970) );
  AOI21_X1 U13559 ( .B1(n11123), .B2(n15514), .A(n10970), .ZN(n10971) );
  INV_X1 U13560 ( .A(n10971), .ZN(P3_U3465) );
  INV_X1 U13561 ( .A(n10972), .ZN(n10973) );
  NAND3_X1 U13562 ( .A1(n10979), .A2(n10976), .A3(n10975), .ZN(n10977) );
  AND2_X1 U13563 ( .A1(n10750), .A2(n10977), .ZN(n10983) );
  OAI21_X1 U13564 ( .B1(n10980), .B2(n10979), .A(n10978), .ZN(n15427) );
  INV_X1 U13565 ( .A(n15422), .ZN(n11247) );
  NAND2_X1 U13566 ( .A1(n15427), .A2(n11247), .ZN(n10982) );
  AOI22_X1 U13567 ( .A1(n13722), .A2(n10801), .B1(n13353), .B2(n13723), .ZN(
        n10981) );
  OAI211_X1 U13568 ( .C1(n10983), .C2(n13701), .A(n10982), .B(n10981), .ZN(
        n15431) );
  NOR2_X1 U13569 ( .A1(n13687), .A2(n15528), .ZN(n10988) );
  OAI211_X1 U13570 ( .C1(n10986), .C2(n7152), .A(n13840), .B(n10985), .ZN(
        n15428) );
  OAI22_X1 U13571 ( .A1(n13549), .A2(n15428), .B1(n13370), .B2(n13683), .ZN(
        n10987) );
  AOI211_X1 U13572 ( .C1(n13687), .C2(n15431), .A(n10988), .B(n10987), .ZN(
        n10992) );
  NOR2_X1 U13573 ( .A1(n13284), .A2(n13666), .ZN(n10989) );
  AND2_X1 U13574 ( .A1(n13687), .A2(n10989), .ZN(n10996) );
  AOI22_X1 U13575 ( .A1(n10996), .A2(n15427), .B1(n13649), .B2(n10805), .ZN(
        n10991) );
  NAND2_X1 U13576 ( .A1(n10992), .A2(n10991), .ZN(P2_U3263) );
  OR2_X1 U13577 ( .A1(n10993), .A2(n11000), .ZN(n10994) );
  NAND2_X1 U13578 ( .A1(n10995), .A2(n10994), .ZN(n15436) );
  INV_X1 U13579 ( .A(n15436), .ZN(n11009) );
  OAI22_X1 U13580 ( .A1(n10997), .A2(n13676), .B1(n11240), .B2(n13678), .ZN(
        n11003) );
  NAND3_X1 U13581 ( .A1(n10749), .A2(n11000), .A3(n10999), .ZN(n11001) );
  AOI21_X1 U13582 ( .B1(n10998), .B2(n11001), .A(n13701), .ZN(n11002) );
  AOI211_X1 U13583 ( .C1(n11247), .C2(n15436), .A(n11003), .B(n11002), .ZN(
        n15433) );
  MUX2_X1 U13584 ( .A(n11004), .B(n15433), .S(n13687), .Z(n11008) );
  OAI211_X1 U13585 ( .C1(n10748), .C2(n7686), .A(n13840), .B(n11064), .ZN(
        n15432) );
  OAI22_X1 U13586 ( .A1(n13549), .A2(n15432), .B1(n11005), .B2(n13683), .ZN(
        n11006) );
  AOI21_X1 U13587 ( .B1(n13649), .B2(n6405), .A(n11006), .ZN(n11007) );
  OAI211_X1 U13588 ( .C1(n11009), .C2(n11256), .A(n11008), .B(n11007), .ZN(
        P2_U3261) );
  AOI21_X1 U13589 ( .B1(n11012), .B2(n11011), .A(n11010), .ZN(n11013) );
  OAI22_X1 U13590 ( .A1(n13049), .A2(n11257), .B1(n11013), .B2(n13089), .ZN(
        n11015) );
  OAI22_X1 U13591 ( .A1(n12994), .A2(n6906), .B1(n9524), .B2(n13081), .ZN(
        n11014) );
  AOI211_X1 U13592 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n11016), .A(n11015), .B(
        n11014), .ZN(n11017) );
  INV_X1 U13593 ( .A(n11017), .ZN(P2_U3194) );
  NAND2_X1 U13594 ( .A1(n11019), .A2(n11018), .ZN(n11175) );
  AND2_X1 U13595 ( .A1(n11179), .A2(n11175), .ZN(n11021) );
  XNOR2_X1 U13596 ( .A(n12293), .B(n11121), .ZN(n11176) );
  XOR2_X1 U13597 ( .A(n12458), .B(n11176), .Z(n11020) );
  NAND2_X1 U13598 ( .A1(n11021), .A2(n11020), .ZN(n11163) );
  OAI211_X1 U13599 ( .C1(n11021), .C2(n11020), .A(n11163), .B(n12439), .ZN(
        n11025) );
  OAI22_X1 U13600 ( .A1(n12448), .A2(n11121), .B1(n6933), .B2(n12429), .ZN(
        n11022) );
  AOI211_X1 U13601 ( .C1(n12427), .C2(n12459), .A(n11023), .B(n11022), .ZN(
        n11024) );
  OAI211_X1 U13602 ( .C1(n11098), .C2(n11433), .A(n11025), .B(n11024), .ZN(
        P3_U3179) );
  XNOR2_X1 U13603 ( .A(n11027), .B(n11026), .ZN(n11033) );
  INV_X1 U13604 ( .A(n13085), .ZN(n13072) );
  INV_X1 U13605 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U13606 ( .A1(n13052), .A2(n13352), .B1(n13083), .B2(n13354), .ZN(
        n11028) );
  NAND2_X1 U13607 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13381) );
  OAI211_X1 U13608 ( .C1(n11029), .C2(n13049), .A(n11028), .B(n13381), .ZN(
        n11030) );
  AOI21_X1 U13609 ( .B1(n13072), .B2(n11031), .A(n11030), .ZN(n11032) );
  OAI21_X1 U13610 ( .B1(n11033), .B2(n13089), .A(n11032), .ZN(P2_U3190) );
  INV_X1 U13611 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11034) );
  OAI22_X1 U13612 ( .A1(n12894), .A2(n11419), .B1(n15510), .B2(n11034), .ZN(
        n11035) );
  INV_X1 U13613 ( .A(n11035), .ZN(n11036) );
  OAI21_X1 U13614 ( .B1(n11037), .B2(n15509), .A(n11036), .ZN(P3_U3411) );
  OAI22_X1 U13615 ( .A1(n12894), .A2(n11406), .B1(n15510), .B2(n7961), .ZN(
        n11038) );
  INV_X1 U13616 ( .A(n11038), .ZN(n11039) );
  OAI21_X1 U13617 ( .B1(n11040), .B2(n15509), .A(n11039), .ZN(P3_U3402) );
  INV_X1 U13618 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11041) );
  OAI22_X1 U13619 ( .A1(n12894), .A2(n11412), .B1(n15510), .B2(n11041), .ZN(
        n11042) );
  INV_X1 U13620 ( .A(n11042), .ZN(n11043) );
  OAI21_X1 U13621 ( .B1(n11044), .B2(n15509), .A(n11043), .ZN(P3_U3399) );
  NAND2_X1 U13622 ( .A1(n15422), .A2(n13666), .ZN(n11045) );
  OR2_X1 U13623 ( .A1(n7148), .A2(n11051), .ZN(n11047) );
  NAND2_X1 U13624 ( .A1(n10803), .A2(n11047), .ZN(n15423) );
  OAI22_X1 U13625 ( .A1(n15423), .A2(n13701), .B1(n6602), .B2(n13678), .ZN(
        n15424) );
  INV_X1 U13626 ( .A(n15424), .ZN(n11049) );
  OAI22_X1 U13627 ( .A1(n6402), .A2(n11049), .B1(n11048), .B2(n13683), .ZN(
        n11050) );
  AOI21_X1 U13628 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n6402), .A(n11050), .ZN(
        n11053) );
  NOR2_X1 U13629 ( .A1(n13549), .A2(n12272), .ZN(n13741) );
  OAI21_X1 U13630 ( .B1(n13741), .B2(n13649), .A(n11051), .ZN(n11052) );
  OAI211_X1 U13631 ( .C1(n13738), .C2(n15423), .A(n11053), .B(n11052), .ZN(
        P2_U3265) );
  OAI21_X1 U13632 ( .B1(n11055), .B2(n13302), .A(n11054), .ZN(n11271) );
  INV_X1 U13633 ( .A(n11271), .ZN(n11072) );
  OAI22_X1 U13634 ( .A1(n11057), .A2(n13676), .B1(n11056), .B2(n13678), .ZN(
        n11062) );
  NAND3_X1 U13635 ( .A1(n10998), .A2(n13302), .A3(n11059), .ZN(n11060) );
  AOI21_X1 U13636 ( .B1(n11058), .B2(n11060), .A(n13701), .ZN(n11061) );
  AOI211_X1 U13637 ( .C1(n11247), .C2(n11271), .A(n11062), .B(n11061), .ZN(
        n11268) );
  MUX2_X1 U13638 ( .A(n11063), .B(n11268), .S(n13687), .Z(n11071) );
  NAND2_X1 U13639 ( .A1(n11064), .A2(n13129), .ZN(n11065) );
  NAND2_X1 U13640 ( .A1(n11065), .A2(n13840), .ZN(n11066) );
  NOR2_X1 U13641 ( .A1(n11249), .A2(n11066), .ZN(n11270) );
  INV_X1 U13642 ( .A(n11270), .ZN(n11068) );
  OAI22_X1 U13643 ( .A1(n13549), .A2(n11068), .B1(n11067), .B2(n13683), .ZN(
        n11069) );
  AOI21_X1 U13644 ( .B1(n13649), .B2(n13129), .A(n11069), .ZN(n11070) );
  OAI211_X1 U13645 ( .C1(n11072), .C2(n11256), .A(n11071), .B(n11070), .ZN(
        P2_U3260) );
  INV_X1 U13646 ( .A(n11073), .ZN(n11080) );
  AOI22_X1 U13647 ( .A1(n13649), .A2(n13119), .B1(n13708), .B2(n11074), .ZN(
        n11079) );
  INV_X1 U13648 ( .A(n13683), .ZN(n13731) );
  AOI21_X1 U13649 ( .B1(n13731), .B2(n11031), .A(n11075), .ZN(n11076) );
  MUX2_X1 U13650 ( .A(n11077), .B(n11076), .S(n13687), .Z(n11078) );
  OAI211_X1 U13651 ( .C1(n11080), .C2(n13738), .A(n11079), .B(n11078), .ZN(
        P2_U3262) );
  NAND2_X1 U13652 ( .A1(n15462), .A2(n11081), .ZN(n11279) );
  NAND2_X1 U13653 ( .A1(n11357), .A2(n11279), .ZN(n15471) );
  NAND2_X1 U13654 ( .A1(n11083), .A2(n11082), .ZN(n11084) );
  XOR2_X1 U13655 ( .A(n11086), .B(n11084), .Z(n11126) );
  INV_X1 U13656 ( .A(n11085), .ZN(n11088) );
  OAI21_X1 U13657 ( .B1(n11088), .B2(n7286), .A(n11087), .ZN(n11089) );
  AOI222_X1 U13658 ( .A1(n12784), .A2(n11089), .B1(n12458), .B2(n15479), .C1(
        n12460), .C2(n12704), .ZN(n11125) );
  MUX2_X1 U13659 ( .A(n11090), .B(n11125), .S(n15472), .Z(n11095) );
  INV_X1 U13660 ( .A(n11091), .ZN(n11092) );
  AOI22_X1 U13661 ( .A1(n12787), .A2(n11093), .B1(n15488), .B2(n11092), .ZN(
        n11094) );
  OAI211_X1 U13662 ( .C1(n12790), .C2(n11126), .A(n11095), .B(n11094), .ZN(
        P3_U3228) );
  MUX2_X1 U13663 ( .A(n11097), .B(n11096), .S(n15493), .Z(n11102) );
  INV_X1 U13664 ( .A(n11098), .ZN(n11099) );
  AOI22_X1 U13665 ( .A1(n12787), .A2(n11100), .B1(n15488), .B2(n11099), .ZN(
        n11101) );
  OAI211_X1 U13666 ( .C1(n11103), .C2(n12790), .A(n11102), .B(n11101), .ZN(
        P3_U3227) );
  XNOR2_X1 U13667 ( .A(n11112), .B(n11104), .ZN(n11153) );
  NAND2_X1 U13668 ( .A1(n11109), .A2(n10770), .ZN(n11150) );
  NAND3_X1 U13669 ( .A1(n11151), .A2(n11153), .A3(n11150), .ZN(n11152) );
  NAND2_X1 U13670 ( .A1(n11112), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11106) );
  MUX2_X1 U13671 ( .A(n8972), .B(P1_REG2_REG_14__SCAN_IN), .S(n11801), .Z(
        n11105) );
  AOI21_X1 U13672 ( .B1(n11152), .B2(n11106), .A(n11105), .ZN(n11800) );
  NAND3_X1 U13673 ( .A1(n11152), .A2(n11106), .A3(n11105), .ZN(n11107) );
  NAND2_X1 U13674 ( .A1(n11107), .A2(n15217), .ZN(n11120) );
  AOI21_X1 U13675 ( .B1(n11110), .B2(n11109), .A(n11108), .ZN(n11156) );
  XOR2_X1 U13676 ( .A(n11112), .B(P1_REG1_REG_13__SCAN_IN), .Z(n11157) );
  NAND2_X1 U13677 ( .A1(n11156), .A2(n11157), .ZN(n11155) );
  XNOR2_X1 U13678 ( .A(n11801), .B(n11111), .ZN(n11113) );
  NAND2_X1 U13679 ( .A1(n11112), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11114) );
  NAND3_X1 U13680 ( .A1(n11155), .A2(n11113), .A3(n11114), .ZN(n11793) );
  INV_X1 U13681 ( .A(n11793), .ZN(n11116) );
  AOI21_X1 U13682 ( .B1(n11155), .B2(n11114), .A(n11113), .ZN(n11115) );
  OAI21_X1 U13683 ( .B1(n11116), .B2(n11115), .A(n15210), .ZN(n11119) );
  INV_X1 U13684 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n11845) );
  NAND2_X1 U13685 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14076)
         );
  OAI21_X1 U13686 ( .B1(n15226), .B2(n11845), .A(n14076), .ZN(n11117) );
  AOI21_X1 U13687 ( .B1(n14654), .B2(n11801), .A(n11117), .ZN(n11118) );
  OAI211_X1 U13688 ( .C1(n11800), .C2(n11120), .A(n11119), .B(n11118), .ZN(
        P1_U3257) );
  OAI22_X1 U13689 ( .A1(n12894), .A2(n11121), .B1(n15510), .B2(n15518), .ZN(
        n11122) );
  AOI21_X1 U13690 ( .B1(n11123), .B2(n15510), .A(n11122), .ZN(n11124) );
  INV_X1 U13691 ( .A(n11124), .ZN(P3_U3408) );
  OAI21_X1 U13692 ( .B1(n12797), .B2(n11126), .A(n11125), .ZN(n11131) );
  OAI22_X1 U13693 ( .A1(n12821), .A2(n11129), .B1(n15514), .B2(n7944), .ZN(
        n11127) );
  AOI21_X1 U13694 ( .B1(n11131), .B2(n15514), .A(n11127), .ZN(n11128) );
  INV_X1 U13695 ( .A(n11128), .ZN(P3_U3464) );
  OAI22_X1 U13696 ( .A1(n12894), .A2(n11129), .B1(n15510), .B2(n7940), .ZN(
        n11130) );
  AOI21_X1 U13697 ( .B1(n11131), .B2(n15510), .A(n11130), .ZN(n11132) );
  INV_X1 U13698 ( .A(n11132), .ZN(P3_U3405) );
  XNOR2_X1 U13699 ( .A(n11608), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11137) );
  NOR2_X1 U13700 ( .A1(n11133), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11134) );
  OR2_X1 U13701 ( .A1(n11135), .A2(n11134), .ZN(n11136) );
  NOR3_X1 U13702 ( .A1(n11135), .A2(n11134), .A3(n11137), .ZN(n11607) );
  AOI211_X1 U13703 ( .C1(n11137), .C2(n11136), .A(n13430), .B(n11607), .ZN(
        n11149) );
  NAND2_X1 U13704 ( .A1(n11138), .A2(n9653), .ZN(n11139) );
  INV_X1 U13705 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11141) );
  MUX2_X1 U13706 ( .A(n11141), .B(P2_REG2_REG_13__SCAN_IN), .S(n11608), .Z(
        n11143) );
  INV_X1 U13707 ( .A(n11603), .ZN(n11142) );
  AOI211_X1 U13708 ( .C1(n11144), .C2(n11143), .A(n11894), .B(n11142), .ZN(
        n11148) );
  NAND2_X1 U13709 ( .A1(n15334), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U13710 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n12117)
         );
  OAI211_X1 U13711 ( .C1(n15395), .C2(n11146), .A(n11145), .B(n12117), .ZN(
        n11147) );
  OR3_X1 U13712 ( .A1(n11149), .A2(n11148), .A3(n11147), .ZN(P2_U3227) );
  AND2_X1 U13713 ( .A1(n11151), .A2(n11150), .ZN(n11154) );
  OAI211_X1 U13714 ( .C1(n11154), .C2(n11153), .A(n15217), .B(n11152), .ZN(
        n11161) );
  NAND2_X1 U13715 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14240)
         );
  OAI211_X1 U13716 ( .C1(n11157), .C2(n11156), .A(n15210), .B(n11155), .ZN(
        n11158) );
  NAND2_X1 U13717 ( .A1(n14240), .A2(n11158), .ZN(n11159) );
  AOI21_X1 U13718 ( .B1(n14653), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11159), 
        .ZN(n11160) );
  OAI211_X1 U13719 ( .C1(n15221), .C2(n11162), .A(n11161), .B(n11160), .ZN(
        P1_U3256) );
  NAND2_X1 U13720 ( .A1(n11176), .A2(n12458), .ZN(n11180) );
  NAND2_X1 U13721 ( .A1(n11163), .A2(n11180), .ZN(n11426) );
  XNOR2_X1 U13722 ( .A(n11426), .B(n11181), .ZN(n11170) );
  INV_X1 U13723 ( .A(n11418), .ZN(n11168) );
  AOI22_X1 U13724 ( .A1(n12427), .A2(n12458), .B1(n12414), .B2(n6932), .ZN(
        n11166) );
  OAI211_X1 U13725 ( .C1(n11353), .C2(n12429), .A(n11166), .B(n11165), .ZN(
        n11167) );
  AOI21_X1 U13726 ( .B1(n11168), .B2(n12441), .A(n11167), .ZN(n11169) );
  OAI21_X1 U13727 ( .B1(n11170), .B2(n12434), .A(n11169), .ZN(P3_U3153) );
  INV_X1 U13728 ( .A(n11171), .ZN(n11173) );
  OAI222_X1 U13729 ( .A1(n7145), .A2(P1_U3086), .B1(n15147), .B2(n11173), .C1(
        n15608), .C2(n15144), .ZN(P1_U3337) );
  INV_X1 U13730 ( .A(n13422), .ZN(n13403) );
  OAI222_X1 U13731 ( .A1(n13403), .A2(P2_U3088), .B1(n13913), .B2(n11173), 
        .C1(n11172), .C2(n13916), .ZN(P2_U3309) );
  XNOR2_X1 U13732 ( .A(n11570), .B(n12293), .ZN(n11304) );
  XNOR2_X1 U13733 ( .A(n11304), .B(n11365), .ZN(n11191) );
  XNOR2_X1 U13734 ( .A(n12293), .B(n11436), .ZN(n11182) );
  XNOR2_X1 U13735 ( .A(n11182), .B(n11353), .ZN(n11427) );
  NOR2_X1 U13736 ( .A1(n11427), .A2(n11177), .ZN(n11178) );
  NAND2_X1 U13737 ( .A1(n11179), .A2(n11178), .ZN(n11187) );
  OAI21_X1 U13738 ( .B1(n11427), .B2(n11180), .A(n11181), .ZN(n11185) );
  INV_X1 U13739 ( .A(n11181), .ZN(n11425) );
  OAI21_X1 U13740 ( .B1(n11427), .B2(n6933), .A(n11425), .ZN(n11184) );
  INV_X1 U13741 ( .A(n11182), .ZN(n11183) );
  AOI22_X1 U13742 ( .A1(n11185), .A2(n11184), .B1(n11183), .B2(n12456), .ZN(
        n11186) );
  INV_X1 U13743 ( .A(n11308), .ZN(n11189) );
  AOI21_X1 U13744 ( .B1(n11191), .B2(n6621), .A(n11189), .ZN(n11197) );
  INV_X1 U13745 ( .A(n11192), .ZN(n11523) );
  AND2_X1 U13746 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11483) );
  NOR2_X1 U13747 ( .A1(n12443), .A2(n11353), .ZN(n11193) );
  AOI211_X1 U13748 ( .C1(n12445), .C2(n12455), .A(n11483), .B(n11193), .ZN(
        n11194) );
  OAI21_X1 U13749 ( .B1(n12448), .B2(n11570), .A(n11194), .ZN(n11195) );
  AOI21_X1 U13750 ( .B1(n11523), .B2(n12441), .A(n11195), .ZN(n11196) );
  OAI21_X1 U13751 ( .B1(n11197), .B2(n12434), .A(n11196), .ZN(P3_U3171) );
  INV_X1 U13752 ( .A(n11198), .ZN(n11200) );
  INV_X1 U13753 ( .A(n14969), .ZN(n11330) );
  OR2_X2 U13754 ( .A1(n15269), .A2(n11201), .ZN(n15262) );
  INV_X1 U13755 ( .A(n15236), .ZN(n15258) );
  AOI22_X1 U13756 ( .A1(n15266), .A2(n11202), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n15258), .ZN(n11203) );
  OAI21_X1 U13757 ( .B1(n11204), .B2(n15262), .A(n11203), .ZN(n11205) );
  AOI21_X1 U13758 ( .B1(n11330), .B2(n14580), .A(n11205), .ZN(n11209) );
  MUX2_X1 U13759 ( .A(n11207), .B(n11206), .S(n14798), .Z(n11208) );
  OAI211_X1 U13760 ( .C1(n11210), .C2(n14978), .A(n11209), .B(n11208), .ZN(
        P1_U3292) );
  XNOR2_X1 U13761 ( .A(n13133), .B(n6425), .ZN(n11219) );
  NAND2_X1 U13762 ( .A1(n13350), .A2(n13542), .ZN(n11218) );
  XNOR2_X1 U13763 ( .A(n11219), .B(n11218), .ZN(n11220) );
  INV_X1 U13764 ( .A(n11211), .ZN(n11212) );
  XOR2_X1 U13765 ( .A(n11221), .B(n11220), .Z(n11214) );
  NAND2_X1 U13766 ( .A1(n11214), .A2(n13042), .ZN(n11217) );
  NOR2_X1 U13767 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9566), .ZN(n15350) );
  OAI22_X1 U13768 ( .A1(n12994), .A2(n11240), .B1(n11239), .B2(n13081), .ZN(
        n11215) );
  AOI211_X1 U13769 ( .C1(n13133), .C2(n13087), .A(n15350), .B(n11215), .ZN(
        n11216) );
  OAI211_X1 U13770 ( .C1(n13085), .C2(n11250), .A(n11217), .B(n11216), .ZN(
        P2_U3211) );
  XNOR2_X1 U13771 ( .A(n13136), .B(n7171), .ZN(n11390) );
  NAND2_X1 U13772 ( .A1(n13349), .A2(n13542), .ZN(n11389) );
  XNOR2_X1 U13773 ( .A(n11390), .B(n11389), .ZN(n11392) );
  XNOR2_X1 U13774 ( .A(n11393), .B(n11392), .ZN(n11228) );
  INV_X1 U13775 ( .A(n11222), .ZN(n11459) );
  NAND2_X1 U13776 ( .A1(n13348), .A2(n13723), .ZN(n11224) );
  NAND2_X1 U13777 ( .A1(n13350), .A2(n13722), .ZN(n11223) );
  AND2_X1 U13778 ( .A1(n11224), .A2(n11223), .ZN(n11299) );
  NAND2_X1 U13779 ( .A1(n13087), .A2(n13136), .ZN(n11225) );
  NAND2_X1 U13780 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15367) );
  OAI211_X1 U13781 ( .C1(n11299), .C2(n13074), .A(n11225), .B(n15367), .ZN(
        n11226) );
  AOI21_X1 U13782 ( .B1(n13072), .B2(n11459), .A(n11226), .ZN(n11227) );
  OAI21_X1 U13783 ( .B1(n11228), .B2(n13089), .A(n11227), .ZN(P2_U3185) );
  AOI22_X1 U13784 ( .A1(n11229), .A2(n15266), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n15258), .ZN(n11230) );
  OAI21_X1 U13785 ( .B1(n8756), .B2(n15262), .A(n11230), .ZN(n11233) );
  MUX2_X1 U13786 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n11231), .S(n14798), .Z(
        n11232) );
  INV_X1 U13787 ( .A(n9734), .ZN(n11236) );
  OAI222_X1 U13788 ( .A1(n13666), .A2(P2_U3088), .B1(n13913), .B2(n11236), 
        .C1(n11234), .C2(n13916), .ZN(P2_U3308) );
  OAI222_X1 U13789 ( .A1(n14934), .A2(P1_U3086), .B1(n15147), .B2(n11236), 
        .C1(n11235), .C2(n15144), .ZN(P1_U3336) );
  OAI21_X1 U13790 ( .B1(n11238), .B2(n11242), .A(n11237), .ZN(n15444) );
  INV_X1 U13791 ( .A(n15444), .ZN(n11254) );
  OAI22_X1 U13792 ( .A1(n11240), .A2(n13676), .B1(n11239), .B2(n13678), .ZN(
        n11246) );
  NAND3_X1 U13793 ( .A1(n11058), .A2(n11242), .A3(n11241), .ZN(n11243) );
  AOI21_X1 U13794 ( .B1(n11244), .B2(n11243), .A(n13701), .ZN(n11245) );
  AOI211_X1 U13795 ( .C1(n11247), .C2(n15444), .A(n11246), .B(n11245), .ZN(
        n15441) );
  MUX2_X1 U13796 ( .A(n11248), .B(n15441), .S(n13687), .Z(n11253) );
  OAI211_X1 U13797 ( .C1(n11249), .C2(n15440), .A(n11296), .B(n13840), .ZN(
        n15438) );
  OAI22_X1 U13798 ( .A1(n13549), .A2(n15438), .B1(n11250), .B2(n13683), .ZN(
        n11251) );
  AOI21_X1 U13799 ( .B1(n13649), .B2(n13133), .A(n11251), .ZN(n11252) );
  OAI211_X1 U13800 ( .C1(n11254), .C2(n11256), .A(n11253), .B(n11252), .ZN(
        P2_U3259) );
  OAI22_X1 U13801 ( .A1(n11257), .A2(n13735), .B1(n11256), .B2(n11255), .ZN(
        n11262) );
  INV_X1 U13802 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13356) );
  OAI22_X1 U13803 ( .A1(n11258), .A2(n6402), .B1(n13356), .B2(n13683), .ZN(
        n11261) );
  OAI22_X1 U13804 ( .A1(n13549), .A2(n11259), .B1(n13687), .B2(n10100), .ZN(
        n11260) );
  OR3_X1 U13805 ( .A1(n11262), .A2(n11261), .A3(n11260), .ZN(P2_U3264) );
  INV_X1 U13806 ( .A(n11263), .ZN(n11266) );
  OAI22_X1 U13807 ( .A1(n11264), .A2(P3_U3151), .B1(SI_22_), .B2(n12941), .ZN(
        n11265) );
  AOI21_X1 U13808 ( .B1(n11266), .B2(n12929), .A(n11265), .ZN(P3_U3273) );
  INV_X1 U13809 ( .A(n11267), .ZN(n15445) );
  INV_X1 U13810 ( .A(n11268), .ZN(n11269) );
  AOI211_X1 U13811 ( .C1(n15445), .C2(n11271), .A(n11270), .B(n11269), .ZN(
        n11277) );
  AOI22_X1 U13812 ( .A1(n13789), .A2(n13129), .B1(n15452), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n11272) );
  OAI21_X1 U13813 ( .B1(n11277), .B2(n15452), .A(n11272), .ZN(P2_U3504) );
  INV_X1 U13814 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11273) );
  OAI22_X1 U13815 ( .A1(n13900), .A2(n11274), .B1(n15448), .B2(n11273), .ZN(
        n11275) );
  INV_X1 U13816 ( .A(n11275), .ZN(n11276) );
  OAI21_X1 U13817 ( .B1(n11277), .B2(n15446), .A(n11276), .ZN(P2_U3445) );
  XNOR2_X1 U13818 ( .A(n11278), .B(n11281), .ZN(n15505) );
  INV_X1 U13819 ( .A(n15505), .ZN(n11293) );
  INV_X1 U13820 ( .A(n11279), .ZN(n11280) );
  NAND2_X1 U13821 ( .A1(n15472), .A2(n11280), .ZN(n15487) );
  INV_X1 U13822 ( .A(n11281), .ZN(n11282) );
  XNOR2_X1 U13823 ( .A(n11283), .B(n11282), .ZN(n11286) );
  INV_X1 U13824 ( .A(n11357), .ZN(n15478) );
  NAND2_X1 U13825 ( .A1(n15505), .A2(n15478), .ZN(n11285) );
  AOI22_X1 U13826 ( .A1(n11365), .A2(n15479), .B1(n12704), .B2(n12457), .ZN(
        n11284) );
  OAI211_X1 U13827 ( .C1(n15484), .C2(n11286), .A(n11285), .B(n11284), .ZN(
        n15508) );
  MUX2_X1 U13828 ( .A(n15508), .B(P3_REG2_REG_8__SCAN_IN), .S(n15493), .Z(
        n11287) );
  INV_X1 U13829 ( .A(n11287), .ZN(n11292) );
  INV_X1 U13830 ( .A(n11432), .ZN(n11290) );
  NAND2_X1 U13831 ( .A1(n11436), .A2(n12829), .ZN(n15503) );
  NOR3_X1 U13832 ( .A1(n11288), .A2(n15462), .A3(n15503), .ZN(n11289) );
  AOI21_X1 U13833 ( .B1(n15488), .B2(n11290), .A(n11289), .ZN(n11291) );
  OAI211_X1 U13834 ( .C1(n11293), .C2(n15487), .A(n11292), .B(n11291), .ZN(
        P3_U3225) );
  OAI21_X1 U13835 ( .B1(n11294), .B2(n11297), .A(n11573), .ZN(n11466) );
  INV_X1 U13836 ( .A(n11577), .ZN(n11295) );
  AOI211_X1 U13837 ( .C1(n13136), .C2(n11296), .A(n13542), .B(n11295), .ZN(
        n11460) );
  XNOR2_X1 U13838 ( .A(n11298), .B(n11297), .ZN(n11300) );
  OAI21_X1 U13839 ( .B1(n11300), .B2(n13701), .A(n11299), .ZN(n11463) );
  AOI211_X1 U13840 ( .C1(n13835), .C2(n11466), .A(n11460), .B(n11463), .ZN(
        n11303) );
  AOI22_X1 U13841 ( .A1(n13881), .A2(n13136), .B1(P2_REG0_REG_7__SCAN_IN), 
        .B2(n15446), .ZN(n11301) );
  OAI21_X1 U13842 ( .B1(n11303), .B2(n15446), .A(n11301), .ZN(P2_U3451) );
  AOI22_X1 U13843 ( .A1(n13789), .A2(n13136), .B1(P2_REG1_REG_7__SCAN_IN), 
        .B2(n15452), .ZN(n11302) );
  OAI21_X1 U13844 ( .B1(n11303), .B2(n15452), .A(n11302), .ZN(P2_U3506) );
  INV_X1 U13845 ( .A(n11304), .ZN(n11305) );
  NAND2_X1 U13846 ( .A1(n11305), .A2(n11431), .ZN(n11306) );
  AND2_X1 U13847 ( .A1(n11308), .A2(n11306), .ZN(n11310) );
  XNOR2_X1 U13848 ( .A(n11677), .B(n12293), .ZN(n11717) );
  XNOR2_X1 U13849 ( .A(n11717), .B(n11352), .ZN(n11309) );
  AND2_X1 U13850 ( .A1(n11309), .A2(n11306), .ZN(n11307) );
  OAI211_X1 U13851 ( .C1(n11310), .C2(n11309), .A(n12439), .B(n11718), .ZN(
        n11315) );
  INV_X1 U13852 ( .A(n11617), .ZN(n11313) );
  AND2_X1 U13853 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11540) );
  AOI21_X1 U13854 ( .B1(n12427), .B2(n11365), .A(n11540), .ZN(n11311) );
  OAI21_X1 U13855 ( .B1(n11908), .B2(n12429), .A(n11311), .ZN(n11312) );
  AOI21_X1 U13856 ( .B1(n11313), .B2(n12441), .A(n11312), .ZN(n11314) );
  OAI211_X1 U13857 ( .C1(n12448), .C2(n11677), .A(n11315), .B(n11314), .ZN(
        P3_U3157) );
  NAND2_X1 U13858 ( .A1(n11317), .A2(n11316), .ZN(n15248) );
  XNOR2_X1 U13859 ( .A(n15250), .B(n15285), .ZN(n14532) );
  XNOR2_X1 U13860 ( .A(n15248), .B(n14532), .ZN(n15288) );
  XNOR2_X1 U13861 ( .A(n11318), .B(n14532), .ZN(n11319) );
  NAND2_X1 U13862 ( .A1(n11319), .A2(n15308), .ZN(n15286) );
  MUX2_X1 U13863 ( .A(n15286), .B(n11320), .S(n15260), .Z(n11326) );
  INV_X1 U13864 ( .A(n15265), .ZN(n11321) );
  AOI211_X1 U13865 ( .C1(n15285), .C2(n11505), .A(n10283), .B(n11321), .ZN(
        n15283) );
  OAI22_X1 U13866 ( .A1(n15262), .A2(n15246), .B1(n11322), .B2(n15236), .ZN(
        n11324) );
  OR2_X1 U13867 ( .A1(n15269), .A2(n15312), .ZN(n14696) );
  OAI22_X1 U13868 ( .A1(n15281), .A2(n14969), .B1(n14696), .B2(n15282), .ZN(
        n11323) );
  AOI211_X1 U13869 ( .C1(n15283), .C2(n15266), .A(n11324), .B(n11323), .ZN(
        n11325) );
  OAI211_X1 U13870 ( .C1(n14978), .C2(n15288), .A(n11326), .B(n11325), .ZN(
        P1_U3289) );
  AOI21_X1 U13871 ( .B1(n15240), .B2(n15266), .A(n14971), .ZN(n11334) );
  OAI22_X1 U13872 ( .A1(n14798), .A2(n11328), .B1(n11327), .B2(n15236), .ZN(
        n11329) );
  AOI21_X1 U13873 ( .B1(n11330), .B2(n9228), .A(n11329), .ZN(n11332) );
  OAI21_X1 U13874 ( .B1(n14879), .B2(n14903), .A(n14525), .ZN(n11331) );
  OAI211_X1 U13875 ( .C1(n11334), .C2(n11333), .A(n11332), .B(n11331), .ZN(
        P1_U3293) );
  OAI21_X1 U13876 ( .B1(n15264), .B2(n15298), .A(n15240), .ZN(n11335) );
  NOR2_X1 U13877 ( .A1(n11335), .A2(n15241), .ZN(n15296) );
  OAI22_X1 U13878 ( .A1(n15262), .A2(n15298), .B1(n11454), .B2(n15236), .ZN(
        n11336) );
  AOI21_X1 U13879 ( .B1(n15296), .B2(n15266), .A(n11336), .ZN(n11346) );
  INV_X1 U13880 ( .A(n14530), .ZN(n11339) );
  XNOR2_X1 U13881 ( .A(n11337), .B(n11339), .ZN(n11343) );
  XNOR2_X1 U13882 ( .A(n11338), .B(n11339), .ZN(n11340) );
  NAND2_X1 U13883 ( .A1(n11340), .A2(n15308), .ZN(n11342) );
  AOI22_X1 U13884 ( .A1(n14576), .A2(n15090), .B1(n15107), .B2(n14578), .ZN(
        n11341) );
  OAI211_X1 U13885 ( .C1(n11343), .C2(n15289), .A(n11342), .B(n11341), .ZN(
        n15299) );
  MUX2_X1 U13886 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n15299), .S(n14798), .Z(
        n11344) );
  INV_X1 U13887 ( .A(n11344), .ZN(n11345) );
  NAND2_X1 U13888 ( .A1(n11346), .A2(n11345), .ZN(P1_U3287) );
  INV_X1 U13889 ( .A(n11347), .ZN(n15504) );
  XNOR2_X1 U13890 ( .A(n11348), .B(n11349), .ZN(n11527) );
  INV_X1 U13891 ( .A(n11527), .ZN(n11358) );
  XNOR2_X1 U13892 ( .A(n11350), .B(n11351), .ZN(n11355) );
  OAI22_X1 U13893 ( .A1(n11353), .A2(n15467), .B1(n11352), .B2(n15469), .ZN(
        n11354) );
  AOI21_X1 U13894 ( .B1(n11355), .B2(n12784), .A(n11354), .ZN(n11356) );
  OAI21_X1 U13895 ( .B1(n11527), .B2(n11357), .A(n11356), .ZN(n11520) );
  AOI21_X1 U13896 ( .B1(n15504), .B2(n11358), .A(n11520), .ZN(n11567) );
  INV_X1 U13897 ( .A(n11570), .ZN(n11524) );
  AOI22_X1 U13898 ( .A1(n12915), .A2(n11524), .B1(n15509), .B2(
        P3_REG0_REG_9__SCAN_IN), .ZN(n11359) );
  OAI21_X1 U13899 ( .B1(n11567), .B2(n15509), .A(n11359), .ZN(P3_U3417) );
  INV_X1 U13900 ( .A(n11360), .ZN(n11361) );
  OAI222_X1 U13901 ( .A1(n12941), .A2(n11363), .B1(P3_U3151), .B2(n11362), 
        .C1(n12948), .C2(n11361), .ZN(P3_U3275) );
  XNOR2_X1 U13902 ( .A(n11364), .B(n11367), .ZN(n11366) );
  AOI222_X1 U13903 ( .A1(n12784), .A2(n11366), .B1(n11955), .B2(n15479), .C1(
        n11365), .C2(n12704), .ZN(n11672) );
  XNOR2_X1 U13904 ( .A(n11368), .B(n11367), .ZN(n11674) );
  INV_X1 U13905 ( .A(n12919), .ZN(n12909) );
  OAI22_X1 U13906 ( .A1(n12894), .A2(n11677), .B1(n15510), .B2(n11369), .ZN(
        n11370) );
  AOI21_X1 U13907 ( .B1(n11674), .B2(n12909), .A(n11370), .ZN(n11371) );
  OAI21_X1 U13908 ( .B1(n11672), .B2(n15509), .A(n11371), .ZN(P3_U3420) );
  INV_X1 U13909 ( .A(n11372), .ZN(n11373) );
  OAI222_X1 U13910 ( .A1(P2_U3088), .A2(n6398), .B1(n13916), .B2(n15584), .C1(
        n13913), .C2(n11373), .ZN(P2_U3307) );
  OAI222_X1 U13911 ( .A1(P1_U3086), .A2(n11375), .B1(n15144), .B2(n11374), 
        .C1(n15147), .C2(n11373), .ZN(P1_U3335) );
  XNOR2_X1 U13912 ( .A(n11376), .B(n14524), .ZN(n15322) );
  INV_X1 U13913 ( .A(n15322), .ZN(n11388) );
  NAND2_X1 U13914 ( .A1(n11378), .A2(n14524), .ZN(n15309) );
  NAND3_X1 U13915 ( .A1(n11377), .A2(n15309), .A3(n14879), .ZN(n11387) );
  NAND2_X1 U13916 ( .A1(n14964), .A2(n14576), .ZN(n11381) );
  INV_X1 U13917 ( .A(n11379), .ZN(n11829) );
  AOI22_X1 U13918 ( .A1(n15260), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n11829), 
        .B2(n15258), .ZN(n11380) );
  OAI211_X1 U13919 ( .C1(n15311), .C2(n14969), .A(n11381), .B(n11380), .ZN(
        n11385) );
  AOI21_X1 U13920 ( .B1(n11382), .B2(n15316), .A(n10283), .ZN(n11383) );
  NAND2_X1 U13921 ( .A1(n11383), .A2(n11646), .ZN(n15317) );
  NOR2_X1 U13922 ( .A1(n15317), .A2(n14974), .ZN(n11384) );
  AOI211_X1 U13923 ( .C1(n14971), .C2(n15316), .A(n11385), .B(n11384), .ZN(
        n11386) );
  OAI211_X1 U13924 ( .C1(n11388), .C2(n14978), .A(n11387), .B(n11386), .ZN(
        P1_U3285) );
  INV_X1 U13925 ( .A(n11389), .ZN(n11391) );
  AND2_X1 U13926 ( .A1(n13348), .A2(n13542), .ZN(n11395) );
  XNOR2_X1 U13927 ( .A(n13145), .B(n7171), .ZN(n11394) );
  NOR2_X1 U13928 ( .A1(n11394), .A2(n11395), .ZN(n11658) );
  AOI21_X1 U13929 ( .B1(n11395), .B2(n11394), .A(n11658), .ZN(n11396) );
  OAI21_X1 U13930 ( .B1(n11397), .B2(n11396), .A(n11660), .ZN(n11398) );
  NAND2_X1 U13931 ( .A1(n11398), .A2(n13042), .ZN(n11404) );
  NAND2_X1 U13932 ( .A1(n13347), .A2(n13723), .ZN(n11400) );
  NAND2_X1 U13933 ( .A1(n13349), .A2(n13722), .ZN(n11399) );
  AND2_X1 U13934 ( .A1(n11400), .A2(n11399), .ZN(n11586) );
  OAI21_X1 U13935 ( .B1(n13074), .B2(n11586), .A(n11401), .ZN(n11402) );
  AOI21_X1 U13936 ( .B1(n13145), .B2(n13087), .A(n11402), .ZN(n11403) );
  OAI211_X1 U13937 ( .C1(n13085), .C2(n11580), .A(n11404), .B(n11403), .ZN(
        P2_U3193) );
  OAI22_X1 U13938 ( .A1(n12726), .A2(n11406), .B1(n11405), .B2(n15460), .ZN(
        n11409) );
  MUX2_X1 U13939 ( .A(n11407), .B(P3_REG2_REG_4__SCAN_IN), .S(n15493), .Z(
        n11408) );
  AOI211_X1 U13940 ( .C1(n12741), .C2(n11410), .A(n11409), .B(n11408), .ZN(
        n11411) );
  INV_X1 U13941 ( .A(n11411), .ZN(P3_U3229) );
  OAI22_X1 U13942 ( .A1(n12726), .A2(n11412), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15460), .ZN(n11415) );
  MUX2_X1 U13943 ( .A(n11413), .B(P3_REG2_REG_3__SCAN_IN), .S(n15493), .Z(
        n11414) );
  AOI211_X1 U13944 ( .C1(n12741), .C2(n11416), .A(n11415), .B(n11414), .ZN(
        n11417) );
  INV_X1 U13945 ( .A(n11417), .ZN(P3_U3230) );
  OAI22_X1 U13946 ( .A1(n12726), .A2(n11419), .B1(n11418), .B2(n15460), .ZN(
        n11422) );
  MUX2_X1 U13947 ( .A(n11420), .B(P3_REG2_REG_7__SCAN_IN), .S(n15493), .Z(
        n11421) );
  AOI211_X1 U13948 ( .C1(n12741), .C2(n11423), .A(n11422), .B(n11421), .ZN(
        n11424) );
  INV_X1 U13949 ( .A(n11424), .ZN(P3_U3226) );
  MUX2_X1 U13950 ( .A(n11426), .B(n12457), .S(n11425), .Z(n11428) );
  XOR2_X1 U13951 ( .A(n11428), .B(n11427), .Z(n11438) );
  AOI21_X1 U13952 ( .B1(n12427), .B2(n12457), .A(n11429), .ZN(n11430) );
  OAI21_X1 U13953 ( .B1(n11431), .B2(n12429), .A(n11430), .ZN(n11435) );
  NOR2_X1 U13954 ( .A1(n11433), .A2(n11432), .ZN(n11434) );
  AOI211_X1 U13955 ( .C1(n11436), .C2(n12414), .A(n11435), .B(n11434), .ZN(
        n11437) );
  OAI21_X1 U13956 ( .B1(n11438), .B2(n12434), .A(n11437), .ZN(P3_U3161) );
  AND2_X1 U13957 ( .A1(n11440), .A2(n11439), .ZN(n11444) );
  INV_X1 U13958 ( .A(n11440), .ZN(n11442) );
  NAND2_X1 U13959 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  NAND2_X1 U13960 ( .A1(n14578), .A2(n14108), .ZN(n11447) );
  NAND2_X1 U13961 ( .A1(n6407), .A2(n10286), .ZN(n11446) );
  NAND2_X1 U13962 ( .A1(n11447), .A2(n11446), .ZN(n14177) );
  OAI22_X1 U13963 ( .A1(n15281), .A2(n14020), .B1(n6406), .B2(n14011), .ZN(
        n11448) );
  XNOR2_X1 U13964 ( .A(n11448), .B(n14111), .ZN(n14178) );
  INV_X1 U13965 ( .A(n14177), .ZN(n11449) );
  NAND2_X1 U13966 ( .A1(n14577), .A2(n10286), .ZN(n11451) );
  OAI21_X1 U13967 ( .B1(n15298), .B2(n14011), .A(n11451), .ZN(n11452) );
  XNOR2_X1 U13968 ( .A(n11452), .B(n14111), .ZN(n11813) );
  INV_X1 U13969 ( .A(n15298), .ZN(n14339) );
  AOI22_X1 U13970 ( .A1(n14339), .A2(n10286), .B1(n14577), .B2(n14108), .ZN(
        n11811) );
  XNOR2_X1 U13971 ( .A(n11813), .B(n11811), .ZN(n11814) );
  XNOR2_X1 U13972 ( .A(n11815), .B(n11814), .ZN(n11458) );
  OAI21_X1 U13973 ( .B1(n14286), .B2(n11454), .A(n11453), .ZN(n11456) );
  OAI22_X1 U13974 ( .A1(n15313), .A2(n14272), .B1(n14227), .B2(n15281), .ZN(
        n11455) );
  AOI211_X1 U13975 ( .C1(n14339), .C2(n14300), .A(n11456), .B(n11455), .ZN(
        n11457) );
  OAI21_X1 U13976 ( .B1(n11458), .B2(n14302), .A(n11457), .ZN(P1_U3239) );
  AOI22_X1 U13977 ( .A1(n11460), .A2(n13708), .B1(n11459), .B2(n13731), .ZN(
        n11461) );
  OAI21_X1 U13978 ( .B1(n11462), .B2(n13735), .A(n11461), .ZN(n11465) );
  MUX2_X1 U13979 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11463), .S(n13687), .Z(
        n11464) );
  AOI211_X1 U13980 ( .C1(n13714), .C2(n11466), .A(n11465), .B(n11464), .ZN(
        n11467) );
  INV_X1 U13981 ( .A(n11467), .ZN(P2_U3258) );
  XNOR2_X1 U13982 ( .A(n11528), .B(P3_REG1_REG_9__SCAN_IN), .ZN(n11490) );
  INV_X1 U13983 ( .A(n11468), .ZN(n11469) );
  INV_X1 U13984 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11522) );
  MUX2_X1 U13985 ( .A(n11522), .B(n11568), .S(n12937), .Z(n11475) );
  INV_X1 U13986 ( .A(n11475), .ZN(n11474) );
  AND2_X1 U13987 ( .A1(n11486), .A2(n11474), .ZN(n11531) );
  INV_X1 U13988 ( .A(n11531), .ZN(n11476) );
  NAND2_X1 U13989 ( .A1(n11529), .A2(n11475), .ZN(n11532) );
  NAND2_X1 U13990 ( .A1(n11476), .A2(n11532), .ZN(n11477) );
  XNOR2_X1 U13991 ( .A(n11533), .B(n11477), .ZN(n11488) );
  OAI21_X1 U13992 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11481), .A(n11538), .ZN(
        n11482) );
  NAND2_X1 U13993 ( .A1(n11482), .A2(n12590), .ZN(n11485) );
  AOI21_X1 U13994 ( .B1(n15455), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11483), .ZN(
        n11484) );
  OAI211_X1 U13995 ( .C1(n12597), .C2(n11486), .A(n11485), .B(n11484), .ZN(
        n11487) );
  AOI21_X1 U13996 ( .B1(n12491), .B2(n11488), .A(n11487), .ZN(n11489) );
  OAI21_X1 U13997 ( .B1(n11490), .B2(n12024), .A(n11489), .ZN(P3_U3191) );
  INV_X1 U13998 ( .A(n11494), .ZN(n11493) );
  OR2_X1 U13999 ( .A1(n11491), .A2(P2_U3088), .ZN(n13334) );
  NAND2_X1 U14000 ( .A1(n13910), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11492) );
  OAI211_X1 U14001 ( .C1(n11493), .C2(n13913), .A(n13334), .B(n11492), .ZN(
        P2_U3304) );
  NAND2_X1 U14002 ( .A1(n11494), .A2(n15139), .ZN(n11495) );
  OAI211_X1 U14003 ( .C1(n11496), .C2(n15144), .A(n11495), .B(n14561), .ZN(
        P1_U3332) );
  INV_X1 U14004 ( .A(n11497), .ZN(n11500) );
  OAI222_X1 U14005 ( .A1(n14307), .A2(P1_U3086), .B1(n15147), .B2(n11500), 
        .C1(n11498), .C2(n15144), .ZN(P1_U3334) );
  OAI222_X1 U14006 ( .A1(n13104), .A2(P2_U3088), .B1(n13913), .B2(n11500), 
        .C1(n11499), .C2(n13916), .ZN(P2_U3306) );
  XNOR2_X1 U14007 ( .A(n11501), .B(n14526), .ZN(n15276) );
  INV_X1 U14008 ( .A(n11502), .ZN(n11504) );
  INV_X1 U14009 ( .A(n14526), .ZN(n14323) );
  AOI21_X1 U14010 ( .B1(n11504), .B2(n14323), .A(n11503), .ZN(n15278) );
  INV_X1 U14011 ( .A(n15278), .ZN(n11514) );
  OAI211_X1 U14012 ( .C1(n11506), .C2(n15275), .A(n11505), .B(n15240), .ZN(
        n15274) );
  INV_X1 U14013 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14014 ( .A1(n14971), .A2(n14094), .B1(n11507), .B2(n15258), .ZN(
        n11512) );
  NAND2_X1 U14015 ( .A1(n14580), .A2(n15107), .ZN(n11509) );
  NAND2_X1 U14016 ( .A1(n15250), .A2(n15090), .ZN(n11508) );
  NAND2_X1 U14017 ( .A1(n11509), .A2(n11508), .ZN(n14095) );
  INV_X1 U14018 ( .A(n14095), .ZN(n15273) );
  MUX2_X1 U14019 ( .A(n15273), .B(n11510), .S(n15260), .Z(n11511) );
  OAI211_X1 U14020 ( .C1(n15274), .C2(n14974), .A(n11512), .B(n11511), .ZN(
        n11513) );
  AOI21_X1 U14021 ( .B1(n11514), .B2(n14903), .A(n11513), .ZN(n11515) );
  OAI21_X1 U14022 ( .B1(n14906), .B2(n15276), .A(n11515), .ZN(P1_U3290) );
  NAND2_X1 U14023 ( .A1(n11516), .A2(n12929), .ZN(n11518) );
  OAI211_X1 U14024 ( .C1(n11519), .C2(n12941), .A(n11518), .B(n11517), .ZN(
        P3_U3272) );
  INV_X1 U14025 ( .A(n11520), .ZN(n11521) );
  MUX2_X1 U14026 ( .A(n11522), .B(n11521), .S(n15472), .Z(n11526) );
  AOI22_X1 U14027 ( .A1(n12787), .A2(n11524), .B1(n15488), .B2(n11523), .ZN(
        n11525) );
  OAI211_X1 U14028 ( .C1(n11527), .C2(n15487), .A(n11526), .B(n11525), .ZN(
        P3_U3224) );
  XOR2_X1 U14029 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11917), .Z(n11914) );
  XOR2_X1 U14030 ( .A(n11914), .B(n11915), .Z(n11546) );
  MUX2_X1 U14031 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12937), .Z(n11530) );
  NOR2_X1 U14032 ( .A1(n11530), .A2(n11917), .ZN(n11920) );
  AOI21_X1 U14033 ( .B1(n11530), .B2(n11917), .A(n11920), .ZN(n11535) );
  AOI21_X1 U14034 ( .B1(n11533), .B2(n11532), .A(n11531), .ZN(n11534) );
  NAND2_X1 U14035 ( .A1(n11534), .A2(n11535), .ZN(n11922) );
  OAI21_X1 U14036 ( .B1(n11535), .B2(n11534), .A(n11922), .ZN(n11544) );
  XNOR2_X1 U14037 ( .A(n11917), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11537) );
  AND3_X1 U14038 ( .A1(n11538), .A2(n11537), .A3(n6941), .ZN(n11539) );
  OAI21_X1 U14039 ( .B1(n11916), .B2(n11539), .A(n12590), .ZN(n11542) );
  AOI21_X1 U14040 ( .B1(n15455), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11540), 
        .ZN(n11541) );
  OAI211_X1 U14041 ( .C1(n12597), .C2(n11917), .A(n11542), .B(n11541), .ZN(
        n11543) );
  AOI21_X1 U14042 ( .B1(n12491), .B2(n11544), .A(n11543), .ZN(n11545) );
  OAI21_X1 U14043 ( .B1(n11546), .B2(n12024), .A(n11545), .ZN(P3_U3192) );
  NAND2_X1 U14044 ( .A1(n11547), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U14045 ( .A1(n11550), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11553) );
  OR2_X1 U14046 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n11551), .ZN(n11552) );
  NAND2_X1 U14047 ( .A1(n11554), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11560) );
  INV_X1 U14048 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11555) );
  NAND2_X1 U14049 ( .A1(n11555), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n11556) );
  AND2_X1 U14050 ( .A1(n11560), .A2(n11556), .ZN(n11558) );
  INV_X1 U14051 ( .A(n11558), .ZN(n11557) );
  XNOR2_X1 U14052 ( .A(n11559), .B(n11557), .ZN(n15159) );
  INV_X1 U14053 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14054 ( .A1(n11561), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n11714) );
  INV_X1 U14055 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n12010) );
  NAND2_X1 U14056 ( .A1(n12010), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11562) );
  AND2_X1 U14057 ( .A1(n11714), .A2(n11562), .ZN(n11712) );
  XNOR2_X1 U14058 ( .A(n11713), .B(n11712), .ZN(n11707) );
  INV_X1 U14059 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n11705) );
  XNOR2_X1 U14060 ( .A(n11706), .B(n11705), .ZN(SUB_1596_U68) );
  INV_X1 U14061 ( .A(n11563), .ZN(n11565) );
  OAI222_X1 U14062 ( .A1(n12941), .A2(n11566), .B1(n12948), .B2(n11565), .C1(
        n11564), .C2(P3_U3151), .ZN(P3_U3274) );
  MUX2_X1 U14063 ( .A(n11568), .B(n11567), .S(n15514), .Z(n11569) );
  OAI21_X1 U14064 ( .B1(n12821), .B2(n11570), .A(n11569), .ZN(P3_U3468) );
  INV_X1 U14065 ( .A(n11571), .ZN(n11572) );
  NAND2_X1 U14066 ( .A1(n11573), .A2(n11572), .ZN(n11576) );
  INV_X1 U14067 ( .A(n11576), .ZN(n11574) );
  NAND2_X1 U14068 ( .A1(n11574), .A2(n13309), .ZN(n11622) );
  INV_X1 U14069 ( .A(n11622), .ZN(n11575) );
  AOI21_X1 U14070 ( .B1(n9830), .B2(n11576), .A(n11575), .ZN(n11638) );
  INV_X1 U14071 ( .A(n11638), .ZN(n11592) );
  NAND2_X1 U14072 ( .A1(n11577), .A2(n13145), .ZN(n11578) );
  NAND2_X1 U14073 ( .A1(n11578), .A2(n13840), .ZN(n11579) );
  NOR2_X1 U14074 ( .A1(n11624), .A2(n11579), .ZN(n11637) );
  OAI22_X1 U14075 ( .A1(n13735), .A2(n11581), .B1(n13683), .B2(n11580), .ZN(
        n11582) );
  AOI21_X1 U14076 ( .B1(n13708), .B2(n11637), .A(n11582), .ZN(n11591) );
  CLKBUF_X1 U14077 ( .A(n11583), .Z(n11585) );
  OAI211_X1 U14078 ( .C1(n11585), .C2(n9830), .A(n11584), .B(n13717), .ZN(
        n11587) );
  NAND2_X1 U14079 ( .A1(n11587), .A2(n11586), .ZN(n11636) );
  INV_X1 U14080 ( .A(n11636), .ZN(n11588) );
  MUX2_X1 U14081 ( .A(n11589), .B(n11588), .S(n13687), .Z(n11590) );
  OAI211_X1 U14082 ( .C1(n11592), .C2(n13738), .A(n11591), .B(n11590), .ZN(
        P2_U3257) );
  XNOR2_X1 U14083 ( .A(n11593), .B(n8087), .ZN(n11594) );
  AOI222_X1 U14084 ( .A1(n12784), .A2(n11594), .B1(n12454), .B2(n15479), .C1(
        n12455), .C2(n12704), .ZN(n11785) );
  NAND2_X1 U14085 ( .A1(n11596), .A2(n11595), .ZN(n11597) );
  NAND2_X1 U14086 ( .A1(n11598), .A2(n11597), .ZN(n11784) );
  OAI22_X1 U14087 ( .A1(n12894), .A2(n11787), .B1(n15510), .B2(n11599), .ZN(
        n11600) );
  AOI21_X1 U14088 ( .B1(n11784), .B2(n12909), .A(n11600), .ZN(n11601) );
  OAI21_X1 U14089 ( .B1(n11785), .B2(n15509), .A(n11601), .ZN(P3_U3423) );
  NAND2_X1 U14090 ( .A1(n11608), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U14091 ( .A1(n11678), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U14092 ( .A1(n11604), .A2(n11687), .ZN(n11605) );
  XNOR2_X1 U14093 ( .A(n11883), .B(n11611), .ZN(n11882) );
  XNOR2_X1 U14094 ( .A(n11882), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n11615) );
  AOI21_X1 U14095 ( .B1(n11608), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11607), 
        .ZN(n11681) );
  XNOR2_X1 U14096 ( .A(n11687), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11680) );
  OAI22_X1 U14097 ( .A1(n11681), .A2(n11680), .B1(n11609), .B2(n13836), .ZN(
        n11886) );
  XOR2_X1 U14098 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n11888), .Z(n11613) );
  NAND2_X1 U14099 ( .A1(n15334), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14100 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13080)
         );
  OAI211_X1 U14101 ( .C1(n15395), .C2(n11611), .A(n11610), .B(n13080), .ZN(
        n11612) );
  AOI21_X1 U14102 ( .B1(n11613), .B2(n15403), .A(n11612), .ZN(n11614) );
  OAI21_X1 U14103 ( .B1(n11615), .B2(n11894), .A(n11614), .ZN(P2_U3229) );
  INV_X1 U14104 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11616) );
  MUX2_X1 U14105 ( .A(n11616), .B(n11672), .S(n15472), .Z(n11620) );
  OAI22_X1 U14106 ( .A1(n12726), .A2(n11677), .B1(n11617), .B2(n15460), .ZN(
        n11618) );
  AOI21_X1 U14107 ( .B1(n11674), .B2(n12741), .A(n11618), .ZN(n11619) );
  NAND2_X1 U14108 ( .A1(n11620), .A2(n11619), .ZN(P3_U3223) );
  NAND2_X1 U14109 ( .A1(n11622), .A2(n11621), .ZN(n11623) );
  XNOR2_X1 U14110 ( .A(n11623), .B(n13310), .ZN(n11734) );
  INV_X1 U14111 ( .A(n11734), .ZN(n11635) );
  INV_X1 U14112 ( .A(n11624), .ZN(n11625) );
  AOI211_X1 U14113 ( .C1(n13148), .C2(n11625), .A(n12272), .B(n11695), .ZN(
        n11733) );
  OAI22_X1 U14114 ( .A1(n13735), .A2(n11626), .B1(n13683), .B2(n11668), .ZN(
        n11627) );
  AOI21_X1 U14115 ( .B1(n11733), .B2(n13708), .A(n11627), .ZN(n11634) );
  OAI211_X1 U14116 ( .C1(n11629), .C2(n13310), .A(n11628), .B(n13717), .ZN(
        n11630) );
  AOI22_X1 U14117 ( .A1(n13722), .A2(n13348), .B1(n13346), .B2(n13723), .ZN(
        n11664) );
  NAND2_X1 U14118 ( .A1(n11630), .A2(n11664), .ZN(n11732) );
  INV_X1 U14119 ( .A(n11732), .ZN(n11631) );
  MUX2_X1 U14120 ( .A(n11632), .B(n11631), .S(n13687), .Z(n11633) );
  OAI211_X1 U14121 ( .C1(n11635), .C2(n13738), .A(n11634), .B(n11633), .ZN(
        P2_U3256) );
  AOI211_X1 U14122 ( .C1(n11638), .C2(n13835), .A(n11637), .B(n11636), .ZN(
        n11641) );
  AOI22_X1 U14123 ( .A1(n13881), .A2(n13145), .B1(P2_REG0_REG_8__SCAN_IN), 
        .B2(n15446), .ZN(n11639) );
  OAI21_X1 U14124 ( .B1(n11641), .B2(n15446), .A(n11639), .ZN(P2_U3454) );
  AOI22_X1 U14125 ( .A1(n13789), .A2(n13145), .B1(P2_REG1_REG_8__SCAN_IN), 
        .B2(n15452), .ZN(n11640) );
  OAI21_X1 U14126 ( .B1(n11641), .B2(n15452), .A(n11640), .ZN(P2_U3507) );
  NAND2_X1 U14127 ( .A1(n11642), .A2(n14535), .ZN(n11643) );
  AOI21_X1 U14128 ( .B1(n11644), .B2(n11643), .A(n15277), .ZN(n11750) );
  INV_X1 U14129 ( .A(n11750), .ZN(n11655) );
  XNOR2_X1 U14130 ( .A(n11645), .B(n14535), .ZN(n11752) );
  AOI21_X1 U14131 ( .B1(n11646), .B2(n14355), .A(n10283), .ZN(n11647) );
  NAND2_X1 U14132 ( .A1(n11647), .A2(n11760), .ZN(n11749) );
  NAND2_X1 U14133 ( .A1(n14964), .A2(n14575), .ZN(n11650) );
  INV_X1 U14134 ( .A(n11648), .ZN(n14219) );
  AOI22_X1 U14135 ( .A1(n15269), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n14219), 
        .B2(n15258), .ZN(n11649) );
  OAI211_X1 U14136 ( .C1(n14360), .C2(n14969), .A(n11650), .B(n11649), .ZN(
        n11651) );
  AOI21_X1 U14137 ( .B1(n14971), .B2(n14355), .A(n11651), .ZN(n11652) );
  OAI21_X1 U14138 ( .B1(n11749), .B2(n14974), .A(n11652), .ZN(n11653) );
  AOI21_X1 U14139 ( .B1(n11752), .B2(n14903), .A(n11653), .ZN(n11654) );
  OAI21_X1 U14140 ( .B1(n11655), .B2(n15260), .A(n11654), .ZN(P1_U3284) );
  AND2_X1 U14141 ( .A1(n13347), .A2(n13542), .ZN(n11657) );
  XNOR2_X1 U14142 ( .A(n13148), .B(n7171), .ZN(n11656) );
  NOR2_X1 U14143 ( .A1(n11656), .A2(n11657), .ZN(n11738) );
  AOI21_X1 U14144 ( .B1(n11657), .B2(n11656), .A(n11738), .ZN(n11662) );
  INV_X1 U14145 ( .A(n11658), .ZN(n11659) );
  OAI21_X1 U14146 ( .B1(n11662), .B2(n11661), .A(n11740), .ZN(n11663) );
  NAND2_X1 U14147 ( .A1(n11663), .A2(n13042), .ZN(n11667) );
  NAND2_X1 U14148 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n15392) );
  OAI21_X1 U14149 ( .B1(n13074), .B2(n11664), .A(n15392), .ZN(n11665) );
  AOI21_X1 U14150 ( .B1(n13148), .B2(n13087), .A(n11665), .ZN(n11666) );
  OAI211_X1 U14151 ( .C1(n13085), .C2(n11668), .A(n11667), .B(n11666), .ZN(
        P2_U3203) );
  INV_X1 U14152 ( .A(n11669), .ZN(n11670) );
  OAI222_X1 U14153 ( .A1(n13916), .A2(n11671), .B1(n13913), .B2(n11670), .C1(
        n9859), .C2(P2_U3088), .ZN(P2_U3305) );
  MUX2_X1 U14154 ( .A(n11673), .B(n11672), .S(n15514), .Z(n11676) );
  NAND2_X1 U14155 ( .A1(n11674), .A2(n12836), .ZN(n11675) );
  OAI211_X1 U14156 ( .C1(n12821), .C2(n11677), .A(n11676), .B(n11675), .ZN(
        P3_U3469) );
  INV_X1 U14157 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n12094) );
  NAND2_X1 U14158 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n12965)
         );
  INV_X1 U14159 ( .A(n12965), .ZN(n11686) );
  XOR2_X1 U14160 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n11678), .Z(n11679) );
  NAND2_X1 U14161 ( .A1(n15405), .A2(n11679), .ZN(n11684) );
  XOR2_X1 U14162 ( .A(n11681), .B(n11680), .Z(n11682) );
  NAND2_X1 U14163 ( .A1(n15403), .A2(n11682), .ZN(n11683) );
  NAND2_X1 U14164 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  AOI211_X1 U14165 ( .C1(n6638), .C2(n11687), .A(n11686), .B(n11685), .ZN(
        n11688) );
  OAI21_X1 U14166 ( .B1(n12094), .B2(n15399), .A(n11688), .ZN(P2_U3228) );
  XNOR2_X1 U14167 ( .A(n11689), .B(n13311), .ZN(n11878) );
  INV_X1 U14168 ( .A(n11878), .ZN(n11704) );
  OAI211_X1 U14169 ( .C1(n11691), .C2(n13311), .A(n11690), .B(n13717), .ZN(
        n11694) );
  OAI22_X1 U14170 ( .A1(n11692), .A2(n13676), .B1(n12045), .B2(n13678), .ZN(
        n11741) );
  INV_X1 U14171 ( .A(n11741), .ZN(n11693) );
  NAND2_X1 U14172 ( .A1(n11694), .A2(n11693), .ZN(n11876) );
  NAND2_X1 U14173 ( .A1(n11876), .A2(n13687), .ZN(n11703) );
  INV_X1 U14174 ( .A(n11695), .ZN(n11697) );
  INV_X1 U14175 ( .A(n11856), .ZN(n11696) );
  AOI211_X1 U14176 ( .C1(n13152), .C2(n11697), .A(n13542), .B(n11696), .ZN(
        n11877) );
  NOR2_X1 U14177 ( .A1(n13735), .A2(n11698), .ZN(n11701) );
  OAI22_X1 U14178 ( .A1(n13687), .A2(n11699), .B1(n11744), .B2(n13683), .ZN(
        n11700) );
  AOI211_X1 U14179 ( .C1(n11877), .C2(n13708), .A(n11701), .B(n11700), .ZN(
        n11702) );
  OAI211_X1 U14180 ( .C1(n13738), .C2(n11704), .A(n11703), .B(n11702), .ZN(
        P2_U3255) );
  NAND2_X1 U14181 ( .A1(n11706), .A2(n11705), .ZN(n11711) );
  INV_X1 U14182 ( .A(n11707), .ZN(n11708) );
  NAND2_X1 U14183 ( .A1(n11709), .A2(n11708), .ZN(n11710) );
  NAND2_X1 U14184 ( .A1(n11711), .A2(n11710), .ZN(n11836) );
  XNOR2_X1 U14185 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n11715) );
  XNOR2_X1 U14186 ( .A(n11841), .B(n11715), .ZN(n11837) );
  XOR2_X1 U14187 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n11837), .Z(n11716) );
  XNOR2_X1 U14188 ( .A(n11836), .B(n11716), .ZN(SUB_1596_U67) );
  XNOR2_X1 U14189 ( .A(n11787), .B(n6610), .ZN(n11771) );
  XNOR2_X1 U14190 ( .A(n11909), .B(n11174), .ZN(n11722) );
  NAND2_X1 U14191 ( .A1(n11722), .A2(n11777), .ZN(n11900) );
  OAI21_X1 U14192 ( .B1(n11771), .B2(n11955), .A(n11900), .ZN(n11719) );
  INV_X1 U14193 ( .A(n11722), .ZN(n11723) );
  NAND2_X1 U14194 ( .A1(n11723), .A2(n12454), .ZN(n11901) );
  XNOR2_X1 U14195 ( .A(n12110), .B(n6610), .ZN(n11865) );
  XNOR2_X1 U14196 ( .A(n11865), .B(n12781), .ZN(n11724) );
  XNOR2_X1 U14197 ( .A(n11868), .B(n11724), .ZN(n11730) );
  NAND2_X1 U14198 ( .A1(n12427), .A2(n12454), .ZN(n11725) );
  NAND2_X1 U14199 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12466)
         );
  OAI211_X1 U14200 ( .C1(n12058), .C2(n12429), .A(n11725), .B(n12466), .ZN(
        n11728) );
  NOR2_X1 U14201 ( .A1(n11726), .A2(n12448), .ZN(n11727) );
  AOI211_X1 U14202 ( .C1(n12109), .C2(n12441), .A(n11728), .B(n11727), .ZN(
        n11729) );
  OAI21_X1 U14203 ( .B1(n11730), .B2(n12434), .A(n11729), .ZN(P3_U3174) );
  NAND2_X1 U14204 ( .A1(n12453), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11731) );
  OAI21_X1 U14205 ( .B1(n12355), .B2(n12453), .A(n11731), .ZN(P3_U3520) );
  AOI211_X1 U14206 ( .C1(n11734), .C2(n13835), .A(n11733), .B(n11732), .ZN(
        n11737) );
  AOI22_X1 U14207 ( .A1(n13789), .A2(n13148), .B1(P2_REG1_REG_9__SCAN_IN), 
        .B2(n15452), .ZN(n11735) );
  OAI21_X1 U14208 ( .B1(n11737), .B2(n15452), .A(n11735), .ZN(P2_U3508) );
  AOI22_X1 U14209 ( .A1(n13881), .A2(n13148), .B1(P2_REG0_REG_9__SCAN_IN), 
        .B2(n15446), .ZN(n11736) );
  OAI21_X1 U14210 ( .B1(n11737), .B2(n15446), .A(n11736), .ZN(P2_U3457) );
  INV_X1 U14211 ( .A(n11738), .ZN(n11739) );
  XNOR2_X1 U14212 ( .A(n13152), .B(n7171), .ZN(n11980) );
  NAND2_X1 U14213 ( .A1(n13346), .A2(n13542), .ZN(n11979) );
  XNOR2_X1 U14214 ( .A(n11980), .B(n11979), .ZN(n11982) );
  XNOR2_X1 U14215 ( .A(n11983), .B(n11982), .ZN(n11747) );
  NAND2_X1 U14216 ( .A1(n13061), .A2(n11741), .ZN(n11742) );
  OAI211_X1 U14217 ( .C1(n13085), .C2(n11744), .A(n11743), .B(n11742), .ZN(
        n11745) );
  AOI21_X1 U14218 ( .B1(n13152), .B2(n13087), .A(n11745), .ZN(n11746) );
  OAI21_X1 U14219 ( .B1(n11747), .B2(n13089), .A(n11746), .ZN(P2_U3189) );
  AOI22_X1 U14220 ( .A1(n14575), .A2(n15107), .B1(n15090), .B2(n14574), .ZN(
        n11748) );
  OAI211_X1 U14221 ( .C1(n7437), .C2(n15302), .A(n11749), .B(n11748), .ZN(
        n11751) );
  AOI211_X1 U14222 ( .C1(n11752), .C2(n15321), .A(n11751), .B(n11750), .ZN(
        n11755) );
  NAND2_X1 U14223 ( .A1(n15323), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11753) );
  OAI21_X1 U14224 ( .B1(n11755), .B2(n15323), .A(n11753), .ZN(P1_U3486) );
  NAND2_X1 U14225 ( .A1(n15331), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11754) );
  OAI21_X1 U14226 ( .B1(n11755), .B2(n15331), .A(n11754), .ZN(P1_U3537) );
  XNOR2_X1 U14227 ( .A(n11756), .B(n11757), .ZN(n15109) );
  INV_X1 U14228 ( .A(n15109), .ZN(n11770) );
  OR2_X1 U14229 ( .A1(n11758), .A2(n14538), .ZN(n15105) );
  NAND3_X1 U14230 ( .A1(n15105), .A2(n14879), .A3(n11759), .ZN(n11769) );
  XNOR2_X1 U14231 ( .A(n11760), .B(n14359), .ZN(n11762) );
  AND2_X1 U14232 ( .A1(n15092), .A2(n15090), .ZN(n11761) );
  AOI21_X1 U14233 ( .B1(n11762), .B2(n15240), .A(n11761), .ZN(n15112) );
  INV_X1 U14234 ( .A(n15112), .ZN(n11767) );
  INV_X1 U14235 ( .A(n15311), .ZN(n15106) );
  OAI22_X1 U14236 ( .A1(n14798), .A2(n11763), .B1(n12181), .B2(n15236), .ZN(
        n11764) );
  AOI21_X1 U14237 ( .B1(n14964), .B2(n15106), .A(n11764), .ZN(n11765) );
  OAI21_X1 U14238 ( .B1(n14359), .B2(n15262), .A(n11765), .ZN(n11766) );
  AOI21_X1 U14239 ( .B1(n11767), .B2(n15266), .A(n11766), .ZN(n11768) );
  OAI211_X1 U14240 ( .C1(n11770), .C2(n14978), .A(n11769), .B(n11768), .ZN(
        P1_U3283) );
  INV_X1 U14241 ( .A(n11772), .ZN(n11774) );
  INV_X1 U14242 ( .A(n11771), .ZN(n11773) );
  OR2_X1 U14243 ( .A1(n11772), .A2(n11771), .ZN(n11902) );
  OAI21_X1 U14244 ( .B1(n11774), .B2(n11773), .A(n11902), .ZN(n11775) );
  NOR2_X1 U14245 ( .A1(n11775), .A2(n11955), .ZN(n11904) );
  AOI21_X1 U14246 ( .B1(n11955), .B2(n11775), .A(n11904), .ZN(n11781) );
  NAND2_X1 U14247 ( .A1(n12427), .A2(n12455), .ZN(n11776) );
  NAND2_X1 U14248 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11926)
         );
  OAI211_X1 U14249 ( .C1(n11777), .C2(n12429), .A(n11776), .B(n11926), .ZN(
        n11779) );
  NOR2_X1 U14250 ( .A1(n11787), .A2(n12448), .ZN(n11778) );
  AOI211_X1 U14251 ( .C1(n11788), .C2(n12441), .A(n11779), .B(n11778), .ZN(
        n11780) );
  OAI21_X1 U14252 ( .B1(n11781), .B2(n12434), .A(n11780), .ZN(P3_U3176) );
  MUX2_X1 U14253 ( .A(n12001), .B(n11785), .S(n15514), .Z(n11783) );
  NAND2_X1 U14254 ( .A1(n11784), .A2(n12836), .ZN(n11782) );
  OAI211_X1 U14255 ( .C1(n12821), .C2(n11787), .A(n11783), .B(n11782), .ZN(
        P3_U3470) );
  INV_X1 U14256 ( .A(n11784), .ZN(n11792) );
  MUX2_X1 U14257 ( .A(n11786), .B(n11785), .S(n15472), .Z(n11791) );
  INV_X1 U14258 ( .A(n11787), .ZN(n11789) );
  AOI22_X1 U14259 ( .A1(n11789), .A2(n12787), .B1(n15488), .B2(n11788), .ZN(
        n11790) );
  OAI211_X1 U14260 ( .C1(n11792), .C2(n12790), .A(n11791), .B(n11790), .ZN(
        P3_U3222) );
  NOR2_X1 U14261 ( .A1(n11972), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11971) );
  INV_X1 U14262 ( .A(n11794), .ZN(n11795) );
  NOR2_X1 U14263 ( .A1(n11795), .A2(n11976), .ZN(n11797) );
  XNOR2_X1 U14264 ( .A(n14636), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11796) );
  INV_X1 U14265 ( .A(n14635), .ZN(n11799) );
  OAI21_X1 U14266 ( .B1(n11971), .B2(n11797), .A(n11796), .ZN(n11798) );
  NAND3_X1 U14267 ( .A1(n11799), .A2(n15210), .A3(n11798), .ZN(n11809) );
  NAND2_X1 U14268 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14171)
         );
  XOR2_X1 U14269 ( .A(n14636), .B(P1_REG2_REG_16__SCAN_IN), .Z(n11805) );
  XNOR2_X1 U14270 ( .A(n11802), .B(n11976), .ZN(n11970) );
  AOI22_X1 U14271 ( .A1(n11970), .A2(n11803), .B1(n11802), .B2(n7072), .ZN(
        n11804) );
  NAND2_X1 U14272 ( .A1(n11804), .A2(n11805), .ZN(n14632) );
  OAI211_X1 U14273 ( .C1(n11805), .C2(n11804), .A(n15217), .B(n14632), .ZN(
        n11806) );
  NAND2_X1 U14274 ( .A1(n14171), .A2(n11806), .ZN(n11807) );
  AOI21_X1 U14275 ( .B1(n14653), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11807), 
        .ZN(n11808) );
  OAI211_X1 U14276 ( .C1(n15221), .C2(n11810), .A(n11809), .B(n11808), .ZN(
        P1_U3259) );
  INV_X1 U14277 ( .A(n11811), .ZN(n11812) );
  NAND2_X1 U14278 ( .A1(n14348), .A2(n10284), .ZN(n11817) );
  OR2_X1 U14279 ( .A1(n15313), .A2(n14020), .ZN(n11816) );
  NAND2_X1 U14280 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  XNOR2_X1 U14281 ( .A(n11818), .B(n14111), .ZN(n11820) );
  OAI22_X1 U14282 ( .A1(n15303), .A2(n14020), .B1(n15313), .B2(n14052), .ZN(
        n11819) );
  XNOR2_X1 U14283 ( .A(n11820), .B(n11819), .ZN(n11938) );
  NAND2_X1 U14284 ( .A1(n15316), .A2(n10284), .ZN(n11822) );
  OR2_X1 U14285 ( .A1(n11933), .A2(n14020), .ZN(n11821) );
  NAND2_X1 U14286 ( .A1(n11822), .A2(n11821), .ZN(n11823) );
  XNOR2_X1 U14287 ( .A(n11823), .B(n14051), .ZN(n11825) );
  AOI22_X1 U14288 ( .A1(n15316), .A2(n10286), .B1(n14108), .B2(n14575), .ZN(
        n11824) );
  NAND2_X1 U14289 ( .A1(n11825), .A2(n11824), .ZN(n12159) );
  OAI21_X1 U14290 ( .B1(n11825), .B2(n11824), .A(n12159), .ZN(n11826) );
  AOI21_X1 U14291 ( .B1(n11827), .B2(n11826), .A(n12161), .ZN(n11834) );
  NAND2_X1 U14292 ( .A1(n14275), .A2(n14576), .ZN(n11831) );
  AOI21_X1 U14293 ( .B1(n14295), .B2(n11829), .A(n11828), .ZN(n11830) );
  OAI211_X1 U14294 ( .C1(n15311), .C2(n14272), .A(n11831), .B(n11830), .ZN(
        n11832) );
  AOI21_X1 U14295 ( .B1(n15316), .B2(n14300), .A(n11832), .ZN(n11833) );
  OAI21_X1 U14296 ( .B1(n11834), .B2(n14302), .A(n11833), .ZN(P1_U3221) );
  NAND2_X1 U14297 ( .A1(n11837), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11835) );
  NAND2_X1 U14298 ( .A1(n11836), .A2(n11835), .ZN(n11839) );
  OR2_X1 U14299 ( .A1(n11837), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U14300 ( .A1(n11839), .A2(n11838), .ZN(n12093) );
  INV_X1 U14301 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12467) );
  NAND2_X1 U14302 ( .A1(n12467), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11840) );
  NAND2_X1 U14303 ( .A1(n11841), .A2(n11840), .ZN(n11844) );
  INV_X1 U14304 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n11842) );
  NAND2_X1 U14305 ( .A1(n11842), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n11843) );
  NAND2_X1 U14306 ( .A1(n11844), .A2(n11843), .ZN(n11848) );
  INV_X1 U14307 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U14308 ( .A1(n12504), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n12097) );
  NAND2_X1 U14309 ( .A1(n11845), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n11846) );
  NAND2_X1 U14310 ( .A1(n12097), .A2(n11846), .ZN(n11847) );
  NAND2_X1 U14311 ( .A1(n11848), .A2(n11847), .ZN(n11849) );
  NAND2_X1 U14312 ( .A1(n12098), .A2(n11849), .ZN(n12095) );
  XNOR2_X1 U14313 ( .A(n12095), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(n11850) );
  XNOR2_X1 U14314 ( .A(n12093), .B(n11850), .ZN(SUB_1596_U66) );
  OAI21_X1 U14315 ( .B1(n6576), .B2(n13315), .A(n11851), .ZN(n11854) );
  INV_X1 U14316 ( .A(n13346), .ZN(n11853) );
  OAI22_X1 U14317 ( .A1(n11853), .A2(n13676), .B1(n11852), .B2(n13678), .ZN(
        n11992) );
  AOI21_X1 U14318 ( .B1(n11854), .B2(n13717), .A(n11992), .ZN(n13853) );
  INV_X1 U14319 ( .A(n12047), .ZN(n11855) );
  AOI211_X1 U14320 ( .C1(n7105), .C2(n11856), .A(n13542), .B(n11855), .ZN(
        n13850) );
  INV_X1 U14321 ( .A(n11989), .ZN(n11857) );
  AOI22_X1 U14322 ( .A1(n6402), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11857), 
        .B2(n13731), .ZN(n11858) );
  OAI21_X1 U14323 ( .B1(n7688), .B2(n13735), .A(n11858), .ZN(n11862) );
  XNOR2_X1 U14324 ( .A(n11860), .B(n11859), .ZN(n13854) );
  NOR2_X1 U14325 ( .A1(n13854), .A2(n13738), .ZN(n11861) );
  AOI211_X1 U14326 ( .C1(n13850), .C2(n13708), .A(n11862), .B(n11861), .ZN(
        n11863) );
  OAI21_X1 U14327 ( .B1(n6402), .B2(n13853), .A(n11863), .ZN(P2_U3254) );
  NAND2_X1 U14328 ( .A1(n11865), .A2(n11864), .ZN(n11867) );
  INV_X1 U14329 ( .A(n11865), .ZN(n11866) );
  XNOR2_X1 U14330 ( .A(n12916), .B(n6610), .ZN(n12055) );
  XNOR2_X1 U14331 ( .A(n12055), .B(n12058), .ZN(n11869) );
  XNOR2_X1 U14332 ( .A(n12054), .B(n11869), .ZN(n11875) );
  NAND2_X1 U14333 ( .A1(n12427), .A2(n12781), .ZN(n11870) );
  NAND2_X1 U14334 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12503)
         );
  OAI211_X1 U14335 ( .C1(n12383), .C2(n12429), .A(n11870), .B(n12503), .ZN(
        n11873) );
  NOR2_X1 U14336 ( .A1(n11871), .A2(n12448), .ZN(n11872) );
  AOI211_X1 U14337 ( .C1(n12786), .C2(n12441), .A(n11873), .B(n11872), .ZN(
        n11874) );
  OAI21_X1 U14338 ( .B1(n11875), .B2(n12434), .A(n11874), .ZN(P3_U3155) );
  AOI211_X1 U14339 ( .C1(n13835), .C2(n11878), .A(n11877), .B(n11876), .ZN(
        n11881) );
  AOI22_X1 U14340 ( .A1(n13881), .A2(n13152), .B1(P2_REG0_REG_10__SCAN_IN), 
        .B2(n15446), .ZN(n11879) );
  OAI21_X1 U14341 ( .B1(n11881), .B2(n15446), .A(n11879), .ZN(P2_U3460) );
  AOI22_X1 U14342 ( .A1(n13789), .A2(n13152), .B1(P2_REG1_REG_10__SCAN_IN), 
        .B2(n15452), .ZN(n11880) );
  OAI21_X1 U14343 ( .B1(n11881), .B2(n15452), .A(n11880), .ZN(P2_U3509) );
  NAND2_X1 U14344 ( .A1(n11882), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11885) );
  NAND2_X1 U14345 ( .A1(n11883), .A2(n11887), .ZN(n11884) );
  NAND2_X1 U14346 ( .A1(n11885), .A2(n11884), .ZN(n13406) );
  INV_X1 U14347 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13669) );
  XNOR2_X1 U14348 ( .A(n13407), .B(n13669), .ZN(n13405) );
  XNOR2_X1 U14349 ( .A(n13406), .B(n13405), .ZN(n11895) );
  NAND2_X1 U14350 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13017)
         );
  XNOR2_X1 U14351 ( .A(n13407), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13399) );
  XOR2_X1 U14352 ( .A(n13400), .B(n13399), .Z(n11889) );
  NAND2_X1 U14353 ( .A1(n15403), .A2(n11889), .ZN(n11890) );
  NAND2_X1 U14354 ( .A1(n13017), .A2(n11890), .ZN(n11892) );
  NOR2_X1 U14355 ( .A1(n15395), .A2(n13398), .ZN(n11891) );
  AOI211_X1 U14356 ( .C1(n15334), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n11892), 
        .B(n11891), .ZN(n11893) );
  OAI21_X1 U14357 ( .B1(n11895), .B2(n11894), .A(n11893), .ZN(P2_U3230) );
  INV_X1 U14358 ( .A(n11896), .ZN(n11898) );
  OAI222_X1 U14359 ( .A1(n12941), .A2(n11899), .B1(n12948), .B2(n11898), .C1(
        P3_U3151), .C2(n11897), .ZN(P3_U3271) );
  NAND2_X1 U14360 ( .A1(n11901), .A2(n11900), .ZN(n11906) );
  INV_X1 U14361 ( .A(n11902), .ZN(n11903) );
  NOR2_X1 U14362 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  XOR2_X1 U14363 ( .A(n11906), .B(n11905), .Z(n11913) );
  NAND2_X1 U14364 ( .A1(n12445), .A2(n12781), .ZN(n11907) );
  NAND2_X1 U14365 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12009)
         );
  OAI211_X1 U14366 ( .C1(n11908), .C2(n12443), .A(n11907), .B(n12009), .ZN(
        n11911) );
  NOR2_X1 U14367 ( .A1(n11909), .A2(n12448), .ZN(n11910) );
  AOI211_X1 U14368 ( .C1(n11961), .C2(n12441), .A(n11911), .B(n11910), .ZN(
        n11912) );
  OAI21_X1 U14369 ( .B1(n11913), .B2(n12434), .A(n11912), .ZN(P3_U3164) );
  XNOR2_X1 U14370 ( .A(n12002), .B(P3_REG1_REG_11__SCAN_IN), .ZN(n11932) );
  OAI21_X1 U14371 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n11918), .A(n12007), 
        .ZN(n11919) );
  NAND2_X1 U14372 ( .A1(n11919), .A2(n12590), .ZN(n11931) );
  INV_X1 U14373 ( .A(n11920), .ZN(n11921) );
  NAND2_X1 U14374 ( .A1(n11922), .A2(n11921), .ZN(n11924) );
  MUX2_X1 U14375 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12937), .Z(n12011) );
  XOR2_X1 U14376 ( .A(n11927), .B(n12011), .Z(n11923) );
  NAND2_X1 U14377 ( .A1(n11924), .A2(n11923), .ZN(n12016) );
  OAI21_X1 U14378 ( .B1(n11924), .B2(n11923), .A(n12016), .ZN(n11929) );
  NAND2_X1 U14379 ( .A1(n15455), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11925) );
  OAI211_X1 U14380 ( .C1(n12597), .C2(n11927), .A(n11926), .B(n11925), .ZN(
        n11928) );
  AOI21_X1 U14381 ( .B1(n11929), .B2(n12491), .A(n11928), .ZN(n11930) );
  OAI211_X1 U14382 ( .C1(n11932), .C2(n12024), .A(n11931), .B(n11930), .ZN(
        P3_U3193) );
  OR2_X1 U14383 ( .A1(n11933), .A2(n15310), .ZN(n11935) );
  NAND2_X1 U14384 ( .A1(n14577), .A2(n15107), .ZN(n11934) );
  NAND2_X1 U14385 ( .A1(n11935), .A2(n11934), .ZN(n15233) );
  NAND2_X1 U14386 ( .A1(n14288), .A2(n15233), .ZN(n11937) );
  OAI211_X1 U14387 ( .C1(n14286), .C2(n15235), .A(n11937), .B(n11936), .ZN(
        n11942) );
  XNOR2_X1 U14388 ( .A(n11939), .B(n11938), .ZN(n11940) );
  NOR2_X1 U14389 ( .A1(n11940), .A2(n14302), .ZN(n11941) );
  AOI211_X1 U14390 ( .C1(n14348), .C2(n14300), .A(n11942), .B(n11941), .ZN(
        n11943) );
  INV_X1 U14391 ( .A(n11943), .ZN(P1_U3213) );
  INV_X1 U14392 ( .A(n11944), .ZN(n11947) );
  OAI222_X1 U14393 ( .A1(P1_U3086), .A2(n11946), .B1(n15144), .B2(n11945), 
        .C1(n15147), .C2(n11947), .ZN(P1_U3329) );
  OAI222_X1 U14394 ( .A1(P2_U3088), .A2(n11949), .B1(n13916), .B2(n11948), 
        .C1(n13913), .C2(n11947), .ZN(P2_U3301) );
  XOR2_X1 U14395 ( .A(n11950), .B(n11951), .Z(n11969) );
  NAND2_X1 U14396 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  NAND2_X1 U14397 ( .A1(n11953), .A2(n12784), .ZN(n11954) );
  OR2_X1 U14398 ( .A1(n6575), .A2(n11954), .ZN(n11957) );
  AOI22_X1 U14399 ( .A1(n11955), .A2(n12704), .B1(n15479), .B2(n12781), .ZN(
        n11956) );
  AND2_X1 U14400 ( .A1(n11957), .A2(n11956), .ZN(n11965) );
  MUX2_X1 U14401 ( .A(n11965), .B(n11958), .S(n9433), .Z(n11960) );
  NAND2_X1 U14402 ( .A1(n11966), .A2(n12840), .ZN(n11959) );
  OAI211_X1 U14403 ( .C1(n12843), .C2(n11969), .A(n11960), .B(n11959), .ZN(
        P3_U3471) );
  MUX2_X1 U14404 ( .A(n11965), .B(n12004), .S(n15493), .Z(n11963) );
  AOI22_X1 U14405 ( .A1(n11966), .A2(n12787), .B1(n15488), .B2(n11961), .ZN(
        n11962) );
  OAI211_X1 U14406 ( .C1(n11969), .C2(n12790), .A(n11963), .B(n11962), .ZN(
        P3_U3221) );
  MUX2_X1 U14407 ( .A(n11965), .B(n11964), .S(n15509), .Z(n11968) );
  NAND2_X1 U14408 ( .A1(n11966), .A2(n12915), .ZN(n11967) );
  OAI211_X1 U14409 ( .C1(n11969), .C2(n12919), .A(n11968), .B(n11967), .ZN(
        P3_U3426) );
  XNOR2_X1 U14410 ( .A(n11970), .B(P1_REG2_REG_15__SCAN_IN), .ZN(n11978) );
  INV_X1 U14411 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15551) );
  NAND2_X1 U14412 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14297)
         );
  OAI21_X1 U14413 ( .B1(n15226), .B2(n15551), .A(n14297), .ZN(n11975) );
  AOI21_X1 U14414 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11972), .A(n11971), 
        .ZN(n11973) );
  NOR2_X1 U14415 ( .A1(n11973), .A2(n14668), .ZN(n11974) );
  AOI211_X1 U14416 ( .C1(n14654), .C2(n11976), .A(n11975), .B(n11974), .ZN(
        n11977) );
  OAI21_X1 U14417 ( .B1(n11978), .B2(n14657), .A(n11977), .ZN(P1_U3258) );
  INV_X1 U14418 ( .A(n11979), .ZN(n11981) );
  AND2_X1 U14419 ( .A1(n13345), .A2(n13542), .ZN(n11985) );
  XNOR2_X1 U14420 ( .A(n7105), .B(n7171), .ZN(n11984) );
  NOR2_X1 U14421 ( .A1(n11984), .A2(n11985), .ZN(n12079) );
  AOI21_X1 U14422 ( .B1(n11985), .B2(n11984), .A(n12079), .ZN(n11986) );
  OAI21_X1 U14423 ( .B1(n11987), .B2(n11986), .A(n12081), .ZN(n11988) );
  NAND2_X1 U14424 ( .A1(n11988), .A2(n13042), .ZN(n11994) );
  NOR2_X1 U14425 ( .A1(n13085), .A2(n11989), .ZN(n11990) );
  AOI211_X1 U14426 ( .C1(n13061), .C2(n11992), .A(n11991), .B(n11990), .ZN(
        n11993) );
  OAI211_X1 U14427 ( .C1(n7688), .C2(n13049), .A(n11994), .B(n11993), .ZN(
        P2_U3208) );
  INV_X1 U14428 ( .A(n11995), .ZN(n11999) );
  OAI222_X1 U14429 ( .A1(n11997), .A2(P2_U3088), .B1(n13913), .B2(n11999), 
        .C1(n11996), .C2(n13916), .ZN(P2_U3303) );
  OAI222_X1 U14430 ( .A1(n15144), .A2(n15647), .B1(n15147), .B2(n11999), .C1(
        P1_U3086), .C2(n11998), .ZN(P1_U3331) );
  XNOR2_X1 U14431 ( .A(n12021), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n12477) );
  XOR2_X1 U14432 ( .A(n12477), .B(n6441), .Z(n12025) );
  INV_X1 U14433 ( .A(n12003), .ZN(n12005) );
  XNOR2_X1 U14434 ( .A(n12021), .B(n12004), .ZN(n12006) );
  AND3_X1 U14435 ( .A1(n12007), .A2(n12006), .A3(n12005), .ZN(n12008) );
  OAI21_X1 U14436 ( .B1(n12462), .B2(n12008), .A(n12590), .ZN(n12023) );
  OAI21_X1 U14437 ( .B1(n12581), .B2(n12010), .A(n12009), .ZN(n12020) );
  INV_X1 U14438 ( .A(n12011), .ZN(n12013) );
  NAND2_X1 U14439 ( .A1(n12013), .A2(n12012), .ZN(n12015) );
  MUX2_X1 U14440 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12937), .Z(n12468) );
  XNOR2_X1 U14441 ( .A(n12468), .B(n12021), .ZN(n12014) );
  NAND3_X1 U14442 ( .A1(n12016), .A2(n12015), .A3(n12014), .ZN(n12472) );
  INV_X1 U14443 ( .A(n12472), .ZN(n12018) );
  AOI21_X1 U14444 ( .B1(n12016), .B2(n12015), .A(n12014), .ZN(n12017) );
  NOR3_X1 U14445 ( .A1(n12018), .A2(n12017), .A3(n12605), .ZN(n12019) );
  AOI211_X1 U14446 ( .C1(n12578), .C2(n12021), .A(n12020), .B(n12019), .ZN(
        n12022) );
  OAI211_X1 U14447 ( .C1(n12025), .C2(n12024), .A(n12023), .B(n12022), .ZN(
        P3_U3194) );
  XNOR2_X1 U14448 ( .A(n12026), .B(n14539), .ZN(n15104) );
  OAI211_X1 U14449 ( .C1(n14539), .C2(n12028), .A(n12027), .B(n15308), .ZN(
        n12031) );
  NAND2_X1 U14450 ( .A1(n14574), .A2(n15107), .ZN(n12030) );
  NAND2_X1 U14451 ( .A1(n14946), .A2(n15090), .ZN(n12029) );
  AND2_X1 U14452 ( .A1(n12030), .A2(n12029), .ZN(n14261) );
  NAND2_X1 U14453 ( .A1(n12031), .A2(n14261), .ZN(n15100) );
  OR2_X1 U14454 ( .A1(n12033), .A2(n14363), .ZN(n12034) );
  AND3_X1 U14455 ( .A1(n12032), .A2(n12034), .A3(n15240), .ZN(n15101) );
  NAND2_X1 U14456 ( .A1(n15101), .A2(n15266), .ZN(n12038) );
  NAND2_X1 U14457 ( .A1(n15260), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n12035) );
  OAI21_X1 U14458 ( .B1(n15236), .B2(n14263), .A(n12035), .ZN(n12036) );
  AOI21_X1 U14459 ( .B1(n7165), .B2(n14971), .A(n12036), .ZN(n12037) );
  NAND2_X1 U14460 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  AOI21_X1 U14461 ( .B1(n15100), .B2(n14798), .A(n12039), .ZN(n12040) );
  OAI21_X1 U14462 ( .B1(n14978), .B2(n15104), .A(n12040), .ZN(P1_U3282) );
  INV_X1 U14463 ( .A(n12044), .ZN(n12042) );
  NAND2_X1 U14464 ( .A1(n12042), .A2(n13313), .ZN(n13694) );
  AOI21_X1 U14465 ( .B1(n12044), .B2(n12043), .A(n13701), .ZN(n12046) );
  OAI22_X1 U14466 ( .A1(n12045), .A2(n13676), .B1(n13695), .B2(n13678), .ZN(
        n12088) );
  AOI21_X1 U14467 ( .B1(n13694), .B2(n12046), .A(n12088), .ZN(n13848) );
  AOI211_X1 U14468 ( .C1(n13846), .C2(n12047), .A(n13542), .B(n13727), .ZN(
        n13845) );
  INV_X1 U14469 ( .A(n12085), .ZN(n12048) );
  AOI22_X1 U14470 ( .A1(n6402), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12048), 
        .B2(n13731), .ZN(n12049) );
  OAI21_X1 U14471 ( .B1(n13735), .B2(n12091), .A(n12049), .ZN(n12052) );
  XNOR2_X1 U14472 ( .A(n12050), .B(n13313), .ZN(n13849) );
  NOR2_X1 U14473 ( .A1(n13849), .A2(n13738), .ZN(n12051) );
  AOI211_X1 U14474 ( .C1(n13845), .C2(n13708), .A(n12052), .B(n12051), .ZN(
        n12053) );
  OAI21_X1 U14475 ( .B1(n6402), .B2(n13848), .A(n12053), .ZN(P2_U3253) );
  XNOR2_X1 U14476 ( .A(n12908), .B(n6610), .ZN(n12295) );
  XNOR2_X1 U14477 ( .A(n12295), .B(n12383), .ZN(n12056) );
  XNOR2_X1 U14478 ( .A(n12294), .B(n12056), .ZN(n12063) );
  NAND2_X1 U14479 ( .A1(n12445), .A2(n12770), .ZN(n12057) );
  NAND2_X1 U14480 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12517)
         );
  OAI211_X1 U14481 ( .C1(n12058), .C2(n12443), .A(n12057), .B(n12517), .ZN(
        n12061) );
  NOR2_X1 U14482 ( .A1(n12059), .A2(n12448), .ZN(n12060) );
  AOI211_X1 U14483 ( .C1(n12773), .C2(n12441), .A(n12061), .B(n12060), .ZN(
        n12062) );
  OAI21_X1 U14484 ( .B1(n12063), .B2(n12434), .A(n12062), .ZN(P3_U3181) );
  INV_X1 U14485 ( .A(n12064), .ZN(n15142) );
  AOI21_X1 U14486 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n13910), .A(n12065), 
        .ZN(n12066) );
  OAI21_X1 U14487 ( .B1(n15142), .B2(n13913), .A(n12066), .ZN(P2_U3300) );
  XNOR2_X1 U14488 ( .A(n12068), .B(n12067), .ZN(n12069) );
  AOI222_X1 U14489 ( .A1(n12784), .A2(n12069), .B1(n12769), .B2(n15479), .C1(
        n12454), .C2(n12704), .ZN(n12108) );
  MUX2_X1 U14490 ( .A(n15554), .B(n12108), .S(n15514), .Z(n12073) );
  XNOR2_X1 U14491 ( .A(n12070), .B(n12071), .ZN(n12107) );
  AOI22_X1 U14492 ( .A1(n12107), .A2(n12836), .B1(n12840), .B2(n12110), .ZN(
        n12072) );
  NAND2_X1 U14493 ( .A1(n12073), .A2(n12072), .ZN(P3_U3472) );
  MUX2_X1 U14494 ( .A(n12074), .B(n12108), .S(n15510), .Z(n12076) );
  AOI22_X1 U14495 ( .A1(n12107), .A2(n12909), .B1(n12915), .B2(n12110), .ZN(
        n12075) );
  NAND2_X1 U14496 ( .A1(n12076), .A2(n12075), .ZN(P3_U3429) );
  AND2_X1 U14497 ( .A1(n13721), .A2(n13542), .ZN(n12078) );
  XNOR2_X1 U14498 ( .A(n13846), .B(n7171), .ZN(n12077) );
  NOR2_X1 U14499 ( .A1(n12077), .A2(n12078), .ZN(n12114) );
  AOI21_X1 U14500 ( .B1(n12078), .B2(n12077), .A(n12114), .ZN(n12083) );
  INV_X1 U14501 ( .A(n12079), .ZN(n12080) );
  OAI21_X1 U14502 ( .B1(n12083), .B2(n12082), .A(n12116), .ZN(n12084) );
  NAND2_X1 U14503 ( .A1(n12084), .A2(n13042), .ZN(n12090) );
  NOR2_X1 U14504 ( .A1(n13085), .A2(n12085), .ZN(n12086) );
  AOI211_X1 U14505 ( .C1(n13061), .C2(n12088), .A(n12087), .B(n12086), .ZN(
        n12089) );
  OAI211_X1 U14506 ( .C1(n12091), .C2(n13049), .A(n12090), .B(n12089), .ZN(
        P2_U3196) );
  OR2_X1 U14507 ( .A1(n12095), .A2(n12094), .ZN(n12092) );
  NAND2_X1 U14508 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  XNOR2_X1 U14509 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n12099) );
  XNOR2_X1 U14510 ( .A(n15163), .B(n12099), .ZN(n12100) );
  NAND2_X1 U14511 ( .A1(n12101), .A2(n12100), .ZN(n15165) );
  INV_X1 U14512 ( .A(n15165), .ZN(n12106) );
  INV_X1 U14513 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n12102) );
  INV_X1 U14514 ( .A(n12103), .ZN(n12104) );
  OAI21_X1 U14515 ( .B1(n12104), .B2(n12106), .A(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n12105) );
  OAI21_X1 U14516 ( .B1(n12106), .B2(n15166), .A(n12105), .ZN(SUB_1596_U65) );
  INV_X1 U14517 ( .A(n12107), .ZN(n12113) );
  INV_X1 U14518 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12465) );
  MUX2_X1 U14519 ( .A(n12465), .B(n12108), .S(n15472), .Z(n12112) );
  AOI22_X1 U14520 ( .A1(n12110), .A2(n12787), .B1(n15488), .B2(n12109), .ZN(
        n12111) );
  OAI211_X1 U14521 ( .C1(n12113), .C2(n12790), .A(n12112), .B(n12111), .ZN(
        P3_U3220) );
  INV_X1 U14522 ( .A(n12114), .ZN(n12115) );
  NAND2_X1 U14523 ( .A1(n13344), .A2(n13542), .ZN(n12211) );
  XNOR2_X1 U14524 ( .A(n13839), .B(n7171), .ZN(n12213) );
  XOR2_X1 U14525 ( .A(n12211), .B(n12213), .Z(n12210) );
  XNOR2_X1 U14526 ( .A(n12209), .B(n12210), .ZN(n12122) );
  NOR2_X1 U14527 ( .A1(n13085), .A2(n13730), .ZN(n12120) );
  NAND2_X1 U14528 ( .A1(n13083), .A2(n13721), .ZN(n12118) );
  OAI211_X1 U14529 ( .C1(n13081), .C2(n13677), .A(n12118), .B(n12117), .ZN(
        n12119) );
  AOI211_X1 U14530 ( .C1(n13839), .C2(n13087), .A(n12120), .B(n12119), .ZN(
        n12121) );
  OAI21_X1 U14531 ( .B1(n12122), .B2(n13089), .A(n12121), .ZN(P2_U3206) );
  INV_X1 U14532 ( .A(n12123), .ZN(n12124) );
  OAI222_X1 U14533 ( .A1(n12941), .A2(n12126), .B1(P3_U3151), .B2(n12125), 
        .C1(n12948), .C2(n12124), .ZN(P3_U3267) );
  INV_X1 U14534 ( .A(n13239), .ZN(n12291) );
  OAI222_X1 U14535 ( .A1(n9480), .A2(P2_U3088), .B1(n13913), .B2(n12291), .C1(
        n13240), .C2(n13916), .ZN(P2_U3298) );
  XNOR2_X1 U14536 ( .A(n12130), .B(n12129), .ZN(n12134) );
  INV_X1 U14537 ( .A(n12135), .ZN(n12136) );
  AOI21_X1 U14538 ( .B1(n7453), .B2(n14449), .A(n10283), .ZN(n12139) );
  INV_X1 U14539 ( .A(n14715), .ZN(n12141) );
  NOR2_X1 U14540 ( .A1(n12143), .A2(n15460), .ZN(n12189) );
  OAI21_X1 U14541 ( .B1(n12844), .B2(n12189), .A(n15472), .ZN(n12609) );
  NAND2_X1 U14542 ( .A1(n15493), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12144) );
  OAI211_X1 U14543 ( .C1(n12848), .C2(n12726), .A(n12609), .B(n12144), .ZN(
        P3_U3203) );
  NAND2_X1 U14544 ( .A1(n12844), .A2(n15514), .ZN(n12791) );
  NAND2_X1 U14545 ( .A1(n9433), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12145) );
  OAI211_X1 U14546 ( .C1(n12848), .C2(n12821), .A(n12791), .B(n12145), .ZN(
        P3_U3489) );
  NAND2_X1 U14547 ( .A1(n12146), .A2(n14545), .ZN(n12147) );
  OAI211_X1 U14548 ( .C1(n12150), .C2(n14545), .A(n12149), .B(n15308), .ZN(
        n12152) );
  OAI22_X1 U14549 ( .A1(n14042), .A2(n15310), .B1(n14251), .B2(n15312), .ZN(
        n14211) );
  INV_X1 U14550 ( .A(n14211), .ZN(n12151) );
  NAND2_X1 U14551 ( .A1(n12152), .A2(n12151), .ZN(n15004) );
  OAI21_X1 U14552 ( .B1(n14777), .B2(n14214), .A(n15240), .ZN(n12153) );
  OR2_X1 U14553 ( .A1(n14747), .A2(n12153), .ZN(n15003) );
  INV_X1 U14554 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n12154) );
  OAI22_X1 U14555 ( .A1(n14209), .A2(n15236), .B1(n12154), .B2(n14798), .ZN(
        n12155) );
  AOI21_X1 U14556 ( .B1(n15006), .B2(n14971), .A(n12155), .ZN(n12156) );
  OAI21_X1 U14557 ( .B1(n15003), .B2(n14974), .A(n12156), .ZN(n12157) );
  AOI21_X1 U14558 ( .B1(n15004), .B2(n14798), .A(n12157), .ZN(n12158) );
  OAI21_X1 U14559 ( .B1(n14978), .B2(n15008), .A(n12158), .ZN(P1_U3269) );
  INV_X1 U14560 ( .A(n14300), .ZN(n14291) );
  INV_X1 U14561 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U14562 ( .A1(n14355), .A2(n10286), .ZN(n12163) );
  OR2_X1 U14563 ( .A1(n15311), .A2(n14052), .ZN(n12162) );
  NAND2_X1 U14564 ( .A1(n12163), .A2(n12162), .ZN(n12172) );
  INV_X1 U14565 ( .A(n12172), .ZN(n12173) );
  NAND2_X1 U14566 ( .A1(n6564), .A2(n12173), .ZN(n12170) );
  OAI21_X1 U14567 ( .B1(n6564), .B2(n12173), .A(n12170), .ZN(n14216) );
  NAND2_X1 U14568 ( .A1(n14355), .A2(n10284), .ZN(n12165) );
  OR2_X1 U14569 ( .A1(n15311), .A2(n14020), .ZN(n12164) );
  NAND2_X1 U14570 ( .A1(n12165), .A2(n12164), .ZN(n12166) );
  XNOR2_X1 U14571 ( .A(n12166), .B(n14111), .ZN(n14217) );
  NOR2_X1 U14572 ( .A1(n14216), .A2(n14217), .ZN(n14215) );
  OAI22_X1 U14573 ( .A1(n14359), .A2(n14011), .B1(n14360), .B2(n14020), .ZN(
        n12167) );
  XNOR2_X1 U14574 ( .A(n12167), .B(n14111), .ZN(n12169) );
  OAI22_X1 U14575 ( .A1(n14359), .A2(n14020), .B1(n14360), .B2(n14052), .ZN(
        n12168) );
  NOR2_X1 U14576 ( .A1(n12169), .A2(n12168), .ZN(n13932) );
  AOI21_X1 U14577 ( .B1(n12169), .B2(n12168), .A(n13932), .ZN(n12175) );
  INV_X1 U14578 ( .A(n12170), .ZN(n12171) );
  NOR3_X1 U14579 ( .A1(n14215), .A2(n12175), .A3(n12171), .ZN(n12179) );
  INV_X1 U14580 ( .A(n14217), .ZN(n12174) );
  INV_X1 U14581 ( .A(n13934), .ZN(n12178) );
  OAI21_X1 U14582 ( .B1(n12179), .B2(n12178), .A(n14281), .ZN(n12185) );
  OAI21_X1 U14583 ( .B1(n14286), .B2(n12181), .A(n12180), .ZN(n12183) );
  NOR2_X1 U14584 ( .A1(n14272), .A2(n14364), .ZN(n12182) );
  AOI211_X1 U14585 ( .C1(n14275), .C2(n15106), .A(n12183), .B(n12182), .ZN(
        n12184) );
  OAI211_X1 U14586 ( .C1(n14359), .C2(n14291), .A(n12185), .B(n12184), .ZN(
        P1_U3217) );
  NAND2_X1 U14587 ( .A1(n12186), .A2(n15472), .ZN(n12191) );
  NOR2_X1 U14588 ( .A1(n12187), .A2(n12726), .ZN(n12188) );
  AOI211_X1 U14589 ( .C1(n15493), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12189), 
        .B(n12188), .ZN(n12190) );
  OAI211_X1 U14590 ( .C1(n12192), .C2(n12790), .A(n12191), .B(n12190), .ZN(
        P3_U3204) );
  INV_X1 U14591 ( .A(n12193), .ZN(n12194) );
  NOR2_X1 U14592 ( .A1(n12194), .A2(SI_29_), .ZN(n12195) );
  MUX2_X1 U14593 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7434), .Z(n12198) );
  NAND2_X1 U14594 ( .A1(n12198), .A2(SI_30_), .ZN(n13257) );
  OAI21_X1 U14595 ( .B1(n12198), .B2(SI_30_), .A(n13257), .ZN(n12201) );
  INV_X1 U14596 ( .A(n12201), .ZN(n12199) );
  NAND2_X1 U14597 ( .A1(n12200), .A2(n12199), .ZN(n13258) );
  INV_X1 U14598 ( .A(n12200), .ZN(n12202) );
  OAI222_X1 U14599 ( .A1(n15147), .A2(n14464), .B1(n12203), .B2(P1_U3086), 
        .C1(n14465), .C2(n15144), .ZN(P1_U3325) );
  OAI222_X1 U14600 ( .A1(n12204), .A2(P2_U3088), .B1(n13913), .B2(n14464), 
        .C1(n15631), .C2(n13916), .ZN(P2_U3297) );
  INV_X1 U14601 ( .A(n12269), .ZN(n13914) );
  INV_X1 U14602 ( .A(n12206), .ZN(n12207) );
  OAI222_X1 U14603 ( .A1(n12941), .A2(n12208), .B1(n12948), .B2(n12207), .C1(
        n7895), .C2(P3_U3151), .ZN(P3_U3265) );
  INV_X1 U14604 ( .A(n12211), .ZN(n12212) );
  NAND2_X1 U14605 ( .A1(n12213), .A2(n12212), .ZN(n12960) );
  XNOR2_X1 U14606 ( .A(n13707), .B(n7171), .ZN(n12216) );
  AND2_X1 U14607 ( .A1(n13724), .A2(n13542), .ZN(n12217) );
  NAND2_X1 U14608 ( .A1(n12216), .A2(n12217), .ZN(n12959) );
  XNOR2_X1 U14609 ( .A(n13180), .B(n7171), .ZN(n12222) );
  AND2_X1 U14610 ( .A1(n13641), .A2(n13542), .ZN(n12221) );
  NOR2_X1 U14611 ( .A1(n12222), .A2(n12221), .ZN(n12215) );
  XNOR2_X1 U14612 ( .A(n13828), .B(n6425), .ZN(n13009) );
  INV_X1 U14613 ( .A(n12215), .ZN(n13013) );
  AND2_X1 U14614 ( .A1(n13343), .A2(n13542), .ZN(n13078) );
  NAND2_X1 U14615 ( .A1(n13013), .A2(n13078), .ZN(n12223) );
  OAI21_X1 U14616 ( .B1(n12215), .B2(n13009), .A(n12223), .ZN(n12220) );
  INV_X1 U14617 ( .A(n12216), .ZN(n12219) );
  INV_X1 U14618 ( .A(n12217), .ZN(n12218) );
  NAND2_X1 U14619 ( .A1(n12219), .A2(n12218), .ZN(n13006) );
  NAND2_X1 U14620 ( .A1(n12222), .A2(n12221), .ZN(n13012) );
  OAI21_X1 U14621 ( .B1(n12223), .B2(n13009), .A(n13012), .ZN(n12224) );
  XNOR2_X1 U14622 ( .A(n13819), .B(n6425), .ZN(n12227) );
  NAND2_X1 U14623 ( .A1(n13342), .A2(n12272), .ZN(n12226) );
  NAND2_X1 U14624 ( .A1(n12227), .A2(n12226), .ZN(n12230) );
  OAI21_X1 U14625 ( .B1(n12227), .B2(n12226), .A(n12230), .ZN(n13025) );
  INV_X1 U14626 ( .A(n13025), .ZN(n12228) );
  NAND2_X1 U14627 ( .A1(n13642), .A2(n12272), .ZN(n12232) );
  XNOR2_X1 U14628 ( .A(n13814), .B(n7171), .ZN(n12231) );
  XOR2_X1 U14629 ( .A(n12232), .B(n12231), .Z(n13058) );
  XNOR2_X1 U14630 ( .A(n13809), .B(n6425), .ZN(n12234) );
  NAND2_X1 U14631 ( .A1(n13598), .A2(n12272), .ZN(n12233) );
  NAND2_X1 U14632 ( .A1(n12234), .A2(n12233), .ZN(n12235) );
  OAI21_X1 U14633 ( .B1(n12234), .B2(n12233), .A(n12235), .ZN(n12984) );
  AND2_X1 U14634 ( .A1(n13341), .A2(n13542), .ZN(n12237) );
  XNOR2_X1 U14635 ( .A(n13804), .B(n7171), .ZN(n12236) );
  NOR2_X1 U14636 ( .A1(n12236), .A2(n12237), .ZN(n12238) );
  AOI21_X1 U14637 ( .B1(n12237), .B2(n12236), .A(n12238), .ZN(n13041) );
  INV_X1 U14638 ( .A(n12238), .ZN(n12239) );
  NAND2_X1 U14639 ( .A1(n13599), .A2(n12272), .ZN(n12240) );
  XNOR2_X1 U14640 ( .A(n13587), .B(n7171), .ZN(n12242) );
  XOR2_X1 U14641 ( .A(n12240), .B(n12242), .Z(n12990) );
  INV_X1 U14642 ( .A(n12240), .ZN(n12241) );
  XNOR2_X1 U14643 ( .A(n13792), .B(n7171), .ZN(n12247) );
  INV_X1 U14644 ( .A(n13051), .ZN(n12245) );
  XNOR2_X1 U14645 ( .A(n13880), .B(n7171), .ZN(n12973) );
  AND2_X1 U14646 ( .A1(n13340), .A2(n13542), .ZN(n12970) );
  OAI21_X1 U14647 ( .B1(n12973), .B2(n13561), .A(n12970), .ZN(n12243) );
  INV_X1 U14648 ( .A(n12243), .ZN(n12244) );
  NAND2_X1 U14649 ( .A1(n12245), .A2(n12244), .ZN(n12253) );
  INV_X1 U14650 ( .A(n12973), .ZN(n12246) );
  AND2_X1 U14651 ( .A1(n13561), .A2(n13542), .ZN(n12249) );
  INV_X1 U14652 ( .A(n12249), .ZN(n12972) );
  NOR2_X1 U14653 ( .A1(n12973), .A2(n12249), .ZN(n12250) );
  XNOR2_X1 U14654 ( .A(n13535), .B(n12214), .ZN(n12256) );
  NAND2_X1 U14655 ( .A1(n13339), .A2(n12272), .ZN(n12254) );
  XNOR2_X1 U14656 ( .A(n12256), .B(n12254), .ZN(n13032) );
  NAND2_X1 U14657 ( .A1(n13031), .A2(n13032), .ZN(n12258) );
  INV_X1 U14658 ( .A(n12254), .ZN(n12255) );
  NAND2_X1 U14659 ( .A1(n12256), .A2(n12255), .ZN(n12257) );
  NAND2_X1 U14660 ( .A1(n12258), .A2(n12257), .ZN(n12998) );
  XNOR2_X1 U14661 ( .A(n13521), .B(n12214), .ZN(n12261) );
  NAND2_X1 U14662 ( .A1(n13338), .A2(n12272), .ZN(n12259) );
  XNOR2_X1 U14663 ( .A(n12261), .B(n12259), .ZN(n12999) );
  INV_X1 U14664 ( .A(n12259), .ZN(n12260) );
  NAND2_X1 U14665 ( .A1(n12261), .A2(n12260), .ZN(n12262) );
  XNOR2_X1 U14666 ( .A(n13771), .B(n6425), .ZN(n12264) );
  NAND2_X1 U14667 ( .A1(n13337), .A2(n12272), .ZN(n12263) );
  NAND2_X1 U14668 ( .A1(n12264), .A2(n12263), .ZN(n12265) );
  OAI21_X1 U14669 ( .B1(n12264), .B2(n12263), .A(n12265), .ZN(n13070) );
  NAND2_X1 U14670 ( .A1(n13449), .A2(n12272), .ZN(n12267) );
  XNOR2_X1 U14671 ( .A(n13491), .B(n12214), .ZN(n12266) );
  XOR2_X1 U14672 ( .A(n12267), .B(n12266), .Z(n12953) );
  INV_X1 U14673 ( .A(n12266), .ZN(n12268) );
  NAND2_X1 U14674 ( .A1(n12269), .A2(n13262), .ZN(n12271) );
  NAND2_X1 U14675 ( .A1(n6400), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U14676 ( .A1(n13456), .A2(n12272), .ZN(n12273) );
  XNOR2_X1 U14677 ( .A(n12273), .B(n12214), .ZN(n12274) );
  XNOR2_X1 U14678 ( .A(n13765), .B(n12274), .ZN(n12275) );
  INV_X1 U14679 ( .A(n12276), .ZN(n13484) );
  NOR2_X1 U14680 ( .A1(n13484), .A2(n13085), .ZN(n12286) );
  INV_X1 U14681 ( .A(n13463), .ZN(n12283) );
  INV_X1 U14682 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13462) );
  NAND2_X1 U14683 ( .A1(n12277), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n12280) );
  NAND2_X1 U14684 ( .A1(n12278), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n12279) );
  OAI211_X1 U14685 ( .C1(n13462), .C2(n9814), .A(n12280), .B(n12279), .ZN(
        n12281) );
  AOI21_X1 U14686 ( .B1(n12283), .B2(n12282), .A(n12281), .ZN(n13477) );
  AOI22_X1 U14687 ( .A1(n13449), .A2(n13083), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12284) );
  OAI21_X1 U14688 ( .B1(n13477), .B2(n13081), .A(n12284), .ZN(n12285) );
  AOI211_X1 U14689 ( .C1(n13765), .C2(n13087), .A(n12286), .B(n12285), .ZN(
        n12287) );
  OAI21_X1 U14690 ( .B1(n12288), .B2(n13089), .A(n12287), .ZN(P2_U3192) );
  OAI222_X1 U14691 ( .A1(n15147), .A2(n12291), .B1(n12290), .B2(P1_U3086), 
        .C1(n12289), .C2(n15144), .ZN(P1_U3326) );
  XNOR2_X1 U14692 ( .A(n12793), .B(n11174), .ZN(n12292) );
  NOR2_X1 U14693 ( .A1(n12292), .A2(n12637), .ZN(n12350) );
  AOI21_X1 U14694 ( .B1(n12292), .B2(n12637), .A(n12350), .ZN(n12322) );
  XNOR2_X1 U14695 ( .A(n12686), .B(n6610), .ZN(n12328) );
  XNOR2_X1 U14696 ( .A(n12902), .B(n6610), .ZN(n12379) );
  INV_X1 U14697 ( .A(n12379), .ZN(n12297) );
  INV_X1 U14698 ( .A(n12295), .ZN(n12296) );
  XNOR2_X1 U14699 ( .A(n12392), .B(n6610), .ZN(n12298) );
  XNOR2_X1 U14700 ( .A(n12298), .B(n12759), .ZN(n12389) );
  XNOR2_X1 U14701 ( .A(n12738), .B(n6610), .ZN(n12299) );
  XNOR2_X1 U14702 ( .A(n12299), .B(n12452), .ZN(n12425) );
  INV_X1 U14703 ( .A(n12299), .ZN(n12300) );
  XNOR2_X1 U14704 ( .A(n12893), .B(n6610), .ZN(n12301) );
  XNOR2_X1 U14705 ( .A(n12301), .B(n12732), .ZN(n12343) );
  INV_X1 U14706 ( .A(n12301), .ZN(n12302) );
  XNOR2_X1 U14707 ( .A(n12884), .B(n6610), .ZN(n12303) );
  XNOR2_X1 U14708 ( .A(n12303), .B(n12694), .ZN(n12409) );
  INV_X1 U14709 ( .A(n12303), .ZN(n12304) );
  XNOR2_X1 U14710 ( .A(n12879), .B(n11174), .ZN(n12305) );
  NOR2_X1 U14711 ( .A1(n12305), .A2(n12705), .ZN(n12306) );
  AOI21_X1 U14712 ( .B1(n12305), .B2(n12705), .A(n12306), .ZN(n12364) );
  INV_X1 U14713 ( .A(n12306), .ZN(n12307) );
  NAND2_X1 U14714 ( .A1(n12362), .A2(n12307), .ZN(n12329) );
  OAI21_X1 U14715 ( .B1(n12419), .B2(n12328), .A(n12329), .ZN(n12311) );
  XNOR2_X1 U14716 ( .A(n12340), .B(n6610), .ZN(n12334) );
  AOI22_X1 U14717 ( .A1(n12334), .A2(n12682), .B1(n12419), .B2(n12328), .ZN(
        n12310) );
  NOR2_X1 U14718 ( .A1(n12334), .A2(n12682), .ZN(n12309) );
  XNOR2_X1 U14719 ( .A(n12406), .B(n6610), .ZN(n12308) );
  NAND2_X1 U14720 ( .A1(n12308), .A2(n12644), .ZN(n12312) );
  OAI21_X1 U14721 ( .B1(n12308), .B2(n12644), .A(n12312), .ZN(n12397) );
  INV_X1 U14722 ( .A(n12312), .ZN(n12372) );
  XNOR2_X1 U14723 ( .A(n12313), .B(n6610), .ZN(n12314) );
  NAND2_X1 U14724 ( .A1(n12314), .A2(n12656), .ZN(n12317) );
  INV_X1 U14725 ( .A(n12314), .ZN(n12315) );
  NAND2_X1 U14726 ( .A1(n12315), .A2(n9352), .ZN(n12316) );
  AND2_X1 U14727 ( .A1(n12317), .A2(n12316), .ZN(n12371) );
  XNOR2_X1 U14728 ( .A(n12449), .B(n6610), .ZN(n12318) );
  NOR2_X1 U14729 ( .A1(n12318), .A2(n12620), .ZN(n12319) );
  AOI21_X1 U14730 ( .B1(n12318), .B2(n12620), .A(n12319), .ZN(n12438) );
  INV_X1 U14731 ( .A(n12319), .ZN(n12320) );
  OAI21_X1 U14732 ( .B1(n12322), .B2(n12321), .A(n12351), .ZN(n12323) );
  NAND2_X1 U14733 ( .A1(n12323), .A2(n12439), .ZN(n12327) );
  AOI22_X1 U14734 ( .A1(n12627), .A2(n12441), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12324) );
  OAI21_X1 U14735 ( .B1(n12645), .B2(n12443), .A(n12324), .ZN(n12325) );
  AOI21_X1 U14736 ( .B1(n12619), .B2(n12445), .A(n12325), .ZN(n12326) );
  OAI211_X1 U14737 ( .C1(n12629), .C2(n12448), .A(n12327), .B(n12326), .ZN(
        P3_U3154) );
  INV_X1 U14738 ( .A(n12328), .ZN(n12331) );
  INV_X1 U14739 ( .A(n12329), .ZN(n12330) );
  AND2_X1 U14740 ( .A1(n12329), .A2(n12328), .ZN(n12332) );
  NAND2_X1 U14741 ( .A1(n12418), .A2(n12419), .ZN(n12417) );
  INV_X1 U14742 ( .A(n12332), .ZN(n12333) );
  NAND2_X1 U14743 ( .A1(n12417), .A2(n12333), .ZN(n12335) );
  NAND2_X1 U14744 ( .A1(n12335), .A2(n12334), .ZN(n12398) );
  AOI22_X1 U14745 ( .A1(n12695), .A2(n12427), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12338) );
  NAND2_X1 U14746 ( .A1(n12671), .A2(n12441), .ZN(n12337) );
  OAI211_X1 U14747 ( .C1(n12644), .C2(n12429), .A(n12338), .B(n12337), .ZN(
        n12339) );
  AOI21_X1 U14748 ( .B1(n12340), .B2(n12414), .A(n12339), .ZN(n12341) );
  OAI21_X1 U14749 ( .B1(n12342), .B2(n12434), .A(n12341), .ZN(P3_U3156) );
  XNOR2_X1 U14750 ( .A(n12344), .B(n12343), .ZN(n12349) );
  NAND2_X1 U14751 ( .A1(n12452), .A2(n12427), .ZN(n12345) );
  NAND2_X1 U14752 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12595)
         );
  OAI211_X1 U14753 ( .C1(n12718), .C2(n12429), .A(n12345), .B(n12595), .ZN(
        n12347) );
  NOR2_X1 U14754 ( .A1(n12893), .A2(n12448), .ZN(n12346) );
  AOI211_X1 U14755 ( .C1(n12724), .C2(n12441), .A(n12347), .B(n12346), .ZN(
        n12348) );
  OAI21_X1 U14756 ( .B1(n12349), .B2(n12434), .A(n12348), .ZN(P3_U3159) );
  XNOR2_X1 U14757 ( .A(n12352), .B(n6610), .ZN(n12353) );
  XNOR2_X1 U14758 ( .A(n12354), .B(n12353), .ZN(n12361) );
  NOR2_X1 U14759 ( .A1(n12355), .A2(n12429), .ZN(n12359) );
  AOI22_X1 U14760 ( .A1(n12613), .A2(n12441), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12356) );
  OAI21_X1 U14761 ( .B1(n12357), .B2(n12443), .A(n12356), .ZN(n12358) );
  AOI211_X1 U14762 ( .C1(n12614), .C2(n12414), .A(n12359), .B(n12358), .ZN(
        n12360) );
  OAI21_X1 U14763 ( .B1(n12361), .B2(n12434), .A(n12360), .ZN(P3_U3160) );
  OAI21_X1 U14764 ( .B1(n12364), .B2(n12363), .A(n12362), .ZN(n12365) );
  NAND2_X1 U14765 ( .A1(n12365), .A2(n12439), .ZN(n12369) );
  AOI22_X1 U14766 ( .A1(n12694), .A2(n12427), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12366) );
  OAI21_X1 U14767 ( .B1(n12419), .B2(n12429), .A(n12366), .ZN(n12367) );
  AOI21_X1 U14768 ( .B1(n12698), .B2(n12441), .A(n12367), .ZN(n12368) );
  OAI211_X1 U14769 ( .C1(n6650), .C2(n12448), .A(n12369), .B(n12368), .ZN(
        P3_U3163) );
  INV_X1 U14770 ( .A(n12370), .ZN(n12374) );
  NOR3_X1 U14771 ( .A1(n12402), .A2(n12372), .A3(n12371), .ZN(n12373) );
  OAI21_X1 U14772 ( .B1(n12374), .B2(n12373), .A(n12439), .ZN(n12378) );
  AOI22_X1 U14773 ( .A1(n12649), .A2(n12441), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12375) );
  OAI21_X1 U14774 ( .B1(n12644), .B2(n12443), .A(n12375), .ZN(n12376) );
  AOI21_X1 U14775 ( .B1(n12620), .B2(n12445), .A(n12376), .ZN(n12377) );
  OAI211_X1 U14776 ( .C1(n12863), .C2(n12448), .A(n12378), .B(n12377), .ZN(
        P3_U3165) );
  XNOR2_X1 U14777 ( .A(n12379), .B(n12748), .ZN(n12380) );
  XNOR2_X1 U14778 ( .A(n12381), .B(n12380), .ZN(n12388) );
  NAND2_X1 U14779 ( .A1(n12759), .A2(n12445), .ZN(n12382) );
  NAND2_X1 U14780 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12545)
         );
  OAI211_X1 U14781 ( .C1(n12383), .C2(n12443), .A(n12382), .B(n12545), .ZN(
        n12386) );
  NOR2_X1 U14782 ( .A1(n12384), .A2(n12448), .ZN(n12385) );
  AOI211_X1 U14783 ( .C1(n12762), .C2(n12441), .A(n12386), .B(n12385), .ZN(
        n12387) );
  OAI21_X1 U14784 ( .B1(n12388), .B2(n12434), .A(n12387), .ZN(P3_U3166) );
  XNOR2_X1 U14785 ( .A(n12390), .B(n12389), .ZN(n12396) );
  NAND2_X1 U14786 ( .A1(n12427), .A2(n12770), .ZN(n12391) );
  NAND2_X1 U14787 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12557)
         );
  OAI211_X1 U14788 ( .C1(n12749), .C2(n12429), .A(n12391), .B(n12557), .ZN(
        n12394) );
  NOR2_X1 U14789 ( .A1(n12392), .A2(n12448), .ZN(n12393) );
  AOI211_X1 U14790 ( .C1(n12750), .C2(n12441), .A(n12394), .B(n12393), .ZN(
        n12395) );
  OAI21_X1 U14791 ( .B1(n12396), .B2(n12434), .A(n12395), .ZN(P3_U3168) );
  INV_X1 U14792 ( .A(n12397), .ZN(n12400) );
  INV_X1 U14793 ( .A(n12398), .ZN(n12399) );
  AOI22_X1 U14794 ( .A1(n9350), .A2(n12427), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12404) );
  NAND2_X1 U14795 ( .A1(n12659), .A2(n12441), .ZN(n12403) );
  OAI211_X1 U14796 ( .C1(n12656), .C2(n12429), .A(n12404), .B(n12403), .ZN(
        n12405) );
  AOI21_X1 U14797 ( .B1(n12406), .B2(n12414), .A(n12405), .ZN(n12407) );
  NAND2_X1 U14798 ( .A1(n12408), .A2(n12407), .ZN(P3_U3169) );
  XNOR2_X1 U14799 ( .A(n12410), .B(n12409), .ZN(n12416) );
  AOI22_X1 U14800 ( .A1(n12732), .A2(n12427), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12412) );
  NAND2_X1 U14801 ( .A1(n12708), .A2(n12441), .ZN(n12411) );
  OAI211_X1 U14802 ( .C1(n12681), .C2(n12429), .A(n12412), .B(n12411), .ZN(
        n12413) );
  AOI21_X1 U14803 ( .B1(n12884), .B2(n12414), .A(n12413), .ZN(n12415) );
  OAI21_X1 U14804 ( .B1(n12416), .B2(n12434), .A(n12415), .ZN(P3_U3173) );
  OAI21_X1 U14805 ( .B1(n12419), .B2(n12418), .A(n12417), .ZN(n12420) );
  NAND2_X1 U14806 ( .A1(n12420), .A2(n12439), .ZN(n12424) );
  AOI22_X1 U14807 ( .A1(n12705), .A2(n12427), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12421) );
  OAI21_X1 U14808 ( .B1(n12682), .B2(n12429), .A(n12421), .ZN(n12422) );
  AOI21_X1 U14809 ( .B1(n12685), .B2(n12441), .A(n12422), .ZN(n12423) );
  OAI211_X1 U14810 ( .C1(n12873), .C2(n12448), .A(n12424), .B(n12423), .ZN(
        P3_U3175) );
  XNOR2_X1 U14811 ( .A(n12426), .B(n12425), .ZN(n12435) );
  NAND2_X1 U14812 ( .A1(n12759), .A2(n12427), .ZN(n12428) );
  NAND2_X1 U14813 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12579)
         );
  OAI211_X1 U14814 ( .C1(n12430), .C2(n12429), .A(n12428), .B(n12579), .ZN(
        n12432) );
  INV_X1 U14815 ( .A(n12738), .ZN(n12826) );
  NOR2_X1 U14816 ( .A1(n12826), .A2(n12448), .ZN(n12431) );
  AOI211_X1 U14817 ( .C1(n12734), .C2(n12441), .A(n12432), .B(n12431), .ZN(
        n12433) );
  OAI21_X1 U14818 ( .B1(n12435), .B2(n12434), .A(n12433), .ZN(P3_U3178) );
  OAI21_X1 U14819 ( .B1(n12438), .B2(n12437), .A(n12436), .ZN(n12440) );
  NAND2_X1 U14820 ( .A1(n12440), .A2(n12439), .ZN(n12447) );
  AOI22_X1 U14821 ( .A1(n12640), .A2(n12441), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12442) );
  OAI21_X1 U14822 ( .B1(n12656), .B2(n12443), .A(n12442), .ZN(n12444) );
  AOI21_X1 U14823 ( .B1(n12637), .B2(n12445), .A(n12444), .ZN(n12446) );
  OAI211_X1 U14824 ( .C1(n12449), .C2(n12448), .A(n12447), .B(n12446), .ZN(
        P3_U3180) );
  MUX2_X1 U14825 ( .A(n12450), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12453), .Z(
        P3_U3522) );
  MUX2_X1 U14826 ( .A(n12451), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12453), .Z(
        P3_U3521) );
  MUX2_X1 U14827 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12619), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14828 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12637), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14829 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12620), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14830 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n9352), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14831 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12668), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14832 ( .A(n9350), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12453), .Z(
        P3_U3514) );
  MUX2_X1 U14833 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12695), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14834 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12705), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14835 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12694), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14836 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12732), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14837 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12452), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14838 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12759), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14839 ( .A(n12770), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12453), .Z(
        P3_U3507) );
  MUX2_X1 U14840 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12782), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14841 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12769), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14842 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12781), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14843 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12454), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14844 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12455), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14845 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12456), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14846 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12457), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14847 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12458), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14848 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12459), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14849 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12460), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14850 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15480), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14851 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12461), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14852 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15481), .S(P3_U3897), .Z(
        P3_U3491) );
  OAI21_X1 U14853 ( .B1(n6415), .B2(n12478), .A(n12463), .ZN(n12464) );
  AOI21_X1 U14854 ( .B1(n12465), .B2(n12464), .A(n12492), .ZN(n12483) );
  OAI21_X1 U14855 ( .B1(n12581), .B2(n12467), .A(n12466), .ZN(n12475) );
  NAND2_X1 U14856 ( .A1(n12468), .A2(n12476), .ZN(n12471) );
  MUX2_X1 U14857 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12937), .Z(n12484) );
  XNOR2_X1 U14858 ( .A(n12484), .B(n12498), .ZN(n12470) );
  AOI21_X1 U14859 ( .B1(n12472), .B2(n12471), .A(n12470), .ZN(n12469) );
  INV_X1 U14860 ( .A(n12469), .ZN(n12473) );
  NAND3_X1 U14861 ( .A1(n12472), .A2(n12471), .A3(n12470), .ZN(n12490) );
  AOI21_X1 U14862 ( .B1(n12473), .B2(n12490), .A(n12605), .ZN(n12474) );
  AOI211_X1 U14863 ( .C1(n12578), .C2(n12498), .A(n12475), .B(n12474), .ZN(
        n12482) );
  NAND2_X1 U14864 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n12479), .ZN(n12499) );
  OAI21_X1 U14865 ( .B1(n12479), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12499), 
        .ZN(n12480) );
  NAND2_X1 U14866 ( .A1(n12480), .A2(n12607), .ZN(n12481) );
  OAI211_X1 U14867 ( .C1(n12483), .C2(n12566), .A(n12482), .B(n12481), .ZN(
        P3_U3195) );
  INV_X1 U14868 ( .A(n12484), .ZN(n12485) );
  NAND2_X1 U14869 ( .A1(n12485), .A2(n12498), .ZN(n12489) );
  NAND2_X1 U14870 ( .A1(n12505), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12518) );
  OR2_X1 U14871 ( .A1(n12505), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12486) );
  AND2_X1 U14872 ( .A1(n12518), .A2(n12486), .ZN(n12493) );
  NAND2_X1 U14873 ( .A1(n12505), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12519) );
  OR2_X1 U14874 ( .A1(n12505), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12487) );
  AND2_X1 U14875 ( .A1(n12519), .A2(n12487), .ZN(n12502) );
  MUX2_X1 U14876 ( .A(n12493), .B(n12502), .S(n12937), .Z(n12488) );
  AOI21_X1 U14877 ( .B1(n12490), .B2(n12489), .A(n12488), .ZN(n12512) );
  NAND3_X1 U14878 ( .A1(n12490), .A2(n12489), .A3(n12488), .ZN(n12521) );
  NAND2_X1 U14879 ( .A1(n12521), .A2(n12491), .ZN(n12511) );
  INV_X1 U14880 ( .A(n12513), .ZN(n12496) );
  NOR3_X1 U14881 ( .A1(n12494), .A2(n12493), .A3(n12492), .ZN(n12495) );
  OAI21_X1 U14882 ( .B1(n12496), .B2(n12495), .A(n12590), .ZN(n12510) );
  OR2_X1 U14883 ( .A1(n12498), .A2(n12497), .ZN(n12500) );
  NAND2_X1 U14884 ( .A1(n12500), .A2(n12499), .ZN(n12501) );
  NAND2_X1 U14885 ( .A1(n12502), .A2(n12501), .ZN(n12515) );
  OAI21_X1 U14886 ( .B1(n12502), .B2(n12501), .A(n12515), .ZN(n12508) );
  OAI21_X1 U14887 ( .B1(n12581), .B2(n12504), .A(n12503), .ZN(n12507) );
  NOR2_X1 U14888 ( .A1(n12597), .A2(n12505), .ZN(n12506) );
  AOI211_X1 U14889 ( .C1(n12607), .C2(n12508), .A(n12507), .B(n12506), .ZN(
        n12509) );
  OAI211_X1 U14890 ( .C1(n12512), .C2(n12511), .A(n12510), .B(n12509), .ZN(
        P3_U3196) );
  INV_X1 U14891 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12772) );
  AOI21_X1 U14892 ( .B1(n12772), .B2(n12514), .A(n6426), .ZN(n12529) );
  NAND2_X1 U14893 ( .A1(n12519), .A2(n12515), .ZN(n12540) );
  XOR2_X1 U14894 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12542), .Z(n12527) );
  NAND2_X1 U14895 ( .A1(n15455), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n12516) );
  OAI211_X1 U14896 ( .C1(n12597), .C2(n12531), .A(n12517), .B(n12516), .ZN(
        n12526) );
  MUX2_X1 U14897 ( .A(n12519), .B(n12518), .S(n11473), .Z(n12520) );
  NAND2_X1 U14898 ( .A1(n12521), .A2(n12520), .ZN(n12530) );
  XNOR2_X1 U14899 ( .A(n12530), .B(n12531), .ZN(n12523) );
  MUX2_X1 U14900 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12937), .Z(n12522) );
  AOI21_X1 U14901 ( .B1(n12523), .B2(n12522), .A(n12532), .ZN(n12524) );
  NOR2_X1 U14902 ( .A1(n12524), .A2(n12605), .ZN(n12525) );
  AOI211_X1 U14903 ( .C1(n12607), .C2(n12527), .A(n12526), .B(n12525), .ZN(
        n12528) );
  OAI21_X1 U14904 ( .B1(n12529), .B2(n12566), .A(n12528), .ZN(P3_U3197) );
  INV_X1 U14905 ( .A(n12530), .ZN(n12533) );
  INV_X1 U14906 ( .A(n12531), .ZN(n12541) );
  INV_X1 U14907 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12761) );
  MUX2_X1 U14908 ( .A(n12761), .B(n12832), .S(n12937), .Z(n12534) );
  NOR2_X1 U14909 ( .A1(n12555), .A2(n12534), .ZN(n12558) );
  NOR2_X1 U14910 ( .A1(n12558), .A2(n6580), .ZN(n12535) );
  XNOR2_X1 U14911 ( .A(n12559), .B(n12535), .ZN(n12551) );
  XNOR2_X1 U14912 ( .A(n12555), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n12537) );
  NOR3_X1 U14913 ( .A1(n6426), .A2(n12538), .A3(n12537), .ZN(n12539) );
  OAI21_X1 U14914 ( .B1(n6490), .B2(n12539), .A(n12590), .ZN(n12550) );
  XNOR2_X1 U14915 ( .A(n12555), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12543) );
  OAI21_X1 U14916 ( .B1(n12544), .B2(n12543), .A(n12554), .ZN(n12548) );
  INV_X1 U14917 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15170) );
  NAND2_X1 U14918 ( .A1(n12578), .A2(n12555), .ZN(n12546) );
  OAI211_X1 U14919 ( .C1(n12581), .C2(n15170), .A(n12546), .B(n12545), .ZN(
        n12547) );
  AOI21_X1 U14920 ( .B1(n12607), .B2(n12548), .A(n12547), .ZN(n12549) );
  OAI211_X1 U14921 ( .C1(n12605), .C2(n12551), .A(n12550), .B(n12549), .ZN(
        P3_U3198) );
  INV_X1 U14922 ( .A(n12574), .ZN(n12552) );
  AOI21_X1 U14923 ( .B1(n12752), .B2(n12553), .A(n12552), .ZN(n12567) );
  XNOR2_X1 U14924 ( .A(n12577), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n12564) );
  NAND2_X1 U14925 ( .A1(n15455), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12556) );
  OAI211_X1 U14926 ( .C1(n12597), .C2(n12576), .A(n12557), .B(n12556), .ZN(
        n12563) );
  MUX2_X1 U14927 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12937), .Z(n12568) );
  XNOR2_X1 U14928 ( .A(n12576), .B(n12568), .ZN(n12561) );
  AOI211_X1 U14929 ( .C1(n12561), .C2(n12560), .A(n12605), .B(n6496), .ZN(
        n12562) );
  AOI211_X1 U14930 ( .C1(n12607), .C2(n12564), .A(n12563), .B(n12562), .ZN(
        n12565) );
  OAI21_X1 U14931 ( .B1(n12567), .B2(n12566), .A(n12565), .ZN(P3_U3199) );
  MUX2_X1 U14932 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12937), .Z(n12570) );
  XNOR2_X1 U14933 ( .A(n12600), .B(n12599), .ZN(n12569) );
  NOR2_X1 U14934 ( .A1(n12569), .A2(n12570), .ZN(n12598) );
  AOI21_X1 U14935 ( .B1(n12570), .B2(n12569), .A(n12598), .ZN(n12586) );
  OR2_X1 U14936 ( .A1(n12599), .A2(n12735), .ZN(n12587) );
  NAND2_X1 U14937 ( .A1(n12599), .A2(n12735), .ZN(n12571) );
  NAND2_X1 U14938 ( .A1(n12587), .A2(n12571), .ZN(n12572) );
  AND3_X1 U14939 ( .A1(n12574), .A2(n12573), .A3(n12572), .ZN(n12575) );
  OAI21_X1 U14940 ( .B1(n12589), .B2(n12575), .A(n12590), .ZN(n12585) );
  XOR2_X1 U14941 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12599), .Z(n12592) );
  XNOR2_X1 U14942 ( .A(n6422), .B(n12592), .ZN(n12583) );
  INV_X1 U14943 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15191) );
  NAND2_X1 U14944 ( .A1(n12578), .A2(n12599), .ZN(n12580) );
  OAI211_X1 U14945 ( .C1(n12581), .C2(n15191), .A(n12580), .B(n12579), .ZN(
        n12582) );
  AOI21_X1 U14946 ( .B1(n12583), .B2(n12607), .A(n12582), .ZN(n12584) );
  OAI211_X1 U14947 ( .C1(n12586), .C2(n12605), .A(n12585), .B(n12584), .ZN(
        P3_U3200) );
  INV_X1 U14948 ( .A(n12587), .ZN(n12588) );
  XNOR2_X1 U14949 ( .A(n12593), .B(n12721), .ZN(n12601) );
  INV_X1 U14950 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12591) );
  XNOR2_X1 U14951 ( .A(n12593), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12602) );
  NAND2_X1 U14952 ( .A1(n15455), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12594) );
  OAI211_X1 U14953 ( .C1(n12597), .C2(n12596), .A(n12595), .B(n12594), .ZN(
        n12606) );
  AOI21_X1 U14954 ( .B1(n12600), .B2(n12599), .A(n12598), .ZN(n12604) );
  MUX2_X1 U14955 ( .A(n12602), .B(n7676), .S(n11473), .Z(n12603) );
  NAND2_X1 U14956 ( .A1(n15493), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12608) );
  OAI211_X1 U14957 ( .C1(n8548), .C2(n12726), .A(n12609), .B(n12608), .ZN(
        P3_U3202) );
  INV_X1 U14958 ( .A(n12610), .ZN(n12611) );
  AOI22_X1 U14959 ( .A1(n12614), .A2(n12787), .B1(n15488), .B2(n12613), .ZN(
        n12615) );
  OAI211_X1 U14960 ( .C1(n12617), .C2(n12790), .A(n12616), .B(n12615), .ZN(
        P3_U3205) );
  AOI21_X1 U14961 ( .B1(n12626), .B2(n12625), .A(n9390), .ZN(n12796) );
  INV_X1 U14962 ( .A(n12796), .ZN(n12631) );
  AOI22_X1 U14963 ( .A1(n12627), .A2(n15488), .B1(n15493), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12628) );
  OAI21_X1 U14964 ( .B1(n12629), .B2(n12726), .A(n12628), .ZN(n12630) );
  AOI21_X1 U14965 ( .B1(n12631), .B2(n12741), .A(n12630), .ZN(n12632) );
  OAI21_X1 U14966 ( .B1(n12795), .B2(n15493), .A(n12632), .ZN(P3_U3206) );
  XNOR2_X1 U14967 ( .A(n12634), .B(n12633), .ZN(n12859) );
  INV_X1 U14968 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12639) );
  XNOR2_X1 U14969 ( .A(n12635), .B(n12636), .ZN(n12638) );
  AOI222_X1 U14970 ( .A1(n12784), .A2(n12638), .B1(n12637), .B2(n15479), .C1(
        n9352), .C2(n12704), .ZN(n12854) );
  MUX2_X1 U14971 ( .A(n12639), .B(n12854), .S(n15472), .Z(n12642) );
  AOI22_X1 U14972 ( .A1(n12856), .A2(n12787), .B1(n15488), .B2(n12640), .ZN(
        n12641) );
  OAI211_X1 U14973 ( .C1(n12859), .C2(n12790), .A(n12642), .B(n12641), .ZN(
        P3_U3207) );
  INV_X1 U14974 ( .A(n12800), .ZN(n12653) );
  OAI21_X1 U14975 ( .B1(n12648), .B2(n12647), .A(n12646), .ZN(n12801) );
  AOI22_X1 U14976 ( .A1(n12649), .A2(n15488), .B1(n15493), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12650) );
  OAI21_X1 U14977 ( .B1(n12863), .B2(n12726), .A(n12650), .ZN(n12651) );
  AOI21_X1 U14978 ( .B1(n12801), .B2(n12741), .A(n12651), .ZN(n12652) );
  OAI21_X1 U14979 ( .B1(n12653), .B2(n15493), .A(n12652), .ZN(P3_U3208) );
  XOR2_X1 U14980 ( .A(n12654), .B(n12658), .Z(n12655) );
  OAI222_X1 U14981 ( .A1(n15469), .A2(n12656), .B1(n15467), .B2(n12682), .C1(
        n12655), .C2(n15484), .ZN(n12803) );
  INV_X1 U14982 ( .A(n12803), .ZN(n12663) );
  OAI21_X1 U14983 ( .B1(n6479), .B2(n12658), .A(n12657), .ZN(n12804) );
  AOI22_X1 U14984 ( .A1(n12659), .A2(n15488), .B1(n15493), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12660) );
  OAI21_X1 U14985 ( .B1(n12867), .B2(n12726), .A(n12660), .ZN(n12661) );
  AOI21_X1 U14986 ( .B1(n12804), .B2(n12741), .A(n12661), .ZN(n12662) );
  OAI21_X1 U14987 ( .B1(n12663), .B2(n15493), .A(n12662), .ZN(P3_U3209) );
  XNOR2_X1 U14988 ( .A(n12664), .B(n12666), .ZN(n12808) );
  INV_X1 U14989 ( .A(n12808), .ZN(n12675) );
  OAI211_X1 U14990 ( .C1(n12667), .C2(n12666), .A(n12665), .B(n12784), .ZN(
        n12670) );
  AOI22_X1 U14991 ( .A1(n12668), .A2(n15479), .B1(n12704), .B2(n12695), .ZN(
        n12669) );
  NAND2_X1 U14992 ( .A1(n12670), .A2(n12669), .ZN(n12807) );
  AOI22_X1 U14993 ( .A1(n12671), .A2(n15488), .B1(n15493), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12672) );
  OAI21_X1 U14994 ( .B1(n12871), .B2(n12726), .A(n12672), .ZN(n12673) );
  AOI21_X1 U14995 ( .B1(n12807), .B2(n15472), .A(n12673), .ZN(n12674) );
  OAI21_X1 U14996 ( .B1(n12675), .B2(n12790), .A(n12674), .ZN(P3_U3210) );
  XNOR2_X1 U14997 ( .A(n12677), .B(n12676), .ZN(n12874) );
  XNOR2_X1 U14998 ( .A(n12679), .B(n12678), .ZN(n12680) );
  OAI222_X1 U14999 ( .A1(n15469), .A2(n12682), .B1(n15467), .B2(n12681), .C1(
        n15484), .C2(n12680), .ZN(n12872) );
  INV_X1 U15000 ( .A(n12872), .ZN(n12683) );
  MUX2_X1 U15001 ( .A(n12684), .B(n12683), .S(n15472), .Z(n12688) );
  AOI22_X1 U15002 ( .A1(n12686), .A2(n12787), .B1(n15488), .B2(n12685), .ZN(
        n12687) );
  OAI211_X1 U15003 ( .C1(n12874), .C2(n12790), .A(n12688), .B(n12687), .ZN(
        P3_U3211) );
  XNOR2_X1 U15004 ( .A(n12690), .B(n12689), .ZN(n12882) );
  OAI21_X1 U15005 ( .B1(n12693), .B2(n12692), .A(n12691), .ZN(n12696) );
  AOI222_X1 U15006 ( .A1(n12784), .A2(n12696), .B1(n12695), .B2(n15479), .C1(
        n12694), .C2(n12704), .ZN(n12877) );
  MUX2_X1 U15007 ( .A(n12697), .B(n12877), .S(n15472), .Z(n12700) );
  AOI22_X1 U15008 ( .A1(n12879), .A2(n12787), .B1(n15488), .B2(n12698), .ZN(
        n12699) );
  OAI211_X1 U15009 ( .C1(n12882), .C2(n12790), .A(n12700), .B(n12699), .ZN(
        P3_U3212) );
  XNOR2_X1 U15010 ( .A(n12701), .B(n12702), .ZN(n12887) );
  XNOR2_X1 U15011 ( .A(n12703), .B(n12702), .ZN(n12706) );
  AOI222_X1 U15012 ( .A1(n12784), .A2(n12706), .B1(n12705), .B2(n15479), .C1(
        n12732), .C2(n12704), .ZN(n12883) );
  MUX2_X1 U15013 ( .A(n12707), .B(n12883), .S(n15472), .Z(n12710) );
  AOI22_X1 U15014 ( .A1(n12884), .A2(n12787), .B1(n15488), .B2(n12708), .ZN(
        n12709) );
  OAI211_X1 U15015 ( .C1(n12887), .C2(n12790), .A(n12710), .B(n12709), .ZN(
        P3_U3213) );
  INV_X1 U15016 ( .A(n12731), .ZN(n12712) );
  NOR2_X1 U15017 ( .A1(n12712), .A2(n12711), .ZN(n12715) );
  INV_X1 U15018 ( .A(n12715), .ZN(n12730) );
  AOI21_X1 U15019 ( .B1(n12730), .B2(n12713), .A(n12722), .ZN(n12717) );
  NOR2_X1 U15020 ( .A1(n12715), .A2(n12714), .ZN(n12716) );
  NOR3_X1 U15021 ( .A1(n12717), .A2(n12716), .A3(n15484), .ZN(n12720) );
  OAI22_X1 U15022 ( .A1(n12718), .A2(n15469), .B1(n12749), .B2(n15467), .ZN(
        n12719) );
  NOR2_X1 U15023 ( .A1(n12720), .A2(n12719), .ZN(n12888) );
  MUX2_X1 U15024 ( .A(n12721), .B(n12888), .S(n15472), .Z(n12729) );
  XNOR2_X1 U15025 ( .A(n12723), .B(n12722), .ZN(n12890) );
  INV_X1 U15026 ( .A(n12724), .ZN(n12725) );
  OAI22_X1 U15027 ( .A1(n12893), .A2(n12726), .B1(n12725), .B2(n15460), .ZN(
        n12727) );
  AOI21_X1 U15028 ( .B1(n12890), .B2(n12741), .A(n12727), .ZN(n12728) );
  NAND2_X1 U15029 ( .A1(n12729), .A2(n12728), .ZN(P3_U3214) );
  OAI21_X1 U15030 ( .B1(n12731), .B2(n12739), .A(n12730), .ZN(n12733) );
  AOI222_X1 U15031 ( .A1(n12784), .A2(n12733), .B1(n12732), .B2(n15479), .C1(
        n12759), .C2(n12704), .ZN(n12825) );
  INV_X1 U15032 ( .A(n12734), .ZN(n12736) );
  OAI22_X1 U15033 ( .A1(n12736), .A2(n15460), .B1(n15472), .B2(n12735), .ZN(
        n12737) );
  AOI21_X1 U15034 ( .B1(n12738), .B2(n12787), .A(n12737), .ZN(n12743) );
  NAND2_X1 U15035 ( .A1(n12740), .A2(n12739), .ZN(n12822) );
  NAND3_X1 U15036 ( .A1(n12823), .A2(n12822), .A3(n12741), .ZN(n12742) );
  OAI211_X1 U15037 ( .C1(n12825), .C2(n15493), .A(n12743), .B(n12742), .ZN(
        P3_U3215) );
  XNOR2_X1 U15038 ( .A(n12744), .B(n12745), .ZN(n12899) );
  XNOR2_X1 U15039 ( .A(n12746), .B(n12745), .ZN(n12747) );
  OAI222_X1 U15040 ( .A1(n15469), .A2(n12749), .B1(n15467), .B2(n12748), .C1(
        n12747), .C2(n15484), .ZN(n12827) );
  NAND2_X1 U15041 ( .A1(n12827), .A2(n15472), .ZN(n12755) );
  NAND2_X1 U15042 ( .A1(n12750), .A2(n15488), .ZN(n12751) );
  OAI21_X1 U15043 ( .B1(n15472), .B2(n12752), .A(n12751), .ZN(n12753) );
  AOI21_X1 U15044 ( .B1(n12828), .B2(n12787), .A(n12753), .ZN(n12754) );
  OAI211_X1 U15045 ( .C1(n12899), .C2(n12790), .A(n12755), .B(n12754), .ZN(
        P3_U3216) );
  XOR2_X1 U15046 ( .A(n12757), .B(n12756), .Z(n12905) );
  XNOR2_X1 U15047 ( .A(n12758), .B(n12757), .ZN(n12760) );
  AOI222_X1 U15048 ( .A1(n12784), .A2(n12760), .B1(n12759), .B2(n15479), .C1(
        n12782), .C2(n12704), .ZN(n12900) );
  MUX2_X1 U15049 ( .A(n12761), .B(n12900), .S(n15472), .Z(n12764) );
  AOI22_X1 U15050 ( .A1(n12902), .A2(n12787), .B1(n15488), .B2(n12762), .ZN(
        n12763) );
  OAI211_X1 U15051 ( .C1(n12905), .C2(n12790), .A(n12764), .B(n12763), .ZN(
        P3_U3217) );
  OAI21_X1 U15052 ( .B1(n12766), .B2(n12767), .A(n12765), .ZN(n12910) );
  INV_X1 U15053 ( .A(n12910), .ZN(n12776) );
  XOR2_X1 U15054 ( .A(n12768), .B(n12767), .Z(n12771) );
  AOI222_X1 U15055 ( .A1(n12784), .A2(n12771), .B1(n12770), .B2(n15479), .C1(
        n12769), .C2(n12704), .ZN(n12906) );
  MUX2_X1 U15056 ( .A(n12772), .B(n12906), .S(n15472), .Z(n12775) );
  AOI22_X1 U15057 ( .A1(n12908), .A2(n12787), .B1(n15488), .B2(n12773), .ZN(
        n12774) );
  OAI211_X1 U15058 ( .C1(n12776), .C2(n12790), .A(n12775), .B(n12774), .ZN(
        P3_U3218) );
  XNOR2_X1 U15059 ( .A(n12777), .B(n12778), .ZN(n12920) );
  INV_X1 U15060 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12785) );
  XNOR2_X1 U15061 ( .A(n12780), .B(n12779), .ZN(n12783) );
  AOI222_X1 U15062 ( .A1(n12784), .A2(n12783), .B1(n12782), .B2(n15479), .C1(
        n12781), .C2(n12704), .ZN(n12913) );
  MUX2_X1 U15063 ( .A(n12785), .B(n12913), .S(n15472), .Z(n12789) );
  AOI22_X1 U15064 ( .A1(n12916), .A2(n12787), .B1(n15488), .B2(n12786), .ZN(
        n12788) );
  OAI211_X1 U15065 ( .C1(n12920), .C2(n12790), .A(n12789), .B(n12788), .ZN(
        P3_U3219) );
  NAND2_X1 U15066 ( .A1(n9433), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12792) );
  OAI211_X1 U15067 ( .C1(n8548), .C2(n12821), .A(n12792), .B(n12791), .ZN(
        P3_U3490) );
  NAND2_X1 U15068 ( .A1(n12793), .A2(n12829), .ZN(n12794) );
  OAI211_X1 U15069 ( .C1(n12797), .C2(n12796), .A(n12795), .B(n12794), .ZN(
        n12853) );
  MUX2_X1 U15070 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12853), .S(n15514), .Z(
        P3_U3486) );
  MUX2_X1 U15071 ( .A(n15617), .B(n12854), .S(n15514), .Z(n12799) );
  NAND2_X1 U15072 ( .A1(n12856), .A2(n12840), .ZN(n12798) );
  OAI211_X1 U15073 ( .C1(n12843), .C2(n12859), .A(n12799), .B(n12798), .ZN(
        P3_U3485) );
  AOI21_X1 U15074 ( .B1(n15501), .B2(n12801), .A(n12800), .ZN(n12860) );
  MUX2_X1 U15075 ( .A(n15575), .B(n12860), .S(n15514), .Z(n12802) );
  OAI21_X1 U15076 ( .B1(n12863), .B2(n12821), .A(n12802), .ZN(P3_U3484) );
  INV_X1 U15077 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12805) );
  AOI21_X1 U15078 ( .B1(n15501), .B2(n12804), .A(n12803), .ZN(n12864) );
  MUX2_X1 U15079 ( .A(n12805), .B(n12864), .S(n15514), .Z(n12806) );
  OAI21_X1 U15080 ( .B1(n12867), .B2(n12821), .A(n12806), .ZN(P3_U3483) );
  INV_X1 U15081 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12809) );
  AOI21_X1 U15082 ( .B1(n15501), .B2(n12808), .A(n12807), .ZN(n12868) );
  MUX2_X1 U15083 ( .A(n12809), .B(n12868), .S(n15514), .Z(n12810) );
  OAI21_X1 U15084 ( .B1(n12871), .B2(n12821), .A(n12810), .ZN(P3_U3482) );
  MUX2_X1 U15085 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n12872), .S(n15514), .Z(
        n12812) );
  OAI22_X1 U15086 ( .A1(n12874), .A2(n12843), .B1(n12873), .B2(n12821), .ZN(
        n12811) );
  OR2_X1 U15087 ( .A1(n12812), .A2(n12811), .ZN(P3_U3481) );
  INV_X1 U15088 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12813) );
  MUX2_X1 U15089 ( .A(n12813), .B(n12877), .S(n15514), .Z(n12815) );
  NAND2_X1 U15090 ( .A1(n12879), .A2(n12840), .ZN(n12814) );
  OAI211_X1 U15091 ( .C1(n12882), .C2(n12843), .A(n12815), .B(n12814), .ZN(
        P3_U3480) );
  MUX2_X1 U15092 ( .A(n15579), .B(n12883), .S(n15514), .Z(n12817) );
  NAND2_X1 U15093 ( .A1(n12884), .A2(n12840), .ZN(n12816) );
  OAI211_X1 U15094 ( .C1(n12887), .C2(n12843), .A(n12817), .B(n12816), .ZN(
        P3_U3479) );
  INV_X1 U15095 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12818) );
  MUX2_X1 U15096 ( .A(n12818), .B(n12888), .S(n15514), .Z(n12820) );
  NAND2_X1 U15097 ( .A1(n12890), .A2(n12836), .ZN(n12819) );
  OAI211_X1 U15098 ( .C1(n12821), .C2(n12893), .A(n12820), .B(n12819), .ZN(
        P3_U3478) );
  NAND3_X1 U15099 ( .A1(n12823), .A2(n12822), .A3(n15501), .ZN(n12824) );
  OAI211_X1 U15100 ( .C1(n12826), .C2(n15475), .A(n12825), .B(n12824), .ZN(
        n12895) );
  MUX2_X1 U15101 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12895), .S(n15514), .Z(
        P3_U3477) );
  INV_X1 U15102 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12830) );
  AOI21_X1 U15103 ( .B1(n12829), .B2(n12828), .A(n12827), .ZN(n12896) );
  MUX2_X1 U15104 ( .A(n12830), .B(n12896), .S(n15514), .Z(n12831) );
  OAI21_X1 U15105 ( .B1(n12843), .B2(n12899), .A(n12831), .ZN(P3_U3476) );
  MUX2_X1 U15106 ( .A(n12832), .B(n12900), .S(n15514), .Z(n12834) );
  NAND2_X1 U15107 ( .A1(n12902), .A2(n12840), .ZN(n12833) );
  OAI211_X1 U15108 ( .C1(n12905), .C2(n12843), .A(n12834), .B(n12833), .ZN(
        P3_U3475) );
  MUX2_X1 U15109 ( .A(n12835), .B(n12906), .S(n15514), .Z(n12838) );
  AOI22_X1 U15110 ( .A1(n12910), .A2(n12836), .B1(n12840), .B2(n12908), .ZN(
        n12837) );
  NAND2_X1 U15111 ( .A1(n12838), .A2(n12837), .ZN(P3_U3474) );
  INV_X1 U15112 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12839) );
  MUX2_X1 U15113 ( .A(n12839), .B(n12913), .S(n15514), .Z(n12842) );
  NAND2_X1 U15114 ( .A1(n12916), .A2(n12840), .ZN(n12841) );
  OAI211_X1 U15115 ( .C1(n12843), .C2(n12920), .A(n12842), .B(n12841), .ZN(
        P3_U3473) );
  NAND2_X1 U15116 ( .A1(n15509), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12845) );
  NAND2_X1 U15117 ( .A1(n12844), .A2(n15510), .ZN(n12847) );
  OAI211_X1 U15118 ( .C1(n8548), .C2(n12894), .A(n12845), .B(n12847), .ZN(
        P3_U3458) );
  NAND2_X1 U15119 ( .A1(n15509), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12846) );
  OAI211_X1 U15120 ( .C1(n12848), .C2(n12894), .A(n12847), .B(n12846), .ZN(
        P3_U3457) );
  NAND2_X1 U15121 ( .A1(n12850), .A2(n12915), .ZN(n12851) );
  NAND2_X1 U15122 ( .A1(n12852), .A2(n12851), .ZN(P3_U3456) );
  MUX2_X1 U15123 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12853), .S(n15510), .Z(
        P3_U3454) );
  INV_X1 U15124 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12855) );
  MUX2_X1 U15125 ( .A(n12855), .B(n12854), .S(n15510), .Z(n12858) );
  NAND2_X1 U15126 ( .A1(n12856), .A2(n12915), .ZN(n12857) );
  OAI211_X1 U15127 ( .C1(n12859), .C2(n12919), .A(n12858), .B(n12857), .ZN(
        P3_U3453) );
  INV_X1 U15128 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12861) );
  MUX2_X1 U15129 ( .A(n12861), .B(n12860), .S(n15510), .Z(n12862) );
  OAI21_X1 U15130 ( .B1(n12863), .B2(n12894), .A(n12862), .ZN(P3_U3452) );
  INV_X1 U15131 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12865) );
  MUX2_X1 U15132 ( .A(n12865), .B(n12864), .S(n15510), .Z(n12866) );
  OAI21_X1 U15133 ( .B1(n12867), .B2(n12894), .A(n12866), .ZN(P3_U3451) );
  INV_X1 U15134 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12869) );
  MUX2_X1 U15135 ( .A(n12869), .B(n12868), .S(n15510), .Z(n12870) );
  OAI21_X1 U15136 ( .B1(n12871), .B2(n12894), .A(n12870), .ZN(P3_U3450) );
  MUX2_X1 U15137 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n12872), .S(n15510), .Z(
        n12876) );
  OAI22_X1 U15138 ( .A1(n12874), .A2(n12919), .B1(n12873), .B2(n12894), .ZN(
        n12875) );
  OR2_X1 U15139 ( .A1(n12876), .A2(n12875), .ZN(P3_U3449) );
  INV_X1 U15140 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12878) );
  MUX2_X1 U15141 ( .A(n12878), .B(n12877), .S(n15510), .Z(n12881) );
  NAND2_X1 U15142 ( .A1(n12879), .A2(n12915), .ZN(n12880) );
  OAI211_X1 U15143 ( .C1(n12882), .C2(n12919), .A(n12881), .B(n12880), .ZN(
        P3_U3448) );
  MUX2_X1 U15144 ( .A(n15630), .B(n12883), .S(n15510), .Z(n12886) );
  NAND2_X1 U15145 ( .A1(n12884), .A2(n12915), .ZN(n12885) );
  OAI211_X1 U15146 ( .C1(n12887), .C2(n12919), .A(n12886), .B(n12885), .ZN(
        P3_U3447) );
  INV_X1 U15147 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12889) );
  MUX2_X1 U15148 ( .A(n12889), .B(n12888), .S(n15510), .Z(n12892) );
  NAND2_X1 U15149 ( .A1(n12890), .A2(n12909), .ZN(n12891) );
  OAI211_X1 U15150 ( .C1(n12894), .C2(n12893), .A(n12892), .B(n12891), .ZN(
        P3_U3446) );
  MUX2_X1 U15151 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12895), .S(n15510), .Z(
        P3_U3444) );
  INV_X1 U15152 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12897) );
  MUX2_X1 U15153 ( .A(n12897), .B(n12896), .S(n15510), .Z(n12898) );
  OAI21_X1 U15154 ( .B1(n12899), .B2(n12919), .A(n12898), .ZN(P3_U3441) );
  INV_X1 U15155 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12901) );
  MUX2_X1 U15156 ( .A(n12901), .B(n12900), .S(n15510), .Z(n12904) );
  NAND2_X1 U15157 ( .A1(n12902), .A2(n12915), .ZN(n12903) );
  OAI211_X1 U15158 ( .C1(n12905), .C2(n12919), .A(n12904), .B(n12903), .ZN(
        P3_U3438) );
  INV_X1 U15159 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12907) );
  MUX2_X1 U15160 ( .A(n12907), .B(n12906), .S(n15510), .Z(n12912) );
  AOI22_X1 U15161 ( .A1(n12910), .A2(n12909), .B1(n12915), .B2(n12908), .ZN(
        n12911) );
  NAND2_X1 U15162 ( .A1(n12912), .A2(n12911), .ZN(P3_U3435) );
  INV_X1 U15163 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12914) );
  MUX2_X1 U15164 ( .A(n12914), .B(n12913), .S(n15510), .Z(n12918) );
  NAND2_X1 U15165 ( .A1(n12916), .A2(n12915), .ZN(n12917) );
  OAI211_X1 U15166 ( .C1(n12920), .C2(n12919), .A(n12918), .B(n12917), .ZN(
        P3_U3432) );
  MUX2_X1 U15167 ( .A(P3_D_REG_1__SCAN_IN), .B(n12921), .S(n12922), .Z(
        P3_U3377) );
  MUX2_X1 U15168 ( .A(P3_D_REG_0__SCAN_IN), .B(n12923), .S(n12922), .Z(
        P3_U3376) );
  NAND3_X1 U15169 ( .A1(n12924), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12926) );
  OAI22_X1 U15170 ( .A1(n12927), .A2(n12926), .B1(n12925), .B2(n12941), .ZN(
        n12928) );
  AOI21_X1 U15171 ( .B1(n12930), .B2(n12929), .A(n12928), .ZN(n12931) );
  INV_X1 U15172 ( .A(n12931), .ZN(P3_U3264) );
  INV_X1 U15173 ( .A(n12932), .ZN(n12934) );
  OAI222_X1 U15174 ( .A1(n12941), .A2(n12935), .B1(n12948), .B2(n12934), .C1(
        n12933), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15175 ( .A(n12936), .ZN(n12938) );
  OAI222_X1 U15176 ( .A1(n12941), .A2(n12939), .B1(n12948), .B2(n12938), .C1(
        n12937), .C2(P3_U3151), .ZN(P3_U3268) );
  INV_X1 U15177 ( .A(n12940), .ZN(n12943) );
  OAI222_X1 U15178 ( .A1(P3_U3151), .A2(n12944), .B1(n12948), .B2(n12943), 
        .C1(n12942), .C2(n12941), .ZN(P3_U3269) );
  INV_X1 U15179 ( .A(n12945), .ZN(n12947) );
  OAI222_X1 U15180 ( .A1(P3_U3151), .A2(n12949), .B1(n12948), .B2(n12947), 
        .C1(n12946), .C2(n12941), .ZN(P3_U3270) );
  MUX2_X1 U15181 ( .A(n12951), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15182 ( .A(n12952), .B(n12953), .ZN(n12958) );
  NOR2_X1 U15183 ( .A1(n13289), .A2(n13081), .ZN(n12956) );
  AOI22_X1 U15184 ( .A1(n13337), .A2(n13083), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12954) );
  OAI21_X1 U15185 ( .B1(n13489), .B2(n13085), .A(n12954), .ZN(n12955) );
  AOI211_X1 U15186 ( .C1(n13491), .C2(n13087), .A(n12956), .B(n12955), .ZN(
        n12957) );
  OAI21_X1 U15187 ( .B1(n12958), .B2(n13089), .A(n12957), .ZN(P2_U3186) );
  NAND2_X1 U15188 ( .A1(n13006), .A2(n12959), .ZN(n12964) );
  NAND2_X1 U15189 ( .A1(n12961), .A2(n12960), .ZN(n12963) );
  INV_X1 U15190 ( .A(n13007), .ZN(n12962) );
  AOI21_X1 U15191 ( .B1(n12964), .B2(n12963), .A(n12962), .ZN(n12969) );
  NOR2_X1 U15192 ( .A1(n13085), .A2(n13709), .ZN(n12967) );
  AOI22_X1 U15193 ( .A1(n13723), .A2(n13343), .B1(n13344), .B2(n13722), .ZN(
        n13700) );
  OAI21_X1 U15194 ( .B1(n13074), .B2(n13700), .A(n12965), .ZN(n12966) );
  AOI211_X1 U15195 ( .C1(n13707), .C2(n13087), .A(n12967), .B(n12966), .ZN(
        n12968) );
  OAI21_X1 U15196 ( .B1(n12969), .B2(n13089), .A(n12968), .ZN(P2_U3187) );
  INV_X1 U15197 ( .A(n12970), .ZN(n13050) );
  OAI21_X1 U15198 ( .B1(n13051), .B2(n13050), .A(n12971), .ZN(n12975) );
  XNOR2_X1 U15199 ( .A(n12973), .B(n12972), .ZN(n12974) );
  XNOR2_X1 U15200 ( .A(n12975), .B(n12974), .ZN(n12981) );
  NAND2_X1 U15201 ( .A1(n13339), .A2(n13723), .ZN(n12977) );
  NAND2_X1 U15202 ( .A1(n13340), .A2(n13722), .ZN(n12976) );
  NAND2_X1 U15203 ( .A1(n12977), .A2(n12976), .ZN(n13553) );
  AOI22_X1 U15204 ( .A1(n13553), .A2(n13061), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12978) );
  OAI21_X1 U15205 ( .B1(n13545), .B2(n13085), .A(n12978), .ZN(n12979) );
  AOI21_X1 U15206 ( .B1(n13880), .B2(n13087), .A(n12979), .ZN(n12980) );
  OAI21_X1 U15207 ( .B1(n12981), .B2(n13089), .A(n12980), .ZN(P2_U3188) );
  INV_X1 U15208 ( .A(n12982), .ZN(n12983) );
  AOI21_X1 U15209 ( .B1(n12985), .B2(n12984), .A(n12983), .ZN(n12989) );
  OAI22_X1 U15210 ( .A1(n13581), .A2(n13678), .B1(n13294), .B2(n13676), .ZN(
        n13613) );
  NAND2_X1 U15211 ( .A1(n13613), .A2(n13061), .ZN(n12986) );
  NAND2_X1 U15212 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13435)
         );
  OAI211_X1 U15213 ( .C1(n13085), .C2(n13616), .A(n12986), .B(n13435), .ZN(
        n12987) );
  AOI21_X1 U15214 ( .B1(n13809), .B2(n13087), .A(n12987), .ZN(n12988) );
  OAI21_X1 U15215 ( .B1(n12989), .B2(n13089), .A(n12988), .ZN(P2_U3191) );
  XNOR2_X1 U15216 ( .A(n12991), .B(n12990), .ZN(n12997) );
  AOI22_X1 U15217 ( .A1(n13052), .A2(n13340), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12993) );
  NAND2_X1 U15218 ( .A1(n13072), .A2(n13588), .ZN(n12992) );
  OAI211_X1 U15219 ( .C1(n13581), .C2(n12994), .A(n12993), .B(n12992), .ZN(
        n12995) );
  AOI21_X1 U15220 ( .B1(n13587), .B2(n13087), .A(n12995), .ZN(n12996) );
  OAI21_X1 U15221 ( .B1(n12997), .B2(n13089), .A(n12996), .ZN(P2_U3195) );
  XNOR2_X1 U15222 ( .A(n12998), .B(n12999), .ZN(n13005) );
  NAND2_X1 U15223 ( .A1(n13337), .A2(n13723), .ZN(n13001) );
  NAND2_X1 U15224 ( .A1(n13339), .A2(n13722), .ZN(n13000) );
  NAND2_X1 U15225 ( .A1(n13001), .A2(n13000), .ZN(n13513) );
  AOI22_X1 U15226 ( .A1(n13513), .A2(n13061), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13002) );
  OAI21_X1 U15227 ( .B1(n13519), .B2(n13085), .A(n13002), .ZN(n13003) );
  AOI21_X1 U15228 ( .B1(n13521), .B2(n13087), .A(n13003), .ZN(n13004) );
  OAI21_X1 U15229 ( .B1(n13005), .B2(n13089), .A(n13004), .ZN(P2_U3197) );
  NAND2_X1 U15230 ( .A1(n13007), .A2(n13006), .ZN(n13008) );
  XOR2_X1 U15231 ( .A(n13009), .B(n13008), .Z(n13079) );
  INV_X1 U15232 ( .A(n13008), .ZN(n13011) );
  INV_X1 U15233 ( .A(n13009), .ZN(n13010) );
  AOI22_X1 U15234 ( .A1(n13079), .A2(n13078), .B1(n13011), .B2(n13010), .ZN(
        n13015) );
  NAND2_X1 U15235 ( .A1(n13013), .A2(n13012), .ZN(n13014) );
  XNOR2_X1 U15236 ( .A(n13015), .B(n13014), .ZN(n13021) );
  NOR2_X1 U15237 ( .A1(n13085), .A2(n13660), .ZN(n13019) );
  AND2_X1 U15238 ( .A1(n13343), .A2(n13722), .ZN(n13016) );
  AOI21_X1 U15239 ( .B1(n13342), .B2(n13723), .A(n13016), .ZN(n13663) );
  OAI21_X1 U15240 ( .B1(n13074), .B2(n13663), .A(n13017), .ZN(n13018) );
  AOI211_X1 U15241 ( .C1(n13180), .C2(n13087), .A(n13019), .B(n13018), .ZN(
        n13020) );
  OAI21_X1 U15242 ( .B1(n13021), .B2(n13089), .A(n13020), .ZN(P2_U3198) );
  INV_X1 U15243 ( .A(n13023), .ZN(n13024) );
  AOI21_X1 U15244 ( .B1(n13022), .B2(n13025), .A(n13024), .ZN(n13030) );
  NAND2_X1 U15245 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15397)
         );
  OAI21_X1 U15246 ( .B1(n13081), .B2(n13294), .A(n15397), .ZN(n13026) );
  AOI21_X1 U15247 ( .B1(n13083), .B2(n13641), .A(n13026), .ZN(n13027) );
  OAI21_X1 U15248 ( .B1(n13646), .B2(n13085), .A(n13027), .ZN(n13028) );
  AOI21_X1 U15249 ( .B1(n13819), .B2(n13087), .A(n13028), .ZN(n13029) );
  OAI21_X1 U15250 ( .B1(n13030), .B2(n13089), .A(n13029), .ZN(P2_U3200) );
  XNOR2_X1 U15251 ( .A(n13031), .B(n13032), .ZN(n13038) );
  AND2_X1 U15252 ( .A1(n13561), .A2(n13722), .ZN(n13033) );
  AOI21_X1 U15253 ( .B1(n13338), .B2(n13723), .A(n13033), .ZN(n13527) );
  OAI22_X1 U15254 ( .A1(n13527), .A2(n13074), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13034), .ZN(n13035) );
  AOI21_X1 U15255 ( .B1(n13534), .B2(n13072), .A(n13035), .ZN(n13037) );
  NAND2_X1 U15256 ( .A1(n13535), .A2(n13087), .ZN(n13036) );
  OAI211_X1 U15257 ( .C1(n13038), .C2(n13089), .A(n13037), .B(n13036), .ZN(
        P2_U3201) );
  OAI21_X1 U15258 ( .B1(n13041), .B2(n13040), .A(n13039), .ZN(n13043) );
  NAND2_X1 U15259 ( .A1(n13043), .A2(n13042), .ZN(n13048) );
  OAI22_X1 U15260 ( .A1(n13081), .A2(n13558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13044), .ZN(n13046) );
  NOR2_X1 U15261 ( .A1(n13085), .A2(n13603), .ZN(n13045) );
  AOI211_X1 U15262 ( .C1(n13083), .C2(n13598), .A(n13046), .B(n13045), .ZN(
        n13047) );
  OAI211_X1 U15263 ( .C1(n13606), .C2(n13049), .A(n13048), .B(n13047), .ZN(
        P2_U3205) );
  XNOR2_X1 U15264 ( .A(n13051), .B(n13050), .ZN(n13057) );
  AOI22_X1 U15265 ( .A1(n13561), .A2(n13052), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13054) );
  NAND2_X1 U15266 ( .A1(n13083), .A2(n13599), .ZN(n13053) );
  OAI211_X1 U15267 ( .C1(n13085), .C2(n13567), .A(n13054), .B(n13053), .ZN(
        n13055) );
  AOI21_X1 U15268 ( .B1(n13792), .B2(n13087), .A(n13055), .ZN(n13056) );
  OAI21_X1 U15269 ( .B1(n13057), .B2(n13089), .A(n13056), .ZN(P2_U3207) );
  XNOR2_X1 U15270 ( .A(n13059), .B(n13058), .ZN(n13066) );
  INV_X1 U15271 ( .A(n13631), .ZN(n13063) );
  NAND2_X1 U15272 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13402)
         );
  OAI22_X1 U15273 ( .A1(n13192), .A2(n13678), .B1(n13060), .B2(n13676), .ZN(
        n13628) );
  NAND2_X1 U15274 ( .A1(n13628), .A2(n13061), .ZN(n13062) );
  OAI211_X1 U15275 ( .C1(n13085), .C2(n13063), .A(n13402), .B(n13062), .ZN(
        n13064) );
  AOI21_X1 U15276 ( .B1(n13814), .B2(n13087), .A(n13064), .ZN(n13065) );
  OAI21_X1 U15277 ( .B1(n13066), .B2(n13089), .A(n13065), .ZN(P2_U3210) );
  INV_X1 U15278 ( .A(n13068), .ZN(n13069) );
  AOI21_X1 U15279 ( .B1(n13067), .B2(n13070), .A(n13069), .ZN(n13077) );
  AND2_X1 U15280 ( .A1(n13338), .A2(n13722), .ZN(n13071) );
  AOI21_X1 U15281 ( .B1(n13449), .B2(n13723), .A(n13071), .ZN(n13499) );
  AOI22_X1 U15282 ( .A1(n13502), .A2(n13072), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13073) );
  OAI21_X1 U15283 ( .B1(n13499), .B2(n13074), .A(n13073), .ZN(n13075) );
  AOI21_X1 U15284 ( .B1(n13771), .B2(n13087), .A(n13075), .ZN(n13076) );
  OAI21_X1 U15285 ( .B1(n13077), .B2(n13089), .A(n13076), .ZN(P2_U3212) );
  XNOR2_X1 U15286 ( .A(n13079), .B(n13078), .ZN(n13090) );
  OAI21_X1 U15287 ( .B1(n13081), .B2(n13679), .A(n13080), .ZN(n13082) );
  AOI21_X1 U15288 ( .B1(n13083), .B2(n13724), .A(n13082), .ZN(n13084) );
  OAI21_X1 U15289 ( .B1(n13684), .B2(n13085), .A(n13084), .ZN(n13086) );
  AOI21_X1 U15290 ( .B1(n13828), .B2(n13087), .A(n13086), .ZN(n13088) );
  OAI21_X1 U15291 ( .B1(n13090), .B2(n13089), .A(n13088), .ZN(P2_U3213) );
  OR2_X1 U15292 ( .A1(n14464), .A2(n13091), .ZN(n13093) );
  OR2_X1 U15293 ( .A1(n13264), .A2(n15631), .ZN(n13092) );
  INV_X1 U15294 ( .A(n13284), .ZN(n13094) );
  INV_X1 U15295 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13098) );
  NAND2_X1 U15296 ( .A1(n9503), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n13097) );
  INV_X1 U15297 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13095) );
  OR2_X1 U15298 ( .A1(n9479), .A2(n13095), .ZN(n13096) );
  OAI211_X1 U15299 ( .C1(n13100), .C2(n13098), .A(n13097), .B(n13096), .ZN(
        n13454) );
  NAND2_X1 U15300 ( .A1(n13099), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13103) );
  INV_X1 U15301 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13745) );
  OR2_X1 U15302 ( .A1(n9479), .A2(n13745), .ZN(n13102) );
  INV_X1 U15303 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13857) );
  OR2_X1 U15304 ( .A1(n13100), .A2(n13857), .ZN(n13101) );
  AND3_X1 U15305 ( .A1(n13103), .A2(n13102), .A3(n13101), .ZN(n13278) );
  AOI211_X1 U15306 ( .C1(n13105), .C2(n6398), .A(n13286), .B(n13104), .ZN(
        n13106) );
  OAI21_X1 U15307 ( .B1(n13278), .B2(n13277), .A(n13106), .ZN(n13107) );
  AOI22_X1 U15308 ( .A1(n13862), .A2(n13277), .B1(n13454), .B2(n13107), .ZN(
        n13276) );
  MUX2_X1 U15309 ( .A(n13454), .B(n13862), .S(n13189), .Z(n13275) );
  NAND2_X1 U15310 ( .A1(n7148), .A2(n15420), .ZN(n13112) );
  NAND2_X1 U15311 ( .A1(n13108), .A2(n13284), .ZN(n13110) );
  NAND2_X1 U15312 ( .A1(n13112), .A2(n13277), .ZN(n13109) );
  OAI211_X1 U15313 ( .C1(n13112), .C2(n13111), .A(n13110), .B(n13109), .ZN(
        n13114) );
  OAI21_X1 U15314 ( .B1(n13354), .B2(n13224), .A(n10805), .ZN(n13118) );
  NAND2_X1 U15315 ( .A1(n13354), .A2(n13224), .ZN(n13116) );
  NAND2_X1 U15316 ( .A1(n13116), .A2(n7152), .ZN(n13117) );
  MUX2_X1 U15317 ( .A(n13353), .B(n13119), .S(n13277), .Z(n13122) );
  NAND2_X1 U15318 ( .A1(n13123), .A2(n13122), .ZN(n13121) );
  MUX2_X1 U15319 ( .A(n13353), .B(n13119), .S(n13189), .Z(n13120) );
  NAND2_X1 U15320 ( .A1(n13121), .A2(n13120), .ZN(n13125) );
  MUX2_X1 U15321 ( .A(n13352), .B(n6405), .S(n13189), .Z(n13128) );
  MUX2_X1 U15322 ( .A(n13352), .B(n6405), .S(n13277), .Z(n13127) );
  MUX2_X1 U15323 ( .A(n13351), .B(n13129), .S(n13277), .Z(n13132) );
  MUX2_X1 U15324 ( .A(n13351), .B(n13129), .S(n13189), .Z(n13130) );
  MUX2_X1 U15325 ( .A(n13350), .B(n13133), .S(n13189), .Z(n13135) );
  MUX2_X1 U15326 ( .A(n13133), .B(n13350), .S(n13189), .Z(n13134) );
  MUX2_X1 U15327 ( .A(n13136), .B(n13349), .S(n13189), .Z(n13140) );
  NAND2_X1 U15328 ( .A1(n13139), .A2(n13140), .ZN(n13138) );
  MUX2_X1 U15329 ( .A(n13349), .B(n13136), .S(n13189), .Z(n13137) );
  NAND2_X1 U15330 ( .A1(n13138), .A2(n13137), .ZN(n13144) );
  INV_X1 U15331 ( .A(n13139), .ZN(n13142) );
  INV_X1 U15332 ( .A(n13140), .ZN(n13141) );
  NAND2_X1 U15333 ( .A1(n13142), .A2(n13141), .ZN(n13143) );
  MUX2_X1 U15334 ( .A(n13348), .B(n13145), .S(n13189), .Z(n13147) );
  MUX2_X1 U15335 ( .A(n13145), .B(n13348), .S(n13189), .Z(n13146) );
  MUX2_X1 U15336 ( .A(n13148), .B(n13347), .S(n13189), .Z(n13150) );
  MUX2_X1 U15337 ( .A(n13148), .B(n13347), .S(n13277), .Z(n13149) );
  MUX2_X1 U15338 ( .A(n13152), .B(n13346), .S(n13277), .Z(n13154) );
  MUX2_X1 U15339 ( .A(n13152), .B(n13346), .S(n13189), .Z(n13153) );
  INV_X1 U15340 ( .A(n13154), .ZN(n13155) );
  MUX2_X1 U15341 ( .A(n13345), .B(n7105), .S(n13277), .Z(n13159) );
  NAND2_X1 U15342 ( .A1(n13158), .A2(n13159), .ZN(n13157) );
  MUX2_X1 U15343 ( .A(n13345), .B(n7105), .S(n13189), .Z(n13156) );
  NAND2_X1 U15344 ( .A1(n13157), .A2(n13156), .ZN(n13163) );
  INV_X1 U15345 ( .A(n13158), .ZN(n13161) );
  INV_X1 U15346 ( .A(n13159), .ZN(n13160) );
  NAND2_X1 U15347 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  MUX2_X1 U15348 ( .A(n13721), .B(n13846), .S(n13189), .Z(n13165) );
  MUX2_X1 U15349 ( .A(n13721), .B(n13846), .S(n13277), .Z(n13164) );
  MUX2_X1 U15350 ( .A(n13344), .B(n13839), .S(n13277), .Z(n13168) );
  NAND2_X1 U15351 ( .A1(n13169), .A2(n13168), .ZN(n13167) );
  MUX2_X1 U15352 ( .A(n13344), .B(n13839), .S(n13189), .Z(n13166) );
  MUX2_X1 U15353 ( .A(n13724), .B(n13707), .S(n13189), .Z(n13172) );
  MUX2_X1 U15354 ( .A(n13707), .B(n13724), .S(n13189), .Z(n13171) );
  MUX2_X1 U15355 ( .A(n13343), .B(n13828), .S(n13277), .Z(n13176) );
  NAND2_X1 U15356 ( .A1(n13175), .A2(n13176), .ZN(n13174) );
  MUX2_X1 U15357 ( .A(n13343), .B(n13828), .S(n13189), .Z(n13173) );
  INV_X1 U15358 ( .A(n13175), .ZN(n13178) );
  INV_X1 U15359 ( .A(n13176), .ZN(n13177) );
  NAND2_X1 U15360 ( .A1(n13178), .A2(n13177), .ZN(n13179) );
  MUX2_X1 U15361 ( .A(n13641), .B(n13180), .S(n13189), .Z(n13182) );
  MUX2_X1 U15362 ( .A(n13641), .B(n13180), .S(n13277), .Z(n13181) );
  INV_X1 U15363 ( .A(n13182), .ZN(n13183) );
  MUX2_X1 U15364 ( .A(n13342), .B(n13819), .S(n13277), .Z(n13185) );
  MUX2_X1 U15365 ( .A(n13342), .B(n13819), .S(n13189), .Z(n13184) );
  INV_X1 U15366 ( .A(n13814), .ZN(n13633) );
  MUX2_X1 U15367 ( .A(n13294), .B(n13633), .S(n13189), .Z(n13191) );
  INV_X1 U15368 ( .A(n13191), .ZN(n13187) );
  MUX2_X1 U15369 ( .A(n13814), .B(n13642), .S(n13189), .Z(n13190) );
  MUX2_X1 U15370 ( .A(n13192), .B(n7696), .S(n13224), .Z(n13212) );
  MUX2_X1 U15371 ( .A(n13598), .B(n13809), .S(n13277), .Z(n13211) );
  INV_X1 U15372 ( .A(n13792), .ZN(n13566) );
  MUX2_X1 U15373 ( .A(n13580), .B(n13566), .S(n13224), .Z(n13202) );
  MUX2_X1 U15374 ( .A(n13340), .B(n13792), .S(n13277), .Z(n13201) );
  NAND2_X1 U15375 ( .A1(n13202), .A2(n13201), .ZN(n13208) );
  MUX2_X1 U15376 ( .A(n13558), .B(n13887), .S(n13224), .Z(n13199) );
  MUX2_X1 U15377 ( .A(n13599), .B(n13587), .S(n13277), .Z(n13198) );
  NAND2_X1 U15378 ( .A1(n13199), .A2(n13198), .ZN(n13193) );
  NAND2_X1 U15379 ( .A1(n13208), .A2(n13193), .ZN(n13205) );
  MUX2_X1 U15380 ( .A(n13581), .B(n13606), .S(n13224), .Z(n13204) );
  MUX2_X1 U15381 ( .A(n13341), .B(n13804), .S(n13277), .Z(n13203) );
  AND2_X1 U15382 ( .A1(n13204), .A2(n13203), .ZN(n13194) );
  OR2_X1 U15383 ( .A1(n13205), .A2(n13194), .ZN(n13210) );
  AOI21_X1 U15384 ( .B1(n13212), .B2(n13211), .A(n13210), .ZN(n13195) );
  INV_X1 U15385 ( .A(n13535), .ZN(n13877) );
  MUX2_X1 U15386 ( .A(n13196), .B(n13877), .S(n13277), .Z(n13227) );
  MUX2_X1 U15387 ( .A(n13339), .B(n13535), .S(n13224), .Z(n13226) );
  MUX2_X1 U15388 ( .A(n13197), .B(n6693), .S(n13224), .Z(n13230) );
  MUX2_X1 U15389 ( .A(n13338), .B(n13521), .S(n13277), .Z(n13229) );
  NOR2_X1 U15390 ( .A1(n13230), .A2(n13229), .ZN(n13228) );
  AOI21_X1 U15391 ( .B1(n13227), .B2(n13226), .A(n13228), .ZN(n13218) );
  NOR2_X1 U15392 ( .A1(n13199), .A2(n13198), .ZN(n13209) );
  INV_X1 U15393 ( .A(n13880), .ZN(n13200) );
  MUX2_X1 U15394 ( .A(n13293), .B(n13200), .S(n13224), .Z(n13220) );
  MUX2_X1 U15395 ( .A(n13561), .B(n13880), .S(n13277), .Z(n13219) );
  OAI22_X1 U15396 ( .A1(n13202), .A2(n13201), .B1(n13220), .B2(n13219), .ZN(
        n13207) );
  NOR3_X1 U15397 ( .A1(n13205), .A2(n13204), .A3(n13203), .ZN(n13206) );
  AOI211_X1 U15398 ( .C1(n13209), .C2(n13208), .A(n13207), .B(n13206), .ZN(
        n13217) );
  INV_X1 U15399 ( .A(n13210), .ZN(n13215) );
  INV_X1 U15400 ( .A(n13211), .ZN(n13214) );
  INV_X1 U15401 ( .A(n13212), .ZN(n13213) );
  NAND3_X1 U15402 ( .A1(n13215), .A2(n13214), .A3(n13213), .ZN(n13216) );
  INV_X1 U15403 ( .A(n13218), .ZN(n13223) );
  INV_X1 U15404 ( .A(n13219), .ZN(n13222) );
  INV_X1 U15405 ( .A(n13220), .ZN(n13221) );
  NOR3_X1 U15406 ( .A1(n13223), .A2(n13222), .A3(n13221), .ZN(n13237) );
  INV_X1 U15407 ( .A(n13765), .ZN(n13457) );
  MUX2_X1 U15408 ( .A(n13289), .B(n13457), .S(n13224), .Z(n13250) );
  MUX2_X1 U15409 ( .A(n13456), .B(n13765), .S(n13277), .Z(n13249) );
  NAND2_X1 U15410 ( .A1(n13250), .A2(n13249), .ZN(n13254) );
  MUX2_X1 U15411 ( .A(n13476), .B(n13869), .S(n13224), .Z(n13248) );
  MUX2_X1 U15412 ( .A(n13449), .B(n13491), .S(n13277), .Z(n13247) );
  NAND2_X1 U15413 ( .A1(n13248), .A2(n13247), .ZN(n13225) );
  NAND2_X1 U15414 ( .A1(n13254), .A2(n13225), .ZN(n13243) );
  NOR3_X1 U15415 ( .A1(n13228), .A2(n13227), .A3(n13226), .ZN(n13236) );
  INV_X1 U15416 ( .A(n13229), .ZN(n13234) );
  INV_X1 U15417 ( .A(n13230), .ZN(n13233) );
  MUX2_X1 U15418 ( .A(n13232), .B(n13231), .S(n13277), .Z(n13245) );
  MUX2_X1 U15419 ( .A(n13337), .B(n13771), .S(n13189), .Z(n13244) );
  OAI22_X1 U15420 ( .A1(n13234), .A2(n13233), .B1(n13245), .B2(n13244), .ZN(
        n13235) );
  NOR4_X1 U15421 ( .A1(n13237), .A2(n13243), .A3(n13236), .A4(n13235), .ZN(
        n13238) );
  NAND2_X1 U15422 ( .A1(n13239), .A2(n13262), .ZN(n13242) );
  OR2_X1 U15423 ( .A1(n13264), .A2(n13240), .ZN(n13241) );
  MUX2_X1 U15424 ( .A(n13477), .B(n13762), .S(n13189), .Z(n13269) );
  INV_X1 U15425 ( .A(n13477), .ZN(n13336) );
  MUX2_X1 U15426 ( .A(n13465), .B(n13336), .S(n13189), .Z(n13268) );
  INV_X1 U15427 ( .A(n13243), .ZN(n13246) );
  NAND3_X1 U15428 ( .A1(n13246), .A2(n13245), .A3(n13244), .ZN(n13256) );
  NOR2_X1 U15429 ( .A1(n13248), .A2(n13247), .ZN(n13253) );
  INV_X1 U15430 ( .A(n13249), .ZN(n13252) );
  INV_X1 U15431 ( .A(n13250), .ZN(n13251) );
  AOI22_X1 U15432 ( .A1(n13254), .A2(n13253), .B1(n13252), .B2(n13251), .ZN(
        n13255) );
  OAI211_X1 U15433 ( .C1(n13269), .C2(n13268), .A(n13256), .B(n13255), .ZN(
        n13267) );
  NAND2_X1 U15434 ( .A1(n13258), .A2(n13257), .ZN(n13261) );
  MUX2_X1 U15435 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7434), .Z(n13259) );
  XNOR2_X1 U15436 ( .A(n13259), .B(SI_31_), .ZN(n13260) );
  NAND2_X1 U15437 ( .A1(n15140), .A2(n13262), .ZN(n13266) );
  INV_X1 U15438 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13263) );
  OR2_X1 U15439 ( .A1(n13264), .A2(n13263), .ZN(n13265) );
  XNOR2_X1 U15440 ( .A(n13437), .B(n13278), .ZN(n13272) );
  INV_X1 U15441 ( .A(n13268), .ZN(n13271) );
  INV_X1 U15442 ( .A(n13269), .ZN(n13270) );
  OAI22_X1 U15443 ( .A1(n13276), .A2(n13275), .B1(n13271), .B2(n13270), .ZN(
        n13273) );
  INV_X1 U15444 ( .A(n13272), .ZN(n13322) );
  INV_X1 U15445 ( .A(n13278), .ZN(n13440) );
  NOR2_X1 U15446 ( .A1(n13440), .A2(n13277), .ZN(n13280) );
  NOR2_X1 U15447 ( .A1(n13278), .A2(n13189), .ZN(n13279) );
  MUX2_X1 U15448 ( .A(n13280), .B(n13279), .S(n13859), .Z(n13281) );
  MUX2_X1 U15449 ( .A(n13331), .B(n13323), .S(n13298), .Z(n13283) );
  NOR2_X1 U15450 ( .A1(n13331), .A2(n13284), .ZN(n13285) );
  AOI211_X1 U15451 ( .C1(n13323), .C2(n13666), .A(n13286), .B(n13285), .ZN(
        n13287) );
  NAND2_X1 U15452 ( .A1(n13765), .A2(n13289), .ZN(n13290) );
  NAND2_X1 U15453 ( .A1(n13292), .A2(n13291), .ZN(n13500) );
  XNOR2_X1 U15454 ( .A(n13880), .B(n13293), .ZN(n13550) );
  XNOR2_X1 U15455 ( .A(n13814), .B(n13294), .ZN(n13626) );
  NAND2_X1 U15456 ( .A1(n13295), .A2(n13557), .ZN(n13608) );
  NAND2_X1 U15457 ( .A1(n13297), .A2(n13296), .ZN(n13622) );
  AND2_X1 U15458 ( .A1(n15423), .A2(n13298), .ZN(n13301) );
  NAND4_X1 U15459 ( .A1(n13300), .A2(n13301), .A3(n13299), .A4(n7079), .ZN(
        n13303) );
  NOR2_X1 U15460 ( .A1(n13303), .A2(n13302), .ZN(n13307) );
  NAND4_X1 U15461 ( .A1(n13307), .A2(n13306), .A3(n13305), .A4(n13304), .ZN(
        n13308) );
  NOR2_X1 U15462 ( .A1(n13309), .A2(n13308), .ZN(n13312) );
  NAND4_X1 U15463 ( .A1(n13313), .A2(n13312), .A3(n13311), .A4(n13310), .ZN(
        n13314) );
  XNOR2_X1 U15464 ( .A(n13839), .B(n13695), .ZN(n13736) );
  NOR2_X1 U15465 ( .A1(n13314), .A2(n13736), .ZN(n13316) );
  NAND4_X1 U15466 ( .A1(n13667), .A2(n13316), .A3(n13315), .A4(n13703), .ZN(
        n13317) );
  NOR2_X1 U15467 ( .A1(n13674), .A2(n13317), .ZN(n13318) );
  NOR4_X1 U15468 ( .A1(n13475), .A2(n13450), .A3(n13515), .A4(n13319), .ZN(
        n13321) );
  XNOR2_X1 U15469 ( .A(n13862), .B(n13454), .ZN(n13320) );
  INV_X1 U15470 ( .A(n13327), .ZN(n13333) );
  OR3_X1 U15471 ( .A1(n13329), .A2(n13328), .A3(n13676), .ZN(n13330) );
  OAI211_X1 U15472 ( .C1(n13331), .C2(n13334), .A(n13330), .B(P2_B_REG_SCAN_IN), .ZN(n13332) );
  OAI211_X1 U15473 ( .C1(n13335), .C2(n13334), .A(n13333), .B(n13332), .ZN(
        P2_U3328) );
  MUX2_X1 U15474 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13440), .S(n6404), .Z(
        P2_U3562) );
  MUX2_X1 U15475 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13454), .S(n6404), .Z(
        P2_U3561) );
  MUX2_X1 U15476 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13336), .S(n6404), .Z(
        P2_U3560) );
  MUX2_X1 U15477 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13456), .S(n6404), .Z(
        P2_U3559) );
  MUX2_X1 U15478 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13449), .S(n6404), .Z(
        P2_U3558) );
  MUX2_X1 U15479 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13337), .S(n6404), .Z(
        P2_U3557) );
  MUX2_X1 U15480 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13338), .S(n6404), .Z(
        P2_U3556) );
  MUX2_X1 U15481 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13339), .S(n6404), .Z(
        P2_U3555) );
  MUX2_X1 U15482 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13561), .S(n6404), .Z(
        P2_U3554) );
  MUX2_X1 U15483 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13340), .S(n6404), .Z(
        P2_U3553) );
  MUX2_X1 U15484 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13599), .S(n6404), .Z(
        P2_U3552) );
  MUX2_X1 U15485 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13341), .S(n6404), .Z(
        P2_U3551) );
  MUX2_X1 U15486 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13598), .S(n6404), .Z(
        P2_U3550) );
  MUX2_X1 U15487 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13642), .S(n6404), .Z(
        P2_U3549) );
  MUX2_X1 U15488 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13342), .S(n6404), .Z(
        P2_U3548) );
  MUX2_X1 U15489 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13641), .S(n6404), .Z(
        P2_U3547) );
  MUX2_X1 U15490 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13343), .S(n6404), .Z(
        P2_U3546) );
  MUX2_X1 U15491 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13724), .S(n6404), .Z(
        P2_U3545) );
  MUX2_X1 U15492 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13344), .S(n6404), .Z(
        P2_U3544) );
  MUX2_X1 U15493 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13721), .S(n6404), .Z(
        P2_U3543) );
  MUX2_X1 U15494 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13345), .S(n6404), .Z(
        P2_U3542) );
  MUX2_X1 U15495 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13346), .S(n6404), .Z(
        P2_U3541) );
  MUX2_X1 U15496 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13347), .S(n6404), .Z(
        P2_U3540) );
  MUX2_X1 U15497 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13348), .S(n6404), .Z(
        P2_U3539) );
  MUX2_X1 U15498 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13349), .S(n6404), .Z(
        P2_U3538) );
  MUX2_X1 U15499 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13350), .S(n6404), .Z(
        P2_U3537) );
  MUX2_X1 U15500 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13351), .S(n6404), .Z(
        P2_U3536) );
  MUX2_X1 U15501 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13352), .S(n6404), .Z(
        P2_U3535) );
  MUX2_X1 U15502 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13353), .S(n6404), .Z(
        P2_U3534) );
  MUX2_X1 U15503 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13354), .S(n6404), .Z(
        P2_U3533) );
  MUX2_X1 U15504 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n10801), .S(n6404), .Z(
        P2_U3532) );
  MUX2_X1 U15505 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7148), .S(n6404), .Z(
        P2_U3531) );
  OAI22_X1 U15506 ( .A1(n15395), .A2(n13362), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13356), .ZN(n13357) );
  AOI21_X1 U15507 ( .B1(n15334), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n13357), .ZN(
        n13369) );
  MUX2_X1 U15508 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10100), .S(n13362), .Z(
        n13358) );
  INV_X1 U15509 ( .A(n13358), .ZN(n13360) );
  OAI211_X1 U15510 ( .C1(n13361), .C2(n13360), .A(n15405), .B(n13359), .ZN(
        n13368) );
  INV_X1 U15511 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13364) );
  MUX2_X1 U15512 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10072), .S(n13362), .Z(
        n13363) );
  OAI21_X1 U15513 ( .B1(n10142), .B2(n13364), .A(n13363), .ZN(n13365) );
  NAND3_X1 U15514 ( .A1(n15403), .A2(n13366), .A3(n13365), .ZN(n13367) );
  NAND3_X1 U15515 ( .A1(n13369), .A2(n13368), .A3(n13367), .ZN(P2_U3215) );
  OAI22_X1 U15516 ( .A1(n15395), .A2(n13372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13370), .ZN(n13371) );
  AOI21_X1 U15517 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n15334), .A(n13371), .ZN(
        n13380) );
  MUX2_X1 U15518 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n15528), .S(n13372), .Z(
        n13373) );
  INV_X1 U15519 ( .A(n13373), .ZN(n13375) );
  OAI211_X1 U15520 ( .C1(n13375), .C2(n13374), .A(n15405), .B(n13385), .ZN(
        n13379) );
  OAI211_X1 U15521 ( .C1(n13377), .C2(n13376), .A(n15403), .B(n13391), .ZN(
        n13378) );
  NAND3_X1 U15522 ( .A1(n13380), .A2(n13379), .A3(n13378), .ZN(P2_U3216) );
  OAI21_X1 U15523 ( .B1(n15395), .B2(n13382), .A(n13381), .ZN(n13383) );
  AOI21_X1 U15524 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15334), .A(n13383), .ZN(
        n13397) );
  MUX2_X1 U15525 ( .A(n11077), .B(P2_REG2_REG_3__SCAN_IN), .S(n13389), .Z(
        n13386) );
  NAND3_X1 U15526 ( .A1(n13386), .A2(n13385), .A3(n13384), .ZN(n13387) );
  NAND3_X1 U15527 ( .A1(n15405), .A2(n13388), .A3(n13387), .ZN(n13396) );
  MUX2_X1 U15528 ( .A(n10077), .B(P2_REG1_REG_3__SCAN_IN), .S(n13389), .Z(
        n13392) );
  NAND3_X1 U15529 ( .A1(n13392), .A2(n13391), .A3(n13390), .ZN(n13393) );
  NAND3_X1 U15530 ( .A1(n15403), .A2(n13394), .A3(n13393), .ZN(n13395) );
  NAND3_X1 U15531 ( .A1(n13397), .A2(n13396), .A3(n13395), .ZN(P2_U3217) );
  INV_X1 U15532 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13401) );
  XNOR2_X1 U15533 ( .A(n13410), .B(n13401), .ZN(n15402) );
  XNOR2_X1 U15534 ( .A(n13420), .B(n13422), .ZN(n13423) );
  XNOR2_X1 U15535 ( .A(n13423), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n13419) );
  OAI21_X1 U15536 ( .B1(n15395), .B2(n13403), .A(n13402), .ZN(n13404) );
  AOI21_X1 U15537 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15334), .A(n13404), 
        .ZN(n13418) );
  NAND2_X1 U15538 ( .A1(n13406), .A2(n13405), .ZN(n13409) );
  NAND2_X1 U15539 ( .A1(n13407), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13408) );
  OR2_X1 U15540 ( .A1(n13410), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U15541 ( .A1(n13410), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13412) );
  AND2_X1 U15542 ( .A1(n13411), .A2(n13412), .ZN(n15407) );
  NAND2_X1 U15543 ( .A1(n15408), .A2(n15407), .ZN(n15406) );
  NAND2_X1 U15544 ( .A1(n15406), .A2(n13412), .ZN(n13413) );
  NAND2_X1 U15545 ( .A1(n13413), .A2(n13422), .ZN(n13414) );
  OAI21_X1 U15546 ( .B1(n6477), .B2(n13415), .A(n13426), .ZN(n13416) );
  NAND2_X1 U15547 ( .A1(n13416), .A2(n15405), .ZN(n13417) );
  OAI211_X1 U15548 ( .C1(n13419), .C2(n13430), .A(n13418), .B(n13417), .ZN(
        P2_U3232) );
  INV_X1 U15549 ( .A(n13420), .ZN(n13421) );
  AOI22_X1 U15550 ( .A1(n13423), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n13422), 
        .B2(n13421), .ZN(n13424) );
  XNOR2_X1 U15551 ( .A(n13424), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13431) );
  NAND2_X1 U15552 ( .A1(n13426), .A2(n13425), .ZN(n13428) );
  INV_X1 U15553 ( .A(n13432), .ZN(n13429) );
  AOI22_X1 U15554 ( .A1(n13431), .A2(n15403), .B1(n15405), .B2(n13429), .ZN(
        n13434) );
  NOR2_X2 U15555 ( .A1(n13461), .A2(n13862), .ZN(n13445) );
  XNOR2_X1 U15556 ( .A(n13445), .B(n13437), .ZN(n13744) );
  NAND2_X1 U15557 ( .A1(n13744), .A2(n13741), .ZN(n13442) );
  NAND2_X1 U15558 ( .A1(n13438), .A2(P2_B_REG_SCAN_IN), .ZN(n13439) );
  AND2_X1 U15559 ( .A1(n13723), .A2(n13439), .ZN(n13455) );
  AND2_X1 U15560 ( .A1(n13440), .A2(n13455), .ZN(n13743) );
  INV_X1 U15561 ( .A(n13743), .ZN(n13747) );
  NOR2_X1 U15562 ( .A1(n6402), .A2(n13747), .ZN(n13446) );
  AOI21_X1 U15563 ( .B1(n6402), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13446), .ZN(
        n13441) );
  OAI211_X1 U15564 ( .C1(n13859), .C2(n13735), .A(n13442), .B(n13441), .ZN(
        P2_U3234) );
  NAND2_X1 U15565 ( .A1(n13461), .A2(n13862), .ZN(n13443) );
  NAND2_X1 U15566 ( .A1(n13443), .A2(n13840), .ZN(n13444) );
  AOI21_X1 U15567 ( .B1(n6402), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13446), .ZN(
        n13448) );
  NAND2_X1 U15568 ( .A1(n13862), .A2(n13649), .ZN(n13447) );
  OAI211_X1 U15569 ( .C1(n13748), .C2(n13549), .A(n13448), .B(n13447), .ZN(
        P2_U3235) );
  AND2_X1 U15570 ( .A1(n13765), .A2(n13456), .ZN(n13751) );
  INV_X1 U15571 ( .A(n13751), .ZN(n13754) );
  OAI21_X1 U15572 ( .B1(n13758), .B2(n13470), .A(n13754), .ZN(n13452) );
  XNOR2_X1 U15573 ( .A(n13452), .B(n13752), .ZN(n13469) );
  AND2_X1 U15574 ( .A1(n13491), .A2(n13476), .ZN(n13472) );
  AOI22_X1 U15575 ( .A1(n13456), .A2(n13722), .B1(n13455), .B2(n13454), .ZN(
        n13460) );
  NAND3_X1 U15576 ( .A1(n13473), .A2(n13752), .A3(n13717), .ZN(n13459) );
  NAND4_X1 U15577 ( .A1(n13752), .A2(n13457), .A3(n13717), .A4(n13456), .ZN(
        n13458) );
  OAI211_X1 U15578 ( .C1(n13481), .C2(n13762), .A(n13840), .B(n13461), .ZN(
        n13761) );
  OAI22_X1 U15579 ( .A1(n13463), .A2(n13683), .B1(n13462), .B2(n13687), .ZN(
        n13464) );
  AOI21_X1 U15580 ( .B1(n13465), .B2(n13649), .A(n13464), .ZN(n13466) );
  OAI21_X1 U15581 ( .B1(n13761), .B2(n13549), .A(n13466), .ZN(n13467) );
  AOI21_X1 U15582 ( .B1(n13760), .B2(n13687), .A(n13467), .ZN(n13468) );
  OAI21_X1 U15583 ( .B1(n13469), .B2(n13738), .A(n13468), .ZN(P2_U3236) );
  AOI211_X1 U15584 ( .C1(n13475), .C2(n13474), .A(n13701), .B(n13473), .ZN(
        n13479) );
  OAI22_X1 U15585 ( .A1(n13477), .A2(n13678), .B1(n13476), .B2(n13676), .ZN(
        n13478) );
  INV_X1 U15586 ( .A(n13480), .ZN(n13482) );
  AOI211_X1 U15587 ( .C1(n13765), .C2(n13482), .A(n13542), .B(n13481), .ZN(
        n13764) );
  NAND2_X1 U15588 ( .A1(n13764), .A2(n13666), .ZN(n13483) );
  OAI211_X1 U15589 ( .C1(n13683), .C2(n13484), .A(n13767), .B(n13483), .ZN(
        n13485) );
  AOI22_X1 U15590 ( .A1(n13765), .A2(n13649), .B1(n6402), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13486) );
  NAND2_X1 U15591 ( .A1(n13487), .A2(n13687), .ZN(n13497) );
  INV_X1 U15592 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13488) );
  OAI22_X1 U15593 ( .A1(n13489), .A2(n13683), .B1(n13488), .B2(n13687), .ZN(
        n13490) );
  AOI21_X1 U15594 ( .B1(n13491), .B2(n13649), .A(n13490), .ZN(n13496) );
  NAND2_X1 U15595 ( .A1(n13492), .A2(n13714), .ZN(n13495) );
  NAND2_X1 U15596 ( .A1(n13493), .A2(n13708), .ZN(n13494) );
  NAND4_X1 U15597 ( .A1(n13497), .A2(n13496), .A3(n13495), .A4(n13494), .ZN(
        P2_U3238) );
  XNOR2_X1 U15598 ( .A(n13501), .B(n13500), .ZN(n13772) );
  NAND2_X1 U15599 ( .A1(n13502), .A2(n13731), .ZN(n13503) );
  OAI21_X1 U15600 ( .B1(n13687), .B2(n13504), .A(n13503), .ZN(n13505) );
  AOI21_X1 U15601 ( .B1(n13771), .B2(n13649), .A(n13505), .ZN(n13509) );
  AOI21_X1 U15602 ( .B1(n13517), .B2(n13771), .A(n13542), .ZN(n13507) );
  AND2_X1 U15603 ( .A1(n13507), .A2(n13506), .ZN(n13770) );
  NAND2_X1 U15604 ( .A1(n13770), .A2(n13708), .ZN(n13508) );
  OAI211_X1 U15605 ( .C1(n13772), .C2(n13738), .A(n13509), .B(n13508), .ZN(
        n13510) );
  AOI21_X1 U15606 ( .B1(n13687), .B2(n13769), .A(n13510), .ZN(n13511) );
  INV_X1 U15607 ( .A(n13511), .ZN(P2_U3239) );
  XNOR2_X1 U15608 ( .A(n13512), .B(n13515), .ZN(n13514) );
  AOI21_X1 U15609 ( .B1(n13514), .B2(n13717), .A(n13513), .ZN(n13776) );
  XNOR2_X1 U15610 ( .A(n13516), .B(n13515), .ZN(n13773) );
  OAI211_X1 U15611 ( .C1(n13532), .C2(n6693), .A(n13840), .B(n13517), .ZN(
        n13774) );
  OAI22_X1 U15612 ( .A1(n13519), .A2(n13683), .B1(n13518), .B2(n13687), .ZN(
        n13520) );
  AOI21_X1 U15613 ( .B1(n13521), .B2(n13649), .A(n13520), .ZN(n13522) );
  OAI21_X1 U15614 ( .B1(n13774), .B2(n13549), .A(n13522), .ZN(n13523) );
  AOI21_X1 U15615 ( .B1(n13773), .B2(n13714), .A(n13523), .ZN(n13524) );
  OAI21_X1 U15616 ( .B1(n13776), .B2(n6402), .A(n13524), .ZN(P2_U3240) );
  XNOR2_X1 U15617 ( .A(n13525), .B(n13526), .ZN(n13529) );
  INV_X1 U15618 ( .A(n13527), .ZN(n13528) );
  AOI21_X1 U15619 ( .B1(n13529), .B2(n13717), .A(n13528), .ZN(n13780) );
  XNOR2_X1 U15620 ( .A(n13530), .B(n6866), .ZN(n13781) );
  INV_X1 U15621 ( .A(n13781), .ZN(n13539) );
  NAND2_X1 U15622 ( .A1(n13543), .A2(n13535), .ZN(n13531) );
  NAND2_X1 U15623 ( .A1(n13531), .A2(n13840), .ZN(n13533) );
  OR2_X1 U15624 ( .A1(n13533), .A2(n13532), .ZN(n13779) );
  AOI22_X1 U15625 ( .A1(n6402), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13534), 
        .B2(n13731), .ZN(n13537) );
  NAND2_X1 U15626 ( .A1(n13535), .A2(n13649), .ZN(n13536) );
  OAI211_X1 U15627 ( .C1(n13779), .C2(n13549), .A(n13537), .B(n13536), .ZN(
        n13538) );
  AOI21_X1 U15628 ( .B1(n13539), .B2(n13714), .A(n13538), .ZN(n13540) );
  OAI21_X1 U15629 ( .B1(n6402), .B2(n13780), .A(n13540), .ZN(P2_U3241) );
  XNOR2_X1 U15630 ( .A(n13541), .B(n6717), .ZN(n13784) );
  AOI21_X1 U15631 ( .B1(n13564), .B2(n13880), .A(n13542), .ZN(n13544) );
  NAND2_X1 U15632 ( .A1(n13544), .A2(n13543), .ZN(n13785) );
  OAI22_X1 U15633 ( .A1(n13687), .A2(n13546), .B1(n13545), .B2(n13683), .ZN(
        n13547) );
  AOI21_X1 U15634 ( .B1(n13880), .B2(n13649), .A(n13547), .ZN(n13548) );
  OAI21_X1 U15635 ( .B1(n13785), .B2(n13549), .A(n13548), .ZN(n13555) );
  XNOR2_X1 U15636 ( .A(n13551), .B(n13550), .ZN(n13552) );
  NAND2_X1 U15637 ( .A1(n13552), .A2(n13717), .ZN(n13786) );
  INV_X1 U15638 ( .A(n13553), .ZN(n13787) );
  AOI21_X1 U15639 ( .B1(n13786), .B2(n13787), .A(n6402), .ZN(n13554) );
  AOI211_X1 U15640 ( .C1(n13714), .C2(n13784), .A(n13555), .B(n13554), .ZN(
        n13556) );
  INV_X1 U15641 ( .A(n13556), .ZN(P2_U3242) );
  AOI21_X1 U15642 ( .B1(n13595), .B2(n13557), .A(n13582), .ZN(n13577) );
  AOI21_X1 U15643 ( .B1(n13558), .B2(n13587), .A(n13577), .ZN(n13560) );
  OAI211_X1 U15644 ( .C1(n13560), .C2(n13571), .A(n13717), .B(n13559), .ZN(
        n13563) );
  AOI22_X1 U15645 ( .A1(n13561), .A2(n13723), .B1(n13722), .B2(n13599), .ZN(
        n13562) );
  AND2_X1 U15646 ( .A1(n13563), .A2(n13562), .ZN(n13797) );
  INV_X1 U15647 ( .A(n13564), .ZN(n13565) );
  AOI211_X1 U15648 ( .C1(n13792), .C2(n13584), .A(n13542), .B(n13565), .ZN(
        n13791) );
  NOR2_X1 U15649 ( .A1(n13566), .A2(n13735), .ZN(n13570) );
  OAI22_X1 U15650 ( .A1(n13687), .A2(n13568), .B1(n13567), .B2(n13683), .ZN(
        n13569) );
  AOI211_X1 U15651 ( .C1(n13791), .C2(n13708), .A(n13570), .B(n13569), .ZN(
        n13574) );
  NAND2_X1 U15652 ( .A1(n13572), .A2(n13571), .ZN(n13793) );
  NAND3_X1 U15653 ( .A1(n13794), .A2(n13793), .A3(n13714), .ZN(n13573) );
  OAI211_X1 U15654 ( .C1(n13797), .C2(n6402), .A(n13574), .B(n13573), .ZN(
        P2_U3243) );
  NOR2_X1 U15655 ( .A1(n13576), .A2(n13575), .ZN(n13578) );
  AOI21_X1 U15656 ( .B1(n13578), .B2(n13595), .A(n13577), .ZN(n13579) );
  OAI222_X1 U15657 ( .A1(n13676), .A2(n13581), .B1(n13678), .B2(n13580), .C1(
        n13701), .C2(n13579), .ZN(n13798) );
  INV_X1 U15658 ( .A(n13798), .ZN(n13593) );
  XNOR2_X1 U15659 ( .A(n13583), .B(n13582), .ZN(n13800) );
  INV_X1 U15660 ( .A(n13601), .ZN(n13586) );
  INV_X1 U15661 ( .A(n13584), .ZN(n13585) );
  AOI211_X1 U15662 ( .C1(n13587), .C2(n13586), .A(n13542), .B(n13585), .ZN(
        n13799) );
  NAND2_X1 U15663 ( .A1(n13799), .A2(n13708), .ZN(n13590) );
  AOI22_X1 U15664 ( .A1(n6402), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13588), 
        .B2(n13731), .ZN(n13589) );
  OAI211_X1 U15665 ( .C1(n13887), .C2(n13735), .A(n13590), .B(n13589), .ZN(
        n13591) );
  AOI21_X1 U15666 ( .B1(n13800), .B2(n13714), .A(n13591), .ZN(n13592) );
  OAI21_X1 U15667 ( .B1(n13593), .B2(n6402), .A(n13592), .ZN(P2_U3244) );
  INV_X1 U15668 ( .A(n13594), .ZN(n13597) );
  INV_X1 U15669 ( .A(n13608), .ZN(n13596) );
  OAI21_X1 U15670 ( .B1(n13597), .B2(n13596), .A(n13595), .ZN(n13600) );
  AOI222_X1 U15671 ( .A1(n13717), .A2(n13600), .B1(n13599), .B2(n13723), .C1(
        n13598), .C2(n13722), .ZN(n13806) );
  INV_X1 U15672 ( .A(n13615), .ZN(n13602) );
  AOI211_X1 U15673 ( .C1(n13804), .C2(n13602), .A(n13542), .B(n13601), .ZN(
        n13803) );
  INV_X1 U15674 ( .A(n13603), .ZN(n13604) );
  AOI22_X1 U15675 ( .A1(n6402), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13604), 
        .B2(n13731), .ZN(n13605) );
  OAI21_X1 U15676 ( .B1(n13606), .B2(n13735), .A(n13605), .ZN(n13610) );
  XOR2_X1 U15677 ( .A(n13607), .B(n13608), .Z(n13807) );
  NOR2_X1 U15678 ( .A1(n13807), .A2(n13738), .ZN(n13609) );
  AOI211_X1 U15679 ( .C1(n13803), .C2(n13708), .A(n13610), .B(n13609), .ZN(
        n13611) );
  OAI21_X1 U15680 ( .B1(n13806), .B2(n6402), .A(n13611), .ZN(P2_U3245) );
  XNOR2_X1 U15681 ( .A(n13612), .B(n13622), .ZN(n13614) );
  AOI21_X1 U15682 ( .B1(n13614), .B2(n13717), .A(n13613), .ZN(n13811) );
  AOI211_X1 U15683 ( .C1(n13809), .C2(n13630), .A(n13542), .B(n13615), .ZN(
        n13808) );
  INV_X1 U15684 ( .A(n13616), .ZN(n13617) );
  AOI22_X1 U15685 ( .A1(n6402), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13617), 
        .B2(n13731), .ZN(n13618) );
  OAI21_X1 U15686 ( .B1(n7696), .B2(n13735), .A(n13618), .ZN(n13624) );
  NAND2_X1 U15687 ( .A1(n13644), .A2(n13619), .ZN(n13635) );
  INV_X1 U15688 ( .A(n13626), .ZN(n13636) );
  NOR2_X1 U15689 ( .A1(n13635), .A2(n13636), .ZN(n13634) );
  NOR2_X1 U15690 ( .A1(n13634), .A2(n13620), .ZN(n13621) );
  XOR2_X1 U15691 ( .A(n13622), .B(n13621), .Z(n13812) );
  NOR2_X1 U15692 ( .A1(n13812), .A2(n13738), .ZN(n13623) );
  AOI211_X1 U15693 ( .C1(n13808), .C2(n13708), .A(n13624), .B(n13623), .ZN(
        n13625) );
  OAI21_X1 U15694 ( .B1(n6402), .B2(n13811), .A(n13625), .ZN(P2_U3246) );
  XNOR2_X1 U15695 ( .A(n13627), .B(n13626), .ZN(n13629) );
  AOI21_X1 U15696 ( .B1(n13629), .B2(n13717), .A(n13628), .ZN(n13816) );
  AOI211_X1 U15697 ( .C1(n13814), .C2(n13652), .A(n13542), .B(n7697), .ZN(
        n13813) );
  AOI22_X1 U15698 ( .A1(n6402), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13631), 
        .B2(n13731), .ZN(n13632) );
  OAI21_X1 U15699 ( .B1(n13633), .B2(n13735), .A(n13632), .ZN(n13638) );
  AOI21_X1 U15700 ( .B1(n13636), .B2(n13635), .A(n13634), .ZN(n13817) );
  NOR2_X1 U15701 ( .A1(n13817), .A2(n13738), .ZN(n13637) );
  AOI211_X1 U15702 ( .C1(n13813), .C2(n13708), .A(n13638), .B(n13637), .ZN(
        n13639) );
  OAI21_X1 U15703 ( .B1(n6402), .B2(n13816), .A(n13639), .ZN(P2_U3247) );
  XNOR2_X1 U15704 ( .A(n13640), .B(n6457), .ZN(n13643) );
  AOI222_X1 U15705 ( .A1(n13717), .A2(n13643), .B1(n13642), .B2(n13723), .C1(
        n13641), .C2(n13722), .ZN(n13821) );
  OAI21_X1 U15706 ( .B1(n13645), .B2(n6457), .A(n13644), .ZN(n13822) );
  OAI22_X1 U15707 ( .A1(n13687), .A2(n13647), .B1(n13646), .B2(n13683), .ZN(
        n13648) );
  AOI21_X1 U15708 ( .B1(n13819), .B2(n13649), .A(n13648), .ZN(n13654) );
  OR2_X1 U15709 ( .A1(n13658), .A2(n13650), .ZN(n13651) );
  AND3_X1 U15710 ( .A1(n13652), .A2(n13651), .A3(n13840), .ZN(n13818) );
  NAND2_X1 U15711 ( .A1(n13818), .A2(n13708), .ZN(n13653) );
  OAI211_X1 U15712 ( .C1(n13822), .C2(n13738), .A(n13654), .B(n13653), .ZN(
        n13655) );
  INV_X1 U15713 ( .A(n13655), .ZN(n13656) );
  OAI21_X1 U15714 ( .B1(n13821), .B2(n6402), .A(n13656), .ZN(P2_U3248) );
  OAI21_X1 U15715 ( .B1(n13657), .B2(n13895), .A(n13840), .ZN(n13659) );
  NOR2_X1 U15716 ( .A1(n13659), .A2(n13658), .ZN(n13824) );
  NOR2_X1 U15717 ( .A1(n13683), .A2(n13660), .ZN(n13665) );
  OAI211_X1 U15718 ( .C1(n13662), .C2(n13667), .A(n13661), .B(n13717), .ZN(
        n13664) );
  NAND2_X1 U15719 ( .A1(n13664), .A2(n13663), .ZN(n13823) );
  AOI211_X1 U15720 ( .C1(n13824), .C2(n13666), .A(n13665), .B(n13823), .ZN(
        n13672) );
  XOR2_X1 U15721 ( .A(n13668), .B(n13667), .Z(n13825) );
  OAI22_X1 U15722 ( .A1(n13895), .A2(n13735), .B1(n13687), .B2(n13669), .ZN(
        n13670) );
  AOI21_X1 U15723 ( .B1(n13825), .B2(n13714), .A(n13670), .ZN(n13671) );
  OAI21_X1 U15724 ( .B1(n13672), .B2(n6402), .A(n13671), .ZN(P2_U3249) );
  XOR2_X1 U15725 ( .A(n13673), .B(n13674), .Z(n13831) );
  AOI21_X1 U15726 ( .B1(n13675), .B2(n13674), .A(n13701), .ZN(n13682) );
  OAI22_X1 U15727 ( .A1(n13679), .A2(n13678), .B1(n13677), .B2(n13676), .ZN(
        n13680) );
  AOI21_X1 U15728 ( .B1(n13682), .B2(n13681), .A(n13680), .ZN(n13830) );
  OAI21_X1 U15729 ( .B1(n13684), .B2(n13683), .A(n13830), .ZN(n13685) );
  NAND2_X1 U15730 ( .A1(n13685), .A2(n13687), .ZN(n13692) );
  XNOR2_X1 U15731 ( .A(n13705), .B(n13828), .ZN(n13686) );
  NOR2_X1 U15732 ( .A1(n13686), .A2(n12272), .ZN(n13827) );
  INV_X1 U15733 ( .A(n13828), .ZN(n13689) );
  INV_X1 U15734 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n13688) );
  OAI22_X1 U15735 ( .A1(n13689), .A2(n13735), .B1(n13688), .B2(n13687), .ZN(
        n13690) );
  AOI21_X1 U15736 ( .B1(n13827), .B2(n13708), .A(n13690), .ZN(n13691) );
  OAI211_X1 U15737 ( .C1(n13831), .C2(n13738), .A(n13692), .B(n13691), .ZN(
        P2_U3250) );
  NAND2_X1 U15738 ( .A1(n13694), .A2(n13693), .ZN(n13720) );
  INV_X1 U15739 ( .A(n13736), .ZN(n13719) );
  NAND2_X1 U15740 ( .A1(n13720), .A2(n13719), .ZN(n13718) );
  OAI21_X1 U15741 ( .B1(n13695), .B2(n13839), .A(n13718), .ZN(n13699) );
  INV_X1 U15742 ( .A(n13703), .ZN(n13698) );
  INV_X1 U15743 ( .A(n13696), .ZN(n13697) );
  AOI21_X1 U15744 ( .B1(n13699), .B2(n13698), .A(n13697), .ZN(n13702) );
  OAI21_X1 U15745 ( .B1(n13702), .B2(n13701), .A(n13700), .ZN(n13832) );
  INV_X1 U15746 ( .A(n13832), .ZN(n13716) );
  XNOR2_X1 U15747 ( .A(n13704), .B(n13703), .ZN(n13834) );
  INV_X1 U15748 ( .A(n13705), .ZN(n13706) );
  AOI211_X1 U15749 ( .C1(n13707), .C2(n13728), .A(n13542), .B(n13706), .ZN(
        n13833) );
  NAND2_X1 U15750 ( .A1(n13833), .A2(n13708), .ZN(n13712) );
  INV_X1 U15751 ( .A(n13709), .ZN(n13710) );
  AOI22_X1 U15752 ( .A1(n6402), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13710), 
        .B2(n13731), .ZN(n13711) );
  OAI211_X1 U15753 ( .C1(n6606), .C2(n13735), .A(n13712), .B(n13711), .ZN(
        n13713) );
  AOI21_X1 U15754 ( .B1(n13834), .B2(n13714), .A(n13713), .ZN(n13715) );
  OAI21_X1 U15755 ( .B1(n13716), .B2(n6402), .A(n13715), .ZN(P2_U3251) );
  OAI211_X1 U15756 ( .C1(n13720), .C2(n13719), .A(n13718), .B(n13717), .ZN(
        n13726) );
  AOI22_X1 U15757 ( .A1(n13724), .A2(n13723), .B1(n13722), .B2(n13721), .ZN(
        n13725) );
  AND2_X1 U15758 ( .A1(n13726), .A2(n13725), .ZN(n13843) );
  INV_X1 U15759 ( .A(n13727), .ZN(n13729) );
  AOI21_X1 U15760 ( .B1(n13839), .B2(n13729), .A(n6607), .ZN(n13841) );
  INV_X1 U15761 ( .A(n13730), .ZN(n13732) );
  AOI22_X1 U15762 ( .A1(n6402), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13732), 
        .B2(n13731), .ZN(n13733) );
  OAI21_X1 U15763 ( .B1(n13735), .B2(n13734), .A(n13733), .ZN(n13740) );
  XNOR2_X1 U15764 ( .A(n13737), .B(n13736), .ZN(n13844) );
  NOR2_X1 U15765 ( .A1(n13844), .A2(n13738), .ZN(n13739) );
  AOI211_X1 U15766 ( .C1(n13841), .C2(n13741), .A(n13740), .B(n13739), .ZN(
        n13742) );
  OAI21_X1 U15767 ( .B1(n6402), .B2(n13843), .A(n13742), .ZN(P2_U3252) );
  AOI21_X1 U15768 ( .B1(n13744), .B2(n13840), .A(n13743), .ZN(n13856) );
  MUX2_X1 U15769 ( .A(n13745), .B(n13856), .S(n15454), .Z(n13746) );
  OAI21_X1 U15770 ( .B1(n13859), .B2(n13838), .A(n13746), .ZN(P2_U3530) );
  NAND2_X1 U15771 ( .A1(n13748), .A2(n13747), .ZN(n13860) );
  AOI21_X1 U15772 ( .B1(n13789), .B2(n13862), .A(n13749), .ZN(n13750) );
  INV_X1 U15773 ( .A(n13750), .ZN(P2_U3529) );
  NOR2_X1 U15774 ( .A1(n13752), .A2(n13751), .ZN(n13757) );
  NAND3_X1 U15775 ( .A1(n13755), .A2(n13470), .A3(n13754), .ZN(n13753) );
  OAI211_X1 U15776 ( .C1(n13755), .C2(n13754), .A(n13753), .B(n13835), .ZN(
        n13756) );
  OAI21_X1 U15777 ( .B1(n13762), .B2(n15439), .A(n13761), .ZN(n13763) );
  AOI21_X1 U15778 ( .B1(n13851), .B2(n13765), .A(n13764), .ZN(n13766) );
  MUX2_X1 U15779 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13870), .S(n15454), .Z(
        P2_U3525) );
  INV_X1 U15780 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13777) );
  NAND2_X1 U15781 ( .A1(n13773), .A2(n13835), .ZN(n13775) );
  AND3_X1 U15782 ( .A1(n13776), .A2(n13775), .A3(n13774), .ZN(n13871) );
  MUX2_X1 U15783 ( .A(n13777), .B(n13871), .S(n15454), .Z(n13778) );
  OAI21_X1 U15784 ( .B1(n6693), .B2(n13838), .A(n13778), .ZN(P2_U3524) );
  OAI211_X1 U15785 ( .C1(n13855), .C2(n13781), .A(n13780), .B(n13779), .ZN(
        n13874) );
  MUX2_X1 U15786 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13874), .S(n15454), .Z(
        n13782) );
  INV_X1 U15787 ( .A(n13782), .ZN(n13783) );
  OAI21_X1 U15788 ( .B1(n13877), .B2(n13838), .A(n13783), .ZN(P2_U3523) );
  MUX2_X1 U15789 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13878), .S(n15454), .Z(
        n13788) );
  AOI21_X1 U15790 ( .B1(n13789), .B2(n13880), .A(n13788), .ZN(n13790) );
  INV_X1 U15791 ( .A(n13790), .ZN(P2_U3522) );
  AOI21_X1 U15792 ( .B1(n13851), .B2(n13792), .A(n13791), .ZN(n13796) );
  NAND3_X1 U15793 ( .A1(n13794), .A2(n13793), .A3(n13835), .ZN(n13795) );
  NAND3_X1 U15794 ( .A1(n13797), .A2(n13796), .A3(n13795), .ZN(n13883) );
  MUX2_X1 U15795 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13883), .S(n15454), .Z(
        P2_U3521) );
  INV_X1 U15796 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13801) );
  AOI211_X1 U15797 ( .C1(n13800), .C2(n13835), .A(n13799), .B(n13798), .ZN(
        n13884) );
  MUX2_X1 U15798 ( .A(n13801), .B(n13884), .S(n15454), .Z(n13802) );
  OAI21_X1 U15799 ( .B1(n13887), .B2(n13838), .A(n13802), .ZN(P2_U3520) );
  AOI21_X1 U15800 ( .B1(n13851), .B2(n13804), .A(n13803), .ZN(n13805) );
  OAI211_X1 U15801 ( .C1(n13855), .C2(n13807), .A(n13806), .B(n13805), .ZN(
        n13888) );
  MUX2_X1 U15802 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13888), .S(n15454), .Z(
        P2_U3519) );
  AOI21_X1 U15803 ( .B1(n13851), .B2(n13809), .A(n13808), .ZN(n13810) );
  OAI211_X1 U15804 ( .C1(n13812), .C2(n13855), .A(n13811), .B(n13810), .ZN(
        n13889) );
  MUX2_X1 U15805 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13889), .S(n15454), .Z(
        P2_U3518) );
  AOI21_X1 U15806 ( .B1(n13851), .B2(n13814), .A(n13813), .ZN(n13815) );
  OAI211_X1 U15807 ( .C1(n13817), .C2(n13855), .A(n13816), .B(n13815), .ZN(
        n13890) );
  MUX2_X1 U15808 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13890), .S(n15454), .Z(
        P2_U3517) );
  AOI21_X1 U15809 ( .B1(n13851), .B2(n13819), .A(n13818), .ZN(n13820) );
  OAI211_X1 U15810 ( .C1(n13855), .C2(n13822), .A(n13821), .B(n13820), .ZN(
        n13891) );
  MUX2_X1 U15811 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13891), .S(n15454), .Z(
        P2_U3516) );
  AOI211_X1 U15812 ( .C1(n13825), .C2(n13835), .A(n13824), .B(n13823), .ZN(
        n13892) );
  MUX2_X1 U15813 ( .A(n15531), .B(n13892), .S(n15454), .Z(n13826) );
  OAI21_X1 U15814 ( .B1(n13895), .B2(n13838), .A(n13826), .ZN(P2_U3515) );
  AOI21_X1 U15815 ( .B1(n13851), .B2(n13828), .A(n13827), .ZN(n13829) );
  OAI211_X1 U15816 ( .C1(n13831), .C2(n13855), .A(n13830), .B(n13829), .ZN(
        n13896) );
  MUX2_X1 U15817 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13896), .S(n15454), .Z(
        P2_U3514) );
  AOI211_X1 U15818 ( .C1(n13835), .C2(n13834), .A(n13833), .B(n13832), .ZN(
        n13897) );
  MUX2_X1 U15819 ( .A(n13836), .B(n13897), .S(n15454), .Z(n13837) );
  OAI21_X1 U15820 ( .B1(n6606), .B2(n13838), .A(n13837), .ZN(P2_U3513) );
  AOI22_X1 U15821 ( .A1(n13841), .A2(n13840), .B1(n13851), .B2(n13839), .ZN(
        n13842) );
  OAI211_X1 U15822 ( .C1(n13855), .C2(n13844), .A(n13843), .B(n13842), .ZN(
        n13901) );
  MUX2_X1 U15823 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13901), .S(n15454), .Z(
        P2_U3512) );
  AOI21_X1 U15824 ( .B1(n13851), .B2(n13846), .A(n13845), .ZN(n13847) );
  OAI211_X1 U15825 ( .C1(n13855), .C2(n13849), .A(n13848), .B(n13847), .ZN(
        n13902) );
  MUX2_X1 U15826 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13902), .S(n15454), .Z(
        P2_U3511) );
  AOI21_X1 U15827 ( .B1(n13851), .B2(n7105), .A(n13850), .ZN(n13852) );
  OAI211_X1 U15828 ( .C1(n13855), .C2(n13854), .A(n13853), .B(n13852), .ZN(
        n13903) );
  MUX2_X1 U15829 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n13903), .S(n15454), .Z(
        P2_U3510) );
  MUX2_X1 U15830 ( .A(n13857), .B(n13856), .S(n15448), .Z(n13858) );
  OAI21_X1 U15831 ( .B1(n13859), .B2(n13900), .A(n13858), .ZN(P2_U3498) );
  INV_X1 U15832 ( .A(n13863), .ZN(P2_U3497) );
  MUX2_X1 U15833 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13865), .S(n15448), .Z(
        P2_U3495) );
  INV_X1 U15834 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13867) );
  OAI21_X1 U15835 ( .B1(n13869), .B2(n13900), .A(n13868), .ZN(P2_U3494) );
  MUX2_X1 U15836 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13870), .S(n15448), .Z(
        P2_U3493) );
  INV_X1 U15837 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13872) );
  MUX2_X1 U15838 ( .A(n13872), .B(n13871), .S(n15448), .Z(n13873) );
  OAI21_X1 U15839 ( .B1(n6693), .B2(n13900), .A(n13873), .ZN(P2_U3492) );
  MUX2_X1 U15840 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13874), .S(n15448), .Z(
        n13875) );
  INV_X1 U15841 ( .A(n13875), .ZN(n13876) );
  OAI21_X1 U15842 ( .B1(n13877), .B2(n13900), .A(n13876), .ZN(P2_U3491) );
  MUX2_X1 U15843 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13878), .S(n15448), .Z(
        n13879) );
  AOI21_X1 U15844 ( .B1(n13881), .B2(n13880), .A(n13879), .ZN(n13882) );
  INV_X1 U15845 ( .A(n13882), .ZN(P2_U3490) );
  MUX2_X1 U15846 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13883), .S(n15448), .Z(
        P2_U3489) );
  INV_X1 U15847 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13885) );
  MUX2_X1 U15848 ( .A(n13885), .B(n13884), .S(n15448), .Z(n13886) );
  OAI21_X1 U15849 ( .B1(n13887), .B2(n13900), .A(n13886), .ZN(P2_U3488) );
  MUX2_X1 U15850 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13888), .S(n15448), .Z(
        P2_U3487) );
  MUX2_X1 U15851 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13889), .S(n15448), .Z(
        P2_U3486) );
  MUX2_X1 U15852 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13890), .S(n15448), .Z(
        P2_U3484) );
  MUX2_X1 U15853 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13891), .S(n15448), .Z(
        P2_U3481) );
  INV_X1 U15854 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n13893) );
  MUX2_X1 U15855 ( .A(n13893), .B(n13892), .S(n15448), .Z(n13894) );
  OAI21_X1 U15856 ( .B1(n13895), .B2(n13900), .A(n13894), .ZN(P2_U3478) );
  MUX2_X1 U15857 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13896), .S(n15448), .Z(
        P2_U3475) );
  MUX2_X1 U15858 ( .A(n13898), .B(n13897), .S(n15448), .Z(n13899) );
  OAI21_X1 U15859 ( .B1(n6606), .B2(n13900), .A(n13899), .ZN(P2_U3472) );
  MUX2_X1 U15860 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13901), .S(n15448), .Z(
        P2_U3469) );
  MUX2_X1 U15861 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n13902), .S(n15448), .Z(
        P2_U3466) );
  MUX2_X1 U15862 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n13903), .S(n15448), .Z(
        P2_U3463) );
  INV_X1 U15863 ( .A(n15140), .ZN(n13909) );
  NOR4_X1 U15864 ( .A1(n13906), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13905), .A4(
        P2_U3088), .ZN(n13907) );
  AOI21_X1 U15865 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13910), .A(n13907), 
        .ZN(n13908) );
  OAI21_X1 U15866 ( .B1(n13909), .B2(n13913), .A(n13908), .ZN(P2_U3296) );
  NAND2_X1 U15867 ( .A1(n13910), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13912) );
  OAI211_X1 U15868 ( .C1(n13914), .C2(n13913), .A(n13912), .B(n13911), .ZN(
        P2_U3299) );
  INV_X1 U15869 ( .A(n13915), .ZN(n15146) );
  OAI222_X1 U15870 ( .A1(n13918), .A2(P2_U3088), .B1(n13913), .B2(n15146), 
        .C1(n13917), .C2(n13916), .ZN(P2_U3302) );
  MUX2_X1 U15871 ( .A(n13919), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15872 ( .A1(n14985), .A2(n10284), .ZN(n13921) );
  NAND2_X1 U15873 ( .A1(n14567), .A2(n10286), .ZN(n13920) );
  NAND2_X1 U15874 ( .A1(n13921), .A2(n13920), .ZN(n13922) );
  XNOR2_X1 U15875 ( .A(n13922), .B(n14051), .ZN(n13925) );
  INV_X1 U15876 ( .A(n13925), .ZN(n13927) );
  AND2_X1 U15877 ( .A1(n14567), .A2(n14108), .ZN(n13923) );
  AOI21_X1 U15878 ( .B1(n14985), .B2(n10286), .A(n13923), .ZN(n13924) );
  INV_X1 U15879 ( .A(n13924), .ZN(n13926) );
  AOI21_X1 U15880 ( .B1(n13927), .B2(n13926), .A(n14122), .ZN(n14058) );
  NAND2_X1 U15881 ( .A1(n15078), .A2(n10284), .ZN(n13929) );
  OR2_X1 U15882 ( .A1(n15082), .A2(n14020), .ZN(n13928) );
  NAND2_X1 U15883 ( .A1(n13929), .A2(n13928), .ZN(n13930) );
  XNOR2_X1 U15884 ( .A(n13930), .B(n14051), .ZN(n13959) );
  NOR2_X1 U15885 ( .A1(n15082), .A2(n14052), .ZN(n13931) );
  AOI21_X1 U15886 ( .B1(n15078), .B2(n10286), .A(n13931), .ZN(n13958) );
  INV_X1 U15887 ( .A(n13932), .ZN(n13933) );
  NAND2_X1 U15888 ( .A1(n7165), .A2(n10286), .ZN(n13936) );
  NAND2_X1 U15889 ( .A1(n15092), .A2(n14108), .ZN(n13935) );
  NAND2_X1 U15890 ( .A1(n13936), .A2(n13935), .ZN(n14068) );
  NAND2_X1 U15891 ( .A1(n7165), .A2(n10284), .ZN(n13938) );
  NAND2_X1 U15892 ( .A1(n15092), .A2(n10286), .ZN(n13937) );
  NAND2_X1 U15893 ( .A1(n13938), .A2(n13937), .ZN(n13939) );
  XNOR2_X1 U15894 ( .A(n13939), .B(n14111), .ZN(n14069) );
  NAND2_X1 U15895 ( .A1(n15086), .A2(n10284), .ZN(n13941) );
  NAND2_X1 U15896 ( .A1(n15091), .A2(n10286), .ZN(n13940) );
  NAND2_X1 U15897 ( .A1(n13941), .A2(n13940), .ZN(n13942) );
  XNOR2_X1 U15898 ( .A(n13942), .B(n14111), .ZN(n13950) );
  NAND2_X1 U15899 ( .A1(n15086), .A2(n10286), .ZN(n13944) );
  NAND2_X1 U15900 ( .A1(n15091), .A2(n14108), .ZN(n13943) );
  NAND2_X1 U15901 ( .A1(n13944), .A2(n13943), .ZN(n13951) );
  AND2_X1 U15902 ( .A1(n13950), .A2(n13951), .ZN(n13949) );
  NAND2_X1 U15903 ( .A1(n14972), .A2(n10284), .ZN(n13946) );
  NAND2_X1 U15904 ( .A1(n14946), .A2(n10286), .ZN(n13945) );
  NAND2_X1 U15905 ( .A1(n13946), .A2(n13945), .ZN(n13947) );
  XNOR2_X1 U15906 ( .A(n13947), .B(n14051), .ZN(n14067) );
  AND2_X1 U15907 ( .A1(n14946), .A2(n14108), .ZN(n13948) );
  AOI21_X1 U15908 ( .B1(n14972), .B2(n10286), .A(n13948), .ZN(n14065) );
  NOR2_X1 U15909 ( .A1(n14067), .A2(n14065), .ZN(n14071) );
  AOI211_X1 U15910 ( .C1(n14068), .C2(n14069), .A(n13949), .B(n14071), .ZN(
        n13957) );
  NOR4_X1 U15911 ( .A1(n14071), .A2(n14069), .A3(n13949), .A4(n14068), .ZN(
        n13956) );
  INV_X1 U15912 ( .A(n13949), .ZN(n14070) );
  NAND3_X1 U15913 ( .A1(n14070), .A2(n14065), .A3(n14067), .ZN(n13954) );
  INV_X1 U15914 ( .A(n13950), .ZN(n13953) );
  INV_X1 U15915 ( .A(n13951), .ZN(n13952) );
  NAND2_X1 U15916 ( .A1(n13953), .A2(n13952), .ZN(n14073) );
  NAND2_X1 U15917 ( .A1(n13954), .A2(n14073), .ZN(n13955) );
  XNOR2_X1 U15918 ( .A(n13959), .B(n13958), .ZN(n14072) );
  NAND2_X1 U15919 ( .A1(n15071), .A2(n10284), .ZN(n13961) );
  OR2_X1 U15920 ( .A1(n15074), .A2(n14020), .ZN(n13960) );
  NAND2_X1 U15921 ( .A1(n13961), .A2(n13960), .ZN(n13962) );
  XNOR2_X1 U15922 ( .A(n13962), .B(n14051), .ZN(n14168) );
  NOR2_X1 U15923 ( .A1(n15074), .A2(n14052), .ZN(n13963) );
  AOI21_X1 U15924 ( .B1(n15071), .B2(n10286), .A(n13963), .ZN(n14292) );
  NAND2_X1 U15925 ( .A1(n15064), .A2(n10284), .ZN(n13965) );
  NAND2_X1 U15926 ( .A1(n14884), .A2(n10286), .ZN(n13964) );
  NAND2_X1 U15927 ( .A1(n13965), .A2(n13964), .ZN(n13966) );
  XNOR2_X1 U15928 ( .A(n13966), .B(n14051), .ZN(n13969) );
  NOR2_X1 U15929 ( .A1(n15053), .A2(n14052), .ZN(n13967) );
  AOI21_X1 U15930 ( .B1(n15064), .B2(n10286), .A(n13967), .ZN(n13968) );
  OR2_X1 U15931 ( .A1(n13969), .A2(n13968), .ZN(n14166) );
  OAI21_X1 U15932 ( .B1(n14168), .B2(n14292), .A(n14166), .ZN(n13971) );
  NAND2_X1 U15933 ( .A1(n13969), .A2(n13968), .ZN(n14191) );
  NAND3_X1 U15934 ( .A1(n14168), .A2(n14166), .A3(n14292), .ZN(n13970) );
  NAND2_X1 U15935 ( .A1(n15057), .A2(n10284), .ZN(n13973) );
  OR2_X1 U15936 ( .A1(n15061), .A2(n14020), .ZN(n13972) );
  NAND2_X1 U15937 ( .A1(n13973), .A2(n13972), .ZN(n13974) );
  XNOR2_X1 U15938 ( .A(n13974), .B(n14051), .ZN(n13977) );
  INV_X1 U15939 ( .A(n13977), .ZN(n13979) );
  NOR2_X1 U15940 ( .A1(n15061), .A2(n14052), .ZN(n13975) );
  AOI21_X1 U15941 ( .B1(n15057), .B2(n10286), .A(n13975), .ZN(n13976) );
  INV_X1 U15942 ( .A(n13976), .ZN(n13978) );
  AND2_X1 U15943 ( .A1(n13977), .A2(n13976), .ZN(n13980) );
  AOI21_X1 U15944 ( .B1(n13979), .B2(n13978), .A(n13980), .ZN(n14192) );
  INV_X1 U15945 ( .A(n13980), .ZN(n13981) );
  OAI22_X1 U15946 ( .A1(n14855), .A2(n14020), .B1(n15054), .B2(n14052), .ZN(
        n13985) );
  NAND2_X1 U15947 ( .A1(n15045), .A2(n10284), .ZN(n13983) );
  OR2_X1 U15948 ( .A1(n15054), .A2(n14020), .ZN(n13982) );
  NAND2_X1 U15949 ( .A1(n13983), .A2(n13982), .ZN(n13984) );
  XNOR2_X1 U15950 ( .A(n13984), .B(n14111), .ZN(n13986) );
  XOR2_X1 U15951 ( .A(n13985), .B(n13986), .Z(n14270) );
  NOR2_X1 U15952 ( .A1(n15043), .A2(n14052), .ZN(n13987) );
  AOI21_X1 U15953 ( .B1(n14850), .B2(n10286), .A(n13987), .ZN(n13992) );
  NAND2_X1 U15954 ( .A1(n14850), .A2(n10284), .ZN(n13989) );
  OR2_X1 U15955 ( .A1(n15043), .A2(n14020), .ZN(n13988) );
  NAND2_X1 U15956 ( .A1(n13989), .A2(n13988), .ZN(n13990) );
  XNOR2_X1 U15957 ( .A(n13990), .B(n14111), .ZN(n13991) );
  XOR2_X1 U15958 ( .A(n13992), .B(n13991), .Z(n14099) );
  INV_X1 U15959 ( .A(n13991), .ZN(n13993) );
  NAND2_X1 U15960 ( .A1(n15030), .A2(n10284), .ZN(n13997) );
  NAND2_X1 U15961 ( .A1(n15035), .A2(n10286), .ZN(n13996) );
  NAND2_X1 U15962 ( .A1(n13997), .A2(n13996), .ZN(n13998) );
  XNOR2_X1 U15963 ( .A(n13998), .B(n14111), .ZN(n14000) );
  AOI22_X1 U15964 ( .A1(n15030), .A2(n10286), .B1(n14108), .B2(n15035), .ZN(
        n13999) );
  XNOR2_X1 U15965 ( .A(n14000), .B(n13999), .ZN(n14225) );
  INV_X1 U15966 ( .A(n13999), .ZN(n14001) );
  NAND2_X1 U15967 ( .A1(n14790), .A2(n10284), .ZN(n14003) );
  NAND2_X1 U15968 ( .A1(n14573), .A2(n10286), .ZN(n14002) );
  NAND2_X1 U15969 ( .A1(n14003), .A2(n14002), .ZN(n14004) );
  XNOR2_X1 U15970 ( .A(n14004), .B(n14051), .ZN(n14007) );
  INV_X1 U15971 ( .A(n14007), .ZN(n14009) );
  NOR2_X1 U15972 ( .A1(n15027), .A2(n14052), .ZN(n14005) );
  AOI21_X1 U15973 ( .B1(n14790), .B2(n10286), .A(n14005), .ZN(n14006) );
  INV_X1 U15974 ( .A(n14006), .ZN(n14008) );
  AOI21_X1 U15975 ( .B1(n14009), .B2(n14008), .A(n14246), .ZN(n14139) );
  OAI22_X1 U15976 ( .A1(n14804), .A2(n14011), .B1(n14010), .B2(n14020), .ZN(
        n14012) );
  XNOR2_X1 U15977 ( .A(n14012), .B(n14051), .ZN(n14015) );
  OR2_X1 U15978 ( .A1(n14804), .A2(n14020), .ZN(n14014) );
  NAND2_X1 U15979 ( .A1(n14572), .A2(n14108), .ZN(n14013) );
  AND2_X1 U15980 ( .A1(n14014), .A2(n14013), .ZN(n14016) );
  NAND2_X1 U15981 ( .A1(n14015), .A2(n14016), .ZN(n14081) );
  INV_X1 U15982 ( .A(n14015), .ZN(n14018) );
  INV_X1 U15983 ( .A(n14016), .ZN(n14017) );
  NAND2_X1 U15984 ( .A1(n14018), .A2(n14017), .ZN(n14019) );
  NAND2_X1 U15985 ( .A1(n15009), .A2(n10284), .ZN(n14022) );
  OR2_X1 U15986 ( .A1(n14251), .A2(n14020), .ZN(n14021) );
  NAND2_X1 U15987 ( .A1(n14022), .A2(n14021), .ZN(n14023) );
  XNOR2_X1 U15988 ( .A(n14023), .B(n14051), .ZN(n14026) );
  NOR2_X1 U15989 ( .A1(n14251), .A2(n14052), .ZN(n14024) );
  AOI21_X1 U15990 ( .B1(n15009), .B2(n10286), .A(n14024), .ZN(n14025) );
  NAND2_X1 U15991 ( .A1(n14026), .A2(n14025), .ZN(n14202) );
  OR2_X1 U15992 ( .A1(n14026), .A2(n14025), .ZN(n14027) );
  AND2_X1 U15993 ( .A1(n14202), .A2(n14027), .ZN(n14082) );
  NAND2_X1 U15994 ( .A1(n14028), .A2(n14082), .ZN(n14083) );
  NAND2_X1 U15995 ( .A1(n14083), .A2(n14202), .ZN(n14038) );
  NAND2_X1 U15996 ( .A1(n15006), .A2(n10284), .ZN(n14030) );
  NAND2_X1 U15997 ( .A1(n14570), .A2(n10286), .ZN(n14029) );
  NAND2_X1 U15998 ( .A1(n14030), .A2(n14029), .ZN(n14031) );
  XNOR2_X1 U15999 ( .A(n14031), .B(n14051), .ZN(n14033) );
  AND2_X1 U16000 ( .A1(n14570), .A2(n14108), .ZN(n14032) );
  AOI21_X1 U16001 ( .B1(n15006), .B2(n10286), .A(n14032), .ZN(n14034) );
  NAND2_X1 U16002 ( .A1(n14033), .A2(n14034), .ZN(n14155) );
  INV_X1 U16003 ( .A(n14033), .ZN(n14036) );
  INV_X1 U16004 ( .A(n14034), .ZN(n14035) );
  NAND2_X1 U16005 ( .A1(n14036), .A2(n14035), .ZN(n14037) );
  NAND2_X1 U16006 ( .A1(n14038), .A2(n14203), .ZN(n14154) );
  NAND2_X1 U16007 ( .A1(n14154), .A2(n14155), .ZN(n14047) );
  NAND2_X1 U16008 ( .A1(n14998), .A2(n10284), .ZN(n14040) );
  NAND2_X1 U16009 ( .A1(n14569), .A2(n10286), .ZN(n14039) );
  NAND2_X1 U16010 ( .A1(n14040), .A2(n14039), .ZN(n14041) );
  XNOR2_X1 U16011 ( .A(n14041), .B(n14051), .ZN(n14045) );
  NOR2_X1 U16012 ( .A1(n14042), .A2(n14052), .ZN(n14043) );
  AOI21_X1 U16013 ( .B1(n14998), .B2(n10286), .A(n14043), .ZN(n14044) );
  NAND2_X1 U16014 ( .A1(n14045), .A2(n14044), .ZN(n14048) );
  OR2_X1 U16015 ( .A1(n14045), .A2(n14044), .ZN(n14046) );
  NAND2_X1 U16016 ( .A1(n14994), .A2(n10284), .ZN(n14050) );
  NAND2_X1 U16017 ( .A1(n14568), .A2(n10286), .ZN(n14049) );
  INV_X1 U16018 ( .A(n14055), .ZN(n14057) );
  NOR2_X1 U16019 ( .A1(n14161), .A2(n14052), .ZN(n14053) );
  AOI21_X1 U16020 ( .B1(n14994), .B2(n10286), .A(n14053), .ZN(n14054) );
  INV_X1 U16021 ( .A(n14054), .ZN(n14056) );
  AOI22_X1 U16022 ( .A1(n14566), .A2(n15090), .B1(n15107), .B2(n14568), .ZN(
        n14721) );
  INV_X1 U16023 ( .A(n14059), .ZN(n14726) );
  AOI22_X1 U16024 ( .A1(n14726), .A2(n14295), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14060) );
  OAI21_X1 U16025 ( .B1(n14721), .B2(n14298), .A(n14060), .ZN(n14061) );
  AOI21_X1 U16026 ( .B1(n14985), .B2(n14300), .A(n14061), .ZN(n14062) );
  NAND2_X1 U16027 ( .A1(n14063), .A2(n14062), .ZN(P1_U3214) );
  XOR2_X1 U16028 ( .A(n14068), .B(n14069), .Z(n14259) );
  NAND2_X1 U16029 ( .A1(n14064), .A2(n14259), .ZN(n14258) );
  INV_X1 U16030 ( .A(n14065), .ZN(n14066) );
  XNOR2_X1 U16031 ( .A(n14067), .B(n14066), .ZN(n14147) );
  OR2_X1 U16032 ( .A1(n14069), .A2(n14068), .ZN(n14146) );
  NAND3_X1 U16033 ( .A1(n14258), .A2(n14147), .A3(n14146), .ZN(n14237) );
  AND2_X1 U16034 ( .A1(n14070), .A2(n14073), .ZN(n14235) );
  INV_X1 U16035 ( .A(n14071), .ZN(n14236) );
  NAND3_X1 U16036 ( .A1(n14237), .A2(n14235), .A3(n14236), .ZN(n14234) );
  AND3_X1 U16037 ( .A1(n14234), .A2(n14073), .A3(n14072), .ZN(n14075) );
  OAI21_X1 U16038 ( .B1(n14075), .B2(n14074), .A(n14281), .ZN(n14080) );
  OAI21_X1 U16039 ( .B1(n14286), .B2(n14936), .A(n14076), .ZN(n14078) );
  NOR2_X1 U16040 ( .A1(n14272), .A2(n15074), .ZN(n14077) );
  AOI211_X1 U16041 ( .C1(n14275), .C2(n15091), .A(n14078), .B(n14077), .ZN(
        n14079) );
  OAI211_X1 U16042 ( .C1(n14932), .C2(n14291), .A(n14080), .B(n14079), .ZN(
        P1_U3215) );
  NOR2_X1 U16043 ( .A1(n6788), .A2(n14082), .ZN(n14084) );
  INV_X1 U16044 ( .A(n14083), .ZN(n14205) );
  AOI21_X1 U16045 ( .B1(n14084), .B2(n14248), .A(n14205), .ZN(n14089) );
  AND2_X1 U16046 ( .A1(n14572), .A2(n15107), .ZN(n14085) );
  AOI21_X1 U16047 ( .B1(n14570), .B2(n15090), .A(n14085), .ZN(n14774) );
  AOI22_X1 U16048 ( .A1(n14778), .A2(n14295), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14086) );
  OAI21_X1 U16049 ( .B1(n14774), .B2(n14298), .A(n14086), .ZN(n14087) );
  AOI21_X1 U16050 ( .B1(n15009), .B2(n14300), .A(n14087), .ZN(n14088) );
  OAI21_X1 U16051 ( .B1(n14089), .B2(n14302), .A(n14088), .ZN(P1_U3216) );
  AOI21_X1 U16052 ( .B1(n14091), .B2(n14090), .A(n14302), .ZN(n14093) );
  NAND2_X1 U16053 ( .A1(n14093), .A2(n14092), .ZN(n14098) );
  AOI22_X1 U16054 ( .A1(n14288), .A2(n14095), .B1(n14094), .B2(n14300), .ZN(
        n14097) );
  MUX2_X1 U16055 ( .A(n14286), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n14096) );
  NAND3_X1 U16056 ( .A1(n14098), .A2(n14097), .A3(n14096), .ZN(P1_U3218) );
  AOI21_X1 U16057 ( .B1(n14100), .B2(n14099), .A(n14302), .ZN(n14102) );
  NAND2_X1 U16058 ( .A1(n14102), .A2(n14101), .ZN(n14107) );
  NOR2_X1 U16059 ( .A1(n14103), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14674) );
  AOI21_X1 U16060 ( .B1(n14845), .B2(n14295), .A(n14674), .ZN(n14104) );
  OAI21_X1 U16061 ( .B1(n14848), .B2(n14272), .A(n14104), .ZN(n14105) );
  AOI21_X1 U16062 ( .B1(n14275), .B2(n15034), .A(n14105), .ZN(n14106) );
  OAI211_X1 U16063 ( .C1(n15038), .C2(n14291), .A(n14107), .B(n14106), .ZN(
        P1_U3219) );
  INV_X1 U16064 ( .A(n14121), .ZN(n14115) );
  NAND2_X1 U16065 ( .A1(n14449), .A2(n10286), .ZN(n14110) );
  NAND2_X1 U16066 ( .A1(n14566), .A2(n14108), .ZN(n14109) );
  NAND2_X1 U16067 ( .A1(n14110), .A2(n14109), .ZN(n14112) );
  XNOR2_X1 U16068 ( .A(n14112), .B(n14111), .ZN(n14114) );
  AOI22_X1 U16069 ( .A1(n14449), .A2(n10284), .B1(n10286), .B2(n14566), .ZN(
        n14113) );
  XNOR2_X1 U16070 ( .A(n14114), .B(n14113), .ZN(n14123) );
  NAND3_X1 U16071 ( .A1(n14115), .A2(n14281), .A3(n14123), .ZN(n14127) );
  NOR2_X1 U16072 ( .A1(n14484), .A2(n14272), .ZN(n14118) );
  AOI22_X1 U16073 ( .A1(n14708), .A2(n14295), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14116) );
  OAI21_X1 U16074 ( .B1(n14311), .B2(n14227), .A(n14116), .ZN(n14117) );
  AOI211_X1 U16075 ( .C1(n14449), .C2(n14300), .A(n14118), .B(n14117), .ZN(
        n14126) );
  INV_X1 U16076 ( .A(n14122), .ZN(n14120) );
  INV_X1 U16077 ( .A(n14123), .ZN(n14119) );
  NAND4_X1 U16078 ( .A1(n14121), .A2(n14281), .A3(n14120), .A4(n14119), .ZN(
        n14125) );
  NAND3_X1 U16079 ( .A1(n14123), .A2(n14122), .A3(n14281), .ZN(n14124) );
  NAND4_X1 U16080 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        P1_U3220) );
  XNOR2_X1 U16081 ( .A(n14128), .B(n14129), .ZN(n14130) );
  NAND2_X1 U16082 ( .A1(n14130), .A2(n14281), .ZN(n14137) );
  AOI22_X1 U16083 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n14132), .B1(n14300), 
        .B2(n14131), .ZN(n14136) );
  NAND2_X1 U16084 ( .A1(n14275), .A2(n14581), .ZN(n14135) );
  NAND2_X1 U16085 ( .A1(n14133), .A2(n14580), .ZN(n14134) );
  NAND4_X1 U16086 ( .A1(n14137), .A2(n14136), .A3(n14135), .A4(n14134), .ZN(
        P1_U3222) );
  OAI21_X1 U16087 ( .B1(n14140), .B2(n14139), .A(n14138), .ZN(n14141) );
  NAND2_X1 U16088 ( .A1(n14141), .A2(n14281), .ZN(n14145) );
  AOI22_X1 U16089 ( .A1(n14572), .A2(n15090), .B1(n15035), .B2(n15107), .ZN(
        n14812) );
  INV_X1 U16090 ( .A(n14812), .ZN(n14143) );
  OAI22_X1 U16091 ( .A1(n14818), .A2(n14286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15581), .ZN(n14142) );
  AOI21_X1 U16092 ( .B1(n14143), .B2(n14288), .A(n14142), .ZN(n14144) );
  OAI211_X1 U16093 ( .C1(n15021), .C2(n14291), .A(n14145), .B(n14144), .ZN(
        P1_U3223) );
  INV_X1 U16094 ( .A(n14972), .ZN(n15095) );
  AND2_X1 U16095 ( .A1(n14258), .A2(n14146), .ZN(n14148) );
  OAI211_X1 U16096 ( .C1(n14148), .C2(n14147), .A(n14281), .B(n14237), .ZN(
        n14153) );
  OAI22_X1 U16097 ( .A1(n14286), .A2(n14965), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14149), .ZN(n14151) );
  NOR2_X1 U16098 ( .A1(n14272), .A2(n15075), .ZN(n14150) );
  AOI211_X1 U16099 ( .C1(n14275), .C2(n15092), .A(n14151), .B(n14150), .ZN(
        n14152) );
  OAI211_X1 U16100 ( .C1(n15095), .C2(n14291), .A(n14153), .B(n14152), .ZN(
        P1_U3224) );
  INV_X1 U16101 ( .A(n14154), .ZN(n14206) );
  INV_X1 U16102 ( .A(n14155), .ZN(n14157) );
  NOR3_X1 U16103 ( .A1(n14206), .A2(n14157), .A3(n14156), .ZN(n14159) );
  OAI21_X1 U16104 ( .B1(n14159), .B2(n6714), .A(n14281), .ZN(n14165) );
  OAI22_X1 U16105 ( .A1(n14161), .A2(n15310), .B1(n14160), .B2(n15312), .ZN(
        n14997) );
  OAI22_X1 U16106 ( .A1(n14753), .A2(n14286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14162), .ZN(n14163) );
  AOI21_X1 U16107 ( .B1(n14997), .B2(n14288), .A(n14163), .ZN(n14164) );
  OAI211_X1 U16108 ( .C1(n14755), .C2(n14291), .A(n14165), .B(n14164), .ZN(
        P1_U3225) );
  NAND2_X1 U16109 ( .A1(n14166), .A2(n14191), .ZN(n14170) );
  XOR2_X1 U16110 ( .A(n14168), .B(n14167), .Z(n14293) );
  OAI22_X1 U16111 ( .A1(n14293), .A2(n14292), .B1(n14168), .B2(n6803), .ZN(
        n14169) );
  NOR2_X1 U16112 ( .A1(n14169), .A2(n14170), .ZN(n14194) );
  AOI21_X1 U16113 ( .B1(n14170), .B2(n14169), .A(n14194), .ZN(n14176) );
  OAI21_X1 U16114 ( .B1(n14286), .B2(n14894), .A(n14171), .ZN(n14173) );
  NOR2_X1 U16115 ( .A1(n14272), .A2(n15061), .ZN(n14172) );
  AOI211_X1 U16116 ( .C1(n14275), .C2(n14897), .A(n14173), .B(n14172), .ZN(
        n14175) );
  NAND2_X1 U16117 ( .A1(n15064), .A2(n14300), .ZN(n14174) );
  OAI211_X1 U16118 ( .C1(n14176), .C2(n14302), .A(n14175), .B(n14174), .ZN(
        P1_U3226) );
  XNOR2_X1 U16119 ( .A(n14178), .B(n14177), .ZN(n14179) );
  XNOR2_X1 U16120 ( .A(n14180), .B(n14179), .ZN(n14181) );
  NAND2_X1 U16121 ( .A1(n14181), .A2(n14281), .ZN(n14190) );
  INV_X1 U16122 ( .A(n14182), .ZN(n14183) );
  AOI21_X1 U16123 ( .B1(n14300), .B2(n6407), .A(n14183), .ZN(n14189) );
  NAND2_X1 U16124 ( .A1(n15250), .A2(n15107), .ZN(n14185) );
  NAND2_X1 U16125 ( .A1(n14577), .A2(n15090), .ZN(n14184) );
  NAND2_X1 U16126 ( .A1(n14185), .A2(n14184), .ZN(n15256) );
  NAND2_X1 U16127 ( .A1(n14288), .A2(n15256), .ZN(n14188) );
  INV_X1 U16128 ( .A(n14186), .ZN(n15259) );
  NAND2_X1 U16129 ( .A1(n14295), .A2(n15259), .ZN(n14187) );
  NAND4_X1 U16130 ( .A1(n14190), .A2(n14189), .A3(n14188), .A4(n14187), .ZN(
        P1_U3227) );
  INV_X1 U16131 ( .A(n15057), .ZN(n14886) );
  INV_X1 U16132 ( .A(n14191), .ZN(n14193) );
  NOR3_X1 U16133 ( .A1(n14194), .A2(n14193), .A3(n14192), .ZN(n14197) );
  INV_X1 U16134 ( .A(n14195), .ZN(n14196) );
  OAI21_X1 U16135 ( .B1(n14197), .B2(n14196), .A(n14281), .ZN(n14201) );
  NAND2_X1 U16136 ( .A1(n14295), .A2(n14881), .ZN(n14198) );
  NAND2_X1 U16137 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14639)
         );
  OAI211_X1 U16138 ( .C1(n15054), .C2(n14272), .A(n14198), .B(n14639), .ZN(
        n14199) );
  AOI21_X1 U16139 ( .B1(n14275), .B2(n14884), .A(n14199), .ZN(n14200) );
  OAI211_X1 U16140 ( .C1(n14886), .C2(n14291), .A(n14201), .B(n14200), .ZN(
        P1_U3228) );
  INV_X1 U16141 ( .A(n14202), .ZN(n14204) );
  NOR3_X1 U16142 ( .A1(n14205), .A2(n14204), .A3(n14203), .ZN(n14207) );
  OAI21_X1 U16143 ( .B1(n14207), .B2(n14206), .A(n14281), .ZN(n14213) );
  OAI22_X1 U16144 ( .A1(n14209), .A2(n14286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14208), .ZN(n14210) );
  AOI21_X1 U16145 ( .B1(n14211), .B2(n14288), .A(n14210), .ZN(n14212) );
  OAI211_X1 U16146 ( .C1(n14214), .C2(n14291), .A(n14213), .B(n14212), .ZN(
        P1_U3229) );
  AOI21_X1 U16147 ( .B1(n14217), .B2(n14216), .A(n14215), .ZN(n14224) );
  NAND2_X1 U16148 ( .A1(n14275), .A2(n14575), .ZN(n14221) );
  AOI21_X1 U16149 ( .B1(n14295), .B2(n14219), .A(n14218), .ZN(n14220) );
  OAI211_X1 U16150 ( .C1(n14360), .C2(n14272), .A(n14221), .B(n14220), .ZN(
        n14222) );
  AOI21_X1 U16151 ( .B1(n14355), .B2(n14300), .A(n14222), .ZN(n14223) );
  OAI21_X1 U16152 ( .B1(n14224), .B2(n14302), .A(n14223), .ZN(P1_U3231) );
  XNOR2_X1 U16153 ( .A(n14226), .B(n14225), .ZN(n14233) );
  NOR2_X1 U16154 ( .A1(n15043), .A2(n14227), .ZN(n14231) );
  INV_X1 U16155 ( .A(n14228), .ZN(n14830) );
  AOI22_X1 U16156 ( .A1(n14830), .A2(n14295), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14229) );
  OAI21_X1 U16157 ( .B1(n15027), .B2(n14272), .A(n14229), .ZN(n14230) );
  AOI211_X1 U16158 ( .C1(n15030), .C2(n14300), .A(n14231), .B(n14230), .ZN(
        n14232) );
  OAI21_X1 U16159 ( .B1(n14233), .B2(n14302), .A(n14232), .ZN(P1_U3233) );
  INV_X1 U16160 ( .A(n14234), .ZN(n14239) );
  AOI21_X1 U16161 ( .B1(n14237), .B2(n14236), .A(n14235), .ZN(n14238) );
  OAI21_X1 U16162 ( .B1(n14239), .B2(n14238), .A(n14281), .ZN(n14244) );
  OAI21_X1 U16163 ( .B1(n14286), .B2(n14947), .A(n14240), .ZN(n14242) );
  NOR2_X1 U16164 ( .A1(n14272), .A2(n15082), .ZN(n14241) );
  AOI211_X1 U16165 ( .C1(n14275), .C2(n14946), .A(n14242), .B(n14241), .ZN(
        n14243) );
  OAI211_X1 U16166 ( .C1(n7446), .C2(n14291), .A(n14244), .B(n14243), .ZN(
        P1_U3234) );
  INV_X1 U16167 ( .A(n14138), .ZN(n14247) );
  NOR3_X1 U16168 ( .A1(n14247), .A2(n14246), .A3(n14245), .ZN(n14250) );
  INV_X1 U16169 ( .A(n14248), .ZN(n14249) );
  OAI21_X1 U16170 ( .B1(n14250), .B2(n14249), .A(n14281), .ZN(n14257) );
  OR2_X1 U16171 ( .A1(n14251), .A2(n15310), .ZN(n14253) );
  NAND2_X1 U16172 ( .A1(n14573), .A2(n15107), .ZN(n14252) );
  NAND2_X1 U16173 ( .A1(n14253), .A2(n14252), .ZN(n14795) );
  OAI22_X1 U16174 ( .A1(n14801), .A2(n14286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14254), .ZN(n14255) );
  AOI21_X1 U16175 ( .B1(n14795), .B2(n14288), .A(n14255), .ZN(n14256) );
  OAI211_X1 U16176 ( .C1(n14291), .C2(n14804), .A(n14257), .B(n14256), .ZN(
        P1_U3235) );
  OAI21_X1 U16177 ( .B1(n14259), .B2(n14064), .A(n14258), .ZN(n14260) );
  NAND2_X1 U16178 ( .A1(n14260), .A2(n14281), .ZN(n14267) );
  INV_X1 U16179 ( .A(n14261), .ZN(n14265) );
  OAI21_X1 U16180 ( .B1(n14286), .B2(n14263), .A(n14262), .ZN(n14264) );
  AOI21_X1 U16181 ( .B1(n14288), .B2(n14265), .A(n14264), .ZN(n14266) );
  OAI211_X1 U16182 ( .C1(n14363), .C2(n14291), .A(n14267), .B(n14266), .ZN(
        P1_U3236) );
  OAI21_X1 U16183 ( .B1(n14270), .B2(n14269), .A(n14268), .ZN(n14271) );
  NAND2_X1 U16184 ( .A1(n14271), .A2(n14281), .ZN(n14277) );
  NAND2_X1 U16185 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14651)
         );
  OAI21_X1 U16186 ( .B1(n14286), .B2(n14859), .A(n14651), .ZN(n14274) );
  NOR2_X1 U16187 ( .A1(n15043), .A2(n14272), .ZN(n14273) );
  AOI211_X1 U16188 ( .C1(n14275), .C2(n14858), .A(n14274), .B(n14273), .ZN(
        n14276) );
  OAI211_X1 U16189 ( .C1(n14855), .C2(n14291), .A(n14277), .B(n14276), .ZN(
        P1_U3238) );
  OAI21_X1 U16190 ( .B1(n14280), .B2(n14279), .A(n14278), .ZN(n14282) );
  NAND2_X1 U16191 ( .A1(n14282), .A2(n14281), .ZN(n14290) );
  NAND2_X1 U16192 ( .A1(n14567), .A2(n15090), .ZN(n14284) );
  NAND2_X1 U16193 ( .A1(n14569), .A2(n15107), .ZN(n14283) );
  NAND2_X1 U16194 ( .A1(n14284), .A2(n14283), .ZN(n14737) );
  OAI22_X1 U16195 ( .A1(n6715), .A2(n14286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14285), .ZN(n14287) );
  AOI21_X1 U16196 ( .B1(n14737), .B2(n14288), .A(n14287), .ZN(n14289) );
  OAI211_X1 U16197 ( .C1(n7452), .C2(n14291), .A(n14290), .B(n14289), .ZN(
        P1_U3240) );
  XNOR2_X1 U16198 ( .A(n14293), .B(n14292), .ZN(n14303) );
  OAI22_X1 U16199 ( .A1(n15053), .A2(n15310), .B1(n15082), .B2(n15312), .ZN(
        n14294) );
  INV_X1 U16200 ( .A(n14294), .ZN(n14913) );
  NAND2_X1 U16201 ( .A1(n14295), .A2(n14919), .ZN(n14296) );
  OAI211_X1 U16202 ( .C1(n14913), .C2(n14298), .A(n14297), .B(n14296), .ZN(
        n14299) );
  AOI21_X1 U16203 ( .B1(n15071), .B2(n14300), .A(n14299), .ZN(n14301) );
  OAI21_X1 U16204 ( .B1(n14303), .B2(n14302), .A(n14301), .ZN(P1_U3241) );
  OR2_X1 U16205 ( .A1(n14304), .A2(n14672), .ZN(n14306) );
  NAND2_X1 U16206 ( .A1(n14309), .A2(n14476), .ZN(n14310) );
  MUX2_X1 U16207 ( .A(n14311), .B(n7451), .S(n14460), .Z(n14447) );
  NAND2_X1 U16208 ( .A1(n14580), .A2(n14448), .ZN(n14312) );
  OAI211_X1 U16209 ( .C1(n14448), .C2(n8756), .A(n9230), .B(n14312), .ZN(
        n14325) );
  NAND2_X1 U16210 ( .A1(n14313), .A2(n14479), .ZN(n14314) );
  NAND2_X1 U16211 ( .A1(n14314), .A2(n10152), .ZN(n14316) );
  NAND2_X1 U16212 ( .A1(n14316), .A2(n14315), .ZN(n14319) );
  NAND4_X1 U16213 ( .A1(n14319), .A2(n14483), .A3(n14318), .A4(n14317), .ZN(
        n14324) );
  NAND2_X1 U16214 ( .A1(n14321), .A2(n14320), .ZN(n14322) );
  NAND4_X1 U16215 ( .A1(n14325), .A2(n14324), .A3(n14323), .A4(n14322), .ZN(
        n14329) );
  MUX2_X1 U16216 ( .A(n14327), .B(n14326), .S(n14448), .Z(n14328) );
  NAND2_X1 U16217 ( .A1(n14329), .A2(n14328), .ZN(n14332) );
  MUX2_X1 U16218 ( .A(n15246), .B(n15247), .S(n14483), .Z(n14331) );
  MUX2_X1 U16219 ( .A(n15250), .B(n15285), .S(n14485), .Z(n14330) );
  NAND2_X1 U16220 ( .A1(n14332), .A2(n14331), .ZN(n14333) );
  MUX2_X1 U16221 ( .A(n14578), .B(n6407), .S(n14485), .Z(n14337) );
  MUX2_X1 U16222 ( .A(n6407), .B(n14578), .S(n14485), .Z(n14335) );
  INV_X1 U16223 ( .A(n14337), .ZN(n14338) );
  MUX2_X1 U16224 ( .A(n14339), .B(n14577), .S(n14485), .Z(n14343) );
  NAND2_X1 U16225 ( .A1(n14342), .A2(n14343), .ZN(n14341) );
  MUX2_X1 U16226 ( .A(n14339), .B(n14577), .S(n14448), .Z(n14340) );
  NAND2_X1 U16227 ( .A1(n14341), .A2(n14340), .ZN(n14347) );
  INV_X1 U16228 ( .A(n14343), .ZN(n14344) );
  NAND2_X1 U16229 ( .A1(n14345), .A2(n14344), .ZN(n14346) );
  MUX2_X1 U16230 ( .A(n14576), .B(n14348), .S(n14485), .Z(n14350) );
  MUX2_X1 U16231 ( .A(n14348), .B(n14576), .S(n14485), .Z(n14349) );
  MUX2_X1 U16232 ( .A(n15316), .B(n14575), .S(n14485), .Z(n14353) );
  MUX2_X1 U16233 ( .A(n14575), .B(n15316), .S(n14485), .Z(n14351) );
  INV_X1 U16234 ( .A(n14353), .ZN(n14354) );
  MUX2_X1 U16235 ( .A(n14355), .B(n15106), .S(n14460), .Z(n14357) );
  MUX2_X1 U16236 ( .A(n7437), .B(n15311), .S(n14485), .Z(n14356) );
  AOI21_X1 U16237 ( .B1(n14358), .B2(n14357), .A(n14356), .ZN(n14362) );
  MUX2_X1 U16238 ( .A(n14360), .B(n14359), .S(n14485), .Z(n14365) );
  MUX2_X1 U16239 ( .A(n15108), .B(n14574), .S(n14485), .Z(n14366) );
  OAI22_X1 U16240 ( .A1(n14362), .A2(n14361), .B1(n14365), .B2(n14366), .ZN(
        n14385) );
  MUX2_X1 U16241 ( .A(n15092), .B(n7165), .S(n14485), .Z(n14374) );
  INV_X1 U16242 ( .A(n14374), .ZN(n14371) );
  MUX2_X1 U16243 ( .A(n14364), .B(n14363), .S(n14460), .Z(n14375) );
  INV_X1 U16244 ( .A(n14375), .ZN(n14370) );
  INV_X1 U16245 ( .A(n14365), .ZN(n14368) );
  INV_X1 U16246 ( .A(n14366), .ZN(n14367) );
  MUX2_X1 U16247 ( .A(n15083), .B(n15095), .S(n14485), .Z(n14377) );
  MUX2_X1 U16248 ( .A(n14946), .B(n14972), .S(n14448), .Z(n14376) );
  NAND2_X1 U16249 ( .A1(n14377), .A2(n14376), .ZN(n14373) );
  OAI21_X1 U16250 ( .B1(n14368), .B2(n14367), .A(n14373), .ZN(n14369) );
  AOI21_X1 U16251 ( .B1(n14371), .B2(n14370), .A(n14369), .ZN(n14384) );
  MUX2_X1 U16252 ( .A(n15091), .B(n15086), .S(n14485), .Z(n14386) );
  NAND2_X1 U16253 ( .A1(n15086), .A2(n14460), .ZN(n14372) );
  OAI211_X1 U16254 ( .C1(n14448), .C2(n15075), .A(n14386), .B(n14372), .ZN(
        n14382) );
  NAND3_X1 U16255 ( .A1(n14375), .A2(n14374), .A3(n14373), .ZN(n14381) );
  INV_X1 U16256 ( .A(n14376), .ZN(n14379) );
  INV_X1 U16257 ( .A(n14377), .ZN(n14378) );
  NAND2_X1 U16258 ( .A1(n14379), .A2(n14378), .ZN(n14380) );
  NAND4_X1 U16259 ( .A1(n14381), .A2(n14382), .A3(n14930), .A4(n14380), .ZN(
        n14383) );
  AOI21_X1 U16260 ( .B1(n14385), .B2(n14384), .A(n14383), .ZN(n14394) );
  INV_X1 U16261 ( .A(n14386), .ZN(n14388) );
  MUX2_X1 U16262 ( .A(n15091), .B(n15086), .S(n14460), .Z(n14387) );
  AND3_X1 U16263 ( .A1(n14930), .A2(n14388), .A3(n14387), .ZN(n14393) );
  AOI21_X1 U16264 ( .B1(n14395), .B2(n14389), .A(n14483), .ZN(n14392) );
  AOI21_X1 U16265 ( .B1(n14872), .B2(n14390), .A(n14448), .ZN(n14391) );
  MUX2_X1 U16266 ( .A(n14395), .B(n14872), .S(n14460), .Z(n14396) );
  MUX2_X1 U16267 ( .A(n14884), .B(n15064), .S(n14485), .Z(n14398) );
  MUX2_X1 U16268 ( .A(n14884), .B(n15064), .S(n14460), .Z(n14397) );
  XNOR2_X1 U16269 ( .A(n15057), .B(n15061), .ZN(n14877) );
  NOR2_X1 U16270 ( .A1(n14399), .A2(n14877), .ZN(n14543) );
  MUX2_X1 U16271 ( .A(n15034), .B(n15045), .S(n14485), .Z(n14400) );
  NAND2_X1 U16272 ( .A1(n7862), .A2(n14400), .ZN(n14407) );
  NOR2_X1 U16273 ( .A1(n15061), .A2(n14448), .ZN(n14402) );
  OAI21_X1 U16274 ( .B1(n14858), .B2(n14483), .A(n15057), .ZN(n14401) );
  OAI21_X1 U16275 ( .B1(n14402), .B2(n15057), .A(n14401), .ZN(n14403) );
  NAND3_X1 U16276 ( .A1(n14405), .A2(n14404), .A3(n14403), .ZN(n14406) );
  NAND2_X1 U16277 ( .A1(n14407), .A2(n14406), .ZN(n14410) );
  NAND3_X1 U16278 ( .A1(n14850), .A2(n15043), .A3(n14448), .ZN(n14409) );
  OR3_X1 U16279 ( .A1(n14850), .A2(n14448), .A3(n15043), .ZN(n14408) );
  OAI211_X1 U16280 ( .C1(n14410), .C2(n14399), .A(n14409), .B(n14408), .ZN(
        n14411) );
  INV_X1 U16281 ( .A(n14411), .ZN(n14412) );
  NAND2_X1 U16282 ( .A1(n14413), .A2(n14412), .ZN(n14416) );
  INV_X1 U16283 ( .A(n15030), .ZN(n14835) );
  MUX2_X1 U16284 ( .A(n14848), .B(n14835), .S(n14485), .Z(n14415) );
  MUX2_X1 U16285 ( .A(n15035), .B(n15030), .S(n14448), .Z(n14414) );
  NAND2_X1 U16286 ( .A1(n14416), .A2(n14415), .ZN(n14417) );
  MUX2_X1 U16287 ( .A(n14573), .B(n14790), .S(n14460), .Z(n14419) );
  MUX2_X1 U16288 ( .A(n14573), .B(n14790), .S(n14485), .Z(n14420) );
  MUX2_X1 U16289 ( .A(n14572), .B(n15017), .S(n14483), .Z(n14422) );
  MUX2_X1 U16290 ( .A(n14572), .B(n15017), .S(n14460), .Z(n14421) );
  INV_X1 U16291 ( .A(n14422), .ZN(n14423) );
  MUX2_X1 U16292 ( .A(n14571), .B(n15009), .S(n14460), .Z(n14425) );
  MUX2_X1 U16293 ( .A(n14571), .B(n15009), .S(n14485), .Z(n14424) );
  INV_X1 U16294 ( .A(n14425), .ZN(n14426) );
  MUX2_X1 U16295 ( .A(n14570), .B(n15006), .S(n14483), .Z(n14430) );
  MUX2_X1 U16296 ( .A(n14570), .B(n15006), .S(n14460), .Z(n14427) );
  NAND2_X1 U16297 ( .A1(n14428), .A2(n14427), .ZN(n14434) );
  INV_X1 U16298 ( .A(n14429), .ZN(n14432) );
  INV_X1 U16299 ( .A(n14430), .ZN(n14431) );
  MUX2_X1 U16300 ( .A(n14569), .B(n14998), .S(n14448), .Z(n14436) );
  MUX2_X1 U16301 ( .A(n14569), .B(n14998), .S(n14485), .Z(n14435) );
  INV_X1 U16302 ( .A(n14436), .ZN(n14437) );
  MUX2_X1 U16303 ( .A(n14568), .B(n14994), .S(n14485), .Z(n14441) );
  MUX2_X1 U16304 ( .A(n14994), .B(n14568), .S(n14483), .Z(n14438) );
  INV_X1 U16305 ( .A(n14440), .ZN(n14443) );
  INV_X1 U16306 ( .A(n14441), .ZN(n14442) );
  NAND2_X1 U16307 ( .A1(n14443), .A2(n14442), .ZN(n14444) );
  MUX2_X1 U16308 ( .A(n14567), .B(n14985), .S(n14485), .Z(n14446) );
  MUX2_X1 U16309 ( .A(n14697), .B(n14710), .S(n14448), .Z(n14488) );
  MUX2_X1 U16310 ( .A(n14566), .B(n14449), .S(n14483), .Z(n14487) );
  NAND2_X1 U16311 ( .A1(n15140), .A2(n6409), .ZN(n14452) );
  INV_X1 U16312 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15136) );
  OR2_X1 U16313 ( .A1(n14466), .A2(n15136), .ZN(n14451) );
  NAND2_X1 U16314 ( .A1(n14453), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n14459) );
  INV_X1 U16315 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14454) );
  OR2_X1 U16316 ( .A1(n14455), .A2(n14454), .ZN(n14458) );
  INV_X1 U16317 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14456) );
  OR2_X1 U16318 ( .A1(n8759), .A2(n14456), .ZN(n14457) );
  AND3_X1 U16319 ( .A1(n14459), .A2(n14458), .A3(n14457), .ZN(n14680) );
  OR2_X1 U16320 ( .A1(n14681), .A2(n14680), .ZN(n14462) );
  NAND2_X1 U16321 ( .A1(n14681), .A2(n14680), .ZN(n14461) );
  OR2_X1 U16322 ( .A1(n14466), .A2(n14465), .ZN(n14467) );
  INV_X1 U16323 ( .A(n14680), .ZN(n14563) );
  INV_X1 U16324 ( .A(n14468), .ZN(n14469) );
  OAI21_X1 U16325 ( .B1(n14563), .B2(n14469), .A(n14564), .ZN(n14470) );
  INV_X1 U16326 ( .A(n14470), .ZN(n14471) );
  MUX2_X1 U16327 ( .A(n14689), .B(n14471), .S(n14483), .Z(n14509) );
  INV_X1 U16328 ( .A(n14509), .ZN(n14482) );
  NAND2_X1 U16329 ( .A1(n14689), .A2(n14483), .ZN(n14475) );
  OAI21_X1 U16330 ( .B1(n14680), .B2(n14483), .A(n14472), .ZN(n14473) );
  NAND2_X1 U16331 ( .A1(n14473), .A2(n14564), .ZN(n14474) );
  NAND2_X1 U16332 ( .A1(n14475), .A2(n14474), .ZN(n14507) );
  OR2_X1 U16333 ( .A1(n14304), .A2(n14476), .ZN(n14477) );
  NAND2_X1 U16334 ( .A1(n14478), .A2(n14477), .ZN(n14481) );
  NAND2_X1 U16335 ( .A1(n14479), .A2(n14672), .ZN(n14480) );
  NAND2_X1 U16336 ( .A1(n14481), .A2(n14480), .ZN(n14506) );
  INV_X1 U16337 ( .A(n14486), .ZN(n14702) );
  MUX2_X1 U16338 ( .A(n14702), .B(n14484), .S(n14483), .Z(n14497) );
  INV_X1 U16339 ( .A(n14484), .ZN(n14565) );
  MUX2_X1 U16340 ( .A(n14565), .B(n14486), .S(n14485), .Z(n14496) );
  NAND2_X1 U16341 ( .A1(n14497), .A2(n14496), .ZN(n14504) );
  INV_X1 U16342 ( .A(n14487), .ZN(n14490) );
  INV_X1 U16343 ( .A(n14488), .ZN(n14489) );
  NAND2_X1 U16344 ( .A1(n14490), .A2(n14489), .ZN(n14521) );
  XNOR2_X1 U16345 ( .A(n14681), .B(n14563), .ZN(n14551) );
  INV_X1 U16346 ( .A(n14507), .ZN(n14493) );
  INV_X1 U16347 ( .A(n14506), .ZN(n14512) );
  AOI21_X1 U16348 ( .B1(n14509), .B2(n14493), .A(n14512), .ZN(n14492) );
  AND2_X1 U16349 ( .A1(n14551), .A2(n14492), .ZN(n14500) );
  INV_X1 U16350 ( .A(n14500), .ZN(n14503) );
  NAND3_X1 U16351 ( .A1(n14509), .A2(n14512), .A3(n14493), .ZN(n14495) );
  INV_X1 U16352 ( .A(n14513), .ZN(n14494) );
  MUX2_X1 U16353 ( .A(n14495), .B(n14512), .S(n14494), .Z(n14502) );
  INV_X1 U16354 ( .A(n14496), .ZN(n14499) );
  INV_X1 U16355 ( .A(n14497), .ZN(n14498) );
  NAND2_X1 U16356 ( .A1(n14499), .A2(n14498), .ZN(n14516) );
  NAND2_X1 U16357 ( .A1(n14500), .A2(n14516), .ZN(n14520) );
  OR2_X1 U16358 ( .A1(n14520), .A2(n6526), .ZN(n14501) );
  OAI211_X1 U16359 ( .C1(n14504), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        n14519) );
  INV_X1 U16360 ( .A(n14505), .ZN(n14517) );
  NAND2_X1 U16361 ( .A1(n14507), .A2(n14506), .ZN(n14508) );
  NOR2_X1 U16362 ( .A1(n14509), .A2(n14508), .ZN(n14510) );
  AOI21_X1 U16363 ( .B1(n14551), .B2(n14510), .A(n14554), .ZN(n14515) );
  INV_X1 U16364 ( .A(n14551), .ZN(n14511) );
  NAND3_X1 U16365 ( .A1(n14513), .A2(n14512), .A3(n14511), .ZN(n14514) );
  OAI211_X1 U16366 ( .C1(n14517), .C2(n14516), .A(n14515), .B(n14514), .ZN(
        n14518) );
  INV_X1 U16367 ( .A(n14520), .ZN(n14522) );
  NAND3_X1 U16368 ( .A1(n14523), .A2(n14522), .A3(n14521), .ZN(n14556) );
  XOR2_X1 U16369 ( .A(n14689), .B(n14564), .Z(n14550) );
  NOR2_X1 U16370 ( .A1(n14526), .A2(n14525), .ZN(n14529) );
  NAND4_X1 U16371 ( .A1(n14529), .A2(n14528), .A3(n15252), .A4(n14527), .ZN(
        n14531) );
  NOR2_X1 U16372 ( .A1(n14531), .A2(n14530), .ZN(n14533) );
  INV_X1 U16373 ( .A(n15227), .ZN(n15229) );
  NAND4_X1 U16374 ( .A1(n8871), .A2(n14533), .A3(n15229), .A4(n14532), .ZN(
        n14534) );
  NOR2_X1 U16375 ( .A1(n14535), .A2(n14534), .ZN(n14537) );
  AND2_X1 U16376 ( .A1(n14944), .A2(n14961), .ZN(n14536) );
  AND4_X1 U16377 ( .A1(n14930), .A2(n14538), .A3(n14537), .A4(n14536), .ZN(
        n14540) );
  NAND4_X1 U16378 ( .A1(n14912), .A2(n14540), .A3(n7050), .A4(n14539), .ZN(
        n14541) );
  XNOR2_X1 U16379 ( .A(n14790), .B(n14573), .ZN(n14815) );
  NAND4_X1 U16380 ( .A1(n7882), .A2(n14543), .A3(n14791), .A4(n14815), .ZN(
        n14544) );
  NOR2_X1 U16381 ( .A1(n14733), .A2(n14544), .ZN(n14546) );
  NAND4_X1 U16382 ( .A1(n14547), .A2(n14546), .A3(n14545), .A4(n14718), .ZN(
        n14548) );
  NOR4_X1 U16383 ( .A1(n14550), .A2(n14549), .A3(n14746), .A4(n14548), .ZN(
        n14552) );
  NAND2_X1 U16384 ( .A1(n14552), .A2(n14551), .ZN(n14553) );
  XNOR2_X1 U16385 ( .A(n14553), .B(n14672), .ZN(n14555) );
  AOI22_X1 U16386 ( .A1(n14557), .A2(n14556), .B1(n14555), .B2(n14554), .ZN(
        n14562) );
  NOR3_X1 U16387 ( .A1(n14558), .A2(n6410), .A3(n15312), .ZN(n14560) );
  OAI21_X1 U16388 ( .B1(n14561), .B2(n14304), .A(P1_B_REG_SCAN_IN), .ZN(n14559) );
  OAI22_X1 U16389 ( .A1(n14562), .A2(n14561), .B1(n14560), .B2(n14559), .ZN(
        P1_U3242) );
  MUX2_X1 U16390 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14563), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16391 ( .A(n14564), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14600), .Z(
        P1_U3590) );
  MUX2_X1 U16392 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14565), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16393 ( .A(n14566), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14600), .Z(
        P1_U3588) );
  MUX2_X1 U16394 ( .A(n14567), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14600), .Z(
        P1_U3587) );
  MUX2_X1 U16395 ( .A(n14568), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14600), .Z(
        P1_U3586) );
  MUX2_X1 U16396 ( .A(n14569), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14600), .Z(
        P1_U3585) );
  MUX2_X1 U16397 ( .A(n14570), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14600), .Z(
        P1_U3584) );
  MUX2_X1 U16398 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14571), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16399 ( .A(n14572), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14600), .Z(
        P1_U3582) );
  MUX2_X1 U16400 ( .A(n14573), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14600), .Z(
        P1_U3581) );
  MUX2_X1 U16401 ( .A(n15035), .B(P1_DATAO_REG_20__SCAN_IN), .S(n14600), .Z(
        P1_U3580) );
  MUX2_X1 U16402 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14833), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16403 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15034), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16404 ( .A(n14858), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14600), .Z(
        P1_U3577) );
  MUX2_X1 U16405 ( .A(n14884), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14600), .Z(
        P1_U3576) );
  MUX2_X1 U16406 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14897), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16407 ( .A(n15091), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14600), .Z(
        P1_U3573) );
  MUX2_X1 U16408 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14946), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16409 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15092), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16410 ( .A(n14574), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14600), .Z(
        P1_U3570) );
  MUX2_X1 U16411 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15106), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16412 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14575), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16413 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14576), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16414 ( .A(n14577), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14600), .Z(
        P1_U3566) );
  MUX2_X1 U16415 ( .A(n14578), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14600), .Z(
        P1_U3565) );
  MUX2_X1 U16416 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15250), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16417 ( .A(n14579), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14600), .Z(
        P1_U3563) );
  MUX2_X1 U16418 ( .A(n14580), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14600), .Z(
        P1_U3562) );
  MUX2_X1 U16419 ( .A(n9228), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14600), .Z(
        P1_U3561) );
  MUX2_X1 U16420 ( .A(n14581), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14600), .Z(
        P1_U3560) );
  OAI22_X1 U16421 ( .A1(n15226), .A2(n14583), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14582), .ZN(n14584) );
  AOI21_X1 U16422 ( .B1(n14654), .B2(n14585), .A(n14584), .ZN(n14595) );
  MUX2_X1 U16423 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10158), .S(n14586), .Z(
        n14587) );
  INV_X1 U16424 ( .A(n14587), .ZN(n14589) );
  OAI211_X1 U16425 ( .C1(n14590), .C2(n14589), .A(n15210), .B(n14588), .ZN(
        n14594) );
  NAND2_X1 U16426 ( .A1(n7069), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14597) );
  OAI211_X1 U16427 ( .C1(n10171), .C2(n14592), .A(n15217), .B(n14591), .ZN(
        n14593) );
  NAND3_X1 U16428 ( .A1(n14595), .A2(n14594), .A3(n14593), .ZN(P1_U3244) );
  MUX2_X1 U16429 ( .A(n14597), .B(n14596), .S(n6410), .Z(n14598) );
  NOR2_X1 U16430 ( .A1(n14598), .A2(n9286), .ZN(n14599) );
  INV_X1 U16431 ( .A(n15223), .ZN(n14614) );
  OAI22_X1 U16432 ( .A1(n15226), .A2(n14602), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8739), .ZN(n14603) );
  AOI21_X1 U16433 ( .B1(n14654), .B2(n14604), .A(n14603), .ZN(n14613) );
  MUX2_X1 U16434 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10160), .S(n14605), .Z(
        n14606) );
  INV_X1 U16435 ( .A(n14606), .ZN(n14608) );
  OAI211_X1 U16436 ( .C1(n14608), .C2(n14607), .A(n15210), .B(n14619), .ZN(
        n14612) );
  OAI211_X1 U16437 ( .C1(n14610), .C2(n14609), .A(n15217), .B(n14624), .ZN(
        n14611) );
  NAND4_X1 U16438 ( .A1(n14614), .A2(n14613), .A3(n14612), .A4(n14611), .ZN(
        P1_U3245) );
  INV_X1 U16439 ( .A(n14621), .ZN(n14616) );
  OAI22_X1 U16440 ( .A1(n15226), .A2(n6881), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11507), .ZN(n14615) );
  AOI21_X1 U16441 ( .B1(n14654), .B2(n14616), .A(n14615), .ZN(n14628) );
  MUX2_X1 U16442 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10162), .S(n14621), .Z(
        n14617) );
  NAND3_X1 U16443 ( .A1(n14619), .A2(n14618), .A3(n14617), .ZN(n14620) );
  NAND3_X1 U16444 ( .A1(n15210), .A2(n15207), .A3(n14620), .ZN(n14627) );
  MUX2_X1 U16445 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11510), .S(n14621), .Z(
        n14622) );
  NAND3_X1 U16446 ( .A1(n14624), .A2(n14623), .A3(n14622), .ZN(n14625) );
  NAND3_X1 U16447 ( .A1(n15217), .A2(n15214), .A3(n14625), .ZN(n14626) );
  NAND3_X1 U16448 ( .A1(n14628), .A2(n14627), .A3(n14626), .ZN(P1_U3246) );
  NAND2_X1 U16449 ( .A1(n14636), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14631) );
  INV_X1 U16450 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14629) );
  MUX2_X1 U16451 ( .A(n14629), .B(P1_REG2_REG_17__SCAN_IN), .S(n14644), .Z(
        n14630) );
  INV_X1 U16452 ( .A(n14643), .ZN(n14634) );
  NAND3_X1 U16453 ( .A1(n14632), .A2(n14631), .A3(n14630), .ZN(n14633) );
  NAND3_X1 U16454 ( .A1(n14634), .A2(n15217), .A3(n14633), .ZN(n14642) );
  AOI21_X1 U16455 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n14636), .A(n14635), 
        .ZN(n14648) );
  XNOR2_X1 U16456 ( .A(n14644), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14647) );
  XOR2_X1 U16457 ( .A(n14648), .B(n14647), .Z(n14637) );
  NAND2_X1 U16458 ( .A1(n15210), .A2(n14637), .ZN(n14638) );
  NAND2_X1 U16459 ( .A1(n14639), .A2(n14638), .ZN(n14640) );
  AOI21_X1 U16460 ( .B1(n14653), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14640), 
        .ZN(n14641) );
  OAI211_X1 U16461 ( .C1(n15221), .C2(n14645), .A(n14642), .B(n14641), .ZN(
        P1_U3260) );
  XNOR2_X1 U16462 ( .A(n14662), .B(n14664), .ZN(n14665) );
  XNOR2_X1 U16463 ( .A(n14665), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14658) );
  INV_X1 U16464 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14646) );
  XOR2_X1 U16465 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14659), .Z(n14649) );
  NAND2_X1 U16466 ( .A1(n15210), .A2(n14649), .ZN(n14650) );
  NAND2_X1 U16467 ( .A1(n14651), .A2(n14650), .ZN(n14652) );
  AOI21_X1 U16468 ( .B1(n14653), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14652), 
        .ZN(n14656) );
  NAND2_X1 U16469 ( .A1(n14654), .A2(n14664), .ZN(n14655) );
  OAI211_X1 U16470 ( .C1(n14658), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        P1_U3261) );
  AOI22_X1 U16471 ( .A1(n14660), .A2(n14664), .B1(P1_REG1_REG_18__SCAN_IN), 
        .B2(n14659), .ZN(n14661) );
  XNOR2_X1 U16472 ( .A(n14661), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14669) );
  INV_X1 U16473 ( .A(n14662), .ZN(n14663) );
  AOI22_X1 U16474 ( .A1(n14665), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14664), 
        .B2(n14663), .ZN(n14666) );
  AOI22_X1 U16475 ( .A1(n14669), .A2(n15210), .B1(n14667), .B2(n15217), .ZN(
        n14673) );
  OAI21_X1 U16476 ( .B1(n14669), .B2(n14668), .A(n15221), .ZN(n14670) );
  INV_X1 U16477 ( .A(n14674), .ZN(n14675) );
  OAI211_X1 U16478 ( .C1(n7901), .C2(n15226), .A(n14676), .B(n14675), .ZN(
        P1_U3262) );
  NAND2_X1 U16479 ( .A1(n14685), .A2(n14983), .ZN(n14684) );
  XOR2_X1 U16480 ( .A(n14681), .B(n14684), .Z(n14677) );
  INV_X1 U16481 ( .A(n14678), .ZN(n14679) );
  OR2_X1 U16482 ( .A1(n14680), .A2(n14679), .ZN(n14981) );
  NOR2_X1 U16483 ( .A1(n15260), .A2(n14981), .ZN(n14687) );
  INV_X1 U16484 ( .A(n14681), .ZN(n14980) );
  NOR2_X1 U16485 ( .A1(n14980), .A2(n15262), .ZN(n14682) );
  AOI211_X1 U16486 ( .C1(n15260), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14687), 
        .B(n14682), .ZN(n14683) );
  OAI21_X1 U16487 ( .B1(n14979), .B2(n14974), .A(n14683), .ZN(P1_U3263) );
  OAI211_X1 U16488 ( .C1(n14685), .C2(n14983), .A(n15240), .B(n14684), .ZN(
        n14982) );
  NOR2_X1 U16489 ( .A1(n14798), .A2(n14686), .ZN(n14688) );
  AOI211_X1 U16490 ( .C1(n14689), .C2(n14971), .A(n14688), .B(n14687), .ZN(
        n14690) );
  OAI21_X1 U16491 ( .B1(n14982), .B2(n14974), .A(n14690), .ZN(P1_U3264) );
  NAND2_X1 U16492 ( .A1(n14692), .A2(n14879), .ZN(n14706) );
  INV_X1 U16493 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n14695) );
  OAI22_X1 U16494 ( .A1(n14798), .A2(n14695), .B1(n14694), .B2(n14693), .ZN(
        n14699) );
  NOR2_X1 U16495 ( .A1(n14697), .A2(n14696), .ZN(n14698) );
  AOI211_X1 U16496 ( .C1(n15258), .C2(n14700), .A(n14699), .B(n14698), .ZN(
        n14701) );
  OAI21_X1 U16497 ( .B1(n14702), .B2(n15262), .A(n14701), .ZN(n14703) );
  AOI21_X1 U16498 ( .B1(n14704), .B2(n15266), .A(n14703), .ZN(n14705) );
  OAI211_X1 U16499 ( .C1(n14707), .C2(n14978), .A(n14706), .B(n14705), .ZN(
        P1_U3356) );
  AOI22_X1 U16500 ( .A1(n14708), .A2(n15258), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15269), .ZN(n14709) );
  OAI21_X1 U16501 ( .B1(n14710), .B2(n15262), .A(n14709), .ZN(n14714) );
  NOR3_X1 U16502 ( .A1(n14712), .A2(n14711), .A3(n14978), .ZN(n14713) );
  XNOR2_X1 U16503 ( .A(n14719), .B(n14718), .ZN(n14720) );
  NAND2_X1 U16504 ( .A1(n14720), .A2(n15308), .ZN(n14722) );
  NAND2_X1 U16505 ( .A1(n14722), .A2(n14721), .ZN(n14989) );
  NAND2_X1 U16506 ( .A1(n14989), .A2(n14798), .ZN(n14730) );
  NAND2_X1 U16507 ( .A1(n14735), .A2(n14985), .ZN(n14723) );
  NAND2_X1 U16508 ( .A1(n14723), .A2(n15240), .ZN(n14724) );
  NOR2_X1 U16509 ( .A1(n14725), .A2(n14724), .ZN(n14984) );
  AOI22_X1 U16510 ( .A1(n14726), .A2(n15258), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15260), .ZN(n14727) );
  OAI21_X1 U16511 ( .B1(n7451), .B2(n15262), .A(n14727), .ZN(n14728) );
  AOI21_X1 U16512 ( .B1(n14984), .B2(n15266), .A(n14728), .ZN(n14729) );
  OAI211_X1 U16513 ( .C1(n14991), .C2(n14978), .A(n14730), .B(n14729), .ZN(
        P1_U3266) );
  NAND2_X1 U16514 ( .A1(n14992), .A2(n14798), .ZN(n14743) );
  INV_X1 U16515 ( .A(n14735), .ZN(n14736) );
  AOI211_X1 U16516 ( .C1(n14994), .C2(n14748), .A(n10283), .B(n14736), .ZN(
        n14738) );
  OR2_X1 U16517 ( .A1(n14738), .A2(n14737), .ZN(n14993) );
  AOI22_X1 U16518 ( .A1(n14739), .A2(n15258), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15260), .ZN(n14740) );
  OAI21_X1 U16519 ( .B1(n7452), .B2(n15262), .A(n14740), .ZN(n14741) );
  AOI21_X1 U16520 ( .B1(n14993), .B2(n15266), .A(n14741), .ZN(n14742) );
  OAI211_X1 U16521 ( .C1(n14995), .C2(n14978), .A(n14743), .B(n14742), .ZN(
        P1_U3267) );
  AOI21_X1 U16522 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(n15002) );
  INV_X1 U16523 ( .A(n14747), .ZN(n14750) );
  INV_X1 U16524 ( .A(n14748), .ZN(n14749) );
  AOI211_X1 U16525 ( .C1(n14998), .C2(n14750), .A(n10283), .B(n14749), .ZN(
        n14996) );
  NAND2_X1 U16526 ( .A1(n14996), .A2(n14934), .ZN(n14752) );
  INV_X1 U16527 ( .A(n14997), .ZN(n14751) );
  OAI211_X1 U16528 ( .C1(n15236), .C2(n14753), .A(n14752), .B(n14751), .ZN(
        n14757) );
  INV_X1 U16529 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14754) );
  OAI22_X1 U16530 ( .A1(n14755), .A2(n15262), .B1(n14754), .B2(n14798), .ZN(
        n14756) );
  AOI21_X1 U16531 ( .B1(n14757), .B2(n14798), .A(n14756), .ZN(n14762) );
  NAND2_X1 U16532 ( .A1(n14760), .A2(n14759), .ZN(n14999) );
  NAND3_X1 U16533 ( .A1(n14758), .A2(n14999), .A3(n14903), .ZN(n14761) );
  OAI211_X1 U16534 ( .C1(n15002), .C2(n14906), .A(n14762), .B(n14761), .ZN(
        P1_U3268) );
  NAND2_X1 U16535 ( .A1(n14763), .A2(n14771), .ZN(n14764) );
  NAND2_X1 U16536 ( .A1(n14765), .A2(n14764), .ZN(n15012) );
  AOI21_X1 U16537 ( .B1(n14766), .B2(n14768), .A(n14767), .ZN(n14792) );
  INV_X1 U16538 ( .A(n14769), .ZN(n14770) );
  OR2_X1 U16539 ( .A1(n14792), .A2(n14770), .ZN(n14772) );
  XNOR2_X1 U16540 ( .A(n14772), .B(n14771), .ZN(n14773) );
  NAND2_X1 U16541 ( .A1(n14773), .A2(n15308), .ZN(n14775) );
  NAND2_X1 U16542 ( .A1(n14775), .A2(n14774), .ZN(n15014) );
  NAND2_X1 U16543 ( .A1(n15014), .A2(n14798), .ZN(n14784) );
  OAI21_X1 U16544 ( .B1(n14799), .B2(n14780), .A(n15240), .ZN(n14776) );
  OR2_X1 U16545 ( .A1(n14777), .A2(n14776), .ZN(n15011) );
  INV_X1 U16546 ( .A(n15011), .ZN(n14782) );
  AOI22_X1 U16547 ( .A1(n14778), .A2(n15258), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15260), .ZN(n14779) );
  OAI21_X1 U16548 ( .B1(n14780), .B2(n15262), .A(n14779), .ZN(n14781) );
  AOI21_X1 U16549 ( .B1(n14782), .B2(n15266), .A(n14781), .ZN(n14783) );
  OAI211_X1 U16550 ( .C1(n15012), .C2(n14978), .A(n14784), .B(n14783), .ZN(
        P1_U3270) );
  NOR2_X1 U16551 ( .A1(n14785), .A2(n14815), .ZN(n14817) );
  NOR2_X1 U16552 ( .A1(n14817), .A2(n14786), .ZN(n14787) );
  XOR2_X1 U16553 ( .A(n14791), .B(n14787), .Z(n15018) );
  INV_X1 U16554 ( .A(n14827), .ZN(n14788) );
  NAND2_X1 U16555 ( .A1(n15025), .A2(n14789), .ZN(n14811) );
  OAI21_X1 U16556 ( .B1(n15027), .B2(n14790), .A(n14810), .ZN(n14794) );
  INV_X1 U16557 ( .A(n14791), .ZN(n14793) );
  INV_X1 U16558 ( .A(n14795), .ZN(n14796) );
  OAI21_X1 U16559 ( .B1(n14797), .B2(n15277), .A(n14796), .ZN(n15015) );
  NAND2_X1 U16560 ( .A1(n15015), .A2(n14798), .ZN(n14807) );
  AOI211_X1 U16561 ( .C1(n15017), .C2(n14800), .A(n10283), .B(n14799), .ZN(
        n15016) );
  INV_X1 U16562 ( .A(n14801), .ZN(n14802) );
  AOI22_X1 U16563 ( .A1(n14802), .A2(n15258), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15260), .ZN(n14803) );
  OAI21_X1 U16564 ( .B1(n14804), .B2(n15262), .A(n14803), .ZN(n14805) );
  AOI21_X1 U16565 ( .B1(n15016), .B2(n15266), .A(n14805), .ZN(n14806) );
  OAI211_X1 U16566 ( .C1(n15018), .C2(n14978), .A(n14807), .B(n14806), .ZN(
        P1_U3271) );
  XNOR2_X1 U16567 ( .A(n7442), .B(n15021), .ZN(n14809) );
  NAND2_X1 U16568 ( .A1(n14809), .A2(n15240), .ZN(n15020) );
  INV_X1 U16569 ( .A(n15020), .ZN(n14814) );
  OAI211_X1 U16570 ( .C1(n14811), .C2(n14815), .A(n14810), .B(n15308), .ZN(
        n14813) );
  NAND2_X1 U16571 ( .A1(n14813), .A2(n14812), .ZN(n15024) );
  AOI21_X1 U16572 ( .B1(n14814), .B2(n14934), .A(n15024), .ZN(n14823) );
  AND2_X1 U16573 ( .A1(n14785), .A2(n14815), .ZN(n14816) );
  OR2_X1 U16574 ( .A1(n14817), .A2(n14816), .ZN(n15019) );
  INV_X1 U16575 ( .A(n14818), .ZN(n14819) );
  AOI22_X1 U16576 ( .A1(n14819), .A2(n15258), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15260), .ZN(n14820) );
  OAI21_X1 U16577 ( .B1(n15021), .B2(n15262), .A(n14820), .ZN(n14821) );
  AOI21_X1 U16578 ( .B1(n15019), .B2(n14903), .A(n14821), .ZN(n14822) );
  OAI21_X1 U16579 ( .B1(n14823), .B2(n15269), .A(n14822), .ZN(P1_U3272) );
  OAI21_X1 U16580 ( .B1(n14824), .B2(n14827), .A(n14825), .ZN(n15033) );
  INV_X1 U16581 ( .A(n14766), .ZN(n14828) );
  NAND2_X1 U16582 ( .A1(n14828), .A2(n14827), .ZN(n15026) );
  NAND3_X1 U16583 ( .A1(n15026), .A2(n14879), .A3(n15025), .ZN(n14838) );
  AOI211_X1 U16584 ( .C1(n15030), .C2(n14829), .A(n10283), .B(n14808), .ZN(
        n15028) );
  AOI22_X1 U16585 ( .A1(n14830), .A2(n15258), .B1(n15269), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14831) );
  OAI21_X1 U16586 ( .B1(n15027), .B2(n14969), .A(n14831), .ZN(n14832) );
  AOI21_X1 U16587 ( .B1(n14964), .B2(n14833), .A(n14832), .ZN(n14834) );
  OAI21_X1 U16588 ( .B1(n14835), .B2(n15262), .A(n14834), .ZN(n14836) );
  AOI21_X1 U16589 ( .B1(n15028), .B2(n15266), .A(n14836), .ZN(n14837) );
  OAI211_X1 U16590 ( .C1(n15033), .C2(n14978), .A(n14838), .B(n14837), .ZN(
        P1_U3273) );
  XOR2_X1 U16591 ( .A(n14399), .B(n14839), .Z(n15042) );
  INV_X1 U16592 ( .A(n14840), .ZN(n14844) );
  INV_X1 U16593 ( .A(n14399), .ZN(n14843) );
  OAI21_X1 U16594 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n15040) );
  OAI211_X1 U16595 ( .C1(n14856), .C2(n15038), .A(n15240), .B(n14829), .ZN(
        n15037) );
  NAND2_X1 U16596 ( .A1(n14964), .A2(n15034), .ZN(n14847) );
  AOI22_X1 U16597 ( .A1(n15269), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14845), 
        .B2(n15258), .ZN(n14846) );
  OAI211_X1 U16598 ( .C1(n14848), .C2(n14969), .A(n14847), .B(n14846), .ZN(
        n14849) );
  AOI21_X1 U16599 ( .B1(n14850), .B2(n14971), .A(n14849), .ZN(n14851) );
  OAI21_X1 U16600 ( .B1(n15037), .B2(n14974), .A(n14851), .ZN(n14852) );
  AOI21_X1 U16601 ( .B1(n15040), .B2(n14879), .A(n14852), .ZN(n14853) );
  OAI21_X1 U16602 ( .B1(n14978), .B2(n15042), .A(n14853), .ZN(P1_U3274) );
  XOR2_X1 U16603 ( .A(n14854), .B(n14865), .Z(n15046) );
  OAI21_X1 U16604 ( .B1(n14880), .B2(n14855), .A(n15240), .ZN(n14857) );
  OR2_X1 U16605 ( .A1(n14857), .A2(n14856), .ZN(n15047) );
  NAND2_X1 U16606 ( .A1(n14964), .A2(n14858), .ZN(n14862) );
  NOR2_X1 U16607 ( .A1(n14859), .A2(n15236), .ZN(n14860) );
  AOI21_X1 U16608 ( .B1(n15269), .B2(P1_REG2_REG_18__SCAN_IN), .A(n14860), 
        .ZN(n14861) );
  OAI211_X1 U16609 ( .C1(n15043), .C2(n14969), .A(n14862), .B(n14861), .ZN(
        n14863) );
  AOI21_X1 U16610 ( .B1(n15045), .B2(n14971), .A(n14863), .ZN(n14864) );
  OAI21_X1 U16611 ( .B1(n15047), .B2(n14974), .A(n14864), .ZN(n14869) );
  OAI211_X1 U16612 ( .C1(n14867), .C2(n9050), .A(n14866), .B(n15308), .ZN(
        n15050) );
  NOR2_X1 U16613 ( .A1(n15050), .A2(n15260), .ZN(n14868) );
  AOI211_X1 U16614 ( .C1(n15046), .C2(n14903), .A(n14869), .B(n14868), .ZN(
        n14870) );
  INV_X1 U16615 ( .A(n14870), .ZN(P1_U3275) );
  XOR2_X1 U16616 ( .A(n14871), .B(n14877), .Z(n15060) );
  NAND2_X1 U16617 ( .A1(n14910), .A2(n14872), .ZN(n14891) );
  NOR2_X1 U16618 ( .A1(n14891), .A2(n14902), .ZN(n14890) );
  INV_X1 U16619 ( .A(n14873), .ZN(n14874) );
  NOR2_X1 U16620 ( .A1(n14890), .A2(n14874), .ZN(n14876) );
  INV_X1 U16621 ( .A(n14877), .ZN(n14875) );
  NAND2_X1 U16622 ( .A1(n14876), .A2(n14875), .ZN(n15052) );
  INV_X1 U16623 ( .A(n14876), .ZN(n14878) );
  NAND2_X1 U16624 ( .A1(n14878), .A2(n14877), .ZN(n15051) );
  NAND3_X1 U16625 ( .A1(n15052), .A2(n14879), .A3(n15051), .ZN(n14889) );
  AOI211_X1 U16626 ( .C1(n15057), .C2(n14892), .A(n10283), .B(n14880), .ZN(
        n15055) );
  AOI22_X1 U16627 ( .A1(n15269), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14881), 
        .B2(n15258), .ZN(n14882) );
  OAI21_X1 U16628 ( .B1(n14969), .B2(n15054), .A(n14882), .ZN(n14883) );
  AOI21_X1 U16629 ( .B1(n14964), .B2(n14884), .A(n14883), .ZN(n14885) );
  OAI21_X1 U16630 ( .B1(n14886), .B2(n15262), .A(n14885), .ZN(n14887) );
  AOI21_X1 U16631 ( .B1(n15055), .B2(n15266), .A(n14887), .ZN(n14888) );
  OAI211_X1 U16632 ( .C1(n15060), .C2(n14978), .A(n14889), .B(n14888), .ZN(
        P1_U3276) );
  AOI21_X1 U16633 ( .B1(n14902), .B2(n14891), .A(n14890), .ZN(n15068) );
  INV_X1 U16634 ( .A(n14892), .ZN(n14893) );
  AOI211_X1 U16635 ( .C1(n15064), .C2(n14916), .A(n10283), .B(n14893), .ZN(
        n15062) );
  NAND2_X1 U16636 ( .A1(n15064), .A2(n14971), .ZN(n14899) );
  OAI22_X1 U16637 ( .A1(n14798), .A2(n14895), .B1(n14894), .B2(n15236), .ZN(
        n14896) );
  AOI21_X1 U16638 ( .B1(n14964), .B2(n14897), .A(n14896), .ZN(n14898) );
  OAI211_X1 U16639 ( .C1(n15061), .C2(n14969), .A(n14899), .B(n14898), .ZN(
        n14900) );
  AOI21_X1 U16640 ( .B1(n15062), .B2(n15266), .A(n14900), .ZN(n14905) );
  XNOR2_X1 U16641 ( .A(n14901), .B(n14902), .ZN(n15065) );
  NAND2_X1 U16642 ( .A1(n15065), .A2(n14903), .ZN(n14904) );
  OAI211_X1 U16643 ( .C1(n15068), .C2(n14906), .A(n14905), .B(n14904), .ZN(
        P1_U3277) );
  NOR2_X1 U16644 ( .A1(n14907), .A2(n14930), .ZN(n14925) );
  NOR2_X1 U16645 ( .A1(n14925), .A2(n14908), .ZN(n14909) );
  XNOR2_X1 U16646 ( .A(n14912), .B(n14909), .ZN(n15073) );
  OAI211_X1 U16647 ( .C1(n14912), .C2(n14911), .A(n14910), .B(n15308), .ZN(
        n14914) );
  NAND2_X1 U16648 ( .A1(n14914), .A2(n14913), .ZN(n15069) );
  NAND2_X1 U16649 ( .A1(n15069), .A2(n14798), .ZN(n14924) );
  INV_X1 U16650 ( .A(n14915), .ZN(n14918) );
  INV_X1 U16651 ( .A(n14916), .ZN(n14917) );
  AOI211_X1 U16652 ( .C1(n15071), .C2(n14918), .A(n10283), .B(n14917), .ZN(
        n15070) );
  AOI22_X1 U16653 ( .A1(n15260), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14919), 
        .B2(n15258), .ZN(n14920) );
  OAI21_X1 U16654 ( .B1(n14921), .B2(n15262), .A(n14920), .ZN(n14922) );
  AOI21_X1 U16655 ( .B1(n15070), .B2(n15266), .A(n14922), .ZN(n14923) );
  OAI211_X1 U16656 ( .C1(n15073), .C2(n14978), .A(n14924), .B(n14923), .ZN(
        P1_U3278) );
  INV_X1 U16657 ( .A(n14907), .ZN(n14928) );
  INV_X1 U16658 ( .A(n14925), .ZN(n14926) );
  OAI21_X1 U16659 ( .B1(n14928), .B2(n14927), .A(n14926), .ZN(n15081) );
  OAI211_X1 U16660 ( .C1(n14931), .C2(n14930), .A(n14929), .B(n15308), .ZN(
        n15080) );
  OAI21_X1 U16661 ( .B1(n14954), .B2(n14932), .A(n15240), .ZN(n14933) );
  NOR2_X1 U16662 ( .A1(n14933), .A2(n14915), .ZN(n15076) );
  NAND2_X1 U16663 ( .A1(n15076), .A2(n14934), .ZN(n14935) );
  OAI211_X1 U16664 ( .C1(n15236), .C2(n14936), .A(n15080), .B(n14935), .ZN(
        n14937) );
  NAND2_X1 U16665 ( .A1(n14937), .A2(n14798), .ZN(n14941) );
  AOI22_X1 U16666 ( .A1(n14964), .A2(n15091), .B1(n15260), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n14938) );
  OAI21_X1 U16667 ( .B1(n15074), .B2(n14969), .A(n14938), .ZN(n14939) );
  AOI21_X1 U16668 ( .B1(n15078), .B2(n14971), .A(n14939), .ZN(n14940) );
  OAI211_X1 U16669 ( .C1(n15081), .C2(n14978), .A(n14941), .B(n14940), .ZN(
        P1_U3279) );
  XNOR2_X1 U16670 ( .A(n14942), .B(n14944), .ZN(n15089) );
  OAI211_X1 U16671 ( .C1(n14945), .C2(n14944), .A(n15308), .B(n14943), .ZN(
        n15088) );
  NAND2_X1 U16672 ( .A1(n14964), .A2(n14946), .ZN(n14950) );
  NOR2_X1 U16673 ( .A1(n15236), .A2(n14947), .ZN(n14948) );
  AOI21_X1 U16674 ( .B1(n15260), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14948), 
        .ZN(n14949) );
  OAI211_X1 U16675 ( .C1(n15082), .C2(n14969), .A(n14950), .B(n14949), .ZN(
        n14951) );
  AOI21_X1 U16676 ( .B1(n15086), .B2(n14971), .A(n14951), .ZN(n14956) );
  NAND2_X1 U16677 ( .A1(n14962), .A2(n15086), .ZN(n14952) );
  NAND2_X1 U16678 ( .A1(n14952), .A2(n15240), .ZN(n14953) );
  NOR2_X1 U16679 ( .A1(n14954), .A2(n14953), .ZN(n15084) );
  NAND2_X1 U16680 ( .A1(n15084), .A2(n15266), .ZN(n14955) );
  OAI211_X1 U16681 ( .C1(n15088), .C2(n15260), .A(n14956), .B(n14955), .ZN(
        n14957) );
  INV_X1 U16682 ( .A(n14957), .ZN(n14958) );
  OAI21_X1 U16683 ( .B1(n14978), .B2(n15089), .A(n14958), .ZN(P1_U3280) );
  XNOR2_X1 U16684 ( .A(n14959), .B(n14961), .ZN(n15099) );
  INV_X1 U16685 ( .A(n15098), .ZN(n14976) );
  AOI21_X1 U16686 ( .B1(n12032), .B2(n14972), .A(n10283), .ZN(n14963) );
  NAND2_X1 U16687 ( .A1(n14963), .A2(n14962), .ZN(n15094) );
  NAND2_X1 U16688 ( .A1(n14964), .A2(n15092), .ZN(n14968) );
  NOR2_X1 U16689 ( .A1(n15236), .A2(n14965), .ZN(n14966) );
  AOI21_X1 U16690 ( .B1(n15269), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14966), 
        .ZN(n14967) );
  OAI211_X1 U16691 ( .C1(n15075), .C2(n14969), .A(n14968), .B(n14967), .ZN(
        n14970) );
  AOI21_X1 U16692 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(n14973) );
  OAI21_X1 U16693 ( .B1(n15094), .B2(n14974), .A(n14973), .ZN(n14975) );
  AOI21_X1 U16694 ( .B1(n14976), .B2(n14798), .A(n14975), .ZN(n14977) );
  OAI21_X1 U16695 ( .B1(n14978), .B2(n15099), .A(n14977), .ZN(P1_U3281) );
  OAI211_X1 U16696 ( .C1(n14980), .C2(n15302), .A(n14979), .B(n14981), .ZN(
        n15114) );
  MUX2_X1 U16697 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15114), .S(n15327), .Z(
        P1_U3559) );
  OAI211_X1 U16698 ( .C1(n14983), .C2(n15302), .A(n14982), .B(n14981), .ZN(
        n15115) );
  MUX2_X1 U16699 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15115), .S(n15327), .Z(
        P1_U3558) );
  MUX2_X1 U16700 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15116), .S(n15327), .Z(
        P1_U3555) );
  MUX2_X1 U16701 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15117), .S(n15327), .Z(
        P1_U3554) );
  AOI211_X1 U16702 ( .C1(n14998), .C2(n15315), .A(n14997), .B(n14996), .ZN(
        n15001) );
  NAND3_X1 U16703 ( .A1(n14758), .A2(n15321), .A3(n14999), .ZN(n15000) );
  OAI211_X1 U16704 ( .C1(n15002), .C2(n15277), .A(n15001), .B(n15000), .ZN(
        n15118) );
  MUX2_X1 U16705 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15118), .S(n15327), .Z(
        P1_U3553) );
  INV_X1 U16706 ( .A(n15003), .ZN(n15005) );
  OAI21_X1 U16707 ( .B1(n15289), .B2(n15008), .A(n15007), .ZN(n15119) );
  MUX2_X1 U16708 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15119), .S(n15327), .Z(
        P1_U3552) );
  NAND2_X1 U16709 ( .A1(n15009), .A2(n15315), .ZN(n15010) );
  OAI211_X1 U16710 ( .C1(n15012), .C2(n15289), .A(n15011), .B(n15010), .ZN(
        n15013) );
  MUX2_X1 U16711 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15120), .S(n15327), .Z(
        P1_U3551) );
  MUX2_X1 U16712 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15121), .S(n15327), .Z(
        P1_U3550) );
  AND2_X1 U16713 ( .A1(n15019), .A2(n15321), .ZN(n15023) );
  OAI21_X1 U16714 ( .B1(n15021), .B2(n15302), .A(n15020), .ZN(n15022) );
  MUX2_X1 U16715 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15122), .S(n15327), .Z(
        P1_U3549) );
  NAND3_X1 U16716 ( .A1(n15026), .A2(n15308), .A3(n15025), .ZN(n15032) );
  OAI22_X1 U16717 ( .A1(n15027), .A2(n15310), .B1(n15043), .B2(n15312), .ZN(
        n15029) );
  AOI211_X1 U16718 ( .C1(n15030), .C2(n15315), .A(n15029), .B(n15028), .ZN(
        n15031) );
  OAI211_X1 U16719 ( .C1(n15289), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        n15123) );
  MUX2_X1 U16720 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15123), .S(n15327), .Z(
        P1_U3548) );
  AOI22_X1 U16721 ( .A1(n15035), .A2(n15090), .B1(n15107), .B2(n15034), .ZN(
        n15036) );
  OAI211_X1 U16722 ( .C1(n15038), .C2(n15302), .A(n15037), .B(n15036), .ZN(
        n15039) );
  AOI21_X1 U16723 ( .B1(n15040), .B2(n15308), .A(n15039), .ZN(n15041) );
  OAI21_X1 U16724 ( .B1(n15289), .B2(n15042), .A(n15041), .ZN(n15124) );
  MUX2_X1 U16725 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15124), .S(n15327), .Z(
        P1_U3547) );
  OAI22_X1 U16726 ( .A1(n15043), .A2(n15310), .B1(n15061), .B2(n15312), .ZN(
        n15044) );
  AOI21_X1 U16727 ( .B1(n15045), .B2(n15315), .A(n15044), .ZN(n15049) );
  NAND2_X1 U16728 ( .A1(n15046), .A2(n15321), .ZN(n15048) );
  NAND4_X1 U16729 ( .A1(n15050), .A2(n15049), .A3(n15048), .A4(n15047), .ZN(
        n15125) );
  MUX2_X1 U16730 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15125), .S(n15327), .Z(
        P1_U3546) );
  NAND3_X1 U16731 ( .A1(n15052), .A2(n15308), .A3(n15051), .ZN(n15059) );
  OAI22_X1 U16732 ( .A1(n15054), .A2(n15310), .B1(n15053), .B2(n15312), .ZN(
        n15056) );
  AOI211_X1 U16733 ( .C1(n15057), .C2(n15315), .A(n15056), .B(n15055), .ZN(
        n15058) );
  OAI211_X1 U16734 ( .C1(n15289), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        n15126) );
  MUX2_X1 U16735 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15126), .S(n15327), .Z(
        P1_U3545) );
  OAI22_X1 U16736 ( .A1(n15061), .A2(n15310), .B1(n15074), .B2(n15312), .ZN(
        n15063) );
  AOI211_X1 U16737 ( .C1(n15064), .C2(n15315), .A(n15063), .B(n15062), .ZN(
        n15067) );
  NAND2_X1 U16738 ( .A1(n15065), .A2(n15321), .ZN(n15066) );
  OAI211_X1 U16739 ( .C1(n15068), .C2(n15277), .A(n15067), .B(n15066), .ZN(
        n15127) );
  MUX2_X1 U16740 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15127), .S(n15327), .Z(
        P1_U3544) );
  AOI211_X1 U16741 ( .C1(n15071), .C2(n15315), .A(n15070), .B(n15069), .ZN(
        n15072) );
  OAI21_X1 U16742 ( .B1(n15289), .B2(n15073), .A(n15072), .ZN(n15128) );
  MUX2_X1 U16743 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15128), .S(n15327), .Z(
        P1_U3543) );
  OAI22_X1 U16744 ( .A1(n15075), .A2(n15312), .B1(n15074), .B2(n15310), .ZN(
        n15077) );
  AOI211_X1 U16745 ( .C1(n15078), .C2(n15315), .A(n15077), .B(n15076), .ZN(
        n15079) );
  OAI211_X1 U16746 ( .C1(n15289), .C2(n15081), .A(n15080), .B(n15079), .ZN(
        n15129) );
  MUX2_X1 U16747 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15129), .S(n15327), .Z(
        P1_U3542) );
  OAI22_X1 U16748 ( .A1(n15083), .A2(n15312), .B1(n15082), .B2(n15310), .ZN(
        n15085) );
  AOI211_X1 U16749 ( .C1(n15086), .C2(n15315), .A(n15085), .B(n15084), .ZN(
        n15087) );
  OAI211_X1 U16750 ( .C1(n15289), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15130) );
  MUX2_X1 U16751 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15130), .S(n15327), .Z(
        P1_U3541) );
  AOI22_X1 U16752 ( .A1(n15107), .A2(n15092), .B1(n15091), .B2(n15090), .ZN(
        n15093) );
  OAI211_X1 U16753 ( .C1(n15095), .C2(n15302), .A(n15094), .B(n15093), .ZN(
        n15096) );
  INV_X1 U16754 ( .A(n15096), .ZN(n15097) );
  OAI211_X1 U16755 ( .C1(n15289), .C2(n15099), .A(n15098), .B(n15097), .ZN(
        n15131) );
  MUX2_X1 U16756 ( .A(n15131), .B(P1_REG1_REG_12__SCAN_IN), .S(n15331), .Z(
        P1_U3540) );
  AOI211_X1 U16757 ( .C1(n7165), .C2(n15315), .A(n15101), .B(n15100), .ZN(
        n15103) );
  OAI21_X1 U16758 ( .B1(n15289), .B2(n15104), .A(n15103), .ZN(n15132) );
  MUX2_X1 U16759 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15132), .S(n15327), .Z(
        P1_U3539) );
  NAND3_X1 U16760 ( .A1(n15105), .A2(n15308), .A3(n11759), .ZN(n15113) );
  AOI22_X1 U16761 ( .A1(n15108), .A2(n15315), .B1(n15107), .B2(n15106), .ZN(
        n15111) );
  NAND2_X1 U16762 ( .A1(n15109), .A2(n15321), .ZN(n15110) );
  NAND4_X1 U16763 ( .A1(n15113), .A2(n15112), .A3(n15111), .A4(n15110), .ZN(
        n15133) );
  MUX2_X1 U16764 ( .A(n15133), .B(P1_REG1_REG_10__SCAN_IN), .S(n15331), .Z(
        P1_U3538) );
  MUX2_X1 U16765 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15114), .S(n6403), .Z(
        P1_U3527) );
  MUX2_X1 U16766 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15115), .S(n6403), .Z(
        P1_U3526) );
  MUX2_X1 U16767 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15116), .S(n6403), .Z(
        P1_U3523) );
  MUX2_X1 U16768 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15118), .S(n6403), .Z(
        P1_U3521) );
  MUX2_X1 U16769 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15119), .S(n6403), .Z(
        P1_U3520) );
  MUX2_X1 U16770 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15120), .S(n6403), .Z(
        P1_U3519) );
  MUX2_X1 U16771 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15122), .S(n6403), .Z(
        P1_U3517) );
  MUX2_X1 U16772 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15123), .S(n6403), .Z(
        P1_U3516) );
  MUX2_X1 U16773 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15124), .S(n6403), .Z(
        P1_U3515) );
  MUX2_X1 U16774 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15125), .S(n6403), .Z(
        P1_U3513) );
  MUX2_X1 U16775 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15126), .S(n6403), .Z(
        P1_U3510) );
  MUX2_X1 U16776 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15127), .S(n6403), .Z(
        P1_U3507) );
  MUX2_X1 U16777 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15128), .S(n6403), .Z(
        P1_U3504) );
  MUX2_X1 U16778 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15129), .S(n6403), .Z(
        P1_U3501) );
  MUX2_X1 U16779 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15130), .S(n6403), .Z(
        P1_U3498) );
  MUX2_X1 U16780 ( .A(n15131), .B(P1_REG0_REG_12__SCAN_IN), .S(n15323), .Z(
        P1_U3495) );
  MUX2_X1 U16781 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15132), .S(n6403), .Z(
        P1_U3492) );
  MUX2_X1 U16782 ( .A(n15133), .B(P1_REG0_REG_10__SCAN_IN), .S(n15323), .Z(
        P1_U3489) );
  NAND3_X1 U16783 ( .A1(n15135), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n15137) );
  OAI22_X1 U16784 ( .A1(n15134), .A2(n15137), .B1(n15136), .B2(n15144), .ZN(
        n15138) );
  AOI21_X1 U16785 ( .B1(n15140), .B2(n15139), .A(n15138), .ZN(n15141) );
  INV_X1 U16786 ( .A(n15141), .ZN(P1_U3324) );
  OAI222_X1 U16787 ( .A1(P1_U3086), .A2(n6410), .B1(n15144), .B2(n15143), .C1(
        n15147), .C2(n15142), .ZN(P1_U3328) );
  OAI222_X1 U16788 ( .A1(n15149), .A2(P1_U3086), .B1(n15147), .B2(n15146), 
        .C1(n15145), .C2(n15144), .ZN(P1_U3330) );
  MUX2_X1 U16789 ( .A(n15150), .B(n14304), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16790 ( .A(n15151), .ZN(n15152) );
  MUX2_X1 U16791 ( .A(n15152), .B(n7069), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  XOR2_X1 U16792 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15153), .Z(SUB_1596_U53) );
  XOR2_X1 U16793 ( .A(n15155), .B(n15154), .Z(SUB_1596_U56) );
  XNOR2_X1 U16794 ( .A(n15156), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(n15157) );
  XOR2_X1 U16795 ( .A(n15158), .B(n15157), .Z(SUB_1596_U54) );
  XNOR2_X1 U16796 ( .A(n15159), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(n15160) );
  XOR2_X1 U16797 ( .A(n15161), .B(n15160), .Z(SUB_1596_U69) );
  INV_X1 U16798 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15162) );
  NAND2_X1 U16799 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15551), .ZN(n15164) );
  XNOR2_X1 U16800 ( .A(n15169), .B(P3_ADDR_REG_16__SCAN_IN), .ZN(n15173) );
  XNOR2_X1 U16801 ( .A(n15173), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(n15167) );
  XNOR2_X1 U16802 ( .A(n15167), .B(n15175), .ZN(SUB_1596_U64) );
  NOR2_X1 U16803 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15168), .ZN(n15172) );
  NOR2_X1 U16804 ( .A1(n15170), .A2(n15169), .ZN(n15171) );
  XNOR2_X1 U16805 ( .A(n15179), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15181) );
  INV_X1 U16806 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15174) );
  OAI21_X1 U16807 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(n15177) );
  NAND2_X1 U16808 ( .A1(n15175), .A2(n15174), .ZN(n15176) );
  XNOR2_X1 U16809 ( .A(n15183), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U16810 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15180) );
  XNOR2_X1 U16811 ( .A(n15190), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(n15185) );
  INV_X1 U16812 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15186) );
  XNOR2_X1 U16813 ( .A(n15185), .B(n15186), .ZN(n15184) );
  INV_X1 U16814 ( .A(n15181), .ZN(n15182) );
  XNOR2_X1 U16815 ( .A(n15184), .B(n15188), .ZN(SUB_1596_U62) );
  NAND2_X1 U16816 ( .A1(n15185), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15189) );
  INV_X1 U16817 ( .A(n15185), .ZN(n15187) );
  INV_X1 U16818 ( .A(n15190), .ZN(n15193) );
  AOI22_X1 U16819 ( .A1(n15193), .A2(P1_ADDR_REG_18__SCAN_IN), .B1(n15192), 
        .B2(n15191), .ZN(n15196) );
  XNOR2_X1 U16820 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15194) );
  XNOR2_X1 U16821 ( .A(n15194), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15195) );
  XNOR2_X1 U16822 ( .A(n15196), .B(n15195), .ZN(n15197) );
  XNOR2_X1 U16823 ( .A(n15198), .B(n15197), .ZN(SUB_1596_U4) );
  AOI21_X1 U16824 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15199) );
  OAI21_X1 U16825 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15199), 
        .ZN(U28) );
  AOI21_X1 U16826 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15200) );
  OAI21_X1 U16827 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15200), 
        .ZN(U29) );
  XOR2_X1 U16828 ( .A(n15202), .B(n15201), .Z(n15203) );
  XNOR2_X1 U16829 ( .A(n15203), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  INV_X1 U16830 ( .A(n15204), .ZN(n15209) );
  NAND3_X1 U16831 ( .A1(n15207), .A2(n15206), .A3(n15205), .ZN(n15208) );
  NAND3_X1 U16832 ( .A1(n15210), .A2(n15209), .A3(n15208), .ZN(n15219) );
  INV_X1 U16833 ( .A(n15211), .ZN(n15216) );
  NAND3_X1 U16834 ( .A1(n15214), .A2(n15213), .A3(n15212), .ZN(n15215) );
  NAND3_X1 U16835 ( .A1(n15217), .A2(n15216), .A3(n15215), .ZN(n15218) );
  OAI211_X1 U16836 ( .C1(n15221), .C2(n15220), .A(n15219), .B(n15218), .ZN(
        n15222) );
  NOR2_X1 U16837 ( .A1(n15223), .A2(n15222), .ZN(n15225) );
  OAI211_X1 U16838 ( .C1(n15226), .C2(n9944), .A(n15225), .B(n15224), .ZN(
        P1_U3247) );
  XNOR2_X1 U16839 ( .A(n15228), .B(n15227), .ZN(n15234) );
  XNOR2_X1 U16840 ( .A(n15230), .B(n15229), .ZN(n15231) );
  NOR2_X1 U16841 ( .A1(n15231), .A2(n15289), .ZN(n15232) );
  AOI211_X1 U16842 ( .C1(n15234), .C2(n15308), .A(n15233), .B(n15232), .ZN(
        n15304) );
  NOR2_X1 U16843 ( .A1(n15236), .A2(n15235), .ZN(n15237) );
  AOI21_X1 U16844 ( .B1(n15260), .B2(P1_REG2_REG_7__SCAN_IN), .A(n15237), .ZN(
        n15238) );
  OAI21_X1 U16845 ( .B1(n15262), .B2(n15303), .A(n15238), .ZN(n15239) );
  INV_X1 U16846 ( .A(n15239), .ZN(n15244) );
  OAI211_X1 U16847 ( .C1(n15241), .C2(n15303), .A(n15240), .B(n11382), .ZN(
        n15301) );
  INV_X1 U16848 ( .A(n15301), .ZN(n15242) );
  NAND2_X1 U16849 ( .A1(n15242), .A2(n15266), .ZN(n15243) );
  OAI211_X1 U16850 ( .C1(n15269), .C2(n15304), .A(n15244), .B(n15243), .ZN(
        P1_U3286) );
  XNOR2_X1 U16851 ( .A(n15245), .B(n15252), .ZN(n15257) );
  INV_X1 U16852 ( .A(n15248), .ZN(n15251) );
  OAI21_X1 U16853 ( .B1(n15248), .B2(n15247), .A(n15246), .ZN(n15249) );
  OAI21_X1 U16854 ( .B1(n15251), .B2(n15250), .A(n15249), .ZN(n15253) );
  XNOR2_X1 U16855 ( .A(n15253), .B(n15252), .ZN(n15254) );
  NOR2_X1 U16856 ( .A1(n15254), .A2(n15289), .ZN(n15255) );
  AOI211_X1 U16857 ( .C1(n15308), .C2(n15257), .A(n15256), .B(n15255), .ZN(
        n15293) );
  AOI22_X1 U16858 ( .A1(n15260), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15259), 
        .B2(n15258), .ZN(n15261) );
  OAI21_X1 U16859 ( .B1(n15262), .B2(n6406), .A(n15261), .ZN(n15263) );
  INV_X1 U16860 ( .A(n15263), .ZN(n15268) );
  AOI211_X1 U16861 ( .C1(n6407), .C2(n15265), .A(n10283), .B(n15264), .ZN(
        n15291) );
  NAND2_X1 U16862 ( .A1(n15291), .A2(n15266), .ZN(n15267) );
  OAI211_X1 U16863 ( .C1(n15269), .C2(n15293), .A(n15268), .B(n15267), .ZN(
        P1_U3288) );
  AND2_X1 U16864 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15270), .ZN(P1_U3294) );
  AND2_X1 U16865 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15270), .ZN(P1_U3295) );
  AND2_X1 U16866 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15270), .ZN(P1_U3296) );
  AND2_X1 U16867 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15270), .ZN(P1_U3297) );
  AND2_X1 U16868 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15270), .ZN(P1_U3298) );
  AND2_X1 U16869 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15270), .ZN(P1_U3299) );
  AND2_X1 U16870 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15270), .ZN(P1_U3300) );
  AND2_X1 U16871 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15270), .ZN(P1_U3301) );
  AND2_X1 U16872 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15270), .ZN(P1_U3302) );
  AND2_X1 U16873 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15270), .ZN(P1_U3303) );
  AND2_X1 U16874 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15270), .ZN(P1_U3304) );
  AND2_X1 U16875 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15270), .ZN(P1_U3305) );
  AND2_X1 U16876 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15270), .ZN(P1_U3306) );
  AND2_X1 U16877 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15270), .ZN(P1_U3307) );
  AND2_X1 U16878 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15270), .ZN(P1_U3308) );
  AND2_X1 U16879 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15270), .ZN(P1_U3309) );
  AND2_X1 U16880 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15270), .ZN(P1_U3310) );
  AND2_X1 U16881 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15270), .ZN(P1_U3311) );
  AND2_X1 U16882 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15270), .ZN(P1_U3312) );
  AND2_X1 U16883 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15270), .ZN(P1_U3313) );
  AND2_X1 U16884 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15270), .ZN(P1_U3314) );
  AND2_X1 U16885 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15270), .ZN(P1_U3315) );
  AND2_X1 U16886 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15270), .ZN(P1_U3316) );
  AND2_X1 U16887 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15270), .ZN(P1_U3317) );
  AND2_X1 U16888 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15270), .ZN(P1_U3318) );
  AND2_X1 U16889 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15270), .ZN(P1_U3319) );
  AND2_X1 U16890 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15270), .ZN(P1_U3320) );
  AND2_X1 U16891 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15270), .ZN(P1_U3321) );
  AND2_X1 U16892 ( .A1(n15270), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3322) );
  AND2_X1 U16893 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15270), .ZN(P1_U3323) );
  INV_X1 U16894 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U16895 ( .A1(n6403), .A2(n15272), .B1(n15271), .B2(n15323), .ZN(
        P1_U3459) );
  OAI211_X1 U16896 ( .C1(n15275), .C2(n15302), .A(n15274), .B(n15273), .ZN(
        n15280) );
  OAI22_X1 U16897 ( .A1(n15278), .A2(n15289), .B1(n15277), .B2(n15276), .ZN(
        n15279) );
  NOR2_X1 U16898 ( .A1(n15280), .A2(n15279), .ZN(n15324) );
  AOI22_X1 U16899 ( .A1(n6403), .A2(n15324), .B1(n8760), .B2(n15323), .ZN(
        P1_U3468) );
  OAI22_X1 U16900 ( .A1(n15282), .A2(n15312), .B1(n15281), .B2(n15310), .ZN(
        n15284) );
  AOI211_X1 U16901 ( .C1(n15285), .C2(n15315), .A(n15284), .B(n15283), .ZN(
        n15287) );
  OAI211_X1 U16902 ( .C1(n15289), .C2(n15288), .A(n15287), .B(n15286), .ZN(
        n15290) );
  INV_X1 U16903 ( .A(n15290), .ZN(n15326) );
  AOI22_X1 U16904 ( .A1(n6403), .A2(n15326), .B1(n8776), .B2(n15323), .ZN(
        P1_U3471) );
  AOI21_X1 U16905 ( .B1(n6407), .B2(n15315), .A(n15291), .ZN(n15294) );
  INV_X1 U16906 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15295) );
  AOI22_X1 U16907 ( .A1(n6403), .A2(n7884), .B1(n15295), .B2(n15323), .ZN(
        P1_U3474) );
  INV_X1 U16908 ( .A(n15296), .ZN(n15297) );
  OAI21_X1 U16909 ( .B1(n15298), .B2(n15302), .A(n15297), .ZN(n15300) );
  NOR2_X1 U16910 ( .A1(n15300), .A2(n15299), .ZN(n15329) );
  AOI22_X1 U16911 ( .A1(n6403), .A2(n15329), .B1(n8819), .B2(n15323), .ZN(
        P1_U3477) );
  OAI21_X1 U16912 ( .B1(n15303), .B2(n15302), .A(n15301), .ZN(n15306) );
  INV_X1 U16913 ( .A(n15304), .ZN(n15305) );
  NOR2_X1 U16914 ( .A1(n15306), .A2(n15305), .ZN(n15330) );
  INV_X1 U16915 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15307) );
  AOI22_X1 U16916 ( .A1(n6403), .A2(n15330), .B1(n15307), .B2(n15323), .ZN(
        P1_U3480) );
  NAND3_X1 U16917 ( .A1(n11377), .A2(n15309), .A3(n15308), .ZN(n15319) );
  OAI22_X1 U16918 ( .A1(n15313), .A2(n15312), .B1(n15311), .B2(n15310), .ZN(
        n15314) );
  AOI21_X1 U16919 ( .B1(n15316), .B2(n15315), .A(n15314), .ZN(n15318) );
  NAND3_X1 U16920 ( .A1(n15319), .A2(n15318), .A3(n15317), .ZN(n15320) );
  AOI21_X1 U16921 ( .B1(n15322), .B2(n15321), .A(n15320), .ZN(n15333) );
  AOI22_X1 U16922 ( .A1(n6403), .A2(n15333), .B1(n8866), .B2(n15323), .ZN(
        P1_U3483) );
  AOI22_X1 U16923 ( .A1(n15327), .A2(n15324), .B1(n10162), .B2(n15331), .ZN(
        P1_U3531) );
  AOI22_X1 U16924 ( .A1(n15327), .A2(n15326), .B1(n15325), .B2(n15331), .ZN(
        P1_U3532) );
  AOI22_X1 U16925 ( .A1(n15327), .A2(n7884), .B1(n8798), .B2(n15331), .ZN(
        P1_U3533) );
  AOI22_X1 U16926 ( .A1(n15327), .A2(n15329), .B1(n15328), .B2(n15331), .ZN(
        P1_U3534) );
  AOI22_X1 U16927 ( .A1(n15327), .A2(n15330), .B1(n8846), .B2(n15331), .ZN(
        P1_U3535) );
  AOI22_X1 U16928 ( .A1(n15327), .A2(n15333), .B1(n15332), .B2(n15331), .ZN(
        P1_U3536) );
  NOR2_X1 U16929 ( .A1(n15334), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16930 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15339) );
  INV_X1 U16931 ( .A(n15335), .ZN(n15338) );
  OR2_X1 U16932 ( .A1(n15395), .A2(n15336), .ZN(n15337) );
  OAI211_X1 U16933 ( .C1(n15399), .C2(n15339), .A(n15338), .B(n15337), .ZN(
        n15340) );
  INV_X1 U16934 ( .A(n15340), .ZN(n15349) );
  OAI211_X1 U16935 ( .C1(n15343), .C2(n15342), .A(n15403), .B(n15341), .ZN(
        n15348) );
  OAI211_X1 U16936 ( .C1(n15346), .C2(n15345), .A(n15405), .B(n15344), .ZN(
        n15347) );
  NAND3_X1 U16937 ( .A1(n15349), .A2(n15348), .A3(n15347), .ZN(P2_U3218) );
  INV_X1 U16938 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15354) );
  INV_X1 U16939 ( .A(n15350), .ZN(n15353) );
  OR2_X1 U16940 ( .A1(n15395), .A2(n15351), .ZN(n15352) );
  OAI211_X1 U16941 ( .C1(n15399), .C2(n15354), .A(n15353), .B(n15352), .ZN(
        n15355) );
  INV_X1 U16942 ( .A(n15355), .ZN(n15364) );
  OAI211_X1 U16943 ( .C1(n15358), .C2(n15357), .A(n15405), .B(n15356), .ZN(
        n15363) );
  OAI211_X1 U16944 ( .C1(n15361), .C2(n15360), .A(n15403), .B(n15359), .ZN(
        n15362) );
  NAND3_X1 U16945 ( .A1(n15364), .A2(n15363), .A3(n15362), .ZN(P2_U3220) );
  OR2_X1 U16946 ( .A1(n15395), .A2(n15365), .ZN(n15366) );
  OAI211_X1 U16947 ( .C1(n15399), .C2(n15368), .A(n15367), .B(n15366), .ZN(
        n15369) );
  INV_X1 U16948 ( .A(n15369), .ZN(n15378) );
  OAI211_X1 U16949 ( .C1(n15372), .C2(n15371), .A(n15405), .B(n15370), .ZN(
        n15377) );
  XOR2_X1 U16950 ( .A(n15374), .B(n15373), .Z(n15375) );
  NAND2_X1 U16951 ( .A1(n15403), .A2(n15375), .ZN(n15376) );
  NAND3_X1 U16952 ( .A1(n15378), .A2(n15377), .A3(n15376), .ZN(P2_U3221) );
  NOR2_X1 U16953 ( .A1(n15380), .A2(n15379), .ZN(n15382) );
  OAI21_X1 U16954 ( .B1(n15382), .B2(n15381), .A(n15403), .ZN(n15389) );
  NAND2_X1 U16955 ( .A1(n15384), .A2(n15383), .ZN(n15385) );
  NAND2_X1 U16956 ( .A1(n15386), .A2(n15385), .ZN(n15387) );
  NAND2_X1 U16957 ( .A1(n15387), .A2(n15405), .ZN(n15388) );
  OAI211_X1 U16958 ( .C1(n15395), .C2(n15390), .A(n15389), .B(n15388), .ZN(
        n15391) );
  INV_X1 U16959 ( .A(n15391), .ZN(n15393) );
  OAI211_X1 U16960 ( .C1(n7095), .C2(n15399), .A(n15393), .B(n15392), .ZN(
        P2_U3223) );
  INV_X1 U16961 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15398) );
  OR2_X1 U16962 ( .A1(n15395), .A2(n15394), .ZN(n15396) );
  OAI211_X1 U16963 ( .C1(n15399), .C2(n15398), .A(n15397), .B(n15396), .ZN(
        n15400) );
  INV_X1 U16964 ( .A(n15400), .ZN(n15411) );
  XOR2_X1 U16965 ( .A(n15402), .B(n15401), .Z(n15404) );
  NAND2_X1 U16966 ( .A1(n15404), .A2(n15403), .ZN(n15410) );
  OAI211_X1 U16967 ( .C1(n15408), .C2(n15407), .A(n15406), .B(n15405), .ZN(
        n15409) );
  NAND3_X1 U16968 ( .A1(n15411), .A2(n15410), .A3(n15409), .ZN(P2_U3231) );
  INV_X1 U16969 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15592) );
  NOR2_X1 U16970 ( .A1(n15413), .A2(n15592), .ZN(P2_U3266) );
  AND2_X1 U16971 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15515), .ZN(P2_U3268) );
  AND2_X1 U16972 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15515), .ZN(P2_U3269) );
  AND2_X1 U16973 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15515), .ZN(P2_U3270) );
  AND2_X1 U16974 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15515), .ZN(P2_U3271) );
  AND2_X1 U16975 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15515), .ZN(P2_U3272) );
  AND2_X1 U16976 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15515), .ZN(P2_U3273) );
  AND2_X1 U16977 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15515), .ZN(P2_U3274) );
  AND2_X1 U16978 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15515), .ZN(P2_U3275) );
  AND2_X1 U16979 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15515), .ZN(P2_U3276) );
  AND2_X1 U16980 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15515), .ZN(P2_U3277) );
  AND2_X1 U16981 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15515), .ZN(P2_U3278) );
  INV_X1 U16982 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15562) );
  NOR2_X1 U16983 ( .A1(n15413), .A2(n15562), .ZN(P2_U3279) );
  AND2_X1 U16984 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15515), .ZN(P2_U3280) );
  AND2_X1 U16985 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15515), .ZN(P2_U3281) );
  AND2_X1 U16986 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15515), .ZN(P2_U3282) );
  AND2_X1 U16987 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15515), .ZN(P2_U3283) );
  AND2_X1 U16988 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15515), .ZN(P2_U3284) );
  AND2_X1 U16989 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15515), .ZN(P2_U3285) );
  AND2_X1 U16990 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15515), .ZN(P2_U3286) );
  AND2_X1 U16991 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15515), .ZN(P2_U3287) );
  AND2_X1 U16992 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15515), .ZN(P2_U3288) );
  AND2_X1 U16993 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15515), .ZN(P2_U3289) );
  AND2_X1 U16994 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15515), .ZN(P2_U3290) );
  AND2_X1 U16995 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15515), .ZN(P2_U3291) );
  AND2_X1 U16996 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15515), .ZN(P2_U3292) );
  AND2_X1 U16997 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15515), .ZN(P2_U3293) );
  AND2_X1 U16998 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15515), .ZN(P2_U3294) );
  AND2_X1 U16999 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15515), .ZN(P2_U3295) );
  AOI22_X1 U17000 ( .A1(n15416), .A2(n15415), .B1(n15414), .B2(n15419), .ZN(
        P2_U3416) );
  AOI21_X1 U17001 ( .B1(n15419), .B2(n15418), .A(n15417), .ZN(P2_U3417) );
  INV_X1 U17002 ( .A(n15423), .ZN(n15426) );
  OAI22_X1 U17003 ( .A1(n15423), .A2(n15422), .B1(n15421), .B2(n15420), .ZN(
        n15425) );
  AOI211_X1 U17004 ( .C1(n15445), .C2(n15426), .A(n15425), .B(n15424), .ZN(
        n15449) );
  AOI22_X1 U17005 ( .A1(n15448), .A2(n15449), .B1(n6895), .B2(n15446), .ZN(
        P2_U3430) );
  NAND2_X1 U17006 ( .A1(n15427), .A2(n15445), .ZN(n15429) );
  OAI211_X1 U17007 ( .C1(n7152), .C2(n15439), .A(n15429), .B(n15428), .ZN(
        n15430) );
  NOR2_X1 U17008 ( .A1(n15431), .A2(n15430), .ZN(n15450) );
  AOI22_X1 U17009 ( .A1(n15448), .A2(n15450), .B1(n9511), .B2(n15446), .ZN(
        P2_U3436) );
  OAI21_X1 U17010 ( .B1(n7686), .B2(n15439), .A(n15432), .ZN(n15435) );
  INV_X1 U17011 ( .A(n15433), .ZN(n15434) );
  AOI211_X1 U17012 ( .C1(n15445), .C2(n15436), .A(n15435), .B(n15434), .ZN(
        n15451) );
  INV_X1 U17013 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15437) );
  AOI22_X1 U17014 ( .A1(n15448), .A2(n15451), .B1(n15437), .B2(n15446), .ZN(
        P2_U3442) );
  OAI21_X1 U17015 ( .B1(n15440), .B2(n15439), .A(n15438), .ZN(n15443) );
  INV_X1 U17016 ( .A(n15441), .ZN(n15442) );
  AOI211_X1 U17017 ( .C1(n15445), .C2(n15444), .A(n15443), .B(n15442), .ZN(
        n15453) );
  INV_X1 U17018 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15447) );
  AOI22_X1 U17019 ( .A1(n15448), .A2(n15453), .B1(n15447), .B2(n15446), .ZN(
        P2_U3448) );
  AOI22_X1 U17020 ( .A1(n15454), .A2(n15449), .B1(n10142), .B2(n15452), .ZN(
        P2_U3499) );
  AOI22_X1 U17021 ( .A1(n15454), .A2(n15450), .B1(n10076), .B2(n15452), .ZN(
        P2_U3501) );
  AOI22_X1 U17022 ( .A1(n15454), .A2(n15451), .B1(n10081), .B2(n15452), .ZN(
        P2_U3503) );
  AOI22_X1 U17023 ( .A1(n15454), .A2(n15453), .B1(n10085), .B2(n15452), .ZN(
        P2_U3505) );
  NOR2_X1 U17024 ( .A1(P3_U3897), .A2(n15455), .ZN(P3_U3150) );
  OAI21_X1 U17025 ( .B1(n15457), .B2(n15464), .A(n15456), .ZN(n15500) );
  NOR2_X1 U17026 ( .A1(n15475), .A2(n15458), .ZN(n15499) );
  INV_X1 U17027 ( .A(n15499), .ZN(n15461) );
  OAI22_X1 U17028 ( .A1(n15462), .A2(n15461), .B1(n15460), .B2(n15459), .ZN(
        n15470) );
  XNOR2_X1 U17029 ( .A(n15463), .B(n15464), .ZN(n15465) );
  OAI222_X1 U17030 ( .A1(n15469), .A2(n15468), .B1(n15467), .B2(n15466), .C1(
        n15484), .C2(n15465), .ZN(n15498) );
  AOI211_X1 U17031 ( .C1(n15471), .C2(n15500), .A(n15470), .B(n15498), .ZN(
        n15473) );
  AOI22_X1 U17032 ( .A1(n15493), .A2(n15474), .B1(n15473), .B2(n15472), .ZN(
        P3_U3231) );
  NOR2_X1 U17033 ( .A1(n15476), .A2(n15475), .ZN(n15495) );
  XNOR2_X1 U17034 ( .A(n9326), .B(n15477), .ZN(n15485) );
  XNOR2_X1 U17035 ( .A(n8425), .B(n9326), .ZN(n15496) );
  NAND2_X1 U17036 ( .A1(n15496), .A2(n15478), .ZN(n15483) );
  AOI22_X1 U17037 ( .A1(n12704), .A2(n15481), .B1(n15480), .B2(n15479), .ZN(
        n15482) );
  OAI211_X1 U17038 ( .C1(n15485), .C2(n15484), .A(n15483), .B(n15482), .ZN(
        n15494) );
  AOI21_X1 U17039 ( .B1(n15495), .B2(n15486), .A(n15494), .ZN(n15492) );
  INV_X1 U17040 ( .A(n15487), .ZN(n15489) );
  AOI22_X1 U17041 ( .A1(n15489), .A2(n15496), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15488), .ZN(n15490) );
  OAI221_X1 U17042 ( .B1(n15493), .B2(n15492), .C1(n15472), .C2(n15491), .A(
        n15490), .ZN(P3_U3232) );
  AOI211_X1 U17043 ( .C1(n15504), .C2(n15496), .A(n15495), .B(n15494), .ZN(
        n15511) );
  INV_X1 U17044 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U17045 ( .A1(n15510), .A2(n15511), .B1(n15497), .B2(n15509), .ZN(
        P3_U3393) );
  AOI211_X1 U17046 ( .C1(n15501), .C2(n15500), .A(n15499), .B(n15498), .ZN(
        n15512) );
  INV_X1 U17047 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U17048 ( .A1(n15510), .A2(n15512), .B1(n15502), .B2(n15509), .ZN(
        P3_U3396) );
  INV_X1 U17049 ( .A(n15503), .ZN(n15507) );
  AND2_X1 U17050 ( .A1(n15505), .A2(n15504), .ZN(n15506) );
  NOR3_X1 U17051 ( .A1(n15508), .A2(n15507), .A3(n15506), .ZN(n15513) );
  AOI22_X1 U17052 ( .A1(n15510), .A2(n15513), .B1(n8017), .B2(n15509), .ZN(
        P3_U3414) );
  AOI22_X1 U17053 ( .A1(n15514), .A2(n15511), .B1(n7907), .B2(n9433), .ZN(
        P3_U3460) );
  AOI22_X1 U17054 ( .A1(n15514), .A2(n15512), .B1(n10329), .B2(n9433), .ZN(
        P3_U3461) );
  AOI22_X1 U17055 ( .A1(n15514), .A2(n15513), .B1(n8020), .B2(n9433), .ZN(
        P3_U3467) );
  NAND2_X1 U17056 ( .A1(n15515), .A2(P2_D_REG_30__SCAN_IN), .ZN(n15663) );
  NAND4_X1 U17057 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(n15630), .A3(n15516), 
        .A4(n15631), .ZN(n15517) );
  NOR3_X1 U17058 ( .A1(n15518), .A2(P1_IR_REG_6__SCAN_IN), .A3(n15517), .ZN(
        n15519) );
  NAND3_X1 U17059 ( .A1(n15519), .A2(P3_IR_REG_29__SCAN_IN), .A3(n15628), .ZN(
        n15523) );
  NAND4_X1 U17060 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), 
        .A3(n15641), .A4(n15640), .ZN(n15522) );
  NAND4_X1 U17061 ( .A1(n15647), .A2(n15520), .A3(n15646), .A4(
        P1_REG1_REG_23__SCAN_IN), .ZN(n15521) );
  NOR3_X1 U17062 ( .A1(n15523), .A2(n15522), .A3(n15521), .ZN(n15661) );
  NAND4_X1 U17063 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), 
        .A3(P2_REG3_REG_7__SCAN_IN), .A4(n9754), .ZN(n15526) );
  NAND4_X1 U17064 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P3_REG1_REG_13__SCAN_IN), 
        .A3(P1_ADDR_REG_15__SCAN_IN), .A4(n15552), .ZN(n15525) );
  NAND3_X1 U17065 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P3_DATAO_REG_9__SCAN_IN), 
        .A3(n10076), .ZN(n15524) );
  NOR4_X1 U17066 ( .A1(P3_D_REG_31__SCAN_IN), .A2(n15526), .A3(n15525), .A4(
        n15524), .ZN(n15546) );
  NAND4_X1 U17067 ( .A1(n15528), .A2(n15527), .A3(n15617), .A4(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n15538) );
  INV_X1 U17068 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15643) );
  AND4_X1 U17069 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .A3(P1_REG3_REG_21__SCAN_IN), .A4(P1_ADDR_REG_16__SCAN_IN), .ZN(n15536) );
  INV_X1 U17070 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15529) );
  NOR4_X1 U17071 ( .A1(P3_REG2_REG_20__SCAN_IN), .A2(SI_12_), .A3(n15529), 
        .A4(n15593), .ZN(n15535) );
  NOR4_X1 U17072 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P3_REG1_REG_7__SCAN_IN), 
        .A3(P1_IR_REG_14__SCAN_IN), .A4(n15530), .ZN(n15534) );
  NOR4_X1 U17073 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .A3(n15532), .A4(n15531), .ZN(n15533) );
  NAND4_X1 U17074 ( .A1(n15536), .A2(n15535), .A3(n15534), .A4(n15533), .ZN(
        n15537) );
  NOR4_X1 U17075 ( .A1(n15538), .A2(n15643), .A3(P2_DATAO_REG_0__SCAN_IN), 
        .A4(n15537), .ZN(n15544) );
  NOR4_X1 U17076 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(n15539), .A3(n15563), .A4(
        n15565), .ZN(n15542) );
  NOR4_X1 U17077 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(P3_REG1_REG_20__SCAN_IN), 
        .A3(n15575), .A4(n15578), .ZN(n15541) );
  NOR3_X1 U17078 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_REG3_REG_26__SCAN_IN), 
        .A3(P3_REG1_REG_0__SCAN_IN), .ZN(n15540) );
  AND4_X1 U17079 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15542), .A3(n15541), .A4(
        n15540), .ZN(n15543) );
  AND4_X1 U17080 ( .A1(n15546), .A2(n15545), .A3(n15544), .A4(n15543), .ZN(
        n15660) );
  AOI22_X1 U17081 ( .A1(n15549), .A2(keyinput10), .B1(n15548), .B2(keyinput1), 
        .ZN(n15547) );
  OAI221_X1 U17082 ( .B1(n15549), .B2(keyinput10), .C1(n15548), .C2(keyinput1), 
        .A(n15547), .ZN(n15560) );
  AOI22_X1 U17083 ( .A1(n15552), .A2(keyinput51), .B1(keyinput44), .B2(n15551), 
        .ZN(n15550) );
  OAI221_X1 U17084 ( .B1(n15552), .B2(keyinput51), .C1(n15551), .C2(keyinput44), .A(n15550), .ZN(n15559) );
  AOI22_X1 U17085 ( .A1(n9754), .A2(keyinput2), .B1(n15554), .B2(keyinput29), 
        .ZN(n15553) );
  OAI221_X1 U17086 ( .B1(n9754), .B2(keyinput2), .C1(n15554), .C2(keyinput29), 
        .A(n15553), .ZN(n15558) );
  XNOR2_X1 U17087 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput0), .ZN(n15556) );
  XNOR2_X1 U17088 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput46), .ZN(n15555) );
  NAND2_X1 U17089 ( .A1(n15556), .A2(n15555), .ZN(n15557) );
  NOR4_X1 U17090 ( .A1(n15560), .A2(n15559), .A3(n15558), .A4(n15557), .ZN(
        n15604) );
  AOI22_X1 U17091 ( .A1(n15563), .A2(keyinput13), .B1(keyinput15), .B2(n15562), 
        .ZN(n15561) );
  OAI221_X1 U17092 ( .B1(n15563), .B2(keyinput13), .C1(n15562), .C2(keyinput15), .A(n15561), .ZN(n15573) );
  AOI22_X1 U17093 ( .A1(n10076), .A2(keyinput23), .B1(keyinput8), .B2(n15565), 
        .ZN(n15564) );
  OAI221_X1 U17094 ( .B1(n10076), .B2(keyinput23), .C1(n15565), .C2(keyinput8), 
        .A(n15564), .ZN(n15572) );
  AOI22_X1 U17095 ( .A1(n15567), .A2(keyinput34), .B1(n7039), .B2(keyinput27), 
        .ZN(n15566) );
  OAI221_X1 U17096 ( .B1(n15567), .B2(keyinput34), .C1(n7039), .C2(keyinput27), 
        .A(n15566), .ZN(n15571) );
  XNOR2_X1 U17097 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput57), .ZN(n15569) );
  XNOR2_X1 U17098 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput28), .ZN(n15568)
         );
  NAND2_X1 U17099 ( .A1(n15569), .A2(n15568), .ZN(n15570) );
  NOR4_X1 U17100 ( .A1(n15573), .A2(n15572), .A3(n15571), .A4(n15570), .ZN(
        n15603) );
  AOI22_X1 U17101 ( .A1(n15576), .A2(keyinput49), .B1(n15575), .B2(keyinput35), 
        .ZN(n15574) );
  OAI221_X1 U17102 ( .B1(n15576), .B2(keyinput49), .C1(n15575), .C2(keyinput35), .A(n15574), .ZN(n15588) );
  AOI22_X1 U17103 ( .A1(n15579), .A2(keyinput22), .B1(keyinput4), .B2(n15578), 
        .ZN(n15577) );
  OAI221_X1 U17104 ( .B1(n15579), .B2(keyinput22), .C1(n15578), .C2(keyinput4), 
        .A(n15577), .ZN(n15587) );
  INV_X1 U17105 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15582) );
  AOI22_X1 U17106 ( .A1(n15582), .A2(keyinput39), .B1(n15581), .B2(keyinput43), 
        .ZN(n15580) );
  OAI221_X1 U17107 ( .B1(n15582), .B2(keyinput39), .C1(n15581), .C2(keyinput43), .A(n15580), .ZN(n15586) );
  AOI22_X1 U17108 ( .A1(n15584), .A2(keyinput31), .B1(keyinput6), .B2(n9566), 
        .ZN(n15583) );
  OAI221_X1 U17109 ( .B1(n15584), .B2(keyinput31), .C1(n9566), .C2(keyinput6), 
        .A(n15583), .ZN(n15585) );
  NOR4_X1 U17110 ( .A1(n15588), .A2(n15587), .A3(n15586), .A4(n15585), .ZN(
        n15602) );
  INV_X1 U17111 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15590) );
  AOI22_X1 U17112 ( .A1(n6700), .A2(keyinput37), .B1(keyinput24), .B2(n15590), 
        .ZN(n15589) );
  OAI221_X1 U17113 ( .B1(n6700), .B2(keyinput37), .C1(n15590), .C2(keyinput24), 
        .A(n15589), .ZN(n15600) );
  AOI22_X1 U17114 ( .A1(n15593), .A2(keyinput59), .B1(n15592), .B2(keyinput3), 
        .ZN(n15591) );
  OAI221_X1 U17115 ( .B1(n15593), .B2(keyinput59), .C1(n15592), .C2(keyinput3), 
        .A(n15591), .ZN(n15599) );
  XOR2_X1 U17116 ( .A(n12707), .B(keyinput16), .Z(n15597) );
  XNOR2_X1 U17117 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput21), .ZN(n15596) );
  XNOR2_X1 U17118 ( .A(P3_REG1_REG_0__SCAN_IN), .B(keyinput20), .ZN(n15595) );
  XNOR2_X1 U17119 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput33), .ZN(n15594) );
  NAND4_X1 U17120 ( .A1(n15597), .A2(n15596), .A3(n15595), .A4(n15594), .ZN(
        n15598) );
  NOR3_X1 U17121 ( .A1(n15600), .A2(n15599), .A3(n15598), .ZN(n15601) );
  NAND4_X1 U17122 ( .A1(n15604), .A2(n15603), .A3(n15602), .A4(n15601), .ZN(
        n15659) );
  AOI22_X1 U17123 ( .A1(n15606), .A2(keyinput61), .B1(keyinput53), .B2(n8983), 
        .ZN(n15605) );
  OAI221_X1 U17124 ( .B1(n15606), .B2(keyinput61), .C1(n8983), .C2(keyinput53), 
        .A(n15605), .ZN(n15615) );
  AOI22_X1 U17125 ( .A1(n8002), .A2(keyinput12), .B1(n15608), .B2(keyinput47), 
        .ZN(n15607) );
  OAI221_X1 U17126 ( .B1(n8002), .B2(keyinput12), .C1(n15608), .C2(keyinput47), 
        .A(n15607), .ZN(n15614) );
  XNOR2_X1 U17127 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput41), .ZN(n15612) );
  XNOR2_X1 U17128 ( .A(P2_REG1_REG_27__SCAN_IN), .B(keyinput32), .ZN(n15611)
         );
  XNOR2_X1 U17129 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(keyinput45), .ZN(n15610)
         );
  XNOR2_X1 U17130 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput50), .ZN(n15609) );
  NAND4_X1 U17131 ( .A1(n15612), .A2(n15611), .A3(n15610), .A4(n15609), .ZN(
        n15613) );
  NOR3_X1 U17132 ( .A1(n15615), .A2(n15614), .A3(n15613), .ZN(n15657) );
  AOI22_X1 U17133 ( .A1(n15528), .A2(keyinput7), .B1(n15617), .B2(keyinput36), 
        .ZN(n15616) );
  OAI221_X1 U17134 ( .B1(n15528), .B2(keyinput7), .C1(n15617), .C2(keyinput36), 
        .A(n15616), .ZN(n15626) );
  XOR2_X1 U17135 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput5), .Z(n15625) );
  XNOR2_X1 U17136 ( .A(n15618), .B(keyinput54), .ZN(n15624) );
  XNOR2_X1 U17137 ( .A(P1_REG0_REG_31__SCAN_IN), .B(keyinput17), .ZN(n15622)
         );
  XNOR2_X1 U17138 ( .A(SI_12_), .B(keyinput40), .ZN(n15621) );
  XNOR2_X1 U17139 ( .A(P2_REG1_REG_16__SCAN_IN), .B(keyinput62), .ZN(n15620)
         );
  XNOR2_X1 U17140 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput9), .ZN(n15619) );
  NAND4_X1 U17141 ( .A1(n15622), .A2(n15621), .A3(n15620), .A4(n15619), .ZN(
        n15623) );
  NOR4_X1 U17142 ( .A1(n15626), .A2(n15625), .A3(n15624), .A4(n15623), .ZN(
        n15656) );
  AOI22_X1 U17143 ( .A1(n7893), .A2(keyinput38), .B1(keyinput56), .B2(n15628), 
        .ZN(n15627) );
  OAI221_X1 U17144 ( .B1(n7893), .B2(keyinput38), .C1(n15628), .C2(keyinput56), 
        .A(n15627), .ZN(n15638) );
  AOI22_X1 U17145 ( .A1(n15631), .A2(keyinput19), .B1(n15630), .B2(keyinput52), 
        .ZN(n15629) );
  OAI221_X1 U17146 ( .B1(n15631), .B2(keyinput19), .C1(n15630), .C2(keyinput52), .A(n15629), .ZN(n15637) );
  XOR2_X1 U17147 ( .A(n15518), .B(keyinput14), .Z(n15635) );
  XNOR2_X1 U17148 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput55), .ZN(n15634) );
  XNOR2_X1 U17149 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput18), .ZN(n15633)
         );
  XNOR2_X1 U17150 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput25), .ZN(n15632) );
  NAND4_X1 U17151 ( .A1(n15635), .A2(n15634), .A3(n15633), .A4(n15632), .ZN(
        n15636) );
  NOR3_X1 U17152 ( .A1(n15638), .A2(n15637), .A3(n15636), .ZN(n15655) );
  AOI22_X1 U17153 ( .A1(n15641), .A2(keyinput30), .B1(keyinput48), .B2(n15640), 
        .ZN(n15639) );
  OAI221_X1 U17154 ( .B1(n15641), .B2(keyinput30), .C1(n15640), .C2(keyinput48), .A(n15639), .ZN(n15653) );
  AOI22_X1 U17155 ( .A1(n15644), .A2(keyinput26), .B1(keyinput60), .B2(n15643), 
        .ZN(n15642) );
  OAI221_X1 U17156 ( .B1(n15644), .B2(keyinput26), .C1(n15643), .C2(keyinput60), .A(n15642), .ZN(n15652) );
  AOI22_X1 U17157 ( .A1(n15647), .A2(keyinput11), .B1(keyinput63), .B2(n15646), 
        .ZN(n15645) );
  OAI221_X1 U17158 ( .B1(n15647), .B2(keyinput11), .C1(n15646), .C2(keyinput63), .A(n15645), .ZN(n15651) );
  XNOR2_X1 U17159 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput42), .ZN(n15649) );
  XNOR2_X1 U17160 ( .A(P1_REG1_REG_23__SCAN_IN), .B(keyinput58), .ZN(n15648)
         );
  NAND2_X1 U17161 ( .A1(n15649), .A2(n15648), .ZN(n15650) );
  NOR4_X1 U17162 ( .A1(n15653), .A2(n15652), .A3(n15651), .A4(n15650), .ZN(
        n15654) );
  NAND4_X1 U17163 ( .A1(n15657), .A2(n15656), .A3(n15655), .A4(n15654), .ZN(
        n15658) );
  AOI211_X1 U17164 ( .C1(n15661), .C2(n15660), .A(n15659), .B(n15658), .ZN(
        n15662) );
  XNOR2_X1 U17165 ( .A(n15663), .B(n15662), .ZN(P2_U3267) );
  AND2_X1 U17166 ( .A1(n15665), .A2(n15664), .ZN(n15666) );
  XOR2_X1 U17167 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15666), .Z(SUB_1596_U60) );
  AOI21_X1 U17168 ( .B1(n15669), .B2(n15668), .A(n15667), .ZN(SUB_1596_U5) );
  NAND2_X1 U9792 ( .A1(n7895), .A2(n12933), .ZN(n7960) );
  OR2_X2 U10017 ( .A1(n7895), .A2(n7896), .ZN(n8390) );
  NAND4_X2 U10401 ( .A1(n7911), .A2(n7910), .A3(n7909), .A4(n7908), .ZN(n12461) );
  INV_X1 U7554 ( .A(n7982), .ZN(n8355) );
  XNOR2_X1 U10381 ( .A(n7894), .B(n7893), .ZN(n12933) );
  INV_X2 U7159 ( .A(n10286), .ZN(n14020) );
  NAND2_X1 U7161 ( .A1(n7918), .A2(n7434), .ZN(n8382) );
  CLKBUF_X1 U7173 ( .A(n12293), .Z(n6610) );
  CLKBUF_X2 U7186 ( .A(n8382), .Z(n6612) );
  CLKBUF_X2 U7194 ( .A(n9536), .Z(n13091) );
  INV_X1 U7205 ( .A(n12203), .ZN(n8633) );
  CLKBUF_X1 U7260 ( .A(n8794), .Z(n14453) );
  NAND2_X1 U7264 ( .A1(n7358), .A2(n7356), .ZN(n14872) );
  CLKBUF_X1 U7354 ( .A(n13126), .Z(n6405) );
  CLKBUF_X1 U7377 ( .A(n15292), .Z(n6407) );
  CLKBUF_X1 U7828 ( .A(n13325), .Z(n6398) );
endmodule

